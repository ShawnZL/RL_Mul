// Benchmark "top" written by ABC on Mon Dec 25 17:56:10 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1922, new_n1923, new_n1924,
    new_n1925, new_n1926, new_n1927, new_n1928, new_n1929, new_n1930,
    new_n1931, new_n1932, new_n1933, new_n1934, new_n1935, new_n1936,
    new_n1937, new_n1938, new_n1939, new_n1940, new_n1941, new_n1942,
    new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948,
    new_n1949, new_n1950, new_n1951, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972,
    new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978,
    new_n1979, new_n1980, new_n1981, new_n1982, new_n1983, new_n1984,
    new_n1985, new_n1986, new_n1987, new_n1988, new_n1989, new_n1990,
    new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996,
    new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2002,
    new_n2003, new_n2004, new_n2005, new_n2006, new_n2007, new_n2008,
    new_n2009, new_n2010, new_n2011, new_n2012, new_n2013, new_n2014,
    new_n2015, new_n2016, new_n2017, new_n2018, new_n2019, new_n2020,
    new_n2021, new_n2022, new_n2023, new_n2024, new_n2025, new_n2026,
    new_n2027, new_n2028, new_n2029, new_n2030, new_n2031, new_n2032,
    new_n2033, new_n2034, new_n2035, new_n2036, new_n2037, new_n2038,
    new_n2039, new_n2040, new_n2041, new_n2042, new_n2043, new_n2044,
    new_n2045, new_n2046, new_n2047, new_n2048, new_n2049, new_n2050,
    new_n2051, new_n2052, new_n2053, new_n2054, new_n2055, new_n2056,
    new_n2057, new_n2058, new_n2059, new_n2060, new_n2061, new_n2062,
    new_n2063, new_n2064, new_n2065, new_n2066, new_n2067, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087,
    new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093,
    new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099,
    new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105,
    new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111,
    new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117,
    new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123,
    new_n2124, new_n2125, new_n2126, new_n2127, new_n2128, new_n2129,
    new_n2130, new_n2131, new_n2132, new_n2133, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141,
    new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2160, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165,
    new_n2166, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171,
    new_n2172, new_n2173, new_n2174, new_n2175, new_n2176, new_n2177,
    new_n2178, new_n2179, new_n2180, new_n2181, new_n2182, new_n2183,
    new_n2184, new_n2185, new_n2186, new_n2187, new_n2188, new_n2189,
    new_n2190, new_n2191, new_n2192, new_n2193, new_n2194, new_n2195,
    new_n2196, new_n2197, new_n2198, new_n2199, new_n2200, new_n2201,
    new_n2202, new_n2203, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431,
    new_n2432, new_n2433, new_n2434, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479,
    new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485,
    new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491,
    new_n2492, new_n2493, new_n2494, new_n2495, new_n2496, new_n2497,
    new_n2498, new_n2499, new_n2500, new_n2501, new_n2502, new_n2503,
    new_n2504, new_n2505, new_n2506, new_n2507, new_n2508, new_n2509,
    new_n2510, new_n2511, new_n2512, new_n2513, new_n2514, new_n2515,
    new_n2516, new_n2517, new_n2518, new_n2519, new_n2520, new_n2521,
    new_n2522, new_n2523, new_n2524, new_n2525, new_n2526, new_n2527,
    new_n2528, new_n2529, new_n2530, new_n2531, new_n2532, new_n2533,
    new_n2534, new_n2535, new_n2536, new_n2537, new_n2538, new_n2539,
    new_n2540, new_n2541, new_n2542, new_n2543, new_n2544, new_n2545,
    new_n2546, new_n2547, new_n2548, new_n2549, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2830, new_n2831, new_n2832, new_n2833, new_n2834, new_n2835,
    new_n2836, new_n2837, new_n2838, new_n2839, new_n2840, new_n2841,
    new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847,
    new_n2848, new_n2849, new_n2850, new_n2851, new_n2852, new_n2853,
    new_n2854, new_n2855, new_n2856, new_n2857, new_n2858, new_n2859,
    new_n2860, new_n2861, new_n2862, new_n2863, new_n2864, new_n2865,
    new_n2866, new_n2867, new_n2868, new_n2869, new_n2870, new_n2871,
    new_n2872, new_n2873, new_n2874, new_n2875, new_n2876, new_n2877,
    new_n2878, new_n2879, new_n2880, new_n2881, new_n2882, new_n2883,
    new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889,
    new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2896, new_n2897, new_n2898, new_n2899, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3095,
    new_n3096, new_n3097, new_n3098, new_n3099, new_n3100, new_n3101,
    new_n3102, new_n3103, new_n3104, new_n3105, new_n3106, new_n3107,
    new_n3108, new_n3109, new_n3110, new_n3111, new_n3112, new_n3113,
    new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239,
    new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269,
    new_n3270, new_n3271, new_n3272, new_n3273, new_n3274, new_n3275,
    new_n3276, new_n3277, new_n3278, new_n3279, new_n3280, new_n3281,
    new_n3282, new_n3283, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502, new_n3503, new_n3504, new_n3505,
    new_n3506, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528, new_n3529,
    new_n3530, new_n3531, new_n3532, new_n3533, new_n3534, new_n3535,
    new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541,
    new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547,
    new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553,
    new_n3554, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561, new_n3562, new_n3563, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595,
    new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601,
    new_n3602, new_n3603, new_n3604, new_n3605, new_n3606, new_n3607,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3615, new_n3616, new_n3617, new_n3618, new_n3619,
    new_n3620, new_n3621, new_n3622, new_n3623, new_n3624, new_n3625,
    new_n3626, new_n3627, new_n3628, new_n3629, new_n3630, new_n3631,
    new_n3632, new_n3633, new_n3634, new_n3635, new_n3636, new_n3637,
    new_n3638, new_n3639, new_n3640, new_n3641, new_n3642, new_n3643,
    new_n3644, new_n3645, new_n3646, new_n3647, new_n3648, new_n3649,
    new_n3650, new_n3651, new_n3652, new_n3653, new_n3654, new_n3655,
    new_n3656, new_n3657, new_n3658, new_n3659, new_n3660, new_n3661,
    new_n3662, new_n3663, new_n3664, new_n3665, new_n3666, new_n3667,
    new_n3668, new_n3669, new_n3670, new_n3671, new_n3672, new_n3673,
    new_n3674, new_n3675, new_n3676, new_n3677, new_n3678, new_n3679,
    new_n3680, new_n3681, new_n3682, new_n3683, new_n3684, new_n3685,
    new_n3686, new_n3687, new_n3688, new_n3689, new_n3690, new_n3691,
    new_n3692, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869, new_n3870, new_n3871, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909, new_n3910, new_n3911, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085, new_n4086, new_n4087, new_n4088, new_n4089,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300,
    new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306,
    new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312,
    new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318,
    new_n4319, new_n4320, new_n4321, new_n4322, new_n4323, new_n4324,
    new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330,
    new_n4331, new_n4332, new_n4333, new_n4334, new_n4335, new_n4336,
    new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342,
    new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873,
    new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879,
    new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915,
    new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921,
    new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927,
    new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4959, new_n4960, new_n4961, new_n4962, new_n4963,
    new_n4964, new_n4965, new_n4966, new_n4967, new_n4968, new_n4969,
    new_n4970, new_n4971, new_n4972, new_n4973, new_n4974, new_n4975,
    new_n4976, new_n4977, new_n4978, new_n4979, new_n4980, new_n4981,
    new_n4982, new_n4983, new_n4984, new_n4985, new_n4986, new_n4987,
    new_n4988, new_n4989, new_n4990, new_n4991, new_n4992, new_n4993,
    new_n4994, new_n4995, new_n4996, new_n4997, new_n4998, new_n4999,
    new_n5000, new_n5001, new_n5002, new_n5003, new_n5004, new_n5005,
    new_n5006, new_n5007, new_n5008, new_n5009, new_n5010, new_n5011,
    new_n5012, new_n5013, new_n5014, new_n5015, new_n5016, new_n5017,
    new_n5018, new_n5019, new_n5020, new_n5021, new_n5022, new_n5023,
    new_n5024, new_n5025, new_n5026, new_n5027, new_n5028, new_n5029,
    new_n5030, new_n5031, new_n5032, new_n5033, new_n5034, new_n5035,
    new_n5036, new_n5037, new_n5038, new_n5039, new_n5040, new_n5041,
    new_n5042, new_n5043, new_n5044, new_n5045, new_n5046, new_n5047,
    new_n5048, new_n5049, new_n5050, new_n5051, new_n5052, new_n5053,
    new_n5054, new_n5055, new_n5056, new_n5057, new_n5058, new_n5059,
    new_n5060, new_n5061, new_n5062, new_n5063, new_n5064, new_n5065,
    new_n5066, new_n5067, new_n5068, new_n5069, new_n5070, new_n5071,
    new_n5072, new_n5073, new_n5074, new_n5075, new_n5076, new_n5077,
    new_n5078, new_n5079, new_n5080, new_n5081, new_n5082, new_n5083,
    new_n5084, new_n5085, new_n5086, new_n5087, new_n5088, new_n5089,
    new_n5090, new_n5091, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162,
    new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168,
    new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174,
    new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180,
    new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189, new_n5190, new_n5191, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198,
    new_n5199, new_n5200, new_n5201, new_n5202, new_n5203, new_n5204,
    new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225, new_n5226, new_n5227, new_n5228,
    new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234,
    new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240,
    new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246,
    new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252,
    new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258,
    new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264,
    new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270,
    new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276,
    new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282,
    new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288,
    new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294,
    new_n5295, new_n5296, new_n5297, new_n5298, new_n5299, new_n5300,
    new_n5301, new_n5302, new_n5303, new_n5304, new_n5305, new_n5306,
    new_n5307, new_n5308, new_n5309, new_n5310, new_n5311, new_n5312,
    new_n5313, new_n5314, new_n5315, new_n5316, new_n5317, new_n5318,
    new_n5319, new_n5320, new_n5321, new_n5322, new_n5323, new_n5324,
    new_n5325, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330,
    new_n5331, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499,
    new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505,
    new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511,
    new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548, new_n5549, new_n5550, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5881, new_n5882, new_n5883, new_n5884, new_n5885,
    new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903,
    new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565,
    new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571,
    new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577,
    new_n6578, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583,
    new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589,
    new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611, new_n6612, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628, new_n6629, new_n6630, new_n6631,
    new_n6632, new_n6633, new_n6634, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652, new_n6653, new_n6654, new_n6655,
    new_n6656, new_n6657, new_n6658, new_n6659, new_n6660, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668, new_n6669, new_n6670, new_n6671, new_n6672, new_n6673,
    new_n6674, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679,
    new_n6680, new_n6681, new_n6682, new_n6683, new_n6684, new_n6685,
    new_n6686, new_n6687, new_n6688, new_n6689, new_n6690, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706, new_n6707, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746,
    new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752,
    new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758,
    new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764,
    new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773, new_n6774, new_n6775, new_n6776,
    new_n6777, new_n6778, new_n6779, new_n6780, new_n6781, new_n6782,
    new_n6783, new_n6784, new_n6785, new_n6786, new_n6787, new_n6788,
    new_n6789, new_n6790, new_n6791, new_n6792, new_n6793, new_n6794,
    new_n6795, new_n6796, new_n6797, new_n6798, new_n6799, new_n6800,
    new_n6801, new_n6802, new_n6803, new_n6804, new_n6805, new_n6806,
    new_n6807, new_n6808, new_n6809, new_n6810, new_n6811, new_n6812,
    new_n6813, new_n6814, new_n6815, new_n6816, new_n6817, new_n6818,
    new_n6819, new_n6820, new_n6821, new_n6822, new_n6823, new_n6824,
    new_n6825, new_n6826, new_n6827, new_n6828, new_n6829, new_n6830,
    new_n6831, new_n6832, new_n6833, new_n6834, new_n6835, new_n6836,
    new_n6837, new_n6838, new_n6839, new_n6840, new_n6841, new_n6842,
    new_n6843, new_n6844, new_n6845, new_n6846, new_n6847, new_n6848,
    new_n6849, new_n6850, new_n6851, new_n6852, new_n6853, new_n6854,
    new_n6855, new_n6856, new_n6857, new_n6858, new_n6859, new_n6860,
    new_n6861, new_n6862, new_n6863, new_n6864, new_n6865, new_n6866,
    new_n6867, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872,
    new_n6873, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878,
    new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884,
    new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890,
    new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896,
    new_n6897, new_n6898, new_n6899, new_n6900, new_n6901, new_n6902,
    new_n6903, new_n6904, new_n6905, new_n6906, new_n6907, new_n6908,
    new_n6909, new_n6910, new_n6911, new_n6912, new_n6913, new_n6914,
    new_n6915, new_n6916, new_n6917, new_n6918, new_n6919, new_n6920,
    new_n6921, new_n6922, new_n6923, new_n6924, new_n6925, new_n6926,
    new_n6927, new_n6928, new_n6929, new_n6930, new_n6931, new_n6932,
    new_n6933, new_n6934, new_n6935, new_n6936, new_n6937, new_n6938,
    new_n6939, new_n6940, new_n6941, new_n6942, new_n6943, new_n6944,
    new_n6945, new_n6946, new_n6947, new_n6948, new_n6949, new_n6950,
    new_n6951, new_n6952, new_n6953, new_n6954, new_n6955, new_n6956,
    new_n6957, new_n6958, new_n6959, new_n6960, new_n6961, new_n6962,
    new_n6963, new_n6964, new_n6965, new_n6966, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7266, new_n7267, new_n7268, new_n7269, new_n7270,
    new_n7271, new_n7272, new_n7273, new_n7274, new_n7275, new_n7276,
    new_n7277, new_n7278, new_n7279, new_n7280, new_n7281, new_n7282,
    new_n7283, new_n7284, new_n7285, new_n7286, new_n7287, new_n7288,
    new_n7289, new_n7290, new_n7291, new_n7292, new_n7293, new_n7294,
    new_n7295, new_n7296, new_n7297, new_n7298, new_n7299, new_n7300,
    new_n7301, new_n7302, new_n7303, new_n7304, new_n7305, new_n7306,
    new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312,
    new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318,
    new_n7319, new_n7320, new_n7321, new_n7322, new_n7323, new_n7324,
    new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330,
    new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336,
    new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342,
    new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348,
    new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354,
    new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414,
    new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420,
    new_n7421, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426,
    new_n7427, new_n7428, new_n7429, new_n7430, new_n7431, new_n7432,
    new_n7433, new_n7434, new_n7435, new_n7436, new_n7437, new_n7438,
    new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730, new_n7731, new_n7732, new_n7733,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8148, new_n8149,
    new_n8150, new_n8151, new_n8152, new_n8153, new_n8154, new_n8155,
    new_n8156, new_n8157, new_n8158, new_n8159, new_n8160, new_n8161,
    new_n8162, new_n8163, new_n8164, new_n8165, new_n8166, new_n8167,
    new_n8168, new_n8169, new_n8170, new_n8171, new_n8172, new_n8173,
    new_n8174, new_n8175, new_n8176, new_n8177, new_n8178, new_n8179,
    new_n8180, new_n8181, new_n8182, new_n8183, new_n8184, new_n8185,
    new_n8186, new_n8187, new_n8188, new_n8189, new_n8190, new_n8191,
    new_n8192, new_n8193, new_n8194, new_n8195, new_n8196, new_n8197,
    new_n8198, new_n8199, new_n8200, new_n8201, new_n8202, new_n8203,
    new_n8204, new_n8205, new_n8206, new_n8207, new_n8208, new_n8209,
    new_n8210, new_n8211, new_n8212, new_n8213, new_n8214, new_n8215,
    new_n8216, new_n8217, new_n8218, new_n8219, new_n8220, new_n8221,
    new_n8222, new_n8223, new_n8224, new_n8225, new_n8226, new_n8227,
    new_n8228, new_n8229, new_n8230, new_n8231, new_n8232, new_n8233,
    new_n8234, new_n8235, new_n8236, new_n8237, new_n8238, new_n8239,
    new_n8240, new_n8241, new_n8242, new_n8243, new_n8244, new_n8245,
    new_n8246, new_n8247, new_n8248, new_n8249, new_n8250, new_n8251,
    new_n8252, new_n8253, new_n8254, new_n8255, new_n8256, new_n8257,
    new_n8258, new_n8259, new_n8260, new_n8261, new_n8262, new_n8263,
    new_n8264, new_n8265, new_n8266, new_n8267, new_n8268, new_n8269,
    new_n8270, new_n8271, new_n8272, new_n8273, new_n8274, new_n8275,
    new_n8276, new_n8277, new_n8278, new_n8279, new_n8280, new_n8281,
    new_n8282, new_n8283, new_n8284, new_n8285, new_n8286, new_n8287,
    new_n8288, new_n8289, new_n8290, new_n8291, new_n8292, new_n8293,
    new_n8294, new_n8295, new_n8296, new_n8297, new_n8298, new_n8299,
    new_n8300, new_n8301, new_n8302, new_n8303, new_n8304, new_n8305,
    new_n8306, new_n8307, new_n8308, new_n8309, new_n8310, new_n8311,
    new_n8312, new_n8313, new_n8314, new_n8315, new_n8316, new_n8317,
    new_n8318, new_n8319, new_n8320, new_n8321, new_n8322, new_n8323,
    new_n8324, new_n8325, new_n8326, new_n8327, new_n8328, new_n8329,
    new_n8330, new_n8331, new_n8332, new_n8333, new_n8334, new_n8335,
    new_n8336, new_n8337, new_n8338, new_n8339, new_n8340, new_n8341,
    new_n8342, new_n8343, new_n8344, new_n8345, new_n8346, new_n8347,
    new_n8348, new_n8349, new_n8350, new_n8351, new_n8352, new_n8353,
    new_n8354, new_n8355, new_n8356, new_n8357, new_n8358, new_n8359,
    new_n8360, new_n8361, new_n8362, new_n8363, new_n8364, new_n8365,
    new_n8366, new_n8367, new_n8368, new_n8369, new_n8370, new_n8371,
    new_n8372, new_n8373, new_n8374, new_n8375, new_n8376, new_n8377,
    new_n8378, new_n8379, new_n8380, new_n8381, new_n8382, new_n8383,
    new_n8384, new_n8385, new_n8386, new_n8387, new_n8388, new_n8389,
    new_n8390, new_n8391, new_n8392, new_n8393, new_n8394, new_n8395,
    new_n8396, new_n8397, new_n8398, new_n8399, new_n8400, new_n8401,
    new_n8402, new_n8403, new_n8404, new_n8405, new_n8406, new_n8407,
    new_n8408, new_n8409, new_n8410, new_n8411, new_n8412, new_n8413,
    new_n8414, new_n8415, new_n8416, new_n8417, new_n8418, new_n8419,
    new_n8420, new_n8421, new_n8422, new_n8423, new_n8424, new_n8425,
    new_n8426, new_n8427, new_n8428, new_n8429, new_n8430, new_n8431,
    new_n8432, new_n8433, new_n8434, new_n8435, new_n8436, new_n8437,
    new_n8438, new_n8439, new_n8440, new_n8441, new_n8442, new_n8443,
    new_n8444, new_n8445, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8777, new_n8778, new_n8779, new_n8780, new_n8781,
    new_n8782, new_n8783, new_n8784, new_n8785, new_n8786, new_n8787,
    new_n8788, new_n8789, new_n8790, new_n8791, new_n8792, new_n8793,
    new_n8794, new_n8795, new_n8796, new_n8797, new_n8798, new_n8799,
    new_n8800, new_n8801, new_n8802, new_n8803, new_n8804, new_n8805,
    new_n8806, new_n8807, new_n8808, new_n8809, new_n8810, new_n8811,
    new_n8812, new_n8813, new_n8814, new_n8815, new_n8816, new_n8817,
    new_n8818, new_n8819, new_n8820, new_n8821, new_n8822, new_n8823,
    new_n8824, new_n8825, new_n8826, new_n8827, new_n8828, new_n8829,
    new_n8830, new_n8831, new_n8832, new_n8833, new_n8834, new_n8835,
    new_n8836, new_n8837, new_n8838, new_n8839, new_n8840, new_n8841,
    new_n8842, new_n8843, new_n8844, new_n8845, new_n8846, new_n8847,
    new_n8848, new_n8849, new_n8850, new_n8851, new_n8852, new_n8853,
    new_n8854, new_n8855, new_n8856, new_n8857, new_n8858, new_n8859,
    new_n8860, new_n8861, new_n8862, new_n8863, new_n8864, new_n8865,
    new_n8866, new_n8867, new_n8868, new_n8869, new_n8870, new_n8871,
    new_n8872, new_n8873, new_n8874, new_n8875, new_n8876, new_n8877,
    new_n8878, new_n8879, new_n8880, new_n8881, new_n8882, new_n8883,
    new_n8884, new_n8885, new_n8886, new_n8887, new_n8888, new_n8889,
    new_n8890, new_n8891, new_n8892, new_n8893, new_n8894, new_n8895,
    new_n8896, new_n8897, new_n8898, new_n8899, new_n8900, new_n8901,
    new_n8902, new_n8903, new_n8904, new_n8905, new_n8906, new_n8907,
    new_n8908, new_n8909, new_n8910, new_n8911, new_n8912, new_n8913,
    new_n8914, new_n8915, new_n8916, new_n8917, new_n8918, new_n8919,
    new_n8920, new_n8921, new_n8922, new_n8923, new_n8924, new_n8925,
    new_n8926, new_n8927, new_n8928, new_n8929, new_n8930, new_n8931,
    new_n8932, new_n8933, new_n8934, new_n8935, new_n8936, new_n8937,
    new_n8938, new_n8939, new_n8940, new_n8941, new_n8942, new_n8943,
    new_n8944, new_n8945, new_n8946, new_n8947, new_n8948, new_n8949,
    new_n8950, new_n8951, new_n8952, new_n8953, new_n8954, new_n8955,
    new_n8956, new_n8957, new_n8958, new_n8959, new_n8960, new_n8961,
    new_n8962, new_n8963, new_n8964, new_n8965, new_n8966, new_n8967,
    new_n8968, new_n8969, new_n8970, new_n8971, new_n8972, new_n8973,
    new_n8974, new_n8975, new_n8976, new_n8977, new_n8978, new_n8979,
    new_n8980, new_n8981, new_n8982, new_n8983, new_n8984, new_n8985,
    new_n8986, new_n8987, new_n8988, new_n8989, new_n8990, new_n8991,
    new_n8992, new_n8993, new_n8994, new_n8995, new_n8996, new_n8997,
    new_n8998, new_n8999, new_n9000, new_n9001, new_n9002, new_n9003,
    new_n9004, new_n9005, new_n9006, new_n9007, new_n9008, new_n9009,
    new_n9010, new_n9011, new_n9012, new_n9013, new_n9014, new_n9015,
    new_n9016, new_n9017, new_n9018, new_n9019, new_n9020, new_n9021,
    new_n9022, new_n9023, new_n9024, new_n9025, new_n9026, new_n9027,
    new_n9028, new_n9029, new_n9030, new_n9031, new_n9032, new_n9033,
    new_n9034, new_n9035, new_n9036, new_n9037, new_n9038, new_n9039,
    new_n9040, new_n9041, new_n9042, new_n9043, new_n9044, new_n9045,
    new_n9046, new_n9047, new_n9048, new_n9049, new_n9050, new_n9051,
    new_n9052, new_n9053, new_n9054, new_n9055, new_n9056, new_n9057,
    new_n9058, new_n9059, new_n9060, new_n9061, new_n9062, new_n9064,
    new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070,
    new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076,
    new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082,
    new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9088,
    new_n9089, new_n9090, new_n9091, new_n9092, new_n9093, new_n9094,
    new_n9095, new_n9096, new_n9097, new_n9098, new_n9099, new_n9100,
    new_n9101, new_n9102, new_n9103, new_n9104, new_n9105, new_n9106,
    new_n9107, new_n9108, new_n9109, new_n9110, new_n9111, new_n9112,
    new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118,
    new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124,
    new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130,
    new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136,
    new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142,
    new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148,
    new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154,
    new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160,
    new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166,
    new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172,
    new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178,
    new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184,
    new_n9185, new_n9186, new_n9187, new_n9188, new_n9189, new_n9190,
    new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202,
    new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208,
    new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214,
    new_n9215, new_n9216, new_n9217, new_n9218, new_n9219, new_n9220,
    new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226,
    new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232,
    new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262,
    new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268,
    new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274,
    new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280,
    new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286,
    new_n9287, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292,
    new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298,
    new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304,
    new_n9305, new_n9306, new_n9307, new_n9308, new_n9309, new_n9310,
    new_n9311, new_n9312, new_n9313, new_n9314, new_n9315, new_n9316,
    new_n9317, new_n9318, new_n9319, new_n9320, new_n9321, new_n9322,
    new_n9323, new_n9324, new_n9325, new_n9326, new_n9327, new_n9328,
    new_n9329, new_n9330, new_n9331, new_n9332, new_n9333, new_n9334,
    new_n9335, new_n9336, new_n9337, new_n9338, new_n9339, new_n9340,
    new_n9341, new_n9342, new_n9343, new_n9344, new_n9345, new_n9346,
    new_n9347, new_n9348, new_n9349, new_n9350, new_n9351, new_n9352,
    new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358,
    new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364,
    new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370,
    new_n9371, new_n9372, new_n9373, new_n9374, new_n9375, new_n9376,
    new_n9377, new_n9378, new_n9379, new_n9380, new_n9381, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912,
    new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9918,
    new_n9919, new_n9920, new_n9921, new_n9922, new_n9923, new_n9924,
    new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930,
    new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936,
    new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942,
    new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948,
    new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954,
    new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960,
    new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966,
    new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972,
    new_n9973, new_n9974, new_n9975, new_n9976, new_n9977, new_n9978,
    new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984,
    new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990,
    new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996,
    new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020,
    new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053, new_n10054, new_n10055, new_n10056, new_n10057,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063,
    new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069,
    new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075,
    new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081,
    new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087,
    new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093,
    new_n10094, new_n10095, new_n10096, new_n10097, new_n10098, new_n10099,
    new_n10100, new_n10101, new_n10102, new_n10103, new_n10104, new_n10105,
    new_n10106, new_n10107, new_n10108, new_n10109, new_n10110, new_n10111,
    new_n10112, new_n10113, new_n10114, new_n10115, new_n10116, new_n10117,
    new_n10118, new_n10119, new_n10120, new_n10121, new_n10122, new_n10123,
    new_n10124, new_n10125, new_n10126, new_n10127, new_n10128, new_n10129,
    new_n10130, new_n10131, new_n10132, new_n10133, new_n10134, new_n10135,
    new_n10136, new_n10137, new_n10138, new_n10139, new_n10140, new_n10141,
    new_n10142, new_n10143, new_n10144, new_n10145, new_n10146, new_n10147,
    new_n10148, new_n10149, new_n10150, new_n10151, new_n10152, new_n10153,
    new_n10154, new_n10155, new_n10156, new_n10157, new_n10158, new_n10159,
    new_n10160, new_n10161, new_n10162, new_n10163, new_n10164, new_n10165,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183,
    new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189,
    new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195,
    new_n10196, new_n10197, new_n10198, new_n10199, new_n10200, new_n10201,
    new_n10202, new_n10203, new_n10204, new_n10205, new_n10206, new_n10207,
    new_n10208, new_n10209, new_n10210, new_n10211, new_n10212, new_n10213,
    new_n10214, new_n10215, new_n10216, new_n10217, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223, new_n10224, new_n10225,
    new_n10226, new_n10227, new_n10228, new_n10229, new_n10230, new_n10231,
    new_n10232, new_n10233, new_n10234, new_n10235, new_n10236, new_n10237,
    new_n10238, new_n10239, new_n10240, new_n10241, new_n10242, new_n10243,
    new_n10244, new_n10245, new_n10246, new_n10247, new_n10248, new_n10249,
    new_n10250, new_n10251, new_n10252, new_n10253, new_n10254, new_n10255,
    new_n10256, new_n10257, new_n10258, new_n10259, new_n10260, new_n10261,
    new_n10262, new_n10263, new_n10264, new_n10265, new_n10266, new_n10267,
    new_n10268, new_n10269, new_n10270, new_n10271, new_n10272, new_n10273,
    new_n10274, new_n10275, new_n10276, new_n10277, new_n10278, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297,
    new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303,
    new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309,
    new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315,
    new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326, new_n10327,
    new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340,
    new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356, new_n10357, new_n10358,
    new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364,
    new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370,
    new_n10371, new_n10372, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385, new_n10386, new_n10387, new_n10388,
    new_n10389, new_n10390, new_n10391, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436,
    new_n10437, new_n10438, new_n10439, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451, new_n10452, new_n10453, new_n10454,
    new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460,
    new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561, new_n10562,
    new_n10563, new_n10564, new_n10565, new_n10566, new_n10567, new_n10568,
    new_n10569, new_n10570, new_n10571, new_n10572, new_n10573, new_n10574,
    new_n10575, new_n10576, new_n10577, new_n10578, new_n10579, new_n10580,
    new_n10581, new_n10582, new_n10583, new_n10584, new_n10585, new_n10586,
    new_n10587, new_n10588, new_n10589, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644, new_n10645, new_n10646,
    new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652,
    new_n10653, new_n10654, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692, new_n10693, new_n10694, new_n10695,
    new_n10696, new_n10697, new_n10698, new_n10699, new_n10700, new_n10701,
    new_n10702, new_n10703, new_n10704, new_n10705, new_n10706, new_n10707,
    new_n10708, new_n10709, new_n10710, new_n10711, new_n10712, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719,
    new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737,
    new_n10738, new_n10739, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756, new_n10757, new_n10758, new_n10759, new_n10760, new_n10761,
    new_n10762, new_n10763, new_n10764, new_n10765, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773,
    new_n10774, new_n10775, new_n10776, new_n10777, new_n10778, new_n10779,
    new_n10780, new_n10781, new_n10782, new_n10783, new_n10784, new_n10785,
    new_n10786, new_n10787, new_n10788, new_n10789, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848, new_n10849, new_n10850, new_n10851,
    new_n10852, new_n10853, new_n10854, new_n10855, new_n10856, new_n10857,
    new_n10858, new_n10859, new_n10860, new_n10861, new_n10862, new_n10863,
    new_n10864, new_n10865, new_n10866, new_n10867, new_n10868, new_n10869,
    new_n10870, new_n10871, new_n10872, new_n10873, new_n10874, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887,
    new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893,
    new_n10894, new_n10895, new_n10896, new_n10897, new_n10898, new_n10899,
    new_n10900, new_n10901, new_n10902, new_n10903, new_n10904, new_n10905,
    new_n10906, new_n10907, new_n10908, new_n10909, new_n10910, new_n10911,
    new_n10912, new_n10913, new_n10914, new_n10915, new_n10916, new_n10917,
    new_n10918, new_n10919, new_n10920, new_n10921, new_n10922, new_n10923,
    new_n10924, new_n10925, new_n10926, new_n10927, new_n10928, new_n10929,
    new_n10930, new_n10931, new_n10932, new_n10933, new_n10934, new_n10935,
    new_n10936, new_n10937, new_n10938, new_n10939, new_n10940, new_n10941,
    new_n10942, new_n10943, new_n10944, new_n10945, new_n10946, new_n10947,
    new_n10948, new_n10949, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961, new_n10962, new_n10963, new_n10964, new_n10965,
    new_n10966, new_n10967, new_n10968, new_n10969, new_n10970, new_n10971,
    new_n10972, new_n10973, new_n10974, new_n10975, new_n10976, new_n10977,
    new_n10978, new_n10979, new_n10980, new_n10981, new_n10982, new_n10983,
    new_n10984, new_n10985, new_n10986, new_n10987, new_n10988, new_n10989,
    new_n10990, new_n10991, new_n10992, new_n10993, new_n10994, new_n10995,
    new_n10996, new_n10997, new_n10998, new_n10999, new_n11000, new_n11001,
    new_n11002, new_n11003, new_n11004, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074,
    new_n11075, new_n11076, new_n11077, new_n11078, new_n11079, new_n11080,
    new_n11081, new_n11082, new_n11083, new_n11084, new_n11085, new_n11086,
    new_n11087, new_n11088, new_n11089, new_n11090, new_n11091, new_n11092,
    new_n11093, new_n11094, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101, new_n11102, new_n11103, new_n11104,
    new_n11105, new_n11106, new_n11107, new_n11108, new_n11109, new_n11110,
    new_n11111, new_n11112, new_n11113, new_n11114, new_n11115, new_n11116,
    new_n11117, new_n11118, new_n11119, new_n11120, new_n11121, new_n11122,
    new_n11123, new_n11124, new_n11125, new_n11126, new_n11127, new_n11128,
    new_n11129, new_n11130, new_n11131, new_n11132, new_n11133, new_n11134,
    new_n11135, new_n11136, new_n11137, new_n11138, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146,
    new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170,
    new_n11171, new_n11172, new_n11173, new_n11174, new_n11175, new_n11176,
    new_n11177, new_n11178, new_n11179, new_n11180, new_n11181, new_n11182,
    new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194,
    new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200,
    new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206,
    new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212,
    new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11218,
    new_n11219, new_n11220, new_n11221, new_n11222, new_n11223, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260,
    new_n11261, new_n11262, new_n11263, new_n11264, new_n11265, new_n11266,
    new_n11267, new_n11268, new_n11269, new_n11270, new_n11271, new_n11272,
    new_n11273, new_n11274, new_n11275, new_n11276, new_n11277, new_n11278,
    new_n11279, new_n11280, new_n11281, new_n11282, new_n11283, new_n11284,
    new_n11285, new_n11286, new_n11287, new_n11288, new_n11289, new_n11290,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311, new_n11312, new_n11313, new_n11314,
    new_n11315, new_n11316, new_n11317, new_n11318, new_n11319, new_n11320,
    new_n11321, new_n11323, new_n11324, new_n11325, new_n11326, new_n11327,
    new_n11328, new_n11329, new_n11330, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347, new_n11348, new_n11349, new_n11350, new_n11351,
    new_n11352, new_n11353, new_n11354, new_n11355, new_n11356, new_n11357,
    new_n11358, new_n11359, new_n11360, new_n11361, new_n11362, new_n11363,
    new_n11364, new_n11365, new_n11366, new_n11367, new_n11368, new_n11369,
    new_n11370, new_n11371, new_n11372, new_n11373, new_n11374, new_n11375,
    new_n11376, new_n11377, new_n11378, new_n11379, new_n11380, new_n11381,
    new_n11382, new_n11383, new_n11384, new_n11385, new_n11386, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391, new_n11392, new_n11393,
    new_n11394, new_n11395, new_n11396, new_n11397, new_n11398, new_n11399,
    new_n11400, new_n11401, new_n11402, new_n11403, new_n11404, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417,
    new_n11418, new_n11419, new_n11420, new_n11421, new_n11422, new_n11423,
    new_n11424, new_n11425, new_n11426, new_n11427, new_n11428, new_n11429,
    new_n11430, new_n11431, new_n11432, new_n11433, new_n11434, new_n11435,
    new_n11436, new_n11437, new_n11438, new_n11439, new_n11440, new_n11441,
    new_n11442, new_n11443, new_n11444, new_n11445, new_n11446, new_n11447,
    new_n11448, new_n11449, new_n11450, new_n11451, new_n11452, new_n11453,
    new_n11454, new_n11455, new_n11456, new_n11457, new_n11458, new_n11459,
    new_n11460, new_n11461, new_n11462, new_n11463, new_n11464, new_n11465,
    new_n11466, new_n11467, new_n11468, new_n11469, new_n11470, new_n11471,
    new_n11472, new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478, new_n11479, new_n11480, new_n11481, new_n11482, new_n11483,
    new_n11484, new_n11485, new_n11486, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496, new_n11497, new_n11498, new_n11499, new_n11500, new_n11501,
    new_n11502, new_n11503, new_n11504, new_n11505, new_n11506, new_n11507,
    new_n11508, new_n11509, new_n11510, new_n11511, new_n11512, new_n11513,
    new_n11514, new_n11515, new_n11516, new_n11517, new_n11518, new_n11519,
    new_n11520, new_n11521, new_n11522, new_n11523, new_n11524, new_n11525,
    new_n11526, new_n11527, new_n11528, new_n11529, new_n11530, new_n11531,
    new_n11532, new_n11533, new_n11534, new_n11535, new_n11536, new_n11537,
    new_n11538, new_n11539, new_n11540, new_n11541, new_n11542, new_n11543,
    new_n11544, new_n11545, new_n11546, new_n11547, new_n11548, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564, new_n11565, new_n11566, new_n11567,
    new_n11568, new_n11569, new_n11570, new_n11571, new_n11572, new_n11573,
    new_n11574, new_n11575, new_n11576, new_n11577, new_n11578, new_n11579,
    new_n11580, new_n11581, new_n11582, new_n11583, new_n11584, new_n11585,
    new_n11586, new_n11587, new_n11588, new_n11589, new_n11590, new_n11591,
    new_n11592, new_n11593, new_n11594, new_n11595, new_n11596, new_n11597,
    new_n11598, new_n11599, new_n11600, new_n11601, new_n11602, new_n11603,
    new_n11604, new_n11605, new_n11606, new_n11607, new_n11608, new_n11609,
    new_n11610, new_n11611, new_n11612, new_n11613, new_n11614, new_n11615,
    new_n11616, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664,
    new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676,
    new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724,
    new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796,
    new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802,
    new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808,
    new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814,
    new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837, new_n11838,
    new_n11839, new_n11840, new_n11841, new_n11842, new_n11843, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922,
    new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928,
    new_n11929, new_n11930, new_n11931, new_n11932, new_n11933, new_n11934,
    new_n11935, new_n11936, new_n11937, new_n11938, new_n11939, new_n11940,
    new_n11941, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971,
    new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980, new_n11981, new_n11982, new_n11983,
    new_n11984, new_n11985, new_n11986, new_n11987, new_n11988, new_n11989,
    new_n11990, new_n11991, new_n11992, new_n11993, new_n11994, new_n11995,
    new_n11996, new_n11997, new_n11998, new_n11999, new_n12000, new_n12001,
    new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025,
    new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031,
    new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037,
    new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043,
    new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049,
    new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055,
    new_n12056, new_n12057, new_n12058, new_n12059, new_n12060, new_n12061,
    new_n12062, new_n12063, new_n12064, new_n12065, new_n12066, new_n12067,
    new_n12068, new_n12069, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076, new_n12077, new_n12078, new_n12079,
    new_n12080, new_n12081, new_n12082, new_n12083, new_n12084, new_n12085,
    new_n12086, new_n12087, new_n12088, new_n12089, new_n12090, new_n12091,
    new_n12092, new_n12093, new_n12094, new_n12095, new_n12096, new_n12097,
    new_n12098, new_n12099, new_n12100, new_n12101, new_n12102, new_n12103,
    new_n12104, new_n12105, new_n12106, new_n12107, new_n12108, new_n12109,
    new_n12110, new_n12111, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146, new_n12147, new_n12148, new_n12149, new_n12150, new_n12151,
    new_n12152, new_n12153, new_n12154, new_n12155, new_n12156, new_n12157,
    new_n12158, new_n12159, new_n12160, new_n12161, new_n12162, new_n12163,
    new_n12164, new_n12165, new_n12166, new_n12167, new_n12168, new_n12169,
    new_n12170, new_n12171, new_n12172, new_n12173, new_n12174, new_n12175,
    new_n12176, new_n12177, new_n12178, new_n12179, new_n12180, new_n12181,
    new_n12182, new_n12183, new_n12184, new_n12185, new_n12186, new_n12187,
    new_n12188, new_n12189, new_n12190, new_n12191, new_n12192, new_n12193,
    new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199,
    new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205,
    new_n12206, new_n12207, new_n12208, new_n12209, new_n12210, new_n12211,
    new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222, new_n12223,
    new_n12224, new_n12225, new_n12226, new_n12227, new_n12228, new_n12229,
    new_n12230, new_n12231, new_n12232, new_n12233, new_n12234, new_n12235,
    new_n12236, new_n12237, new_n12238, new_n12239, new_n12240, new_n12241,
    new_n12242, new_n12243, new_n12244, new_n12245, new_n12246, new_n12247,
    new_n12248, new_n12249, new_n12250, new_n12251, new_n12252, new_n12253,
    new_n12254, new_n12255, new_n12256, new_n12257, new_n12258, new_n12259,
    new_n12260, new_n12261, new_n12262, new_n12263, new_n12264, new_n12265,
    new_n12266, new_n12267, new_n12268, new_n12269, new_n12270, new_n12271,
    new_n12272, new_n12273, new_n12274, new_n12275, new_n12276, new_n12277,
    new_n12278, new_n12279, new_n12280, new_n12281, new_n12282, new_n12283,
    new_n12284, new_n12285, new_n12286, new_n12287, new_n12288, new_n12289,
    new_n12290, new_n12291, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299, new_n12300, new_n12301, new_n12302,
    new_n12303, new_n12304, new_n12305, new_n12306, new_n12307, new_n12308,
    new_n12309, new_n12310, new_n12311, new_n12312, new_n12313, new_n12314,
    new_n12315, new_n12316, new_n12317, new_n12318, new_n12319, new_n12320,
    new_n12321, new_n12322, new_n12323, new_n12324, new_n12325, new_n12326,
    new_n12327, new_n12328, new_n12329, new_n12330, new_n12331, new_n12332,
    new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346, new_n12347, new_n12348, new_n12349, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380,
    new_n12381, new_n12382, new_n12383, new_n12384, new_n12385, new_n12386,
    new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464,
    new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470,
    new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476,
    new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494,
    new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500,
    new_n12501, new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507, new_n12508, new_n12509, new_n12510, new_n12511, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542,
    new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566,
    new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572,
    new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578,
    new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584,
    new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590,
    new_n12591, new_n12592, new_n12593, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607, new_n12608,
    new_n12609, new_n12610, new_n12611, new_n12612, new_n12613, new_n12614,
    new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648, new_n12649, new_n12650, new_n12651,
    new_n12652, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675,
    new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681,
    new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687,
    new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693,
    new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704, new_n12705,
    new_n12706, new_n12707, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725, new_n12726, new_n12727, new_n12728, new_n12729,
    new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735,
    new_n12736, new_n12737, new_n12738, new_n12739, new_n12740, new_n12741,
    new_n12742, new_n12743, new_n12744, new_n12745, new_n12746, new_n12747,
    new_n12748, new_n12749, new_n12750, new_n12751, new_n12752, new_n12753,
    new_n12754, new_n12755, new_n12756, new_n12757, new_n12758, new_n12759,
    new_n12760, new_n12761, new_n12762, new_n12763, new_n12764, new_n12765,
    new_n12766, new_n12767, new_n12768, new_n12769, new_n12770, new_n12771,
    new_n12772, new_n12773, new_n12774, new_n12775, new_n12776, new_n12777,
    new_n12778, new_n12779, new_n12780, new_n12781, new_n12782, new_n12783,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800, new_n12801,
    new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842, new_n12843,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860, new_n12861,
    new_n12862, new_n12863, new_n12864, new_n12865, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870, new_n12871, new_n12872, new_n12873,
    new_n12874, new_n12875, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897,
    new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903,
    new_n12904, new_n12905, new_n12906, new_n12907, new_n12908, new_n12909,
    new_n12910, new_n12911, new_n12912, new_n12913, new_n12914, new_n12915,
    new_n12916, new_n12917, new_n12918, new_n12919, new_n12920, new_n12921,
    new_n12922, new_n12923, new_n12924, new_n12925, new_n12926, new_n12927,
    new_n12928, new_n12929, new_n12930, new_n12931, new_n12932, new_n12933,
    new_n12934, new_n12935, new_n12936, new_n12937, new_n12938, new_n12939,
    new_n12940, new_n12941, new_n12942, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956, new_n12957,
    new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963,
    new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969,
    new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975,
    new_n12976, new_n12977, new_n12978, new_n12979, new_n12980, new_n12982,
    new_n12983, new_n12984, new_n12985, new_n12986, new_n12987, new_n12988,
    new_n12989, new_n12990, new_n12991, new_n12992, new_n12993, new_n12994,
    new_n12995, new_n12996, new_n12997, new_n12998, new_n12999, new_n13000,
    new_n13001, new_n13002, new_n13003, new_n13004, new_n13005, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030,
    new_n13031, new_n13032, new_n13033, new_n13034, new_n13035, new_n13036,
    new_n13037, new_n13038, new_n13039, new_n13040, new_n13041, new_n13042,
    new_n13043, new_n13044, new_n13045, new_n13046, new_n13047, new_n13048,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053, new_n13054,
    new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126,
    new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132,
    new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138,
    new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144,
    new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150,
    new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156,
    new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162,
    new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264,
    new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270,
    new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13292, new_n13293, new_n13294, new_n13295,
    new_n13296, new_n13297, new_n13298, new_n13299, new_n13300, new_n13301,
    new_n13302, new_n13303, new_n13304, new_n13305, new_n13306, new_n13307,
    new_n13308, new_n13309, new_n13310, new_n13311, new_n13312, new_n13313,
    new_n13314, new_n13315, new_n13316, new_n13317, new_n13318, new_n13319,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333, new_n13334, new_n13335, new_n13336, new_n13337,
    new_n13338, new_n13339, new_n13340, new_n13341, new_n13342, new_n13343,
    new_n13344, new_n13345, new_n13346, new_n13347, new_n13348, new_n13349,
    new_n13350, new_n13351, new_n13352, new_n13353, new_n13354, new_n13355,
    new_n13356, new_n13357, new_n13358, new_n13359, new_n13360, new_n13361,
    new_n13362, new_n13363, new_n13364, new_n13365, new_n13366, new_n13367,
    new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373,
    new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407, new_n13408, new_n13409,
    new_n13410, new_n13411, new_n13412, new_n13413, new_n13414, new_n13415,
    new_n13416, new_n13417, new_n13418, new_n13419, new_n13420, new_n13421,
    new_n13422, new_n13423, new_n13424, new_n13425, new_n13426, new_n13427,
    new_n13428, new_n13429, new_n13430, new_n13431, new_n13432, new_n13433,
    new_n13434, new_n13435, new_n13436, new_n13437, new_n13438, new_n13439,
    new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445,
    new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451,
    new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457,
    new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481,
    new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487,
    new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493,
    new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511,
    new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517,
    new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523,
    new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529,
    new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559,
    new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565,
    new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571,
    new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577,
    new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583,
    new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589,
    new_n13590, new_n13591, new_n13592, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602,
    new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608,
    new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614,
    new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620,
    new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626,
    new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632,
    new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638,
    new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053,
    new_n14054, new_n14055, new_n14056, new_n14057, new_n14058, new_n14059,
    new_n14060, new_n14061, new_n14062, new_n14063, new_n14064, new_n14065,
    new_n14066, new_n14067, new_n14068, new_n14069, new_n14070, new_n14071,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083,
    new_n14084, new_n14085, new_n14086, new_n14087, new_n14088, new_n14089,
    new_n14090, new_n14091, new_n14092, new_n14093, new_n14094, new_n14095,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106, new_n14107,
    new_n14108, new_n14109, new_n14110, new_n14111, new_n14112, new_n14113,
    new_n14114, new_n14115, new_n14116, new_n14117, new_n14118, new_n14119,
    new_n14120, new_n14121, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126, new_n14127, new_n14128, new_n14129, new_n14130, new_n14131,
    new_n14132, new_n14133, new_n14134, new_n14135, new_n14136, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147, new_n14148, new_n14149,
    new_n14150, new_n14151, new_n14152, new_n14153, new_n14154, new_n14155,
    new_n14156, new_n14157, new_n14158, new_n14159, new_n14160, new_n14161,
    new_n14162, new_n14163, new_n14164, new_n14165, new_n14166, new_n14167,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211, new_n14212, new_n14213, new_n14214, new_n14215, new_n14216,
    new_n14217, new_n14218, new_n14219, new_n14220, new_n14221, new_n14222,
    new_n14223, new_n14224, new_n14225, new_n14226, new_n14227, new_n14228,
    new_n14229, new_n14230, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267, new_n14268, new_n14269, new_n14270,
    new_n14271, new_n14272, new_n14273, new_n14274, new_n14275, new_n14276,
    new_n14277, new_n14278, new_n14279, new_n14280, new_n14281, new_n14282,
    new_n14283, new_n14284, new_n14285, new_n14286, new_n14287, new_n14288,
    new_n14289, new_n14290, new_n14291, new_n14292, new_n14293, new_n14294,
    new_n14295, new_n14296, new_n14297, new_n14298, new_n14299, new_n14300,
    new_n14301, new_n14302, new_n14303, new_n14304, new_n14305, new_n14306,
    new_n14307, new_n14308, new_n14309, new_n14310, new_n14311, new_n14312,
    new_n14313, new_n14314, new_n14315, new_n14316, new_n14317, new_n14318,
    new_n14319, new_n14320, new_n14321, new_n14322, new_n14323, new_n14324,
    new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336,
    new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342,
    new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366,
    new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372,
    new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378,
    new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384,
    new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390,
    new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396,
    new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402,
    new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408,
    new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426,
    new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432,
    new_n14433, new_n14434, new_n14435, new_n14436, new_n14437, new_n14438,
    new_n14439, new_n14440, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457, new_n14458, new_n14459, new_n14460, new_n14461, new_n14462,
    new_n14463, new_n14464, new_n14466, new_n14467, new_n14468, new_n14469,
    new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475,
    new_n14476, new_n14477, new_n14478, new_n14479, new_n14480, new_n14481,
    new_n14482, new_n14483, new_n14484, new_n14485, new_n14486, new_n14487,
    new_n14488, new_n14489, new_n14490, new_n14491, new_n14492, new_n14493,
    new_n14494, new_n14495, new_n14496, new_n14497, new_n14498, new_n14499,
    new_n14500, new_n14501, new_n14502, new_n14503, new_n14504, new_n14505,
    new_n14506, new_n14507, new_n14508, new_n14509, new_n14510, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540, new_n14541,
    new_n14542, new_n14543, new_n14544, new_n14545, new_n14546, new_n14547,
    new_n14548, new_n14549, new_n14550, new_n14551, new_n14552, new_n14553,
    new_n14554, new_n14555, new_n14556, new_n14557, new_n14558, new_n14559,
    new_n14560, new_n14561, new_n14562, new_n14563, new_n14564, new_n14565,
    new_n14566, new_n14567, new_n14568, new_n14569, new_n14570, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575, new_n14576, new_n14577,
    new_n14578, new_n14579, new_n14580, new_n14581, new_n14582, new_n14583,
    new_n14584, new_n14585, new_n14586, new_n14587, new_n14588, new_n14589,
    new_n14590, new_n14591, new_n14592, new_n14593, new_n14594, new_n14595,
    new_n14596, new_n14597, new_n14598, new_n14599, new_n14600, new_n14601,
    new_n14602, new_n14603, new_n14604, new_n14605, new_n14606, new_n14607,
    new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613,
    new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619,
    new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633, new_n14634, new_n14635, new_n14636, new_n14637,
    new_n14638, new_n14639, new_n14640, new_n14641, new_n14642, new_n14643,
    new_n14644, new_n14645, new_n14646, new_n14647, new_n14648, new_n14649,
    new_n14650, new_n14651, new_n14652, new_n14653, new_n14654, new_n14655,
    new_n14656, new_n14657, new_n14658, new_n14659, new_n14660, new_n14661,
    new_n14662, new_n14663, new_n14664, new_n14665, new_n14666, new_n14667,
    new_n14668, new_n14669, new_n14670, new_n14671, new_n14672, new_n14673,
    new_n14674, new_n14675, new_n14676, new_n14677, new_n14678, new_n14679,
    new_n14680, new_n14681, new_n14682, new_n14683, new_n14684, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692, new_n14693, new_n14694, new_n14695, new_n14696, new_n14697,
    new_n14698, new_n14699, new_n14700, new_n14701, new_n14702, new_n14703,
    new_n14704, new_n14705, new_n14706, new_n14707, new_n14708, new_n14709,
    new_n14710, new_n14711, new_n14712, new_n14713, new_n14714, new_n14715,
    new_n14716, new_n14717, new_n14718, new_n14719, new_n14720, new_n14721,
    new_n14722, new_n14723, new_n14724, new_n14725, new_n14726, new_n14727,
    new_n14728, new_n14729, new_n14730, new_n14731, new_n14732, new_n14733,
    new_n14734, new_n14735, new_n14736, new_n14737, new_n14738, new_n14739,
    new_n14740, new_n14741, new_n14742, new_n14743, new_n14744, new_n14745,
    new_n14746, new_n14747, new_n14748, new_n14749, new_n14750, new_n14751,
    new_n14752, new_n14753, new_n14754, new_n14755, new_n14756, new_n14757,
    new_n14758, new_n14759, new_n14760, new_n14761, new_n14762, new_n14764,
    new_n14765, new_n14766, new_n14767, new_n14768, new_n14769, new_n14770,
    new_n14771, new_n14772, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801, new_n14802, new_n14803, new_n14804, new_n14805, new_n14806,
    new_n14807, new_n14808, new_n14809, new_n14810, new_n14811, new_n14812,
    new_n14813, new_n14814, new_n14815, new_n14816, new_n14817, new_n14818,
    new_n14819, new_n14820, new_n14821, new_n14822, new_n14823, new_n14824,
    new_n14825, new_n14826, new_n14827, new_n14828, new_n14829, new_n14830,
    new_n14831, new_n14832, new_n14833, new_n14834, new_n14835, new_n14836,
    new_n14837, new_n14838, new_n14839, new_n14840, new_n14841, new_n14842,
    new_n14843, new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849, new_n14850, new_n14851, new_n14852, new_n14853, new_n14854,
    new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860,
    new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866,
    new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872,
    new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878,
    new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884,
    new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890,
    new_n14891, new_n14892, new_n14893, new_n14894, new_n14895, new_n14896,
    new_n14897, new_n14898, new_n14899, new_n14900, new_n14901, new_n14902,
    new_n14903, new_n14904, new_n14905, new_n14906, new_n14907, new_n14908,
    new_n14909, new_n14910, new_n14911, new_n14912, new_n14913, new_n14914,
    new_n14915, new_n14916, new_n14917, new_n14918, new_n14919, new_n14920,
    new_n14921, new_n14922, new_n14923, new_n14924, new_n14925, new_n14926,
    new_n14927, new_n14928, new_n14929, new_n14930, new_n14931, new_n14932,
    new_n14933, new_n14934, new_n14935, new_n14936, new_n14937, new_n14938,
    new_n14939, new_n14940, new_n14941, new_n14942, new_n14943, new_n14944,
    new_n14945, new_n14946, new_n14947, new_n14948, new_n14949, new_n14950,
    new_n14951, new_n14952, new_n14953, new_n14954, new_n14955, new_n14956,
    new_n14957, new_n14958, new_n14959, new_n14960, new_n14961, new_n14962,
    new_n14963, new_n14964, new_n14965, new_n14966, new_n14967, new_n14968,
    new_n14969, new_n14970, new_n14971, new_n14972, new_n14973, new_n14974,
    new_n14975, new_n14976, new_n14977, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002, new_n15003, new_n15004,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011, new_n15012, new_n15013, new_n15014, new_n15015, new_n15016,
    new_n15017, new_n15018, new_n15019, new_n15020, new_n15021, new_n15022,
    new_n15023, new_n15024, new_n15025, new_n15026, new_n15027, new_n15028,
    new_n15029, new_n15030, new_n15032, new_n15033, new_n15034, new_n15035,
    new_n15036, new_n15037, new_n15038, new_n15039, new_n15040, new_n15041,
    new_n15042, new_n15043, new_n15044, new_n15045, new_n15046, new_n15047,
    new_n15048, new_n15049, new_n15050, new_n15051, new_n15052, new_n15053,
    new_n15054, new_n15055, new_n15056, new_n15057, new_n15058, new_n15059,
    new_n15060, new_n15061, new_n15062, new_n15063, new_n15064, new_n15065,
    new_n15066, new_n15067, new_n15068, new_n15069, new_n15070, new_n15071,
    new_n15072, new_n15073, new_n15074, new_n15075, new_n15076, new_n15077,
    new_n15078, new_n15079, new_n15080, new_n15081, new_n15082, new_n15083,
    new_n15084, new_n15085, new_n15086, new_n15087, new_n15088, new_n15089,
    new_n15090, new_n15091, new_n15092, new_n15093, new_n15094, new_n15095,
    new_n15096, new_n15097, new_n15098, new_n15099, new_n15100, new_n15101,
    new_n15102, new_n15103, new_n15104, new_n15105, new_n15106, new_n15107,
    new_n15108, new_n15109, new_n15110, new_n15111, new_n15112, new_n15113,
    new_n15114, new_n15115, new_n15116, new_n15117, new_n15118, new_n15119,
    new_n15120, new_n15121, new_n15122, new_n15123, new_n15124, new_n15125,
    new_n15126, new_n15127, new_n15128, new_n15129, new_n15130, new_n15131,
    new_n15132, new_n15133, new_n15134, new_n15135, new_n15136, new_n15137,
    new_n15138, new_n15139, new_n15140, new_n15141, new_n15142, new_n15143,
    new_n15144, new_n15145, new_n15146, new_n15147, new_n15148, new_n15149,
    new_n15150, new_n15151, new_n15152, new_n15153, new_n15154, new_n15155,
    new_n15156, new_n15157, new_n15158, new_n15159, new_n15160, new_n15161,
    new_n15162, new_n15163, new_n15164, new_n15165, new_n15166, new_n15167,
    new_n15168, new_n15169, new_n15170, new_n15171, new_n15172, new_n15173,
    new_n15174, new_n15175, new_n15176, new_n15177, new_n15178, new_n15179,
    new_n15180, new_n15181, new_n15182, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205, new_n15206, new_n15207, new_n15208, new_n15209,
    new_n15210, new_n15211, new_n15212, new_n15213, new_n15214, new_n15215,
    new_n15216, new_n15217, new_n15218, new_n15219, new_n15220, new_n15221,
    new_n15222, new_n15223, new_n15224, new_n15225, new_n15226, new_n15227,
    new_n15228, new_n15229, new_n15230, new_n15231, new_n15232, new_n15233,
    new_n15234, new_n15235, new_n15236, new_n15237, new_n15238, new_n15239,
    new_n15240, new_n15241, new_n15242, new_n15243, new_n15244, new_n15245,
    new_n15246, new_n15247, new_n15248, new_n15249, new_n15250, new_n15251,
    new_n15252, new_n15253, new_n15254, new_n15255, new_n15256, new_n15257,
    new_n15258, new_n15259, new_n15260, new_n15261, new_n15262, new_n15263,
    new_n15264, new_n15265, new_n15266, new_n15267, new_n15268, new_n15269,
    new_n15270, new_n15271, new_n15272, new_n15273, new_n15274, new_n15275,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289, new_n15290, new_n15291, new_n15292, new_n15293,
    new_n15294, new_n15295, new_n15296, new_n15297, new_n15298, new_n15299,
    new_n15300, new_n15301, new_n15302, new_n15303, new_n15304, new_n15305,
    new_n15306, new_n15307, new_n15308, new_n15309, new_n15310, new_n15311,
    new_n15312, new_n15313, new_n15314, new_n15315, new_n15316, new_n15317,
    new_n15318, new_n15319, new_n15320, new_n15321, new_n15322, new_n15323,
    new_n15324, new_n15325, new_n15326, new_n15327, new_n15328, new_n15329,
    new_n15330, new_n15331, new_n15332, new_n15333, new_n15334, new_n15335,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345, new_n15346, new_n15347, new_n15348,
    new_n15349, new_n15350, new_n15351, new_n15352, new_n15353, new_n15354,
    new_n15355, new_n15356, new_n15357, new_n15358, new_n15359, new_n15360,
    new_n15361, new_n15362, new_n15363, new_n15364, new_n15365, new_n15366,
    new_n15367, new_n15368, new_n15369, new_n15370, new_n15371, new_n15372,
    new_n15373, new_n15374, new_n15375, new_n15376, new_n15377, new_n15378,
    new_n15379, new_n15380, new_n15381, new_n15382, new_n15383, new_n15384,
    new_n15385, new_n15386, new_n15387, new_n15388, new_n15389, new_n15390,
    new_n15391, new_n15392, new_n15393, new_n15394, new_n15395, new_n15396,
    new_n15397, new_n15398, new_n15399, new_n15400, new_n15401, new_n15402,
    new_n15403, new_n15404, new_n15405, new_n15406, new_n15407, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424, new_n15425, new_n15426,
    new_n15427, new_n15428, new_n15429, new_n15430, new_n15431, new_n15432,
    new_n15433, new_n15434, new_n15435, new_n15436, new_n15437, new_n15438,
    new_n15439, new_n15440, new_n15441, new_n15442, new_n15443, new_n15444,
    new_n15445, new_n15446, new_n15447, new_n15448, new_n15449, new_n15450,
    new_n15451, new_n15452, new_n15453, new_n15454, new_n15455, new_n15456,
    new_n15457, new_n15458, new_n15459, new_n15460, new_n15461, new_n15462,
    new_n15463, new_n15464, new_n15465, new_n15466, new_n15467, new_n15468,
    new_n15469, new_n15470, new_n15471, new_n15472, new_n15473, new_n15474,
    new_n15475, new_n15476, new_n15477, new_n15478, new_n15479, new_n15480,
    new_n15481, new_n15482, new_n15483, new_n15484, new_n15485, new_n15486,
    new_n15487, new_n15488, new_n15489, new_n15490, new_n15491, new_n15492,
    new_n15493, new_n15494, new_n15495, new_n15496, new_n15497, new_n15498,
    new_n15499, new_n15500, new_n15501, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506, new_n15507, new_n15508, new_n15509, new_n15510,
    new_n15511, new_n15512, new_n15513, new_n15514, new_n15515, new_n15516,
    new_n15517, new_n15518, new_n15519, new_n15520, new_n15521, new_n15522,
    new_n15523, new_n15524, new_n15525, new_n15526, new_n15527, new_n15528,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539, new_n15540,
    new_n15541, new_n15542, new_n15543, new_n15544, new_n15545, new_n15546,
    new_n15547, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552,
    new_n15553, new_n15554, new_n15555, new_n15556, new_n15557, new_n15558,
    new_n15559, new_n15560, new_n15561, new_n15562, new_n15563, new_n15564,
    new_n15565, new_n15566, new_n15567, new_n15568, new_n15569, new_n15570,
    new_n15571, new_n15572, new_n15573, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587, new_n15588,
    new_n15589, new_n15590, new_n15591, new_n15592, new_n15593, new_n15594,
    new_n15595, new_n15596, new_n15597, new_n15598, new_n15599, new_n15600,
    new_n15601, new_n15602, new_n15603, new_n15604, new_n15605, new_n15606,
    new_n15607, new_n15608, new_n15609, new_n15610, new_n15611, new_n15612,
    new_n15613, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15620, new_n15621, new_n15622, new_n15623, new_n15624, new_n15625,
    new_n15626, new_n15627, new_n15628, new_n15629, new_n15630, new_n15631,
    new_n15632, new_n15633, new_n15634, new_n15635, new_n15636, new_n15637,
    new_n15638, new_n15639, new_n15640, new_n15641, new_n15642, new_n15643,
    new_n15644, new_n15645, new_n15646, new_n15647, new_n15648, new_n15649,
    new_n15650, new_n15651, new_n15652, new_n15653, new_n15654, new_n15655,
    new_n15656, new_n15657, new_n15658, new_n15659, new_n15660, new_n15661,
    new_n15662, new_n15663, new_n15664, new_n15665, new_n15666, new_n15667,
    new_n15668, new_n15669, new_n15670, new_n15671, new_n15672, new_n15673,
    new_n15674, new_n15675, new_n15676, new_n15677, new_n15678, new_n15679,
    new_n15680, new_n15681, new_n15682, new_n15683, new_n15684, new_n15685,
    new_n15686, new_n15687, new_n15688, new_n15689, new_n15690, new_n15691,
    new_n15692, new_n15693, new_n15694, new_n15695, new_n15696, new_n15697,
    new_n15698, new_n15699, new_n15700, new_n15701, new_n15702, new_n15703,
    new_n15704, new_n15705, new_n15706, new_n15707, new_n15708, new_n15709,
    new_n15710, new_n15711, new_n15712, new_n15713, new_n15714, new_n15715,
    new_n15716, new_n15717, new_n15718, new_n15719, new_n15720, new_n15721,
    new_n15722, new_n15723, new_n15724, new_n15725, new_n15726, new_n15727,
    new_n15728, new_n15729, new_n15730, new_n15731, new_n15732, new_n15733,
    new_n15734, new_n15735, new_n15736, new_n15737, new_n15738, new_n15739,
    new_n15740, new_n15741, new_n15742, new_n15743, new_n15744, new_n15745,
    new_n15746, new_n15747, new_n15748, new_n15749, new_n15750, new_n15751,
    new_n15752, new_n15753, new_n15754, new_n15755, new_n15756, new_n15757,
    new_n15758, new_n15759, new_n15760, new_n15761, new_n15762, new_n15763,
    new_n15764, new_n15765, new_n15766, new_n15767, new_n15768, new_n15769,
    new_n15770, new_n15771, new_n15772, new_n15773, new_n15774, new_n15775,
    new_n15776, new_n15777, new_n15778, new_n15779, new_n15780, new_n15781,
    new_n15782, new_n15783, new_n15784, new_n15785, new_n15786, new_n15787,
    new_n15788, new_n15789, new_n15790, new_n15791, new_n15792, new_n15793,
    new_n15794, new_n15795, new_n15796, new_n15797, new_n15798, new_n15799,
    new_n15800, new_n15801, new_n15802, new_n15803, new_n15804, new_n15805,
    new_n15806, new_n15807, new_n15808, new_n15809, new_n15810, new_n15811,
    new_n15812, new_n15813, new_n15814, new_n15815, new_n15816, new_n15817,
    new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823,
    new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829,
    new_n15830, new_n15831, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15842, new_n15843, new_n15844, new_n15845, new_n15846, new_n15847,
    new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853,
    new_n15854, new_n15855, new_n15856, new_n15857, new_n15858, new_n15859,
    new_n15860, new_n15861, new_n15862, new_n15863, new_n15864, new_n15865,
    new_n15866, new_n15867, new_n15868, new_n15869, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884, new_n15885, new_n15886, new_n15887, new_n15888, new_n15889,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917, new_n15918, new_n15919,
    new_n15920, new_n15921, new_n15922, new_n15923, new_n15924, new_n15926,
    new_n15927, new_n15928, new_n15929, new_n15930, new_n15931, new_n15932,
    new_n15933, new_n15934, new_n15935, new_n15936, new_n15937, new_n15938,
    new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944,
    new_n15945, new_n15946, new_n15947, new_n15948, new_n15949, new_n15950,
    new_n15951, new_n15952, new_n15953, new_n15954, new_n15955, new_n15956,
    new_n15957, new_n15958, new_n15959, new_n15960, new_n15961, new_n15962,
    new_n15963, new_n15964, new_n15965, new_n15966, new_n15967, new_n15968,
    new_n15969, new_n15970, new_n15971, new_n15972, new_n15973, new_n15974,
    new_n15975, new_n15976, new_n15977, new_n15978, new_n15979, new_n15980,
    new_n15981, new_n15982, new_n15983, new_n15984, new_n15985, new_n15986,
    new_n15987, new_n15988, new_n15989, new_n15990, new_n15991, new_n15992,
    new_n15993, new_n15994, new_n15995, new_n15996, new_n15997, new_n15998,
    new_n15999, new_n16000, new_n16001, new_n16002, new_n16003, new_n16004,
    new_n16005, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010,
    new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016,
    new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022,
    new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034,
    new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040,
    new_n16041, new_n16042, new_n16043, new_n16044, new_n16045, new_n16046,
    new_n16047, new_n16048, new_n16049, new_n16050, new_n16051, new_n16052,
    new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058,
    new_n16059, new_n16060, new_n16061, new_n16062, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068, new_n16069, new_n16070,
    new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076,
    new_n16077, new_n16078, new_n16079, new_n16080, new_n16081, new_n16082,
    new_n16083, new_n16084, new_n16085, new_n16086, new_n16087, new_n16088,
    new_n16089, new_n16090, new_n16091, new_n16092, new_n16093, new_n16094,
    new_n16095, new_n16096, new_n16097, new_n16098, new_n16099, new_n16100,
    new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106,
    new_n16107, new_n16108, new_n16109, new_n16110, new_n16111, new_n16112,
    new_n16113, new_n16114, new_n16115, new_n16116, new_n16117, new_n16118,
    new_n16119, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124,
    new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16218, new_n16219, new_n16220, new_n16221,
    new_n16222, new_n16223, new_n16224, new_n16225, new_n16226, new_n16227,
    new_n16228, new_n16229, new_n16230, new_n16231, new_n16232, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239,
    new_n16240, new_n16241, new_n16242, new_n16243, new_n16244, new_n16245,
    new_n16246, new_n16247, new_n16248, new_n16249, new_n16250, new_n16251,
    new_n16252, new_n16253, new_n16254, new_n16255, new_n16256, new_n16257,
    new_n16258, new_n16259, new_n16260, new_n16261, new_n16262, new_n16263,
    new_n16264, new_n16265, new_n16266, new_n16267, new_n16268, new_n16269,
    new_n16270, new_n16271, new_n16272, new_n16273, new_n16274, new_n16275,
    new_n16276, new_n16277, new_n16278, new_n16279, new_n16280, new_n16281,
    new_n16282, new_n16283, new_n16284, new_n16285, new_n16286, new_n16287,
    new_n16288, new_n16289, new_n16290, new_n16291, new_n16292, new_n16293,
    new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311,
    new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317,
    new_n16318, new_n16319, new_n16320, new_n16321, new_n16322, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350, new_n16351, new_n16352, new_n16353,
    new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359,
    new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365,
    new_n16366, new_n16367, new_n16368, new_n16369, new_n16370, new_n16371,
    new_n16372, new_n16373, new_n16374, new_n16375, new_n16376, new_n16377,
    new_n16378, new_n16379, new_n16380, new_n16381, new_n16382, new_n16383,
    new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389,
    new_n16390, new_n16391, new_n16392, new_n16393, new_n16394, new_n16395,
    new_n16396, new_n16397, new_n16398, new_n16399, new_n16400, new_n16401,
    new_n16402, new_n16403, new_n16404, new_n16405, new_n16406, new_n16407,
    new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413,
    new_n16414, new_n16415, new_n16416, new_n16417, new_n16418, new_n16419,
    new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425,
    new_n16426, new_n16427, new_n16428, new_n16429, new_n16430, new_n16431,
    new_n16432, new_n16433, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439, new_n16440, new_n16441, new_n16442, new_n16443,
    new_n16444, new_n16445, new_n16446, new_n16447, new_n16448, new_n16449,
    new_n16450, new_n16451, new_n16452, new_n16453, new_n16454, new_n16455,
    new_n16456, new_n16457, new_n16458, new_n16459, new_n16460, new_n16461,
    new_n16462, new_n16463, new_n16464, new_n16465, new_n16466, new_n16467,
    new_n16468, new_n16469, new_n16470, new_n16471, new_n16472, new_n16473,
    new_n16474, new_n16475, new_n16476, new_n16477, new_n16478, new_n16479,
    new_n16480, new_n16481, new_n16482, new_n16483, new_n16484, new_n16485,
    new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491,
    new_n16492, new_n16493, new_n16494, new_n16495, new_n16496, new_n16497,
    new_n16498, new_n16499, new_n16500, new_n16501, new_n16502, new_n16503,
    new_n16504, new_n16505, new_n16506, new_n16507, new_n16508, new_n16509,
    new_n16510, new_n16511, new_n16512, new_n16513, new_n16514, new_n16515,
    new_n16516, new_n16517, new_n16518, new_n16519, new_n16520, new_n16521,
    new_n16522, new_n16523, new_n16525, new_n16526, new_n16527, new_n16528,
    new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534,
    new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540,
    new_n16541, new_n16542, new_n16543, new_n16544, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583, new_n16584, new_n16585, new_n16586, new_n16587, new_n16588,
    new_n16589, new_n16590, new_n16591, new_n16592, new_n16593, new_n16594,
    new_n16595, new_n16596, new_n16597, new_n16598, new_n16599, new_n16600,
    new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606,
    new_n16607, new_n16608, new_n16609, new_n16610, new_n16611, new_n16612,
    new_n16613, new_n16614, new_n16615, new_n16616, new_n16617, new_n16618,
    new_n16619, new_n16620, new_n16621, new_n16622, new_n16623, new_n16624,
    new_n16625, new_n16626, new_n16627, new_n16628, new_n16629, new_n16630,
    new_n16631, new_n16632, new_n16633, new_n16634, new_n16635, new_n16636,
    new_n16637, new_n16638, new_n16639, new_n16640, new_n16641, new_n16642,
    new_n16643, new_n16644, new_n16645, new_n16646, new_n16647, new_n16648,
    new_n16649, new_n16650, new_n16651, new_n16652, new_n16653, new_n16654,
    new_n16655, new_n16656, new_n16657, new_n16658, new_n16659, new_n16660,
    new_n16661, new_n16662, new_n16663, new_n16664, new_n16665, new_n16666,
    new_n16667, new_n16668, new_n16669, new_n16670, new_n16671, new_n16672,
    new_n16673, new_n16674, new_n16675, new_n16676, new_n16677, new_n16678,
    new_n16679, new_n16680, new_n16681, new_n16682, new_n16683, new_n16684,
    new_n16685, new_n16686, new_n16687, new_n16688, new_n16689, new_n16690,
    new_n16691, new_n16692, new_n16693, new_n16694, new_n16695, new_n16696,
    new_n16697, new_n16698, new_n16699, new_n16700, new_n16701, new_n16702,
    new_n16703, new_n16704, new_n16705, new_n16706, new_n16707, new_n16708,
    new_n16709, new_n16710, new_n16711, new_n16712, new_n16713, new_n16714,
    new_n16715, new_n16716, new_n16717, new_n16718, new_n16719, new_n16720,
    new_n16721, new_n16722, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733, new_n16734, new_n16735, new_n16736, new_n16737, new_n16738,
    new_n16739, new_n16740, new_n16741, new_n16742, new_n16743, new_n16744,
    new_n16745, new_n16746, new_n16747, new_n16748, new_n16749, new_n16750,
    new_n16751, new_n16752, new_n16753, new_n16754, new_n16755, new_n16756,
    new_n16757, new_n16758, new_n16759, new_n16760, new_n16761, new_n16762,
    new_n16763, new_n16764, new_n16765, new_n16766, new_n16767, new_n16768,
    new_n16769, new_n16770, new_n16771, new_n16772, new_n16773, new_n16774,
    new_n16775, new_n16776, new_n16777, new_n16778, new_n16779, new_n16780,
    new_n16781, new_n16782, new_n16783, new_n16784, new_n16785, new_n16786,
    new_n16787, new_n16788, new_n16789, new_n16790, new_n16791, new_n16792,
    new_n16793, new_n16794, new_n16795, new_n16796, new_n16797, new_n16799,
    new_n16800, new_n16801, new_n16802, new_n16803, new_n16804, new_n16805,
    new_n16806, new_n16807, new_n16808, new_n16809, new_n16810, new_n16811,
    new_n16812, new_n16813, new_n16814, new_n16815, new_n16816, new_n16817,
    new_n16818, new_n16819, new_n16820, new_n16821, new_n16822, new_n16823,
    new_n16824, new_n16825, new_n16826, new_n16827, new_n16828, new_n16829,
    new_n16830, new_n16831, new_n16832, new_n16833, new_n16834, new_n16835,
    new_n16836, new_n16837, new_n16838, new_n16839, new_n16840, new_n16841,
    new_n16842, new_n16843, new_n16844, new_n16845, new_n16846, new_n16847,
    new_n16848, new_n16849, new_n16850, new_n16851, new_n16852, new_n16853,
    new_n16854, new_n16855, new_n16856, new_n16857, new_n16858, new_n16859,
    new_n16860, new_n16861, new_n16862, new_n16863, new_n16864, new_n16865,
    new_n16866, new_n16867, new_n16868, new_n16869, new_n16870, new_n16871,
    new_n16872, new_n16873, new_n16874, new_n16875, new_n16876, new_n16877,
    new_n16878, new_n16879, new_n16880, new_n16881, new_n16882, new_n16883,
    new_n16884, new_n16885, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895,
    new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901,
    new_n16902, new_n16903, new_n16904, new_n16905, new_n16906, new_n16907,
    new_n16908, new_n16909, new_n16910, new_n16911, new_n16912, new_n16913,
    new_n16914, new_n16915, new_n16916, new_n16917, new_n16918, new_n16919,
    new_n16920, new_n16921, new_n16922, new_n16923, new_n16924, new_n16925,
    new_n16926, new_n16927, new_n16928, new_n16929, new_n16930, new_n16931,
    new_n16932, new_n16933, new_n16934, new_n16935, new_n16936, new_n16937,
    new_n16938, new_n16939, new_n16940, new_n16941, new_n16942, new_n16943,
    new_n16944, new_n16945, new_n16946, new_n16947, new_n16948, new_n16949,
    new_n16950, new_n16951, new_n16952, new_n16953, new_n16954, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968, new_n16969, new_n16970, new_n16971, new_n16972, new_n16973,
    new_n16974, new_n16975, new_n16976, new_n16977, new_n16978, new_n16979,
    new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985,
    new_n16986, new_n16987, new_n16988, new_n16989, new_n16990, new_n16991,
    new_n16992, new_n16993, new_n16994, new_n16995, new_n16996, new_n16997,
    new_n16998, new_n16999, new_n17000, new_n17001, new_n17002, new_n17003,
    new_n17004, new_n17005, new_n17006, new_n17007, new_n17008, new_n17009,
    new_n17010, new_n17011, new_n17012, new_n17013, new_n17014, new_n17015,
    new_n17016, new_n17017, new_n17018, new_n17019, new_n17020, new_n17021,
    new_n17022, new_n17023, new_n17024, new_n17025, new_n17026, new_n17027,
    new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033,
    new_n17034, new_n17035, new_n17036, new_n17037, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057,
    new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063,
    new_n17064, new_n17065, new_n17066, new_n17067, new_n17068, new_n17069,
    new_n17070, new_n17071, new_n17072, new_n17073, new_n17074, new_n17075,
    new_n17076, new_n17077, new_n17078, new_n17080, new_n17081, new_n17082,
    new_n17083, new_n17084, new_n17085, new_n17086, new_n17087, new_n17088,
    new_n17089, new_n17090, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095, new_n17096, new_n17097, new_n17098, new_n17099, new_n17100,
    new_n17101, new_n17102, new_n17103, new_n17104, new_n17105, new_n17106,
    new_n17107, new_n17108, new_n17109, new_n17110, new_n17111, new_n17112,
    new_n17113, new_n17114, new_n17115, new_n17116, new_n17117, new_n17118,
    new_n17119, new_n17120, new_n17121, new_n17122, new_n17123, new_n17124,
    new_n17125, new_n17126, new_n17127, new_n17128, new_n17129, new_n17130,
    new_n17131, new_n17132, new_n17133, new_n17134, new_n17135, new_n17136,
    new_n17137, new_n17138, new_n17139, new_n17140, new_n17141, new_n17142,
    new_n17143, new_n17144, new_n17145, new_n17146, new_n17147, new_n17148,
    new_n17149, new_n17150, new_n17151, new_n17152, new_n17153, new_n17154,
    new_n17155, new_n17156, new_n17157, new_n17158, new_n17159, new_n17160,
    new_n17161, new_n17162, new_n17163, new_n17164, new_n17165, new_n17166,
    new_n17167, new_n17168, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201, new_n17202,
    new_n17203, new_n17204, new_n17205, new_n17206, new_n17207, new_n17208,
    new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214,
    new_n17215, new_n17216, new_n17217, new_n17218, new_n17219, new_n17220,
    new_n17221, new_n17222, new_n17223, new_n17224, new_n17225, new_n17226,
    new_n17227, new_n17228, new_n17229, new_n17230, new_n17231, new_n17232,
    new_n17233, new_n17234, new_n17235, new_n17236, new_n17237, new_n17238,
    new_n17239, new_n17240, new_n17241, new_n17242, new_n17243, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249, new_n17250,
    new_n17251, new_n17252, new_n17253, new_n17254, new_n17255, new_n17256,
    new_n17257, new_n17258, new_n17259, new_n17260, new_n17261, new_n17262,
    new_n17263, new_n17264, new_n17265, new_n17266, new_n17267, new_n17268,
    new_n17269, new_n17270, new_n17271, new_n17272, new_n17273, new_n17274,
    new_n17275, new_n17276, new_n17277, new_n17278, new_n17279, new_n17280,
    new_n17281, new_n17282, new_n17283, new_n17284, new_n17285, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17292,
    new_n17293, new_n17294, new_n17295, new_n17296, new_n17297, new_n17298,
    new_n17299, new_n17300, new_n17301, new_n17302, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320, new_n17321, new_n17323,
    new_n17324, new_n17325, new_n17326, new_n17327, new_n17328, new_n17329,
    new_n17330, new_n17331, new_n17332, new_n17333, new_n17334, new_n17335,
    new_n17336, new_n17337, new_n17338, new_n17339, new_n17340, new_n17341,
    new_n17342, new_n17343, new_n17344, new_n17345, new_n17346, new_n17347,
    new_n17348, new_n17349, new_n17350, new_n17351, new_n17352, new_n17353,
    new_n17354, new_n17355, new_n17356, new_n17357, new_n17358, new_n17359,
    new_n17360, new_n17361, new_n17362, new_n17363, new_n17364, new_n17365,
    new_n17366, new_n17367, new_n17368, new_n17369, new_n17370, new_n17371,
    new_n17372, new_n17373, new_n17374, new_n17375, new_n17376, new_n17377,
    new_n17378, new_n17379, new_n17380, new_n17381, new_n17382, new_n17383,
    new_n17384, new_n17385, new_n17386, new_n17387, new_n17388, new_n17389,
    new_n17390, new_n17391, new_n17392, new_n17393, new_n17394, new_n17395,
    new_n17396, new_n17397, new_n17398, new_n17399, new_n17400, new_n17401,
    new_n17402, new_n17403, new_n17404, new_n17405, new_n17406, new_n17407,
    new_n17408, new_n17409, new_n17410, new_n17411, new_n17412, new_n17413,
    new_n17414, new_n17415, new_n17416, new_n17417, new_n17418, new_n17419,
    new_n17420, new_n17421, new_n17422, new_n17423, new_n17424, new_n17425,
    new_n17426, new_n17427, new_n17428, new_n17429, new_n17430, new_n17431,
    new_n17432, new_n17433, new_n17434, new_n17435, new_n17436, new_n17437,
    new_n17438, new_n17439, new_n17440, new_n17441, new_n17442, new_n17443,
    new_n17444, new_n17445, new_n17446, new_n17447, new_n17448, new_n17449,
    new_n17450, new_n17451, new_n17452, new_n17453, new_n17454, new_n17455,
    new_n17456, new_n17457, new_n17458, new_n17459, new_n17460, new_n17461,
    new_n17462, new_n17463, new_n17464, new_n17465, new_n17466, new_n17467,
    new_n17468, new_n17469, new_n17470, new_n17471, new_n17472, new_n17473,
    new_n17474, new_n17475, new_n17476, new_n17477, new_n17478, new_n17479,
    new_n17480, new_n17481, new_n17482, new_n17483, new_n17484, new_n17485,
    new_n17486, new_n17487, new_n17488, new_n17489, new_n17490, new_n17491,
    new_n17492, new_n17493, new_n17494, new_n17495, new_n17496, new_n17497,
    new_n17498, new_n17499, new_n17500, new_n17501, new_n17502, new_n17503,
    new_n17504, new_n17505, new_n17506, new_n17507, new_n17508, new_n17509,
    new_n17510, new_n17511, new_n17512, new_n17513, new_n17514, new_n17515,
    new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521,
    new_n17522, new_n17523, new_n17524, new_n17525, new_n17526, new_n17527,
    new_n17528, new_n17529, new_n17530, new_n17531, new_n17532, new_n17533,
    new_n17534, new_n17535, new_n17536, new_n17537, new_n17538, new_n17539,
    new_n17540, new_n17541, new_n17542, new_n17543, new_n17544, new_n17545,
    new_n17546, new_n17547, new_n17548, new_n17549, new_n17550, new_n17551,
    new_n17552, new_n17553, new_n17554, new_n17555, new_n17556, new_n17557,
    new_n17558, new_n17559, new_n17560, new_n17561, new_n17562, new_n17563,
    new_n17564, new_n17565, new_n17566, new_n17567, new_n17568, new_n17569,
    new_n17570, new_n17571, new_n17573, new_n17574, new_n17575, new_n17576,
    new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583, new_n17584, new_n17585, new_n17586, new_n17587, new_n17588,
    new_n17589, new_n17590, new_n17591, new_n17592, new_n17593, new_n17594,
    new_n17595, new_n17596, new_n17597, new_n17598, new_n17599, new_n17600,
    new_n17601, new_n17602, new_n17603, new_n17604, new_n17605, new_n17606,
    new_n17607, new_n17608, new_n17609, new_n17610, new_n17611, new_n17612,
    new_n17613, new_n17614, new_n17615, new_n17616, new_n17617, new_n17618,
    new_n17619, new_n17620, new_n17621, new_n17622, new_n17623, new_n17624,
    new_n17625, new_n17626, new_n17627, new_n17628, new_n17629, new_n17630,
    new_n17631, new_n17632, new_n17633, new_n17634, new_n17635, new_n17636,
    new_n17637, new_n17638, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648,
    new_n17649, new_n17650, new_n17651, new_n17652, new_n17653, new_n17654,
    new_n17655, new_n17656, new_n17657, new_n17658, new_n17659, new_n17660,
    new_n17661, new_n17662, new_n17663, new_n17664, new_n17665, new_n17666,
    new_n17667, new_n17668, new_n17669, new_n17670, new_n17671, new_n17672,
    new_n17673, new_n17674, new_n17675, new_n17676, new_n17677, new_n17678,
    new_n17679, new_n17680, new_n17681, new_n17682, new_n17683, new_n17684,
    new_n17685, new_n17686, new_n17687, new_n17688, new_n17689, new_n17690,
    new_n17691, new_n17692, new_n17693, new_n17694, new_n17695, new_n17696,
    new_n17697, new_n17698, new_n17699, new_n17700, new_n17701, new_n17702,
    new_n17703, new_n17704, new_n17705, new_n17706, new_n17707, new_n17708,
    new_n17709, new_n17710, new_n17711, new_n17712, new_n17713, new_n17714,
    new_n17715, new_n17716, new_n17717, new_n17718, new_n17719, new_n17720,
    new_n17721, new_n17722, new_n17723, new_n17724, new_n17725, new_n17726,
    new_n17727, new_n17728, new_n17729, new_n17730, new_n17731, new_n17732,
    new_n17733, new_n17734, new_n17735, new_n17736, new_n17737, new_n17738,
    new_n17739, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744,
    new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17807, new_n17808, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820, new_n17821, new_n17822, new_n17823,
    new_n17824, new_n17825, new_n17826, new_n17827, new_n17828, new_n17829,
    new_n17830, new_n17831, new_n17832, new_n17833, new_n17834, new_n17835,
    new_n17836, new_n17837, new_n17838, new_n17839, new_n17840, new_n17841,
    new_n17842, new_n17843, new_n17844, new_n17845, new_n17846, new_n17847,
    new_n17848, new_n17849, new_n17850, new_n17851, new_n17852, new_n17853,
    new_n17854, new_n17855, new_n17856, new_n17857, new_n17858, new_n17859,
    new_n17860, new_n17861, new_n17862, new_n17863, new_n17864, new_n17865,
    new_n17866, new_n17867, new_n17868, new_n17869, new_n17870, new_n17871,
    new_n17872, new_n17873, new_n17874, new_n17875, new_n17876, new_n17877,
    new_n17878, new_n17879, new_n17880, new_n17881, new_n17882, new_n17883,
    new_n17884, new_n17885, new_n17886, new_n17887, new_n17888, new_n17889,
    new_n17890, new_n17891, new_n17892, new_n17893, new_n17894, new_n17895,
    new_n17896, new_n17897, new_n17898, new_n17899, new_n17900, new_n17901,
    new_n17902, new_n17903, new_n17904, new_n17905, new_n17906, new_n17907,
    new_n17908, new_n17909, new_n17910, new_n17911, new_n17912, new_n17913,
    new_n17914, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919,
    new_n17920, new_n17921, new_n17922, new_n17923, new_n17924, new_n17925,
    new_n17926, new_n17927, new_n17928, new_n17929, new_n17930, new_n17931,
    new_n17932, new_n17933, new_n17934, new_n17935, new_n17936, new_n17937,
    new_n17938, new_n17939, new_n17940, new_n17941, new_n17942, new_n17943,
    new_n17944, new_n17945, new_n17946, new_n17947, new_n17948, new_n17949,
    new_n17950, new_n17951, new_n17952, new_n17953, new_n17954, new_n17955,
    new_n17956, new_n17957, new_n17958, new_n17959, new_n17960, new_n17961,
    new_n17962, new_n17963, new_n17964, new_n17965, new_n17966, new_n17967,
    new_n17968, new_n17969, new_n17970, new_n17971, new_n17972, new_n17973,
    new_n17974, new_n17975, new_n17976, new_n17977, new_n17978, new_n17979,
    new_n17980, new_n17981, new_n17982, new_n17983, new_n17984, new_n17985,
    new_n17986, new_n17987, new_n17988, new_n17989, new_n17990, new_n17991,
    new_n17992, new_n17993, new_n17994, new_n17995, new_n17996, new_n17997,
    new_n17998, new_n17999, new_n18000, new_n18001, new_n18002, new_n18003,
    new_n18004, new_n18005, new_n18006, new_n18007, new_n18008, new_n18009,
    new_n18010, new_n18011, new_n18012, new_n18013, new_n18014, new_n18015,
    new_n18016, new_n18017, new_n18018, new_n18019, new_n18020, new_n18021,
    new_n18022, new_n18023, new_n18024, new_n18025, new_n18026, new_n18027,
    new_n18028, new_n18029, new_n18030, new_n18031, new_n18032, new_n18033,
    new_n18034, new_n18035, new_n18036, new_n18037, new_n18038, new_n18039,
    new_n18040, new_n18041, new_n18042, new_n18043, new_n18044, new_n18045,
    new_n18047, new_n18048, new_n18049, new_n18050, new_n18051, new_n18052,
    new_n18053, new_n18054, new_n18055, new_n18056, new_n18057, new_n18058,
    new_n18059, new_n18060, new_n18061, new_n18062, new_n18063, new_n18064,
    new_n18065, new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071, new_n18072, new_n18073, new_n18074, new_n18075, new_n18076,
    new_n18077, new_n18078, new_n18079, new_n18080, new_n18081, new_n18082,
    new_n18083, new_n18084, new_n18085, new_n18086, new_n18087, new_n18088,
    new_n18089, new_n18090, new_n18091, new_n18092, new_n18093, new_n18094,
    new_n18095, new_n18096, new_n18097, new_n18098, new_n18099, new_n18100,
    new_n18101, new_n18102, new_n18103, new_n18104, new_n18105, new_n18106,
    new_n18107, new_n18108, new_n18109, new_n18110, new_n18111, new_n18112,
    new_n18113, new_n18114, new_n18115, new_n18116, new_n18117, new_n18118,
    new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124,
    new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130,
    new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136,
    new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143, new_n18144, new_n18145, new_n18146, new_n18147, new_n18148,
    new_n18149, new_n18150, new_n18151, new_n18152, new_n18153, new_n18154,
    new_n18155, new_n18156, new_n18157, new_n18158, new_n18159, new_n18160,
    new_n18161, new_n18162, new_n18163, new_n18164, new_n18165, new_n18166,
    new_n18167, new_n18168, new_n18169, new_n18170, new_n18171, new_n18172,
    new_n18173, new_n18174, new_n18175, new_n18176, new_n18177, new_n18178,
    new_n18179, new_n18180, new_n18181, new_n18182, new_n18183, new_n18184,
    new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190,
    new_n18191, new_n18192, new_n18193, new_n18194, new_n18195, new_n18196,
    new_n18197, new_n18198, new_n18199, new_n18200, new_n18201, new_n18202,
    new_n18203, new_n18204, new_n18205, new_n18206, new_n18207, new_n18208,
    new_n18209, new_n18210, new_n18211, new_n18212, new_n18213, new_n18214,
    new_n18215, new_n18216, new_n18217, new_n18218, new_n18219, new_n18220,
    new_n18221, new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227, new_n18228, new_n18229, new_n18230, new_n18231, new_n18232,
    new_n18233, new_n18234, new_n18235, new_n18236, new_n18237, new_n18238,
    new_n18239, new_n18240, new_n18241, new_n18242, new_n18243, new_n18244,
    new_n18245, new_n18246, new_n18247, new_n18248, new_n18249, new_n18250,
    new_n18251, new_n18252, new_n18253, new_n18254, new_n18255, new_n18256,
    new_n18257, new_n18258, new_n18259, new_n18260, new_n18261, new_n18262,
    new_n18263, new_n18264, new_n18265, new_n18266, new_n18267, new_n18268,
    new_n18269, new_n18270, new_n18271, new_n18272, new_n18273, new_n18274,
    new_n18275, new_n18276, new_n18278, new_n18279, new_n18280, new_n18281,
    new_n18282, new_n18283, new_n18284, new_n18285, new_n18286, new_n18287,
    new_n18288, new_n18289, new_n18290, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301, new_n18302, new_n18303, new_n18304, new_n18305,
    new_n18306, new_n18307, new_n18308, new_n18309, new_n18310, new_n18311,
    new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317,
    new_n18318, new_n18319, new_n18320, new_n18321, new_n18322, new_n18323,
    new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329,
    new_n18330, new_n18331, new_n18332, new_n18333, new_n18334, new_n18335,
    new_n18336, new_n18337, new_n18338, new_n18339, new_n18340, new_n18341,
    new_n18342, new_n18343, new_n18344, new_n18345, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362, new_n18363, new_n18364, new_n18365,
    new_n18366, new_n18367, new_n18368, new_n18369, new_n18370, new_n18371,
    new_n18372, new_n18373, new_n18374, new_n18375, new_n18376, new_n18377,
    new_n18378, new_n18379, new_n18380, new_n18381, new_n18382, new_n18383,
    new_n18384, new_n18385, new_n18386, new_n18387, new_n18388, new_n18389,
    new_n18390, new_n18391, new_n18392, new_n18393, new_n18394, new_n18395,
    new_n18396, new_n18397, new_n18398, new_n18399, new_n18400, new_n18401,
    new_n18402, new_n18403, new_n18404, new_n18405, new_n18406, new_n18407,
    new_n18408, new_n18409, new_n18410, new_n18411, new_n18412, new_n18413,
    new_n18414, new_n18415, new_n18416, new_n18417, new_n18418, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436, new_n18437,
    new_n18438, new_n18439, new_n18440, new_n18441, new_n18442, new_n18443,
    new_n18444, new_n18445, new_n18446, new_n18447, new_n18448, new_n18449,
    new_n18450, new_n18451, new_n18452, new_n18453, new_n18454, new_n18455,
    new_n18456, new_n18457, new_n18458, new_n18459, new_n18460, new_n18461,
    new_n18462, new_n18463, new_n18464, new_n18465, new_n18466, new_n18467,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482, new_n18483, new_n18484, new_n18485,
    new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491,
    new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497,
    new_n18499, new_n18500, new_n18501, new_n18502, new_n18503, new_n18504,
    new_n18505, new_n18506, new_n18507, new_n18508, new_n18509, new_n18510,
    new_n18511, new_n18512, new_n18513, new_n18514, new_n18515, new_n18516,
    new_n18517, new_n18518, new_n18519, new_n18520, new_n18521, new_n18522,
    new_n18523, new_n18524, new_n18525, new_n18526, new_n18527, new_n18528,
    new_n18529, new_n18530, new_n18531, new_n18532, new_n18533, new_n18534,
    new_n18535, new_n18536, new_n18537, new_n18538, new_n18539, new_n18540,
    new_n18541, new_n18542, new_n18543, new_n18544, new_n18545, new_n18546,
    new_n18547, new_n18548, new_n18549, new_n18550, new_n18551, new_n18552,
    new_n18553, new_n18554, new_n18555, new_n18556, new_n18557, new_n18558,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18570,
    new_n18571, new_n18572, new_n18573, new_n18574, new_n18575, new_n18576,
    new_n18577, new_n18578, new_n18579, new_n18580, new_n18581, new_n18582,
    new_n18583, new_n18584, new_n18585, new_n18586, new_n18587, new_n18588,
    new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594,
    new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600,
    new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18606,
    new_n18607, new_n18608, new_n18609, new_n18610, new_n18611, new_n18612,
    new_n18613, new_n18614, new_n18615, new_n18616, new_n18617, new_n18618,
    new_n18619, new_n18620, new_n18621, new_n18622, new_n18623, new_n18624,
    new_n18625, new_n18626, new_n18627, new_n18628, new_n18629, new_n18630,
    new_n18631, new_n18632, new_n18633, new_n18634, new_n18635, new_n18636,
    new_n18637, new_n18638, new_n18639, new_n18640, new_n18641, new_n18642,
    new_n18643, new_n18644, new_n18645, new_n18646, new_n18647, new_n18648,
    new_n18649, new_n18650, new_n18651, new_n18652, new_n18653, new_n18654,
    new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18711, new_n18712, new_n18713, new_n18714, new_n18715,
    new_n18716, new_n18717, new_n18718, new_n18719, new_n18720, new_n18721,
    new_n18722, new_n18723, new_n18724, new_n18725, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18734, new_n18735, new_n18736, new_n18737, new_n18738, new_n18739,
    new_n18740, new_n18741, new_n18742, new_n18743, new_n18744, new_n18745,
    new_n18746, new_n18747, new_n18748, new_n18749, new_n18750, new_n18751,
    new_n18752, new_n18753, new_n18754, new_n18755, new_n18756, new_n18757,
    new_n18758, new_n18759, new_n18760, new_n18761, new_n18762, new_n18763,
    new_n18764, new_n18765, new_n18766, new_n18767, new_n18768, new_n18769,
    new_n18770, new_n18771, new_n18772, new_n18773, new_n18774, new_n18775,
    new_n18776, new_n18777, new_n18778, new_n18779, new_n18780, new_n18781,
    new_n18782, new_n18783, new_n18784, new_n18785, new_n18786, new_n18787,
    new_n18788, new_n18789, new_n18790, new_n18791, new_n18792, new_n18793,
    new_n18794, new_n18795, new_n18796, new_n18797, new_n18798, new_n18799,
    new_n18800, new_n18801, new_n18802, new_n18803, new_n18804, new_n18805,
    new_n18806, new_n18807, new_n18808, new_n18809, new_n18810, new_n18811,
    new_n18812, new_n18813, new_n18814, new_n18815, new_n18816, new_n18817,
    new_n18818, new_n18819, new_n18820, new_n18821, new_n18822, new_n18823,
    new_n18824, new_n18825, new_n18826, new_n18827, new_n18828, new_n18829,
    new_n18830, new_n18831, new_n18832, new_n18833, new_n18834, new_n18835,
    new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843, new_n18844, new_n18845, new_n18846, new_n18847,
    new_n18848, new_n18849, new_n18850, new_n18851, new_n18852, new_n18853,
    new_n18854, new_n18855, new_n18856, new_n18857, new_n18858, new_n18859,
    new_n18860, new_n18861, new_n18862, new_n18863, new_n18864, new_n18865,
    new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871,
    new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877,
    new_n18878, new_n18879, new_n18880, new_n18881, new_n18882, new_n18883,
    new_n18884, new_n18885, new_n18886, new_n18887, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900, new_n18901,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906, new_n18907,
    new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18913,
    new_n18914, new_n18915, new_n18916, new_n18917, new_n18918, new_n18919,
    new_n18920, new_n18921, new_n18922, new_n18923, new_n18924, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962,
    new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968,
    new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004,
    new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010,
    new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016,
    new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022,
    new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028,
    new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058,
    new_n19059, new_n19060, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112,
    new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130,
    new_n19132, new_n19133, new_n19134, new_n19135, new_n19136, new_n19137,
    new_n19138, new_n19139, new_n19140, new_n19141, new_n19142, new_n19143,
    new_n19144, new_n19145, new_n19146, new_n19147, new_n19148, new_n19149,
    new_n19150, new_n19151, new_n19152, new_n19153, new_n19154, new_n19155,
    new_n19156, new_n19157, new_n19158, new_n19159, new_n19160, new_n19161,
    new_n19162, new_n19163, new_n19164, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174, new_n19175, new_n19176, new_n19177, new_n19178, new_n19179,
    new_n19180, new_n19181, new_n19182, new_n19183, new_n19184, new_n19185,
    new_n19186, new_n19187, new_n19188, new_n19189, new_n19190, new_n19191,
    new_n19192, new_n19193, new_n19194, new_n19195, new_n19196, new_n19197,
    new_n19198, new_n19199, new_n19200, new_n19201, new_n19202, new_n19203,
    new_n19204, new_n19205, new_n19206, new_n19207, new_n19208, new_n19209,
    new_n19210, new_n19211, new_n19212, new_n19213, new_n19214, new_n19215,
    new_n19216, new_n19217, new_n19218, new_n19219, new_n19220, new_n19221,
    new_n19222, new_n19223, new_n19224, new_n19225, new_n19226, new_n19227,
    new_n19228, new_n19229, new_n19230, new_n19231, new_n19232, new_n19233,
    new_n19234, new_n19235, new_n19236, new_n19237, new_n19238, new_n19239,
    new_n19240, new_n19241, new_n19242, new_n19243, new_n19244, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263,
    new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270, new_n19271, new_n19272, new_n19273, new_n19274, new_n19275,
    new_n19276, new_n19277, new_n19278, new_n19279, new_n19280, new_n19281,
    new_n19282, new_n19283, new_n19284, new_n19285, new_n19286, new_n19287,
    new_n19288, new_n19289, new_n19290, new_n19291, new_n19292, new_n19293,
    new_n19294, new_n19295, new_n19296, new_n19297, new_n19298, new_n19299,
    new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305,
    new_n19306, new_n19307, new_n19308, new_n19309, new_n19310, new_n19311,
    new_n19312, new_n19313, new_n19314, new_n19315, new_n19316, new_n19317,
    new_n19318, new_n19319, new_n19320, new_n19321, new_n19322, new_n19323,
    new_n19324, new_n19325, new_n19326, new_n19327, new_n19328, new_n19329,
    new_n19330, new_n19331, new_n19332, new_n19334, new_n19335, new_n19336,
    new_n19337, new_n19338, new_n19339, new_n19340, new_n19341, new_n19342,
    new_n19343, new_n19344, new_n19345, new_n19346, new_n19347, new_n19348,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353, new_n19354,
    new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360,
    new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367, new_n19368, new_n19369, new_n19370, new_n19371, new_n19372,
    new_n19373, new_n19374, new_n19375, new_n19376, new_n19377, new_n19378,
    new_n19379, new_n19380, new_n19381, new_n19382, new_n19383, new_n19384,
    new_n19385, new_n19386, new_n19387, new_n19388, new_n19389, new_n19390,
    new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396,
    new_n19397, new_n19398, new_n19399, new_n19400, new_n19401, new_n19402,
    new_n19403, new_n19404, new_n19405, new_n19406, new_n19407, new_n19408,
    new_n19409, new_n19410, new_n19411, new_n19412, new_n19413, new_n19414,
    new_n19415, new_n19416, new_n19417, new_n19418, new_n19419, new_n19420,
    new_n19421, new_n19422, new_n19423, new_n19424, new_n19425, new_n19426,
    new_n19427, new_n19428, new_n19429, new_n19430, new_n19431, new_n19432,
    new_n19433, new_n19434, new_n19435, new_n19436, new_n19437, new_n19438,
    new_n19439, new_n19440, new_n19441, new_n19442, new_n19443, new_n19444,
    new_n19445, new_n19446, new_n19447, new_n19448, new_n19449, new_n19450,
    new_n19451, new_n19452, new_n19453, new_n19454, new_n19455, new_n19456,
    new_n19457, new_n19458, new_n19459, new_n19460, new_n19461, new_n19462,
    new_n19463, new_n19464, new_n19465, new_n19466, new_n19467, new_n19468,
    new_n19469, new_n19470, new_n19471, new_n19472, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477, new_n19478, new_n19479, new_n19480,
    new_n19481, new_n19482, new_n19483, new_n19484, new_n19485, new_n19486,
    new_n19487, new_n19488, new_n19489, new_n19490, new_n19491, new_n19492,
    new_n19493, new_n19494, new_n19495, new_n19496, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19514, new_n19515, new_n19516,
    new_n19517, new_n19518, new_n19519, new_n19520, new_n19521, new_n19522,
    new_n19523, new_n19524, new_n19525, new_n19526, new_n19527, new_n19528,
    new_n19529, new_n19530, new_n19531, new_n19532, new_n19533, new_n19534,
    new_n19535, new_n19536, new_n19537, new_n19538, new_n19539, new_n19540,
    new_n19541, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547,
    new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553,
    new_n19554, new_n19555, new_n19556, new_n19557, new_n19558, new_n19559,
    new_n19560, new_n19561, new_n19562, new_n19563, new_n19564, new_n19565,
    new_n19566, new_n19567, new_n19568, new_n19569, new_n19570, new_n19571,
    new_n19572, new_n19573, new_n19574, new_n19575, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584, new_n19585, new_n19586, new_n19587, new_n19588, new_n19589,
    new_n19590, new_n19591, new_n19592, new_n19593, new_n19594, new_n19595,
    new_n19596, new_n19597, new_n19598, new_n19599, new_n19600, new_n19601,
    new_n19602, new_n19603, new_n19604, new_n19605, new_n19606, new_n19607,
    new_n19608, new_n19609, new_n19610, new_n19611, new_n19612, new_n19613,
    new_n19614, new_n19615, new_n19616, new_n19617, new_n19618, new_n19619,
    new_n19620, new_n19621, new_n19622, new_n19623, new_n19624, new_n19625,
    new_n19626, new_n19627, new_n19628, new_n19629, new_n19630, new_n19631,
    new_n19632, new_n19633, new_n19634, new_n19635, new_n19636, new_n19637,
    new_n19638, new_n19639, new_n19640, new_n19641, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648, new_n19649,
    new_n19650, new_n19651, new_n19652, new_n19653, new_n19654, new_n19655,
    new_n19656, new_n19657, new_n19658, new_n19659, new_n19660, new_n19661,
    new_n19662, new_n19663, new_n19664, new_n19665, new_n19666, new_n19667,
    new_n19668, new_n19669, new_n19670, new_n19671, new_n19672, new_n19673,
    new_n19674, new_n19675, new_n19676, new_n19677, new_n19678, new_n19679,
    new_n19680, new_n19681, new_n19682, new_n19683, new_n19684, new_n19685,
    new_n19686, new_n19687, new_n19688, new_n19689, new_n19690, new_n19691,
    new_n19692, new_n19693, new_n19694, new_n19695, new_n19696, new_n19697,
    new_n19698, new_n19699, new_n19700, new_n19701, new_n19702, new_n19703,
    new_n19704, new_n19705, new_n19706, new_n19707, new_n19708, new_n19709,
    new_n19710, new_n19711, new_n19712, new_n19713, new_n19714, new_n19715,
    new_n19716, new_n19717, new_n19718, new_n19719, new_n19720, new_n19721,
    new_n19722, new_n19723, new_n19724, new_n19725, new_n19726, new_n19727,
    new_n19728, new_n19729, new_n19730, new_n19731, new_n19732, new_n19734,
    new_n19735, new_n19736, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749, new_n19750, new_n19751, new_n19752,
    new_n19753, new_n19754, new_n19755, new_n19756, new_n19757, new_n19758,
    new_n19759, new_n19760, new_n19761, new_n19762, new_n19763, new_n19764,
    new_n19765, new_n19766, new_n19767, new_n19768, new_n19769, new_n19770,
    new_n19771, new_n19772, new_n19773, new_n19774, new_n19775, new_n19776,
    new_n19777, new_n19778, new_n19779, new_n19780, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789, new_n19790, new_n19791, new_n19792, new_n19793, new_n19794,
    new_n19795, new_n19796, new_n19797, new_n19798, new_n19799, new_n19800,
    new_n19801, new_n19802, new_n19803, new_n19804, new_n19805, new_n19806,
    new_n19807, new_n19808, new_n19809, new_n19810, new_n19811, new_n19812,
    new_n19813, new_n19814, new_n19815, new_n19816, new_n19817, new_n19818,
    new_n19819, new_n19820, new_n19821, new_n19822, new_n19823, new_n19824,
    new_n19825, new_n19826, new_n19827, new_n19828, new_n19829, new_n19830,
    new_n19831, new_n19832, new_n19833, new_n19834, new_n19835, new_n19836,
    new_n19837, new_n19838, new_n19839, new_n19840, new_n19841, new_n19842,
    new_n19843, new_n19844, new_n19845, new_n19846, new_n19847, new_n19848,
    new_n19849, new_n19850, new_n19851, new_n19852, new_n19853, new_n19854,
    new_n19855, new_n19856, new_n19857, new_n19858, new_n19859, new_n19860,
    new_n19861, new_n19862, new_n19863, new_n19864, new_n19865, new_n19866,
    new_n19867, new_n19868, new_n19869, new_n19870, new_n19871, new_n19872,
    new_n19873, new_n19874, new_n19875, new_n19876, new_n19877, new_n19878,
    new_n19879, new_n19880, new_n19881, new_n19882, new_n19883, new_n19884,
    new_n19885, new_n19886, new_n19887, new_n19888, new_n19889, new_n19890,
    new_n19891, new_n19892, new_n19893, new_n19894, new_n19895, new_n19896,
    new_n19897, new_n19898, new_n19899, new_n19900, new_n19901, new_n19902,
    new_n19903, new_n19904, new_n19905, new_n19906, new_n19907, new_n19908,
    new_n19909, new_n19910, new_n19911, new_n19912, new_n19914, new_n19915,
    new_n19916, new_n19917, new_n19918, new_n19919, new_n19920, new_n19921,
    new_n19922, new_n19923, new_n19924, new_n19925, new_n19926, new_n19927,
    new_n19928, new_n19929, new_n19930, new_n19931, new_n19932, new_n19933,
    new_n19934, new_n19935, new_n19936, new_n19937, new_n19938, new_n19939,
    new_n19940, new_n19941, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951,
    new_n19952, new_n19953, new_n19954, new_n19955, new_n19956, new_n19957,
    new_n19958, new_n19959, new_n19960, new_n19961, new_n19962, new_n19963,
    new_n19964, new_n19965, new_n19966, new_n19967, new_n19968, new_n19969,
    new_n19970, new_n19971, new_n19972, new_n19973, new_n19974, new_n19975,
    new_n19976, new_n19977, new_n19978, new_n19979, new_n19980, new_n19981,
    new_n19982, new_n19983, new_n19984, new_n19985, new_n19986, new_n19987,
    new_n19988, new_n19989, new_n19990, new_n19991, new_n19992, new_n19993,
    new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999,
    new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005,
    new_n20006, new_n20007, new_n20008, new_n20009, new_n20010, new_n20011,
    new_n20012, new_n20013, new_n20014, new_n20015, new_n20016, new_n20017,
    new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023,
    new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029,
    new_n20030, new_n20031, new_n20032, new_n20033, new_n20034, new_n20035,
    new_n20036, new_n20037, new_n20038, new_n20039, new_n20040, new_n20041,
    new_n20042, new_n20043, new_n20044, new_n20045, new_n20046, new_n20047,
    new_n20048, new_n20049, new_n20050, new_n20051, new_n20052, new_n20053,
    new_n20054, new_n20055, new_n20056, new_n20057, new_n20058, new_n20059,
    new_n20060, new_n20061, new_n20062, new_n20063, new_n20064, new_n20065,
    new_n20066, new_n20067, new_n20068, new_n20069, new_n20070, new_n20071,
    new_n20072, new_n20073, new_n20074, new_n20075, new_n20076, new_n20077,
    new_n20078, new_n20079, new_n20080, new_n20081, new_n20082, new_n20083,
    new_n20084, new_n20085, new_n20086, new_n20087, new_n20088, new_n20089,
    new_n20090, new_n20091, new_n20092, new_n20093, new_n20094, new_n20095,
    new_n20096, new_n20097, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162,
    new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169, new_n20170, new_n20171, new_n20172, new_n20173, new_n20174,
    new_n20175, new_n20176, new_n20177, new_n20178, new_n20179, new_n20180,
    new_n20181, new_n20182, new_n20183, new_n20184, new_n20185, new_n20186,
    new_n20187, new_n20188, new_n20189, new_n20190, new_n20191, new_n20192,
    new_n20193, new_n20194, new_n20195, new_n20196, new_n20197, new_n20198,
    new_n20199, new_n20200, new_n20201, new_n20202, new_n20203, new_n20204,
    new_n20205, new_n20206, new_n20207, new_n20208, new_n20209, new_n20210,
    new_n20211, new_n20212, new_n20213, new_n20214, new_n20215, new_n20216,
    new_n20217, new_n20218, new_n20219, new_n20220, new_n20221, new_n20222,
    new_n20223, new_n20224, new_n20225, new_n20226, new_n20227, new_n20228,
    new_n20229, new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235, new_n20236, new_n20237, new_n20238, new_n20239, new_n20240,
    new_n20241, new_n20242, new_n20243, new_n20244, new_n20245, new_n20246,
    new_n20247, new_n20248, new_n20249, new_n20250, new_n20251, new_n20252,
    new_n20253, new_n20254, new_n20255, new_n20256, new_n20257, new_n20258,
    new_n20259, new_n20260, new_n20261, new_n20262, new_n20263, new_n20264,
    new_n20265, new_n20266, new_n20267, new_n20268, new_n20269, new_n20270,
    new_n20271, new_n20272, new_n20273, new_n20274, new_n20275, new_n20276,
    new_n20277, new_n20278, new_n20279, new_n20280, new_n20281, new_n20282,
    new_n20283, new_n20284, new_n20285, new_n20287, new_n20288, new_n20289,
    new_n20290, new_n20291, new_n20292, new_n20293, new_n20294, new_n20295,
    new_n20296, new_n20297, new_n20298, new_n20299, new_n20300, new_n20301,
    new_n20302, new_n20303, new_n20304, new_n20305, new_n20306, new_n20307,
    new_n20308, new_n20309, new_n20310, new_n20311, new_n20312, new_n20313,
    new_n20314, new_n20315, new_n20316, new_n20317, new_n20318, new_n20319,
    new_n20320, new_n20321, new_n20322, new_n20323, new_n20324, new_n20325,
    new_n20326, new_n20327, new_n20328, new_n20329, new_n20330, new_n20331,
    new_n20332, new_n20333, new_n20334, new_n20335, new_n20336, new_n20337,
    new_n20338, new_n20339, new_n20340, new_n20341, new_n20342, new_n20343,
    new_n20344, new_n20345, new_n20346, new_n20347, new_n20348, new_n20349,
    new_n20350, new_n20351, new_n20352, new_n20353, new_n20354, new_n20355,
    new_n20356, new_n20357, new_n20358, new_n20359, new_n20360, new_n20361,
    new_n20362, new_n20363, new_n20364, new_n20365, new_n20366, new_n20367,
    new_n20368, new_n20369, new_n20370, new_n20371, new_n20372, new_n20373,
    new_n20374, new_n20375, new_n20376, new_n20377, new_n20378, new_n20379,
    new_n20380, new_n20381, new_n20382, new_n20383, new_n20384, new_n20385,
    new_n20386, new_n20387, new_n20388, new_n20389, new_n20390, new_n20391,
    new_n20392, new_n20393, new_n20394, new_n20395, new_n20396, new_n20397,
    new_n20398, new_n20399, new_n20400, new_n20401, new_n20402, new_n20403,
    new_n20404, new_n20405, new_n20406, new_n20407, new_n20408, new_n20409,
    new_n20410, new_n20411, new_n20412, new_n20413, new_n20414, new_n20415,
    new_n20416, new_n20417, new_n20418, new_n20419, new_n20420, new_n20421,
    new_n20422, new_n20423, new_n20424, new_n20425, new_n20426, new_n20427,
    new_n20428, new_n20429, new_n20430, new_n20431, new_n20432, new_n20433,
    new_n20434, new_n20435, new_n20436, new_n20437, new_n20438, new_n20439,
    new_n20440, new_n20441, new_n20442, new_n20443, new_n20444, new_n20445,
    new_n20446, new_n20447, new_n20448, new_n20449, new_n20450, new_n20451,
    new_n20452, new_n20453, new_n20454, new_n20455, new_n20456, new_n20457,
    new_n20458, new_n20459, new_n20460, new_n20461, new_n20462, new_n20463,
    new_n20464, new_n20465, new_n20466, new_n20467, new_n20468, new_n20469,
    new_n20470, new_n20471, new_n20472, new_n20473, new_n20474, new_n20475,
    new_n20477, new_n20478, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489, new_n20490, new_n20491, new_n20492, new_n20493, new_n20494,
    new_n20495, new_n20496, new_n20497, new_n20498, new_n20499, new_n20500,
    new_n20501, new_n20502, new_n20503, new_n20504, new_n20505, new_n20506,
    new_n20507, new_n20508, new_n20509, new_n20510, new_n20511, new_n20512,
    new_n20513, new_n20514, new_n20515, new_n20516, new_n20517, new_n20518,
    new_n20519, new_n20520, new_n20521, new_n20522, new_n20523, new_n20524,
    new_n20525, new_n20526, new_n20527, new_n20528, new_n20529, new_n20530,
    new_n20531, new_n20532, new_n20533, new_n20534, new_n20535, new_n20536,
    new_n20537, new_n20538, new_n20539, new_n20540, new_n20541, new_n20542,
    new_n20543, new_n20544, new_n20545, new_n20546, new_n20547, new_n20548,
    new_n20549, new_n20550, new_n20551, new_n20552, new_n20553, new_n20554,
    new_n20555, new_n20556, new_n20557, new_n20558, new_n20559, new_n20560,
    new_n20561, new_n20562, new_n20563, new_n20564, new_n20565, new_n20566,
    new_n20567, new_n20568, new_n20569, new_n20570, new_n20571, new_n20572,
    new_n20573, new_n20574, new_n20575, new_n20576, new_n20577, new_n20578,
    new_n20579, new_n20580, new_n20581, new_n20582, new_n20583, new_n20584,
    new_n20585, new_n20586, new_n20587, new_n20588, new_n20589, new_n20590,
    new_n20591, new_n20592, new_n20593, new_n20594, new_n20595, new_n20596,
    new_n20597, new_n20598, new_n20599, new_n20600, new_n20601, new_n20602,
    new_n20603, new_n20604, new_n20605, new_n20606, new_n20607, new_n20608,
    new_n20609, new_n20610, new_n20611, new_n20612, new_n20613, new_n20614,
    new_n20615, new_n20616, new_n20617, new_n20618, new_n20619, new_n20620,
    new_n20621, new_n20622, new_n20623, new_n20624, new_n20625, new_n20626,
    new_n20627, new_n20628, new_n20629, new_n20630, new_n20631, new_n20632,
    new_n20633, new_n20634, new_n20635, new_n20636, new_n20637, new_n20638,
    new_n20639, new_n20640, new_n20641, new_n20642, new_n20643, new_n20644,
    new_n20645, new_n20646, new_n20647, new_n20648, new_n20649, new_n20650,
    new_n20651, new_n20652, new_n20653, new_n20655, new_n20656, new_n20657,
    new_n20658, new_n20659, new_n20660, new_n20661, new_n20662, new_n20663,
    new_n20664, new_n20665, new_n20666, new_n20667, new_n20668, new_n20669,
    new_n20670, new_n20671, new_n20672, new_n20673, new_n20674, new_n20675,
    new_n20676, new_n20677, new_n20678, new_n20679, new_n20680, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685, new_n20686, new_n20687,
    new_n20688, new_n20689, new_n20690, new_n20691, new_n20692, new_n20693,
    new_n20694, new_n20695, new_n20696, new_n20697, new_n20698, new_n20699,
    new_n20700, new_n20701, new_n20702, new_n20703, new_n20704, new_n20705,
    new_n20706, new_n20707, new_n20708, new_n20709, new_n20710, new_n20711,
    new_n20712, new_n20713, new_n20714, new_n20715, new_n20716, new_n20717,
    new_n20718, new_n20719, new_n20720, new_n20721, new_n20722, new_n20723,
    new_n20724, new_n20725, new_n20726, new_n20727, new_n20728, new_n20729,
    new_n20730, new_n20731, new_n20732, new_n20733, new_n20734, new_n20735,
    new_n20736, new_n20737, new_n20738, new_n20739, new_n20740, new_n20741,
    new_n20742, new_n20743, new_n20744, new_n20745, new_n20746, new_n20747,
    new_n20748, new_n20749, new_n20750, new_n20751, new_n20752, new_n20753,
    new_n20754, new_n20755, new_n20756, new_n20757, new_n20758, new_n20759,
    new_n20760, new_n20761, new_n20762, new_n20763, new_n20764, new_n20765,
    new_n20766, new_n20767, new_n20768, new_n20769, new_n20770, new_n20771,
    new_n20772, new_n20773, new_n20774, new_n20775, new_n20776, new_n20777,
    new_n20778, new_n20779, new_n20780, new_n20781, new_n20782, new_n20783,
    new_n20784, new_n20785, new_n20786, new_n20787, new_n20788, new_n20789,
    new_n20790, new_n20791, new_n20792, new_n20793, new_n20794, new_n20795,
    new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801,
    new_n20802, new_n20803, new_n20804, new_n20805, new_n20806, new_n20807,
    new_n20808, new_n20809, new_n20810, new_n20811, new_n20812, new_n20813,
    new_n20814, new_n20815, new_n20816, new_n20817, new_n20818, new_n20819,
    new_n20820, new_n20821, new_n20822, new_n20823, new_n20824, new_n20825,
    new_n20826, new_n20827, new_n20828, new_n20829, new_n20830, new_n20831,
    new_n20832, new_n20833, new_n20834, new_n20836, new_n20837, new_n20838,
    new_n20839, new_n20840, new_n20841, new_n20842, new_n20843, new_n20844,
    new_n20845, new_n20846, new_n20847, new_n20848, new_n20849, new_n20850,
    new_n20851, new_n20852, new_n20853, new_n20854, new_n20855, new_n20856,
    new_n20857, new_n20858, new_n20859, new_n20860, new_n20861, new_n20862,
    new_n20863, new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869, new_n20870, new_n20871, new_n20872, new_n20873, new_n20874,
    new_n20875, new_n20876, new_n20877, new_n20878, new_n20879, new_n20880,
    new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898,
    new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904,
    new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910,
    new_n20911, new_n20912, new_n20913, new_n20914, new_n20915, new_n20916,
    new_n20917, new_n20918, new_n20919, new_n20920, new_n20921, new_n20922,
    new_n20923, new_n20924, new_n20925, new_n20926, new_n20927, new_n20928,
    new_n20929, new_n20930, new_n20931, new_n20932, new_n20933, new_n20934,
    new_n20935, new_n20936, new_n20937, new_n20938, new_n20939, new_n20940,
    new_n20941, new_n20942, new_n20943, new_n20944, new_n20945, new_n20946,
    new_n20947, new_n20948, new_n20949, new_n20950, new_n20951, new_n20952,
    new_n20953, new_n20954, new_n20955, new_n20956, new_n20957, new_n20958,
    new_n20959, new_n20960, new_n20961, new_n20962, new_n20963, new_n20964,
    new_n20965, new_n20966, new_n20967, new_n20968, new_n20969, new_n20970,
    new_n20971, new_n20972, new_n20973, new_n20974, new_n20975, new_n20976,
    new_n20977, new_n20978, new_n20979, new_n20980, new_n20981, new_n20982,
    new_n20983, new_n20984, new_n20985, new_n20986, new_n20987, new_n20988,
    new_n20989, new_n20990, new_n20991, new_n20992, new_n20993, new_n20994,
    new_n20995, new_n20996, new_n20997, new_n20998, new_n20999, new_n21000,
    new_n21001, new_n21002, new_n21003, new_n21004, new_n21006, new_n21007,
    new_n21008, new_n21009, new_n21010, new_n21011, new_n21012, new_n21013,
    new_n21014, new_n21015, new_n21016, new_n21017, new_n21018, new_n21019,
    new_n21020, new_n21021, new_n21022, new_n21023, new_n21024, new_n21025,
    new_n21026, new_n21027, new_n21028, new_n21029, new_n21030, new_n21031,
    new_n21032, new_n21033, new_n21034, new_n21035, new_n21036, new_n21037,
    new_n21038, new_n21039, new_n21040, new_n21041, new_n21042, new_n21043,
    new_n21044, new_n21045, new_n21046, new_n21047, new_n21048, new_n21049,
    new_n21050, new_n21051, new_n21052, new_n21053, new_n21054, new_n21055,
    new_n21056, new_n21057, new_n21058, new_n21059, new_n21060, new_n21061,
    new_n21062, new_n21063, new_n21064, new_n21065, new_n21066, new_n21067,
    new_n21068, new_n21069, new_n21070, new_n21071, new_n21072, new_n21073,
    new_n21074, new_n21075, new_n21076, new_n21077, new_n21078, new_n21079,
    new_n21080, new_n21081, new_n21082, new_n21083, new_n21084, new_n21085,
    new_n21086, new_n21087, new_n21088, new_n21089, new_n21090, new_n21091,
    new_n21092, new_n21093, new_n21094, new_n21095, new_n21096, new_n21097,
    new_n21098, new_n21099, new_n21100, new_n21101, new_n21102, new_n21103,
    new_n21104, new_n21105, new_n21106, new_n21107, new_n21108, new_n21109,
    new_n21110, new_n21111, new_n21112, new_n21113, new_n21114, new_n21115,
    new_n21116, new_n21117, new_n21118, new_n21119, new_n21120, new_n21121,
    new_n21122, new_n21123, new_n21124, new_n21125, new_n21126, new_n21127,
    new_n21128, new_n21129, new_n21130, new_n21131, new_n21132, new_n21133,
    new_n21134, new_n21135, new_n21136, new_n21137, new_n21138, new_n21139,
    new_n21140, new_n21141, new_n21142, new_n21143, new_n21144, new_n21145,
    new_n21146, new_n21147, new_n21148, new_n21149, new_n21150, new_n21151,
    new_n21152, new_n21153, new_n21154, new_n21155, new_n21156, new_n21157,
    new_n21158, new_n21159, new_n21160, new_n21161, new_n21162, new_n21163,
    new_n21164, new_n21165, new_n21167, new_n21168, new_n21169, new_n21170,
    new_n21171, new_n21172, new_n21173, new_n21174, new_n21175, new_n21176,
    new_n21177, new_n21178, new_n21179, new_n21180, new_n21181, new_n21182,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203, new_n21204, new_n21205, new_n21206,
    new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212,
    new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218,
    new_n21219, new_n21220, new_n21221, new_n21222, new_n21223, new_n21224,
    new_n21225, new_n21226, new_n21227, new_n21228, new_n21229, new_n21230,
    new_n21231, new_n21232, new_n21233, new_n21234, new_n21235, new_n21236,
    new_n21237, new_n21238, new_n21239, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248,
    new_n21249, new_n21250, new_n21251, new_n21252, new_n21253, new_n21254,
    new_n21255, new_n21256, new_n21257, new_n21258, new_n21259, new_n21260,
    new_n21261, new_n21262, new_n21263, new_n21264, new_n21265, new_n21266,
    new_n21267, new_n21268, new_n21269, new_n21270, new_n21271, new_n21272,
    new_n21273, new_n21274, new_n21275, new_n21276, new_n21277, new_n21278,
    new_n21279, new_n21280, new_n21281, new_n21282, new_n21283, new_n21284,
    new_n21285, new_n21286, new_n21287, new_n21288, new_n21289, new_n21290,
    new_n21291, new_n21292, new_n21293, new_n21294, new_n21295, new_n21296,
    new_n21297, new_n21298, new_n21299, new_n21300, new_n21301, new_n21302,
    new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308,
    new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314,
    new_n21315, new_n21316, new_n21317, new_n21318, new_n21319, new_n21320,
    new_n21321, new_n21322, new_n21323, new_n21324, new_n21325, new_n21326,
    new_n21328, new_n21329, new_n21330, new_n21331, new_n21332, new_n21333,
    new_n21334, new_n21335, new_n21336, new_n21337, new_n21338, new_n21339,
    new_n21340, new_n21341, new_n21342, new_n21343, new_n21344, new_n21345,
    new_n21346, new_n21347, new_n21348, new_n21349, new_n21350, new_n21351,
    new_n21352, new_n21353, new_n21354, new_n21355, new_n21356, new_n21357,
    new_n21358, new_n21359, new_n21360, new_n21361, new_n21362, new_n21363,
    new_n21364, new_n21365, new_n21366, new_n21367, new_n21368, new_n21369,
    new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375,
    new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381,
    new_n21382, new_n21383, new_n21384, new_n21385, new_n21386, new_n21387,
    new_n21388, new_n21389, new_n21390, new_n21391, new_n21392, new_n21393,
    new_n21394, new_n21395, new_n21396, new_n21397, new_n21398, new_n21399,
    new_n21400, new_n21401, new_n21402, new_n21403, new_n21404, new_n21405,
    new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411,
    new_n21412, new_n21413, new_n21414, new_n21415, new_n21416, new_n21417,
    new_n21418, new_n21419, new_n21420, new_n21421, new_n21422, new_n21423,
    new_n21424, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21444, new_n21445, new_n21446, new_n21447,
    new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453,
    new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459,
    new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21465,
    new_n21466, new_n21467, new_n21468, new_n21469, new_n21470, new_n21471,
    new_n21472, new_n21473, new_n21474, new_n21475, new_n21476, new_n21477,
    new_n21478, new_n21479, new_n21481, new_n21482, new_n21483, new_n21484,
    new_n21485, new_n21486, new_n21487, new_n21488, new_n21489, new_n21490,
    new_n21491, new_n21492, new_n21493, new_n21494, new_n21495, new_n21496,
    new_n21497, new_n21498, new_n21499, new_n21500, new_n21501, new_n21502,
    new_n21503, new_n21504, new_n21505, new_n21506, new_n21507, new_n21508,
    new_n21509, new_n21510, new_n21511, new_n21512, new_n21513, new_n21514,
    new_n21515, new_n21516, new_n21517, new_n21518, new_n21519, new_n21520,
    new_n21521, new_n21522, new_n21523, new_n21524, new_n21525, new_n21526,
    new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532,
    new_n21533, new_n21534, new_n21535, new_n21536, new_n21537, new_n21538,
    new_n21539, new_n21540, new_n21541, new_n21542, new_n21543, new_n21544,
    new_n21545, new_n21546, new_n21547, new_n21548, new_n21549, new_n21550,
    new_n21551, new_n21552, new_n21553, new_n21554, new_n21555, new_n21556,
    new_n21557, new_n21558, new_n21559, new_n21560, new_n21561, new_n21562,
    new_n21563, new_n21564, new_n21565, new_n21566, new_n21567, new_n21568,
    new_n21569, new_n21570, new_n21571, new_n21572, new_n21573, new_n21574,
    new_n21575, new_n21576, new_n21577, new_n21578, new_n21579, new_n21580,
    new_n21581, new_n21582, new_n21583, new_n21584, new_n21585, new_n21586,
    new_n21587, new_n21588, new_n21589, new_n21590, new_n21591, new_n21592,
    new_n21593, new_n21594, new_n21595, new_n21596, new_n21597, new_n21598,
    new_n21599, new_n21600, new_n21601, new_n21602, new_n21603, new_n21604,
    new_n21605, new_n21606, new_n21607, new_n21608, new_n21609, new_n21610,
    new_n21611, new_n21612, new_n21613, new_n21614, new_n21615, new_n21616,
    new_n21617, new_n21618, new_n21619, new_n21620, new_n21621, new_n21622,
    new_n21623, new_n21624, new_n21625, new_n21626, new_n21627, new_n21628,
    new_n21629, new_n21630, new_n21631, new_n21632, new_n21634, new_n21635,
    new_n21636, new_n21637, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645, new_n21646, new_n21647,
    new_n21648, new_n21649, new_n21650, new_n21651, new_n21652, new_n21653,
    new_n21654, new_n21655, new_n21656, new_n21657, new_n21658, new_n21659,
    new_n21660, new_n21661, new_n21662, new_n21663, new_n21664, new_n21665,
    new_n21666, new_n21667, new_n21668, new_n21669, new_n21670, new_n21671,
    new_n21672, new_n21673, new_n21674, new_n21675, new_n21676, new_n21677,
    new_n21678, new_n21679, new_n21680, new_n21681, new_n21682, new_n21683,
    new_n21684, new_n21685, new_n21686, new_n21687, new_n21688, new_n21689,
    new_n21690, new_n21691, new_n21692, new_n21693, new_n21694, new_n21695,
    new_n21696, new_n21697, new_n21698, new_n21699, new_n21700, new_n21701,
    new_n21702, new_n21703, new_n21704, new_n21705, new_n21706, new_n21707,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21714, new_n21715, new_n21716, new_n21717, new_n21718, new_n21719,
    new_n21720, new_n21721, new_n21722, new_n21723, new_n21724, new_n21725,
    new_n21726, new_n21727, new_n21728, new_n21729, new_n21730, new_n21731,
    new_n21732, new_n21733, new_n21734, new_n21735, new_n21736, new_n21737,
    new_n21738, new_n21739, new_n21740, new_n21741, new_n21742, new_n21743,
    new_n21744, new_n21745, new_n21746, new_n21747, new_n21748, new_n21749,
    new_n21750, new_n21751, new_n21752, new_n21753, new_n21754, new_n21755,
    new_n21756, new_n21757, new_n21758, new_n21759, new_n21760, new_n21761,
    new_n21762, new_n21763, new_n21764, new_n21765, new_n21766, new_n21767,
    new_n21768, new_n21769, new_n21770, new_n21771, new_n21772, new_n21773,
    new_n21774, new_n21775, new_n21777, new_n21778, new_n21779, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784, new_n21785, new_n21786,
    new_n21787, new_n21788, new_n21789, new_n21790, new_n21791, new_n21792,
    new_n21793, new_n21794, new_n21795, new_n21796, new_n21797, new_n21798,
    new_n21799, new_n21800, new_n21801, new_n21802, new_n21803, new_n21804,
    new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810,
    new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816,
    new_n21817, new_n21818, new_n21819, new_n21820, new_n21821, new_n21822,
    new_n21823, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828,
    new_n21829, new_n21830, new_n21831, new_n21832, new_n21833, new_n21834,
    new_n21835, new_n21836, new_n21837, new_n21838, new_n21839, new_n21840,
    new_n21841, new_n21842, new_n21843, new_n21844, new_n21845, new_n21846,
    new_n21847, new_n21848, new_n21849, new_n21850, new_n21851, new_n21852,
    new_n21853, new_n21854, new_n21855, new_n21856, new_n21857, new_n21858,
    new_n21859, new_n21860, new_n21861, new_n21862, new_n21863, new_n21864,
    new_n21865, new_n21866, new_n21867, new_n21868, new_n21869, new_n21870,
    new_n21871, new_n21872, new_n21873, new_n21874, new_n21875, new_n21876,
    new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882,
    new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888,
    new_n21889, new_n21890, new_n21891, new_n21892, new_n21893, new_n21894,
    new_n21895, new_n21896, new_n21897, new_n21898, new_n21899, new_n21900,
    new_n21901, new_n21902, new_n21903, new_n21904, new_n21905, new_n21906,
    new_n21907, new_n21908, new_n21909, new_n21910, new_n21911, new_n21912,
    new_n21913, new_n21914, new_n21915, new_n21917, new_n21918, new_n21919,
    new_n21920, new_n21921, new_n21922, new_n21923, new_n21924, new_n21925,
    new_n21926, new_n21927, new_n21928, new_n21929, new_n21930, new_n21931,
    new_n21932, new_n21933, new_n21934, new_n21935, new_n21936, new_n21937,
    new_n21938, new_n21939, new_n21940, new_n21941, new_n21942, new_n21943,
    new_n21944, new_n21945, new_n21946, new_n21947, new_n21948, new_n21949,
    new_n21950, new_n21951, new_n21952, new_n21953, new_n21954, new_n21955,
    new_n21956, new_n21957, new_n21958, new_n21959, new_n21960, new_n21961,
    new_n21962, new_n21963, new_n21964, new_n21965, new_n21966, new_n21967,
    new_n21968, new_n21969, new_n21970, new_n21971, new_n21972, new_n21973,
    new_n21974, new_n21975, new_n21976, new_n21977, new_n21978, new_n21979,
    new_n21980, new_n21981, new_n21982, new_n21983, new_n21984, new_n21985,
    new_n21986, new_n21987, new_n21988, new_n21989, new_n21990, new_n21991,
    new_n21992, new_n21993, new_n21994, new_n21995, new_n21996, new_n21997,
    new_n21998, new_n21999, new_n22000, new_n22001, new_n22002, new_n22003,
    new_n22004, new_n22005, new_n22006, new_n22007, new_n22008, new_n22009,
    new_n22010, new_n22011, new_n22012, new_n22013, new_n22014, new_n22015,
    new_n22016, new_n22017, new_n22018, new_n22019, new_n22020, new_n22021,
    new_n22022, new_n22023, new_n22024, new_n22025, new_n22026, new_n22027,
    new_n22028, new_n22029, new_n22030, new_n22031, new_n22032, new_n22033,
    new_n22034, new_n22035, new_n22036, new_n22037, new_n22038, new_n22039,
    new_n22040, new_n22041, new_n22042, new_n22043, new_n22044, new_n22045,
    new_n22047, new_n22048, new_n22049, new_n22050, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058,
    new_n22059, new_n22060, new_n22061, new_n22062, new_n22063, new_n22064,
    new_n22065, new_n22066, new_n22067, new_n22068, new_n22069, new_n22070,
    new_n22071, new_n22072, new_n22073, new_n22074, new_n22075, new_n22076,
    new_n22077, new_n22078, new_n22079, new_n22080, new_n22081, new_n22082,
    new_n22083, new_n22084, new_n22085, new_n22086, new_n22087, new_n22088,
    new_n22089, new_n22090, new_n22091, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107, new_n22108, new_n22109, new_n22110, new_n22111, new_n22112,
    new_n22113, new_n22114, new_n22115, new_n22116, new_n22117, new_n22118,
    new_n22119, new_n22120, new_n22121, new_n22122, new_n22123, new_n22124,
    new_n22125, new_n22126, new_n22127, new_n22128, new_n22129, new_n22130,
    new_n22131, new_n22132, new_n22133, new_n22134, new_n22135, new_n22136,
    new_n22137, new_n22138, new_n22139, new_n22140, new_n22141, new_n22142,
    new_n22143, new_n22144, new_n22145, new_n22146, new_n22147, new_n22148,
    new_n22149, new_n22150, new_n22151, new_n22152, new_n22153, new_n22154,
    new_n22155, new_n22156, new_n22157, new_n22158, new_n22159, new_n22160,
    new_n22161, new_n22162, new_n22163, new_n22164, new_n22165, new_n22166,
    new_n22167, new_n22168, new_n22169, new_n22170, new_n22171, new_n22172,
    new_n22173, new_n22174, new_n22175, new_n22176, new_n22177, new_n22179,
    new_n22180, new_n22181, new_n22182, new_n22183, new_n22184, new_n22185,
    new_n22186, new_n22187, new_n22188, new_n22189, new_n22190, new_n22191,
    new_n22192, new_n22193, new_n22194, new_n22195, new_n22196, new_n22197,
    new_n22198, new_n22199, new_n22200, new_n22201, new_n22202, new_n22203,
    new_n22204, new_n22205, new_n22206, new_n22207, new_n22208, new_n22209,
    new_n22210, new_n22211, new_n22212, new_n22213, new_n22214, new_n22215,
    new_n22216, new_n22217, new_n22218, new_n22219, new_n22220, new_n22221,
    new_n22222, new_n22223, new_n22224, new_n22225, new_n22226, new_n22227,
    new_n22228, new_n22229, new_n22230, new_n22231, new_n22232, new_n22233,
    new_n22234, new_n22235, new_n22236, new_n22237, new_n22238, new_n22239,
    new_n22240, new_n22241, new_n22242, new_n22243, new_n22244, new_n22245,
    new_n22246, new_n22247, new_n22248, new_n22249, new_n22250, new_n22251,
    new_n22252, new_n22253, new_n22254, new_n22255, new_n22256, new_n22257,
    new_n22258, new_n22259, new_n22260, new_n22261, new_n22262, new_n22263,
    new_n22264, new_n22265, new_n22266, new_n22267, new_n22268, new_n22269,
    new_n22270, new_n22271, new_n22272, new_n22273, new_n22274, new_n22275,
    new_n22276, new_n22277, new_n22278, new_n22279, new_n22280, new_n22281,
    new_n22282, new_n22283, new_n22284, new_n22285, new_n22286, new_n22287,
    new_n22288, new_n22289, new_n22290, new_n22291, new_n22292, new_n22293,
    new_n22294, new_n22295, new_n22296, new_n22297, new_n22298, new_n22299,
    new_n22300, new_n22301, new_n22302, new_n22303, new_n22304, new_n22306,
    new_n22307, new_n22308, new_n22309, new_n22310, new_n22311, new_n22312,
    new_n22313, new_n22314, new_n22315, new_n22316, new_n22317, new_n22318,
    new_n22319, new_n22320, new_n22321, new_n22322, new_n22323, new_n22324,
    new_n22325, new_n22326, new_n22327, new_n22328, new_n22329, new_n22330,
    new_n22331, new_n22332, new_n22333, new_n22334, new_n22335, new_n22336,
    new_n22337, new_n22338, new_n22339, new_n22340, new_n22341, new_n22342,
    new_n22343, new_n22344, new_n22345, new_n22346, new_n22347, new_n22348,
    new_n22349, new_n22350, new_n22351, new_n22352, new_n22353, new_n22354,
    new_n22355, new_n22356, new_n22357, new_n22358, new_n22359, new_n22360,
    new_n22361, new_n22362, new_n22363, new_n22364, new_n22365, new_n22366,
    new_n22367, new_n22368, new_n22369, new_n22370, new_n22371, new_n22372,
    new_n22373, new_n22374, new_n22375, new_n22376, new_n22377, new_n22378,
    new_n22379, new_n22380, new_n22381, new_n22382, new_n22383, new_n22384,
    new_n22385, new_n22386, new_n22387, new_n22388, new_n22389, new_n22390,
    new_n22391, new_n22392, new_n22393, new_n22394, new_n22395, new_n22396,
    new_n22397, new_n22398, new_n22399, new_n22400, new_n22401, new_n22402,
    new_n22403, new_n22404, new_n22405, new_n22406, new_n22407, new_n22408,
    new_n22409, new_n22410, new_n22411, new_n22412, new_n22413, new_n22414,
    new_n22415, new_n22416, new_n22417, new_n22418, new_n22419, new_n22420,
    new_n22421, new_n22422, new_n22423, new_n22425, new_n22426, new_n22427,
    new_n22428, new_n22429, new_n22430, new_n22431, new_n22432, new_n22433,
    new_n22434, new_n22435, new_n22436, new_n22437, new_n22438, new_n22439,
    new_n22440, new_n22441, new_n22442, new_n22443, new_n22444, new_n22445,
    new_n22446, new_n22447, new_n22448, new_n22449, new_n22450, new_n22451,
    new_n22452, new_n22453, new_n22454, new_n22455, new_n22456, new_n22457,
    new_n22458, new_n22459, new_n22460, new_n22461, new_n22462, new_n22463,
    new_n22464, new_n22465, new_n22466, new_n22467, new_n22468, new_n22469,
    new_n22470, new_n22471, new_n22472, new_n22473, new_n22474, new_n22475,
    new_n22476, new_n22477, new_n22478, new_n22479, new_n22480, new_n22481,
    new_n22482, new_n22483, new_n22484, new_n22485, new_n22486, new_n22487,
    new_n22488, new_n22489, new_n22490, new_n22491, new_n22492, new_n22493,
    new_n22494, new_n22495, new_n22496, new_n22497, new_n22498, new_n22499,
    new_n22500, new_n22501, new_n22502, new_n22503, new_n22504, new_n22505,
    new_n22506, new_n22507, new_n22508, new_n22509, new_n22510, new_n22511,
    new_n22512, new_n22513, new_n22514, new_n22515, new_n22516, new_n22517,
    new_n22518, new_n22519, new_n22520, new_n22521, new_n22522, new_n22523,
    new_n22524, new_n22525, new_n22526, new_n22527, new_n22528, new_n22529,
    new_n22530, new_n22531, new_n22532, new_n22533, new_n22534, new_n22535,
    new_n22536, new_n22537, new_n22538, new_n22539, new_n22540, new_n22541,
    new_n22542, new_n22543, new_n22544, new_n22546, new_n22547, new_n22548,
    new_n22549, new_n22550, new_n22551, new_n22552, new_n22553, new_n22554,
    new_n22555, new_n22556, new_n22557, new_n22558, new_n22559, new_n22560,
    new_n22561, new_n22562, new_n22563, new_n22564, new_n22565, new_n22566,
    new_n22567, new_n22568, new_n22569, new_n22570, new_n22571, new_n22572,
    new_n22573, new_n22574, new_n22575, new_n22576, new_n22577, new_n22578,
    new_n22579, new_n22580, new_n22581, new_n22582, new_n22583, new_n22584,
    new_n22585, new_n22586, new_n22587, new_n22588, new_n22589, new_n22590,
    new_n22591, new_n22592, new_n22593, new_n22594, new_n22595, new_n22596,
    new_n22597, new_n22598, new_n22599, new_n22600, new_n22601, new_n22602,
    new_n22603, new_n22604, new_n22605, new_n22606, new_n22607, new_n22608,
    new_n22609, new_n22610, new_n22611, new_n22612, new_n22613, new_n22614,
    new_n22615, new_n22616, new_n22617, new_n22618, new_n22619, new_n22620,
    new_n22621, new_n22622, new_n22623, new_n22624, new_n22625, new_n22626,
    new_n22627, new_n22628, new_n22629, new_n22630, new_n22631, new_n22632,
    new_n22633, new_n22634, new_n22635, new_n22636, new_n22637, new_n22638,
    new_n22639, new_n22640, new_n22641, new_n22642, new_n22643, new_n22644,
    new_n22645, new_n22646, new_n22647, new_n22648, new_n22649, new_n22651,
    new_n22652, new_n22653, new_n22654, new_n22655, new_n22656, new_n22657,
    new_n22658, new_n22659, new_n22660, new_n22661, new_n22662, new_n22663,
    new_n22664, new_n22665, new_n22666, new_n22667, new_n22668, new_n22669,
    new_n22670, new_n22671, new_n22672, new_n22673, new_n22674, new_n22675,
    new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681,
    new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687,
    new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22693,
    new_n22694, new_n22695, new_n22696, new_n22697, new_n22698, new_n22699,
    new_n22700, new_n22701, new_n22702, new_n22703, new_n22704, new_n22705,
    new_n22706, new_n22707, new_n22708, new_n22709, new_n22710, new_n22711,
    new_n22712, new_n22713, new_n22714, new_n22715, new_n22716, new_n22717,
    new_n22718, new_n22719, new_n22720, new_n22721, new_n22722, new_n22723,
    new_n22724, new_n22725, new_n22726, new_n22727, new_n22728, new_n22729,
    new_n22730, new_n22731, new_n22732, new_n22733, new_n22734, new_n22735,
    new_n22736, new_n22737, new_n22738, new_n22739, new_n22740, new_n22741,
    new_n22742, new_n22743, new_n22744, new_n22745, new_n22746, new_n22747,
    new_n22748, new_n22750, new_n22751, new_n22752, new_n22753, new_n22754,
    new_n22755, new_n22756, new_n22757, new_n22758, new_n22759, new_n22760,
    new_n22761, new_n22762, new_n22763, new_n22764, new_n22765, new_n22766,
    new_n22767, new_n22768, new_n22769, new_n22770, new_n22771, new_n22772,
    new_n22773, new_n22774, new_n22775, new_n22776, new_n22777, new_n22778,
    new_n22779, new_n22780, new_n22781, new_n22782, new_n22783, new_n22784,
    new_n22785, new_n22786, new_n22787, new_n22788, new_n22789, new_n22790,
    new_n22791, new_n22792, new_n22793, new_n22794, new_n22795, new_n22796,
    new_n22797, new_n22798, new_n22799, new_n22800, new_n22801, new_n22802,
    new_n22803, new_n22804, new_n22805, new_n22806, new_n22807, new_n22808,
    new_n22809, new_n22810, new_n22811, new_n22812, new_n22813, new_n22814,
    new_n22815, new_n22816, new_n22817, new_n22818, new_n22819, new_n22820,
    new_n22821, new_n22822, new_n22823, new_n22824, new_n22825, new_n22826,
    new_n22827, new_n22828, new_n22829, new_n22830, new_n22831, new_n22832,
    new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22838,
    new_n22839, new_n22840, new_n22841, new_n22842, new_n22843, new_n22844,
    new_n22845, new_n22846, new_n22847, new_n22848, new_n22849, new_n22850,
    new_n22851, new_n22853, new_n22854, new_n22855, new_n22856, new_n22857,
    new_n22858, new_n22859, new_n22860, new_n22861, new_n22862, new_n22863,
    new_n22864, new_n22865, new_n22866, new_n22867, new_n22868, new_n22869,
    new_n22870, new_n22871, new_n22872, new_n22873, new_n22874, new_n22875,
    new_n22876, new_n22877, new_n22878, new_n22879, new_n22880, new_n22881,
    new_n22882, new_n22883, new_n22884, new_n22885, new_n22886, new_n22887,
    new_n22888, new_n22889, new_n22890, new_n22891, new_n22892, new_n22893,
    new_n22894, new_n22895, new_n22896, new_n22897, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903, new_n22904, new_n22905,
    new_n22906, new_n22907, new_n22908, new_n22909, new_n22910, new_n22911,
    new_n22912, new_n22913, new_n22914, new_n22915, new_n22916, new_n22917,
    new_n22918, new_n22919, new_n22920, new_n22921, new_n22922, new_n22923,
    new_n22924, new_n22925, new_n22926, new_n22927, new_n22928, new_n22929,
    new_n22930, new_n22931, new_n22932, new_n22933, new_n22934, new_n22935,
    new_n22936, new_n22937, new_n22938, new_n22939, new_n22940, new_n22941,
    new_n22942, new_n22943, new_n22944, new_n22946, new_n22947, new_n22948,
    new_n22949, new_n22950, new_n22951, new_n22952, new_n22953, new_n22954,
    new_n22955, new_n22956, new_n22957, new_n22958, new_n22959, new_n22960,
    new_n22961, new_n22962, new_n22963, new_n22964, new_n22965, new_n22966,
    new_n22967, new_n22968, new_n22969, new_n22970, new_n22971, new_n22972,
    new_n22973, new_n22974, new_n22975, new_n22976, new_n22977, new_n22978,
    new_n22979, new_n22980, new_n22981, new_n22982, new_n22983, new_n22984,
    new_n22985, new_n22986, new_n22987, new_n22988, new_n22989, new_n22990,
    new_n22991, new_n22992, new_n22993, new_n22994, new_n22995, new_n22996,
    new_n22997, new_n22998, new_n22999, new_n23000, new_n23001, new_n23002,
    new_n23003, new_n23004, new_n23005, new_n23006, new_n23007, new_n23008,
    new_n23009, new_n23010, new_n23011, new_n23012, new_n23013, new_n23014,
    new_n23015, new_n23016, new_n23017, new_n23018, new_n23019, new_n23020,
    new_n23021, new_n23022, new_n23023, new_n23024, new_n23025, new_n23026,
    new_n23027, new_n23028, new_n23029, new_n23030, new_n23031, new_n23032,
    new_n23033, new_n23034, new_n23035, new_n23036, new_n23038, new_n23039,
    new_n23040, new_n23041, new_n23042, new_n23043, new_n23044, new_n23045,
    new_n23046, new_n23047, new_n23048, new_n23049, new_n23050, new_n23051,
    new_n23052, new_n23053, new_n23054, new_n23055, new_n23056, new_n23057,
    new_n23058, new_n23059, new_n23060, new_n23061, new_n23062, new_n23063,
    new_n23064, new_n23065, new_n23066, new_n23067, new_n23068, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23074, new_n23075,
    new_n23076, new_n23077, new_n23078, new_n23079, new_n23080, new_n23081,
    new_n23082, new_n23083, new_n23084, new_n23085, new_n23086, new_n23087,
    new_n23088, new_n23089, new_n23090, new_n23091, new_n23092, new_n23093,
    new_n23094, new_n23095, new_n23096, new_n23097, new_n23098, new_n23099,
    new_n23100, new_n23101, new_n23102, new_n23103, new_n23104, new_n23105,
    new_n23106, new_n23107, new_n23108, new_n23109, new_n23110, new_n23111,
    new_n23112, new_n23113, new_n23114, new_n23115, new_n23116, new_n23117,
    new_n23118, new_n23120, new_n23121, new_n23122, new_n23123, new_n23124,
    new_n23125, new_n23126, new_n23127, new_n23128, new_n23129, new_n23130,
    new_n23131, new_n23132, new_n23133, new_n23134, new_n23135, new_n23136,
    new_n23137, new_n23138, new_n23139, new_n23140, new_n23141, new_n23142,
    new_n23143, new_n23144, new_n23145, new_n23146, new_n23147, new_n23148,
    new_n23149, new_n23150, new_n23151, new_n23152, new_n23153, new_n23154,
    new_n23155, new_n23156, new_n23157, new_n23158, new_n23159, new_n23160,
    new_n23161, new_n23162, new_n23163, new_n23164, new_n23165, new_n23166,
    new_n23167, new_n23168, new_n23169, new_n23170, new_n23171, new_n23172,
    new_n23173, new_n23174, new_n23175, new_n23176, new_n23177, new_n23178,
    new_n23179, new_n23180, new_n23181, new_n23182, new_n23183, new_n23184,
    new_n23185, new_n23186, new_n23187, new_n23188, new_n23189, new_n23190,
    new_n23191, new_n23192, new_n23193, new_n23194, new_n23195, new_n23196,
    new_n23197, new_n23198, new_n23199, new_n23200, new_n23202, new_n23203,
    new_n23204, new_n23205, new_n23206, new_n23207, new_n23208, new_n23209,
    new_n23210, new_n23211, new_n23212, new_n23213, new_n23214, new_n23215,
    new_n23216, new_n23217, new_n23218, new_n23219, new_n23220, new_n23221,
    new_n23222, new_n23223, new_n23224, new_n23225, new_n23226, new_n23227,
    new_n23228, new_n23229, new_n23230, new_n23231, new_n23232, new_n23233,
    new_n23234, new_n23235, new_n23236, new_n23237, new_n23238, new_n23239,
    new_n23240, new_n23241, new_n23242, new_n23243, new_n23244, new_n23245,
    new_n23246, new_n23247, new_n23248, new_n23249, new_n23250, new_n23251,
    new_n23252, new_n23253, new_n23254, new_n23255, new_n23256, new_n23257,
    new_n23258, new_n23259, new_n23260, new_n23261, new_n23262, new_n23263,
    new_n23264, new_n23265, new_n23266, new_n23267, new_n23268, new_n23269,
    new_n23270, new_n23271, new_n23272, new_n23273, new_n23275, new_n23276,
    new_n23277, new_n23278, new_n23279, new_n23280, new_n23281, new_n23282,
    new_n23283, new_n23284, new_n23285, new_n23286, new_n23287, new_n23288,
    new_n23289, new_n23290, new_n23291, new_n23292, new_n23293, new_n23294,
    new_n23295, new_n23296, new_n23297, new_n23298, new_n23299, new_n23300,
    new_n23301, new_n23302, new_n23303, new_n23304, new_n23305, new_n23306,
    new_n23307, new_n23308, new_n23309, new_n23310, new_n23311, new_n23312,
    new_n23313, new_n23314, new_n23315, new_n23316, new_n23317, new_n23318,
    new_n23319, new_n23320, new_n23321, new_n23322, new_n23323, new_n23324,
    new_n23325, new_n23326, new_n23327, new_n23328, new_n23329, new_n23330,
    new_n23331, new_n23332, new_n23334, new_n23335, new_n23336, new_n23337,
    new_n23338, new_n23339, new_n23340, new_n23341, new_n23342, new_n23343,
    new_n23344, new_n23345, new_n23346, new_n23347, new_n23348, new_n23349,
    new_n23350, new_n23351, new_n23352, new_n23353, new_n23354, new_n23355,
    new_n23356, new_n23357, new_n23358, new_n23359, new_n23360, new_n23361,
    new_n23362, new_n23363, new_n23364, new_n23365, new_n23366, new_n23367,
    new_n23368, new_n23369, new_n23370, new_n23371, new_n23372, new_n23373,
    new_n23374, new_n23375, new_n23376, new_n23377, new_n23378, new_n23379,
    new_n23380, new_n23381, new_n23382, new_n23383, new_n23384, new_n23385,
    new_n23386, new_n23387, new_n23388, new_n23389, new_n23390, new_n23391,
    new_n23392, new_n23393, new_n23394, new_n23395, new_n23396, new_n23397,
    new_n23399, new_n23400, new_n23401, new_n23402, new_n23403, new_n23404,
    new_n23405, new_n23406, new_n23407, new_n23408, new_n23409, new_n23410,
    new_n23411, new_n23412, new_n23413, new_n23414, new_n23415, new_n23416,
    new_n23417, new_n23418, new_n23419, new_n23420, new_n23421, new_n23422,
    new_n23423, new_n23424, new_n23425, new_n23426, new_n23427, new_n23428,
    new_n23429, new_n23430, new_n23431, new_n23432, new_n23433, new_n23434,
    new_n23435, new_n23436, new_n23437, new_n23438, new_n23439, new_n23440,
    new_n23441, new_n23442, new_n23443, new_n23444, new_n23445, new_n23446,
    new_n23447, new_n23448, new_n23449, new_n23450, new_n23451, new_n23452,
    new_n23453, new_n23454, new_n23455, new_n23456, new_n23458, new_n23459,
    new_n23460, new_n23461, new_n23462, new_n23463, new_n23464, new_n23465,
    new_n23466, new_n23467, new_n23468, new_n23469, new_n23470, new_n23471,
    new_n23472, new_n23473, new_n23474, new_n23475, new_n23476, new_n23477,
    new_n23478, new_n23479, new_n23480, new_n23481, new_n23482, new_n23483,
    new_n23484, new_n23485, new_n23486, new_n23487, new_n23488, new_n23489,
    new_n23490, new_n23491, new_n23492, new_n23493, new_n23494, new_n23495,
    new_n23496, new_n23497, new_n23498, new_n23499, new_n23500, new_n23501,
    new_n23502, new_n23503, new_n23504, new_n23505, new_n23506, new_n23507,
    new_n23508, new_n23509, new_n23510, new_n23512, new_n23513, new_n23514,
    new_n23515, new_n23516, new_n23517, new_n23518, new_n23519, new_n23520,
    new_n23521, new_n23522, new_n23523, new_n23524, new_n23525, new_n23526,
    new_n23527, new_n23528, new_n23529, new_n23530, new_n23531, new_n23532,
    new_n23533, new_n23534, new_n23535, new_n23536, new_n23537, new_n23538,
    new_n23539, new_n23540, new_n23541, new_n23542, new_n23543, new_n23544,
    new_n23545, new_n23546, new_n23547, new_n23548, new_n23549, new_n23550,
    new_n23551, new_n23552, new_n23553, new_n23554, new_n23555, new_n23556,
    new_n23558, new_n23559, new_n23560, new_n23561, new_n23562, new_n23563,
    new_n23564, new_n23565, new_n23566, new_n23567, new_n23568, new_n23569,
    new_n23570, new_n23571, new_n23572, new_n23573, new_n23574, new_n23575,
    new_n23576, new_n23577, new_n23578, new_n23579, new_n23580, new_n23581,
    new_n23582, new_n23583, new_n23584, new_n23585, new_n23586, new_n23587,
    new_n23588, new_n23589, new_n23590, new_n23591, new_n23592, new_n23593,
    new_n23594, new_n23595, new_n23596, new_n23597, new_n23598, new_n23599,
    new_n23600, new_n23602, new_n23603, new_n23604, new_n23605, new_n23606,
    new_n23607, new_n23608, new_n23609, new_n23610, new_n23611, new_n23612,
    new_n23613, new_n23614, new_n23615, new_n23616, new_n23617, new_n23618,
    new_n23619, new_n23620, new_n23621, new_n23622, new_n23623, new_n23624,
    new_n23625, new_n23626, new_n23627, new_n23628, new_n23629, new_n23630,
    new_n23631, new_n23632, new_n23633, new_n23634, new_n23635, new_n23636,
    new_n23637, new_n23638, new_n23639, new_n23640, new_n23642, new_n23643,
    new_n23644, new_n23645, new_n23646, new_n23647, new_n23648, new_n23649,
    new_n23650, new_n23651, new_n23652, new_n23653, new_n23654, new_n23655,
    new_n23656, new_n23657, new_n23658, new_n23659, new_n23660, new_n23661,
    new_n23662, new_n23663, new_n23664, new_n23665, new_n23666, new_n23667,
    new_n23668, new_n23669, new_n23670, new_n23671, new_n23672, new_n23673,
    new_n23674, new_n23675, new_n23676, new_n23678, new_n23679, new_n23680,
    new_n23681, new_n23682, new_n23683, new_n23684, new_n23685, new_n23686,
    new_n23687, new_n23688, new_n23689, new_n23690, new_n23691, new_n23692,
    new_n23693, new_n23694, new_n23695, new_n23696, new_n23697, new_n23698,
    new_n23699, new_n23700, new_n23701, new_n23702, new_n23703, new_n23705,
    new_n23706, new_n23707, new_n23708, new_n23709, new_n23710, new_n23711,
    new_n23712, new_n23713, new_n23714, new_n23715, new_n23716, new_n23717,
    new_n23718, new_n23719, new_n23720, new_n23721, new_n23722, new_n23723,
    new_n23724, new_n23725, new_n23726, new_n23727, new_n23728, new_n23729,
    new_n23730, new_n23731, new_n23733, new_n23734, new_n23735, new_n23736,
    new_n23737, new_n23738, new_n23739, new_n23740, new_n23741, new_n23742,
    new_n23743, new_n23744, new_n23746, new_n23747, new_n23748, new_n23749,
    new_n23750, new_n23751, new_n23752, new_n23753;
  INVx1_ASAP7_75t_L         g00000(.A(\a[2] ), .Y(new_n257));
  AOI21xp33_ASAP7_75t_L     g00001(.A1(\a[0] ), .A2(\b[0] ), .B(new_n257), .Y(new_n258));
  AOI21xp33_ASAP7_75t_L     g00002(.A1(\a[0] ), .A2(\b[0] ), .B(\a[2] ), .Y(new_n259));
  NOR2xp33_ASAP7_75t_L      g00003(.A(new_n259), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00004(.A(\b[0] ), .B(\a[0] ), .Y(new_n261));
  INVx1_ASAP7_75t_L         g00005(.A(\b[1] ), .Y(new_n262));
  INVx1_ASAP7_75t_L         g00006(.A(\a[1] ), .Y(new_n263));
  NOR2xp33_ASAP7_75t_L      g00007(.A(\a[0] ), .B(new_n263), .Y(new_n264));
  NAND2xp33_ASAP7_75t_L     g00008(.A(\b[0] ), .B(new_n264), .Y(new_n265));
  NOR2xp33_ASAP7_75t_L      g00009(.A(\a[1] ), .B(new_n257), .Y(new_n266));
  NOR2xp33_ASAP7_75t_L      g00010(.A(\a[2] ), .B(new_n263), .Y(new_n267));
  NOR2xp33_ASAP7_75t_L      g00011(.A(new_n266), .B(new_n267), .Y(new_n268));
  NAND2xp33_ASAP7_75t_L     g00012(.A(\a[0] ), .B(new_n268), .Y(new_n269));
  OAI21xp33_ASAP7_75t_L     g00013(.A1(new_n262), .A2(new_n269), .B(new_n265), .Y(new_n270));
  INVx1_ASAP7_75t_L         g00014(.A(new_n270), .Y(new_n271));
  INVx1_ASAP7_75t_L         g00015(.A(\a[0] ), .Y(new_n272));
  NOR2xp33_ASAP7_75t_L      g00016(.A(new_n272), .B(new_n268), .Y(new_n273));
  XNOR2x2_ASAP7_75t_L       g00017(.A(\b[1] ), .B(\b[0] ), .Y(new_n274));
  INVx1_ASAP7_75t_L         g00018(.A(new_n274), .Y(new_n275));
  NAND2xp33_ASAP7_75t_L     g00019(.A(new_n275), .B(new_n273), .Y(new_n276));
  AND4x1_ASAP7_75t_L        g00020(.A(new_n276), .B(new_n271), .C(new_n261), .D(\a[2] ), .Y(new_n277));
  A2O1A1Ixp33_ASAP7_75t_L   g00021(.A1(new_n273), .A2(new_n275), .B(new_n270), .C(\a[2] ), .Y(new_n278));
  INVx1_ASAP7_75t_L         g00022(.A(new_n273), .Y(new_n279));
  O2A1O1Ixp33_ASAP7_75t_L   g00023(.A1(new_n279), .A2(new_n274), .B(new_n271), .C(\a[2] ), .Y(new_n280));
  O2A1O1Ixp33_ASAP7_75t_L   g00024(.A1(new_n261), .A2(new_n278), .B(\a[2] ), .C(new_n280), .Y(new_n281));
  NOR2xp33_ASAP7_75t_L      g00025(.A(new_n277), .B(new_n281), .Y(\f[1] ));
  INVx1_ASAP7_75t_L         g00026(.A(new_n269), .Y(new_n283));
  INVx1_ASAP7_75t_L         g00027(.A(\b[0] ), .Y(new_n284));
  INVx1_ASAP7_75t_L         g00028(.A(new_n264), .Y(new_n285));
  NOR3xp33_ASAP7_75t_L      g00029(.A(new_n257), .B(\a[1] ), .C(\a[0] ), .Y(new_n286));
  INVx1_ASAP7_75t_L         g00030(.A(new_n286), .Y(new_n287));
  OAI22xp33_ASAP7_75t_L     g00031(.A1(new_n287), .A2(new_n284), .B1(new_n262), .B2(new_n285), .Y(new_n288));
  INVx1_ASAP7_75t_L         g00032(.A(\b[2] ), .Y(new_n289));
  NAND3xp33_ASAP7_75t_L     g00033(.A(new_n289), .B(\b[1] ), .C(\b[0] ), .Y(new_n290));
  NAND2xp33_ASAP7_75t_L     g00034(.A(\b[1] ), .B(new_n289), .Y(new_n291));
  NAND2xp33_ASAP7_75t_L     g00035(.A(\b[2] ), .B(new_n262), .Y(new_n292));
  OAI211xp5_ASAP7_75t_L     g00036(.A1(new_n262), .A2(new_n284), .B(new_n291), .C(new_n292), .Y(new_n293));
  AND2x2_ASAP7_75t_L        g00037(.A(new_n290), .B(new_n293), .Y(new_n294));
  AOI221xp5_ASAP7_75t_L     g00038(.A1(new_n294), .A2(new_n273), .B1(\b[2] ), .B2(new_n283), .C(new_n288), .Y(new_n295));
  XNOR2x2_ASAP7_75t_L       g00039(.A(\a[2] ), .B(new_n295), .Y(new_n296));
  NAND2xp33_ASAP7_75t_L     g00040(.A(new_n277), .B(new_n296), .Y(new_n297));
  INVx1_ASAP7_75t_L         g00041(.A(new_n297), .Y(new_n298));
  A2O1A1O1Ixp25_ASAP7_75t_L g00042(.A1(new_n278), .A2(\a[2] ), .B(new_n280), .C(new_n258), .D(new_n296), .Y(new_n299));
  NOR2xp33_ASAP7_75t_L      g00043(.A(new_n299), .B(new_n298), .Y(\f[2] ));
  INVx1_ASAP7_75t_L         g00044(.A(\b[3] ), .Y(new_n301));
  AOI22xp33_ASAP7_75t_L     g00045(.A1(new_n264), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n286), .Y(new_n302));
  OAI21xp33_ASAP7_75t_L     g00046(.A1(new_n301), .A2(new_n269), .B(new_n302), .Y(new_n303));
  NOR2xp33_ASAP7_75t_L      g00047(.A(\b[2] ), .B(\b[3] ), .Y(new_n304));
  INVx1_ASAP7_75t_L         g00048(.A(new_n304), .Y(new_n305));
  NAND2xp33_ASAP7_75t_L     g00049(.A(\b[3] ), .B(\b[2] ), .Y(new_n306));
  NAND2xp33_ASAP7_75t_L     g00050(.A(new_n306), .B(new_n305), .Y(new_n307));
  O2A1O1Ixp33_ASAP7_75t_L   g00051(.A1(new_n262), .A2(new_n289), .B(new_n290), .C(new_n307), .Y(new_n308));
  INVx1_ASAP7_75t_L         g00052(.A(new_n306), .Y(new_n309));
  NOR2xp33_ASAP7_75t_L      g00053(.A(new_n304), .B(new_n309), .Y(new_n310));
  O2A1O1Ixp33_ASAP7_75t_L   g00054(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n310), .Y(new_n311));
  NOR2xp33_ASAP7_75t_L      g00055(.A(new_n311), .B(new_n308), .Y(new_n312));
  A2O1A1Ixp33_ASAP7_75t_L   g00056(.A1(new_n312), .A2(new_n273), .B(new_n303), .C(\a[2] ), .Y(new_n313));
  INVx1_ASAP7_75t_L         g00057(.A(new_n303), .Y(new_n314));
  OAI21xp33_ASAP7_75t_L     g00058(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n315));
  INVx1_ASAP7_75t_L         g00059(.A(new_n315), .Y(new_n316));
  NAND2xp33_ASAP7_75t_L     g00060(.A(new_n316), .B(new_n310), .Y(new_n317));
  A2O1A1Ixp33_ASAP7_75t_L   g00061(.A1(new_n289), .A2(new_n284), .B(new_n262), .C(new_n307), .Y(new_n318));
  NAND2xp33_ASAP7_75t_L     g00062(.A(new_n317), .B(new_n318), .Y(new_n319));
  O2A1O1Ixp33_ASAP7_75t_L   g00063(.A1(new_n319), .A2(new_n279), .B(new_n314), .C(\a[2] ), .Y(new_n320));
  INVx1_ASAP7_75t_L         g00064(.A(\a[3] ), .Y(new_n321));
  NAND2xp33_ASAP7_75t_L     g00065(.A(\a[2] ), .B(new_n321), .Y(new_n322));
  NAND2xp33_ASAP7_75t_L     g00066(.A(\a[3] ), .B(new_n257), .Y(new_n323));
  NAND2xp33_ASAP7_75t_L     g00067(.A(new_n323), .B(new_n322), .Y(new_n324));
  NAND2xp33_ASAP7_75t_L     g00068(.A(\b[0] ), .B(new_n324), .Y(new_n325));
  INVx1_ASAP7_75t_L         g00069(.A(new_n325), .Y(new_n326));
  A2O1A1Ixp33_ASAP7_75t_L   g00070(.A1(new_n313), .A2(\a[2] ), .B(new_n320), .C(new_n326), .Y(new_n327));
  AOI21xp33_ASAP7_75t_L     g00071(.A1(new_n313), .A2(\a[2] ), .B(new_n320), .Y(new_n328));
  A2O1A1Ixp33_ASAP7_75t_L   g00072(.A1(new_n322), .A2(new_n323), .B(new_n284), .C(new_n328), .Y(new_n329));
  NAND2xp33_ASAP7_75t_L     g00073(.A(new_n327), .B(new_n329), .Y(new_n330));
  XNOR2x2_ASAP7_75t_L       g00074(.A(new_n298), .B(new_n330), .Y(\f[3] ));
  INVx1_ASAP7_75t_L         g00075(.A(\b[4] ), .Y(new_n332));
  NAND2xp33_ASAP7_75t_L     g00076(.A(\b[2] ), .B(new_n286), .Y(new_n333));
  OAI221xp5_ASAP7_75t_L     g00077(.A1(new_n285), .A2(new_n301), .B1(new_n332), .B2(new_n269), .C(new_n333), .Y(new_n334));
  NOR2xp33_ASAP7_75t_L      g00078(.A(\b[3] ), .B(\b[4] ), .Y(new_n335));
  NOR2xp33_ASAP7_75t_L      g00079(.A(new_n301), .B(new_n332), .Y(new_n336));
  NOR2xp33_ASAP7_75t_L      g00080(.A(new_n335), .B(new_n336), .Y(new_n337));
  A2O1A1Ixp33_ASAP7_75t_L   g00081(.A1(new_n305), .A2(new_n316), .B(new_n309), .C(new_n337), .Y(new_n338));
  INVx1_ASAP7_75t_L         g00082(.A(new_n338), .Y(new_n339));
  OAI21xp33_ASAP7_75t_L     g00083(.A1(new_n304), .A2(new_n315), .B(new_n306), .Y(new_n340));
  NOR2xp33_ASAP7_75t_L      g00084(.A(new_n340), .B(new_n337), .Y(new_n341));
  NOR2xp33_ASAP7_75t_L      g00085(.A(new_n341), .B(new_n339), .Y(new_n342));
  A2O1A1Ixp33_ASAP7_75t_L   g00086(.A1(new_n342), .A2(new_n273), .B(new_n334), .C(\a[2] ), .Y(new_n343));
  A2O1A1Ixp33_ASAP7_75t_L   g00087(.A1(new_n342), .A2(new_n273), .B(new_n334), .C(new_n257), .Y(new_n344));
  INVx1_ASAP7_75t_L         g00088(.A(new_n344), .Y(new_n345));
  INVx1_ASAP7_75t_L         g00089(.A(\a[5] ), .Y(new_n346));
  AND2x2_ASAP7_75t_L        g00090(.A(new_n322), .B(new_n323), .Y(new_n347));
  XNOR2x2_ASAP7_75t_L       g00091(.A(\a[4] ), .B(\a[3] ), .Y(new_n348));
  NOR2xp33_ASAP7_75t_L      g00092(.A(new_n348), .B(new_n324), .Y(new_n349));
  INVx1_ASAP7_75t_L         g00093(.A(new_n349), .Y(new_n350));
  INVx1_ASAP7_75t_L         g00094(.A(\a[4] ), .Y(new_n351));
  NAND2xp33_ASAP7_75t_L     g00095(.A(\a[5] ), .B(new_n351), .Y(new_n352));
  NAND2xp33_ASAP7_75t_L     g00096(.A(\a[4] ), .B(new_n346), .Y(new_n353));
  NAND2xp33_ASAP7_75t_L     g00097(.A(new_n353), .B(new_n352), .Y(new_n354));
  OAI32xp33_ASAP7_75t_L     g00098(.A1(new_n262), .A2(new_n354), .A3(new_n347), .B1(new_n350), .B2(new_n284), .Y(new_n355));
  NAND2xp33_ASAP7_75t_L     g00099(.A(new_n354), .B(new_n324), .Y(new_n356));
  NOR2xp33_ASAP7_75t_L      g00100(.A(new_n274), .B(new_n356), .Y(new_n357));
  NOR4xp25_ASAP7_75t_L      g00101(.A(new_n355), .B(new_n346), .C(new_n357), .D(new_n326), .Y(new_n358));
  INVx1_ASAP7_75t_L         g00102(.A(new_n356), .Y(new_n359));
  A2O1A1Ixp33_ASAP7_75t_L   g00103(.A1(new_n359), .A2(new_n275), .B(new_n355), .C(\a[5] ), .Y(new_n360));
  NOR2xp33_ASAP7_75t_L      g00104(.A(new_n354), .B(new_n347), .Y(new_n361));
  AOI221xp5_ASAP7_75t_L     g00105(.A1(\b[1] ), .A2(new_n361), .B1(new_n349), .B2(\b[0] ), .C(new_n357), .Y(new_n362));
  NOR2xp33_ASAP7_75t_L      g00106(.A(\a[5] ), .B(new_n362), .Y(new_n363));
  O2A1O1Ixp33_ASAP7_75t_L   g00107(.A1(new_n325), .A2(new_n360), .B(\a[5] ), .C(new_n363), .Y(new_n364));
  NOR2xp33_ASAP7_75t_L      g00108(.A(new_n358), .B(new_n364), .Y(new_n365));
  A2O1A1Ixp33_ASAP7_75t_L   g00109(.A1(\a[2] ), .A2(new_n343), .B(new_n345), .C(new_n365), .Y(new_n366));
  AO21x2_ASAP7_75t_L        g00110(.A1(\a[2] ), .A2(new_n343), .B(new_n345), .Y(new_n367));
  NOR3xp33_ASAP7_75t_L      g00111(.A(new_n367), .B(new_n364), .C(new_n358), .Y(new_n368));
  A2O1A1O1Ixp25_ASAP7_75t_L g00112(.A1(new_n343), .A2(\a[2] ), .B(new_n345), .C(new_n366), .D(new_n368), .Y(new_n369));
  O2A1O1Ixp33_ASAP7_75t_L   g00113(.A1(new_n297), .A2(new_n330), .B(new_n327), .C(new_n369), .Y(new_n370));
  MAJIxp5_ASAP7_75t_L       g00114(.A(new_n297), .B(new_n328), .C(new_n325), .Y(new_n371));
  AOI211xp5_ASAP7_75t_L     g00115(.A1(new_n366), .A2(new_n367), .B(new_n371), .C(new_n368), .Y(new_n372));
  NOR2xp33_ASAP7_75t_L      g00116(.A(new_n372), .B(new_n370), .Y(\f[4] ));
  NAND2xp33_ASAP7_75t_L     g00117(.A(\b[2] ), .B(new_n361), .Y(new_n374));
  NAND3xp33_ASAP7_75t_L     g00118(.A(new_n347), .B(new_n348), .C(new_n354), .Y(new_n375));
  OAI221xp5_ASAP7_75t_L     g00119(.A1(new_n350), .A2(new_n262), .B1(new_n375), .B2(new_n284), .C(new_n374), .Y(new_n376));
  AOI21xp33_ASAP7_75t_L     g00120(.A1(new_n359), .A2(new_n294), .B(new_n376), .Y(new_n377));
  NAND4xp25_ASAP7_75t_L     g00121(.A(new_n377), .B(\a[5] ), .C(new_n325), .D(new_n362), .Y(new_n378));
  INVx1_ASAP7_75t_L         g00122(.A(new_n358), .Y(new_n379));
  NAND2xp33_ASAP7_75t_L     g00123(.A(\a[5] ), .B(new_n377), .Y(new_n380));
  A2O1A1Ixp33_ASAP7_75t_L   g00124(.A1(new_n294), .A2(new_n359), .B(new_n376), .C(new_n346), .Y(new_n381));
  NAND3xp33_ASAP7_75t_L     g00125(.A(new_n380), .B(new_n379), .C(new_n381), .Y(new_n382));
  NAND2xp33_ASAP7_75t_L     g00126(.A(new_n378), .B(new_n382), .Y(new_n383));
  INVx1_ASAP7_75t_L         g00127(.A(\b[5] ), .Y(new_n384));
  NOR2xp33_ASAP7_75t_L      g00128(.A(new_n301), .B(new_n287), .Y(new_n385));
  INVx1_ASAP7_75t_L         g00129(.A(new_n385), .Y(new_n386));
  OAI221xp5_ASAP7_75t_L     g00130(.A1(new_n285), .A2(new_n332), .B1(new_n384), .B2(new_n269), .C(new_n386), .Y(new_n387));
  NOR2xp33_ASAP7_75t_L      g00131(.A(\b[4] ), .B(\b[5] ), .Y(new_n388));
  NOR2xp33_ASAP7_75t_L      g00132(.A(new_n332), .B(new_n384), .Y(new_n389));
  NOR2xp33_ASAP7_75t_L      g00133(.A(new_n388), .B(new_n389), .Y(new_n390));
  A2O1A1Ixp33_ASAP7_75t_L   g00134(.A1(new_n337), .A2(new_n340), .B(new_n336), .C(new_n390), .Y(new_n391));
  A2O1A1O1Ixp25_ASAP7_75t_L g00135(.A1(new_n305), .A2(new_n316), .B(new_n309), .C(new_n337), .D(new_n336), .Y(new_n392));
  OAI21xp33_ASAP7_75t_L     g00136(.A1(new_n388), .A2(new_n389), .B(new_n392), .Y(new_n393));
  AND2x2_ASAP7_75t_L        g00137(.A(new_n391), .B(new_n393), .Y(new_n394));
  A2O1A1Ixp33_ASAP7_75t_L   g00138(.A1(new_n394), .A2(new_n273), .B(new_n387), .C(\a[2] ), .Y(new_n395));
  INVx1_ASAP7_75t_L         g00139(.A(new_n395), .Y(new_n396));
  A2O1A1Ixp33_ASAP7_75t_L   g00140(.A1(new_n394), .A2(new_n273), .B(new_n387), .C(new_n257), .Y(new_n397));
  O2A1O1Ixp33_ASAP7_75t_L   g00141(.A1(new_n396), .A2(new_n257), .B(new_n397), .C(new_n383), .Y(new_n398));
  INVx1_ASAP7_75t_L         g00142(.A(new_n397), .Y(new_n399));
  A2O1A1Ixp33_ASAP7_75t_L   g00143(.A1(\a[2] ), .A2(new_n395), .B(new_n399), .C(new_n383), .Y(new_n400));
  MAJIxp5_ASAP7_75t_L       g00144(.A(new_n371), .B(new_n367), .C(new_n365), .Y(new_n401));
  O2A1O1Ixp33_ASAP7_75t_L   g00145(.A1(new_n383), .A2(new_n398), .B(new_n400), .C(new_n401), .Y(new_n402));
  OA211x2_ASAP7_75t_L       g00146(.A1(new_n383), .A2(new_n398), .B(new_n400), .C(new_n401), .Y(new_n403));
  NOR2xp33_ASAP7_75t_L      g00147(.A(new_n402), .B(new_n403), .Y(\f[5] ));
  NOR2xp33_ASAP7_75t_L      g00148(.A(new_n257), .B(new_n396), .Y(new_n405));
  A2O1A1O1Ixp25_ASAP7_75t_L g00149(.A1(new_n273), .A2(new_n394), .B(new_n387), .C(new_n395), .D(new_n405), .Y(new_n406));
  MAJIxp5_ASAP7_75t_L       g00150(.A(new_n401), .B(new_n383), .C(new_n406), .Y(new_n407));
  AND4x1_ASAP7_75t_L        g00151(.A(new_n377), .B(new_n362), .C(new_n325), .D(\a[5] ), .Y(new_n408));
  INVx1_ASAP7_75t_L         g00152(.A(\a[6] ), .Y(new_n409));
  NAND2xp33_ASAP7_75t_L     g00153(.A(\a[5] ), .B(new_n409), .Y(new_n410));
  NAND2xp33_ASAP7_75t_L     g00154(.A(\a[6] ), .B(new_n346), .Y(new_n411));
  A2O1A1Ixp33_ASAP7_75t_L   g00155(.A1(new_n410), .A2(new_n411), .B(new_n284), .C(new_n408), .Y(new_n412));
  AND2x2_ASAP7_75t_L        g00156(.A(new_n410), .B(new_n411), .Y(new_n413));
  NOR2xp33_ASAP7_75t_L      g00157(.A(new_n284), .B(new_n413), .Y(new_n414));
  A2O1A1Ixp33_ASAP7_75t_L   g00158(.A1(new_n380), .A2(new_n381), .B(new_n379), .C(new_n414), .Y(new_n415));
  NAND2xp33_ASAP7_75t_L     g00159(.A(\b[3] ), .B(new_n361), .Y(new_n416));
  OAI221xp5_ASAP7_75t_L     g00160(.A1(new_n350), .A2(new_n289), .B1(new_n262), .B2(new_n375), .C(new_n416), .Y(new_n417));
  NOR2xp33_ASAP7_75t_L      g00161(.A(new_n356), .B(new_n319), .Y(new_n418));
  A2O1A1Ixp33_ASAP7_75t_L   g00162(.A1(new_n312), .A2(new_n359), .B(new_n417), .C(\a[5] ), .Y(new_n419));
  NOR3xp33_ASAP7_75t_L      g00163(.A(new_n417), .B(new_n418), .C(new_n346), .Y(new_n420));
  O2A1O1Ixp33_ASAP7_75t_L   g00164(.A1(new_n417), .A2(new_n418), .B(new_n419), .C(new_n420), .Y(new_n421));
  INVx1_ASAP7_75t_L         g00165(.A(new_n421), .Y(new_n422));
  AO21x2_ASAP7_75t_L        g00166(.A1(new_n415), .A2(new_n412), .B(new_n422), .Y(new_n423));
  NAND3xp33_ASAP7_75t_L     g00167(.A(new_n412), .B(new_n415), .C(new_n422), .Y(new_n424));
  NOR2xp33_ASAP7_75t_L      g00168(.A(new_n332), .B(new_n287), .Y(new_n425));
  AOI221xp5_ASAP7_75t_L     g00169(.A1(\b[5] ), .A2(new_n264), .B1(\b[6] ), .B2(new_n283), .C(new_n425), .Y(new_n426));
  INVx1_ASAP7_75t_L         g00170(.A(\b[6] ), .Y(new_n427));
  NAND2xp33_ASAP7_75t_L     g00171(.A(new_n427), .B(new_n384), .Y(new_n428));
  NAND2xp33_ASAP7_75t_L     g00172(.A(\b[6] ), .B(\b[5] ), .Y(new_n429));
  NAND2xp33_ASAP7_75t_L     g00173(.A(new_n429), .B(new_n428), .Y(new_n430));
  O2A1O1Ixp33_ASAP7_75t_L   g00174(.A1(new_n332), .A2(new_n384), .B(new_n391), .C(new_n430), .Y(new_n431));
  INVx1_ASAP7_75t_L         g00175(.A(new_n389), .Y(new_n432));
  AND3x1_ASAP7_75t_L        g00176(.A(new_n391), .B(new_n430), .C(new_n432), .Y(new_n433));
  OR2x4_ASAP7_75t_L         g00177(.A(new_n431), .B(new_n433), .Y(new_n434));
  O2A1O1Ixp33_ASAP7_75t_L   g00178(.A1(new_n279), .A2(new_n434), .B(new_n426), .C(new_n257), .Y(new_n435));
  OAI21xp33_ASAP7_75t_L     g00179(.A1(new_n279), .A2(new_n434), .B(new_n426), .Y(new_n436));
  NAND2xp33_ASAP7_75t_L     g00180(.A(new_n257), .B(new_n436), .Y(new_n437));
  OA21x2_ASAP7_75t_L        g00181(.A1(new_n257), .A2(new_n435), .B(new_n437), .Y(new_n438));
  AOI21xp33_ASAP7_75t_L     g00182(.A1(new_n423), .A2(new_n424), .B(new_n438), .Y(new_n439));
  INVx1_ASAP7_75t_L         g00183(.A(new_n439), .Y(new_n440));
  NAND3xp33_ASAP7_75t_L     g00184(.A(new_n423), .B(new_n424), .C(new_n438), .Y(new_n441));
  AND3x1_ASAP7_75t_L        g00185(.A(new_n440), .B(new_n441), .C(new_n407), .Y(new_n442));
  AOI21xp33_ASAP7_75t_L     g00186(.A1(new_n440), .A2(new_n441), .B(new_n407), .Y(new_n443));
  NOR2xp33_ASAP7_75t_L      g00187(.A(new_n443), .B(new_n442), .Y(\f[6] ));
  O2A1O1Ixp33_ASAP7_75t_L   g00188(.A1(new_n398), .A2(new_n402), .B(new_n441), .C(new_n439), .Y(new_n445));
  NOR2xp33_ASAP7_75t_L      g00189(.A(new_n384), .B(new_n287), .Y(new_n446));
  AOI221xp5_ASAP7_75t_L     g00190(.A1(\b[6] ), .A2(new_n264), .B1(\b[7] ), .B2(new_n283), .C(new_n446), .Y(new_n447));
  INVx1_ASAP7_75t_L         g00191(.A(\b[7] ), .Y(new_n448));
  NAND2xp33_ASAP7_75t_L     g00192(.A(new_n448), .B(new_n427), .Y(new_n449));
  NAND2xp33_ASAP7_75t_L     g00193(.A(\b[7] ), .B(\b[6] ), .Y(new_n450));
  NAND2xp33_ASAP7_75t_L     g00194(.A(new_n450), .B(new_n449), .Y(new_n451));
  A2O1A1O1Ixp25_ASAP7_75t_L g00195(.A1(new_n432), .A2(new_n391), .B(new_n430), .C(new_n429), .D(new_n451), .Y(new_n452));
  INVx1_ASAP7_75t_L         g00196(.A(new_n452), .Y(new_n453));
  A2O1A1O1Ixp25_ASAP7_75t_L g00197(.A1(new_n340), .A2(new_n337), .B(new_n336), .C(new_n390), .D(new_n389), .Y(new_n454));
  OAI211xp5_ASAP7_75t_L     g00198(.A1(new_n430), .A2(new_n454), .B(new_n429), .C(new_n451), .Y(new_n455));
  NAND2xp33_ASAP7_75t_L     g00199(.A(new_n455), .B(new_n453), .Y(new_n456));
  OAI21xp33_ASAP7_75t_L     g00200(.A1(new_n279), .A2(new_n456), .B(new_n447), .Y(new_n457));
  NOR2xp33_ASAP7_75t_L      g00201(.A(new_n257), .B(new_n457), .Y(new_n458));
  O2A1O1Ixp33_ASAP7_75t_L   g00202(.A1(new_n279), .A2(new_n456), .B(new_n447), .C(\a[2] ), .Y(new_n459));
  NOR2xp33_ASAP7_75t_L      g00203(.A(new_n459), .B(new_n458), .Y(new_n460));
  NAND2xp33_ASAP7_75t_L     g00204(.A(\b[4] ), .B(new_n361), .Y(new_n461));
  OAI221xp5_ASAP7_75t_L     g00205(.A1(new_n350), .A2(new_n301), .B1(new_n289), .B2(new_n375), .C(new_n461), .Y(new_n462));
  A2O1A1Ixp33_ASAP7_75t_L   g00206(.A1(new_n342), .A2(new_n359), .B(new_n462), .C(\a[5] ), .Y(new_n463));
  AOI211xp5_ASAP7_75t_L     g00207(.A1(new_n359), .A2(new_n342), .B(new_n346), .C(new_n462), .Y(new_n464));
  A2O1A1O1Ixp25_ASAP7_75t_L g00208(.A1(new_n342), .A2(new_n359), .B(new_n462), .C(new_n463), .D(new_n464), .Y(new_n465));
  INVx1_ASAP7_75t_L         g00209(.A(\a[8] ), .Y(new_n466));
  A2O1A1Ixp33_ASAP7_75t_L   g00210(.A1(new_n410), .A2(new_n411), .B(new_n284), .C(\a[8] ), .Y(new_n467));
  NAND2xp33_ASAP7_75t_L     g00211(.A(new_n411), .B(new_n410), .Y(new_n468));
  XNOR2x2_ASAP7_75t_L       g00212(.A(\a[7] ), .B(\a[6] ), .Y(new_n469));
  NOR2xp33_ASAP7_75t_L      g00213(.A(new_n469), .B(new_n468), .Y(new_n470));
  INVx1_ASAP7_75t_L         g00214(.A(\a[7] ), .Y(new_n471));
  NAND2xp33_ASAP7_75t_L     g00215(.A(\a[8] ), .B(new_n471), .Y(new_n472));
  NAND2xp33_ASAP7_75t_L     g00216(.A(\a[7] ), .B(new_n466), .Y(new_n473));
  NAND2xp33_ASAP7_75t_L     g00217(.A(new_n473), .B(new_n472), .Y(new_n474));
  NOR2xp33_ASAP7_75t_L      g00218(.A(new_n474), .B(new_n413), .Y(new_n475));
  AOI22xp33_ASAP7_75t_L     g00219(.A1(new_n470), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n475), .Y(new_n476));
  NAND2xp33_ASAP7_75t_L     g00220(.A(new_n474), .B(new_n468), .Y(new_n477));
  O2A1O1Ixp33_ASAP7_75t_L   g00221(.A1(new_n477), .A2(new_n274), .B(new_n476), .C(new_n466), .Y(new_n478));
  O2A1O1Ixp33_ASAP7_75t_L   g00222(.A1(new_n477), .A2(new_n274), .B(new_n476), .C(\a[8] ), .Y(new_n479));
  INVx1_ASAP7_75t_L         g00223(.A(new_n479), .Y(new_n480));
  O2A1O1Ixp33_ASAP7_75t_L   g00224(.A1(new_n478), .A2(new_n466), .B(new_n480), .C(new_n467), .Y(new_n481));
  INVx1_ASAP7_75t_L         g00225(.A(new_n414), .Y(new_n482));
  INVx1_ASAP7_75t_L         g00226(.A(new_n477), .Y(new_n483));
  NAND2xp33_ASAP7_75t_L     g00227(.A(new_n275), .B(new_n483), .Y(new_n484));
  AND3x1_ASAP7_75t_L        g00228(.A(new_n484), .B(new_n476), .C(\a[8] ), .Y(new_n485));
  AOI211xp5_ASAP7_75t_L     g00229(.A1(new_n482), .A2(\a[8] ), .B(new_n479), .C(new_n485), .Y(new_n486));
  NOR3xp33_ASAP7_75t_L      g00230(.A(new_n465), .B(new_n486), .C(new_n481), .Y(new_n487));
  AND2x2_ASAP7_75t_L        g00231(.A(new_n476), .B(new_n484), .Y(new_n488));
  NAND3xp33_ASAP7_75t_L     g00232(.A(new_n488), .B(new_n482), .C(\a[8] ), .Y(new_n489));
  A2O1A1Ixp33_ASAP7_75t_L   g00233(.A1(new_n414), .A2(new_n478), .B(new_n466), .C(new_n480), .Y(new_n490));
  INVx1_ASAP7_75t_L         g00234(.A(new_n464), .Y(new_n491));
  A2O1A1Ixp33_ASAP7_75t_L   g00235(.A1(new_n342), .A2(new_n359), .B(new_n462), .C(new_n346), .Y(new_n492));
  NAND4xp25_ASAP7_75t_L     g00236(.A(new_n490), .B(new_n491), .C(new_n492), .D(new_n489), .Y(new_n493));
  MAJIxp5_ASAP7_75t_L       g00237(.A(new_n422), .B(new_n414), .C(new_n408), .Y(new_n494));
  O2A1O1Ixp33_ASAP7_75t_L   g00238(.A1(new_n465), .A2(new_n487), .B(new_n493), .C(new_n494), .Y(new_n495));
  INVx1_ASAP7_75t_L         g00239(.A(new_n492), .Y(new_n496));
  OAI22xp33_ASAP7_75t_L     g00240(.A1(new_n481), .A2(new_n486), .B1(new_n496), .B2(new_n464), .Y(new_n497));
  NAND2xp33_ASAP7_75t_L     g00241(.A(new_n493), .B(new_n497), .Y(new_n498));
  MAJIxp5_ASAP7_75t_L       g00242(.A(new_n421), .B(new_n482), .C(new_n378), .Y(new_n499));
  NOR2xp33_ASAP7_75t_L      g00243(.A(new_n499), .B(new_n498), .Y(new_n500));
  NOR3xp33_ASAP7_75t_L      g00244(.A(new_n495), .B(new_n500), .C(new_n460), .Y(new_n501));
  INVx1_ASAP7_75t_L         g00245(.A(new_n501), .Y(new_n502));
  OAI21xp33_ASAP7_75t_L     g00246(.A1(new_n500), .A2(new_n495), .B(new_n460), .Y(new_n503));
  NAND2xp33_ASAP7_75t_L     g00247(.A(new_n503), .B(new_n502), .Y(new_n504));
  XOR2x2_ASAP7_75t_L        g00248(.A(new_n445), .B(new_n504), .Y(\f[7] ));
  NAND3xp33_ASAP7_75t_L     g00249(.A(new_n413), .B(new_n469), .C(new_n474), .Y(new_n506));
  NOR2xp33_ASAP7_75t_L      g00250(.A(new_n284), .B(new_n506), .Y(new_n507));
  AOI221xp5_ASAP7_75t_L     g00251(.A1(\b[2] ), .A2(new_n475), .B1(new_n470), .B2(\b[1] ), .C(new_n507), .Y(new_n508));
  NAND2xp33_ASAP7_75t_L     g00252(.A(new_n290), .B(new_n293), .Y(new_n509));
  NOR2xp33_ASAP7_75t_L      g00253(.A(new_n477), .B(new_n509), .Y(new_n510));
  INVx1_ASAP7_75t_L         g00254(.A(new_n510), .Y(new_n511));
  NAND3xp33_ASAP7_75t_L     g00255(.A(new_n508), .B(\a[8] ), .C(new_n511), .Y(new_n512));
  OR2x4_ASAP7_75t_L         g00256(.A(new_n469), .B(new_n468), .Y(new_n513));
  NAND2xp33_ASAP7_75t_L     g00257(.A(\b[2] ), .B(new_n475), .Y(new_n514));
  OAI221xp5_ASAP7_75t_L     g00258(.A1(new_n513), .A2(new_n262), .B1(new_n506), .B2(new_n284), .C(new_n514), .Y(new_n515));
  A2O1A1Ixp33_ASAP7_75t_L   g00259(.A1(new_n294), .A2(new_n483), .B(new_n515), .C(new_n466), .Y(new_n516));
  NAND3xp33_ASAP7_75t_L     g00260(.A(new_n489), .B(new_n512), .C(new_n516), .Y(new_n517));
  NAND5xp2_ASAP7_75t_L      g00261(.A(\a[8] ), .B(new_n488), .C(new_n511), .D(new_n508), .E(new_n482), .Y(new_n518));
  NAND2xp33_ASAP7_75t_L     g00262(.A(\b[5] ), .B(new_n361), .Y(new_n519));
  OAI221xp5_ASAP7_75t_L     g00263(.A1(new_n350), .A2(new_n332), .B1(new_n301), .B2(new_n375), .C(new_n519), .Y(new_n520));
  A2O1A1Ixp33_ASAP7_75t_L   g00264(.A1(new_n394), .A2(new_n359), .B(new_n520), .C(\a[5] ), .Y(new_n521));
  NAND2xp33_ASAP7_75t_L     g00265(.A(\a[5] ), .B(new_n521), .Y(new_n522));
  A2O1A1Ixp33_ASAP7_75t_L   g00266(.A1(new_n394), .A2(new_n359), .B(new_n520), .C(new_n346), .Y(new_n523));
  NAND4xp25_ASAP7_75t_L     g00267(.A(new_n517), .B(new_n522), .C(new_n523), .D(new_n518), .Y(new_n524));
  AO22x1_ASAP7_75t_L        g00268(.A1(new_n523), .A2(new_n522), .B1(new_n518), .B2(new_n517), .Y(new_n525));
  AOI21xp33_ASAP7_75t_L     g00269(.A1(new_n498), .A2(new_n499), .B(new_n487), .Y(new_n526));
  NAND3xp33_ASAP7_75t_L     g00270(.A(new_n526), .B(new_n525), .C(new_n524), .Y(new_n527));
  NAND2xp33_ASAP7_75t_L     g00271(.A(new_n524), .B(new_n525), .Y(new_n528));
  A2O1A1Ixp33_ASAP7_75t_L   g00272(.A1(new_n498), .A2(new_n499), .B(new_n487), .C(new_n528), .Y(new_n529));
  NAND2xp33_ASAP7_75t_L     g00273(.A(new_n529), .B(new_n527), .Y(new_n530));
  NOR2xp33_ASAP7_75t_L      g00274(.A(new_n427), .B(new_n287), .Y(new_n531));
  AOI221xp5_ASAP7_75t_L     g00275(.A1(\b[7] ), .A2(new_n264), .B1(\b[8] ), .B2(new_n283), .C(new_n531), .Y(new_n532));
  NOR2xp33_ASAP7_75t_L      g00276(.A(\b[7] ), .B(\b[8] ), .Y(new_n533));
  INVx1_ASAP7_75t_L         g00277(.A(\b[8] ), .Y(new_n534));
  NOR2xp33_ASAP7_75t_L      g00278(.A(new_n448), .B(new_n534), .Y(new_n535));
  NOR2xp33_ASAP7_75t_L      g00279(.A(new_n533), .B(new_n535), .Y(new_n536));
  A2O1A1Ixp33_ASAP7_75t_L   g00280(.A1(\b[7] ), .A2(\b[6] ), .B(new_n452), .C(new_n536), .Y(new_n537));
  INVx1_ASAP7_75t_L         g00281(.A(new_n536), .Y(new_n538));
  NAND3xp33_ASAP7_75t_L     g00282(.A(new_n453), .B(new_n450), .C(new_n538), .Y(new_n539));
  NAND2xp33_ASAP7_75t_L     g00283(.A(new_n537), .B(new_n539), .Y(new_n540));
  O2A1O1Ixp33_ASAP7_75t_L   g00284(.A1(new_n279), .A2(new_n540), .B(new_n532), .C(new_n257), .Y(new_n541));
  NOR2xp33_ASAP7_75t_L      g00285(.A(new_n257), .B(new_n541), .Y(new_n542));
  O2A1O1Ixp33_ASAP7_75t_L   g00286(.A1(new_n279), .A2(new_n540), .B(new_n532), .C(\a[2] ), .Y(new_n543));
  NOR2xp33_ASAP7_75t_L      g00287(.A(new_n543), .B(new_n542), .Y(new_n544));
  XNOR2x2_ASAP7_75t_L       g00288(.A(new_n544), .B(new_n530), .Y(new_n545));
  O2A1O1Ixp33_ASAP7_75t_L   g00289(.A1(new_n445), .A2(new_n504), .B(new_n502), .C(new_n545), .Y(new_n546));
  A2O1A1O1Ixp25_ASAP7_75t_L g00290(.A1(new_n441), .A2(new_n407), .B(new_n439), .C(new_n503), .D(new_n501), .Y(new_n547));
  AND2x2_ASAP7_75t_L        g00291(.A(new_n547), .B(new_n545), .Y(new_n548));
  NOR2xp33_ASAP7_75t_L      g00292(.A(new_n546), .B(new_n548), .Y(\f[8] ));
  INVx1_ASAP7_75t_L         g00293(.A(\a[9] ), .Y(new_n550));
  NAND2xp33_ASAP7_75t_L     g00294(.A(\a[8] ), .B(new_n550), .Y(new_n551));
  NAND2xp33_ASAP7_75t_L     g00295(.A(\a[9] ), .B(new_n466), .Y(new_n552));
  AND2x2_ASAP7_75t_L        g00296(.A(new_n551), .B(new_n552), .Y(new_n553));
  NOR2xp33_ASAP7_75t_L      g00297(.A(new_n284), .B(new_n553), .Y(new_n554));
  A2O1A1Ixp33_ASAP7_75t_L   g00298(.A1(new_n512), .A2(new_n516), .B(new_n489), .C(new_n554), .Y(new_n555));
  NAND2xp33_ASAP7_75t_L     g00299(.A(new_n476), .B(new_n484), .Y(new_n556));
  NOR5xp2_ASAP7_75t_L       g00300(.A(new_n556), .B(new_n515), .C(new_n510), .D(new_n414), .E(new_n466), .Y(new_n557));
  A2O1A1Ixp33_ASAP7_75t_L   g00301(.A1(new_n551), .A2(new_n552), .B(new_n284), .C(new_n557), .Y(new_n558));
  NAND2xp33_ASAP7_75t_L     g00302(.A(\b[3] ), .B(new_n475), .Y(new_n559));
  INVx1_ASAP7_75t_L         g00303(.A(new_n506), .Y(new_n560));
  NAND2xp33_ASAP7_75t_L     g00304(.A(\b[1] ), .B(new_n560), .Y(new_n561));
  NAND2xp33_ASAP7_75t_L     g00305(.A(\b[2] ), .B(new_n470), .Y(new_n562));
  NAND2xp33_ASAP7_75t_L     g00306(.A(new_n483), .B(new_n312), .Y(new_n563));
  NAND5xp2_ASAP7_75t_L      g00307(.A(new_n563), .B(new_n562), .C(new_n561), .D(new_n559), .E(\a[8] ), .Y(new_n564));
  OAI211xp5_ASAP7_75t_L     g00308(.A1(new_n506), .A2(new_n262), .B(new_n559), .C(new_n562), .Y(new_n565));
  A2O1A1Ixp33_ASAP7_75t_L   g00309(.A1(new_n312), .A2(new_n483), .B(new_n565), .C(new_n466), .Y(new_n566));
  AND2x2_ASAP7_75t_L        g00310(.A(new_n564), .B(new_n566), .Y(new_n567));
  AO21x2_ASAP7_75t_L        g00311(.A1(new_n555), .A2(new_n558), .B(new_n567), .Y(new_n568));
  NAND3xp33_ASAP7_75t_L     g00312(.A(new_n558), .B(new_n555), .C(new_n567), .Y(new_n569));
  NOR2xp33_ASAP7_75t_L      g00313(.A(new_n332), .B(new_n375), .Y(new_n570));
  AOI221xp5_ASAP7_75t_L     g00314(.A1(\b[6] ), .A2(new_n361), .B1(new_n349), .B2(\b[5] ), .C(new_n570), .Y(new_n571));
  O2A1O1Ixp33_ASAP7_75t_L   g00315(.A1(new_n356), .A2(new_n434), .B(new_n571), .C(new_n346), .Y(new_n572));
  OAI21xp33_ASAP7_75t_L     g00316(.A1(new_n356), .A2(new_n434), .B(new_n571), .Y(new_n573));
  NAND2xp33_ASAP7_75t_L     g00317(.A(new_n346), .B(new_n573), .Y(new_n574));
  OA21x2_ASAP7_75t_L        g00318(.A1(new_n346), .A2(new_n572), .B(new_n574), .Y(new_n575));
  NAND3xp33_ASAP7_75t_L     g00319(.A(new_n575), .B(new_n568), .C(new_n569), .Y(new_n576));
  AO21x2_ASAP7_75t_L        g00320(.A1(new_n568), .A2(new_n569), .B(new_n575), .Y(new_n577));
  NAND2xp33_ASAP7_75t_L     g00321(.A(new_n576), .B(new_n577), .Y(new_n578));
  NAND2xp33_ASAP7_75t_L     g00322(.A(new_n518), .B(new_n517), .Y(new_n579));
  INVx1_ASAP7_75t_L         g00323(.A(new_n522), .Y(new_n580));
  A2O1A1O1Ixp25_ASAP7_75t_L g00324(.A1(new_n394), .A2(new_n359), .B(new_n520), .C(new_n521), .D(new_n580), .Y(new_n581));
  MAJIxp5_ASAP7_75t_L       g00325(.A(new_n526), .B(new_n579), .C(new_n581), .Y(new_n582));
  NOR2xp33_ASAP7_75t_L      g00326(.A(new_n578), .B(new_n582), .Y(new_n583));
  NAND2xp33_ASAP7_75t_L     g00327(.A(new_n569), .B(new_n568), .Y(new_n584));
  O2A1O1Ixp33_ASAP7_75t_L   g00328(.A1(new_n572), .A2(new_n346), .B(new_n574), .C(new_n584), .Y(new_n585));
  INVx1_ASAP7_75t_L         g00329(.A(new_n521), .Y(new_n586));
  O2A1O1Ixp33_ASAP7_75t_L   g00330(.A1(new_n586), .A2(new_n346), .B(new_n523), .C(new_n579), .Y(new_n587));
  A2O1A1O1Ixp25_ASAP7_75t_L g00331(.A1(new_n498), .A2(new_n499), .B(new_n487), .C(new_n528), .D(new_n587), .Y(new_n588));
  O2A1O1Ixp33_ASAP7_75t_L   g00332(.A1(new_n575), .A2(new_n585), .B(new_n576), .C(new_n588), .Y(new_n589));
  INVx1_ASAP7_75t_L         g00333(.A(\b[9] ), .Y(new_n590));
  NAND2xp33_ASAP7_75t_L     g00334(.A(\b[7] ), .B(new_n286), .Y(new_n591));
  OAI221xp5_ASAP7_75t_L     g00335(.A1(new_n285), .A2(new_n534), .B1(new_n590), .B2(new_n269), .C(new_n591), .Y(new_n592));
  INVx1_ASAP7_75t_L         g00336(.A(new_n535), .Y(new_n593));
  NOR2xp33_ASAP7_75t_L      g00337(.A(\b[8] ), .B(\b[9] ), .Y(new_n594));
  NOR2xp33_ASAP7_75t_L      g00338(.A(new_n534), .B(new_n590), .Y(new_n595));
  NOR2xp33_ASAP7_75t_L      g00339(.A(new_n594), .B(new_n595), .Y(new_n596));
  INVx1_ASAP7_75t_L         g00340(.A(new_n596), .Y(new_n597));
  A2O1A1O1Ixp25_ASAP7_75t_L g00341(.A1(new_n450), .A2(new_n453), .B(new_n533), .C(new_n593), .D(new_n597), .Y(new_n598));
  A2O1A1O1Ixp25_ASAP7_75t_L g00342(.A1(\b[7] ), .A2(\b[6] ), .B(new_n452), .C(new_n536), .D(new_n535), .Y(new_n599));
  NAND2xp33_ASAP7_75t_L     g00343(.A(new_n597), .B(new_n599), .Y(new_n600));
  INVx1_ASAP7_75t_L         g00344(.A(new_n600), .Y(new_n601));
  NOR2xp33_ASAP7_75t_L      g00345(.A(new_n598), .B(new_n601), .Y(new_n602));
  A2O1A1Ixp33_ASAP7_75t_L   g00346(.A1(new_n602), .A2(new_n273), .B(new_n592), .C(\a[2] ), .Y(new_n603));
  AOI211xp5_ASAP7_75t_L     g00347(.A1(new_n602), .A2(new_n273), .B(new_n592), .C(new_n257), .Y(new_n604));
  A2O1A1O1Ixp25_ASAP7_75t_L g00348(.A1(new_n273), .A2(new_n602), .B(new_n592), .C(new_n603), .D(new_n604), .Y(new_n605));
  INVx1_ASAP7_75t_L         g00349(.A(new_n605), .Y(new_n606));
  NOR3xp33_ASAP7_75t_L      g00350(.A(new_n583), .B(new_n589), .C(new_n606), .Y(new_n607));
  NAND3xp33_ASAP7_75t_L     g00351(.A(new_n588), .B(new_n577), .C(new_n576), .Y(new_n608));
  NOR2xp33_ASAP7_75t_L      g00352(.A(new_n486), .B(new_n481), .Y(new_n609));
  A2O1A1Ixp33_ASAP7_75t_L   g00353(.A1(\a[5] ), .A2(new_n463), .B(new_n496), .C(new_n609), .Y(new_n610));
  A2O1A1Ixp33_ASAP7_75t_L   g00354(.A1(new_n493), .A2(new_n497), .B(new_n494), .C(new_n610), .Y(new_n611));
  A2O1A1Ixp33_ASAP7_75t_L   g00355(.A1(new_n528), .A2(new_n611), .B(new_n587), .C(new_n578), .Y(new_n612));
  AOI21xp33_ASAP7_75t_L     g00356(.A1(new_n612), .A2(new_n608), .B(new_n605), .Y(new_n613));
  MAJIxp5_ASAP7_75t_L       g00357(.A(new_n547), .B(new_n544), .C(new_n530), .Y(new_n614));
  OAI21xp33_ASAP7_75t_L     g00358(.A1(new_n607), .A2(new_n613), .B(new_n614), .Y(new_n615));
  INVx1_ASAP7_75t_L         g00359(.A(new_n615), .Y(new_n616));
  NOR3xp33_ASAP7_75t_L      g00360(.A(new_n614), .B(new_n613), .C(new_n607), .Y(new_n617));
  NOR2xp33_ASAP7_75t_L      g00361(.A(new_n617), .B(new_n616), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g00362(.A(new_n589), .B(new_n583), .Y(new_n619));
  NAND2xp33_ASAP7_75t_L     g00363(.A(new_n606), .B(new_n619), .Y(new_n620));
  INVx1_ASAP7_75t_L         g00364(.A(new_n620), .Y(new_n621));
  O2A1O1Ixp33_ASAP7_75t_L   g00365(.A1(new_n606), .A2(new_n607), .B(new_n614), .C(new_n621), .Y(new_n622));
  INVx1_ASAP7_75t_L         g00366(.A(new_n554), .Y(new_n623));
  MAJIxp5_ASAP7_75t_L       g00367(.A(new_n567), .B(new_n623), .C(new_n518), .Y(new_n624));
  NAND2xp33_ASAP7_75t_L     g00368(.A(\b[4] ), .B(new_n475), .Y(new_n625));
  OAI221xp5_ASAP7_75t_L     g00369(.A1(new_n513), .A2(new_n301), .B1(new_n289), .B2(new_n506), .C(new_n625), .Y(new_n626));
  A2O1A1Ixp33_ASAP7_75t_L   g00370(.A1(new_n342), .A2(new_n483), .B(new_n626), .C(\a[8] ), .Y(new_n627));
  AOI211xp5_ASAP7_75t_L     g00371(.A1(new_n342), .A2(new_n483), .B(new_n466), .C(new_n626), .Y(new_n628));
  A2O1A1O1Ixp25_ASAP7_75t_L g00372(.A1(new_n483), .A2(new_n342), .B(new_n626), .C(new_n627), .D(new_n628), .Y(new_n629));
  NAND2xp33_ASAP7_75t_L     g00373(.A(new_n552), .B(new_n551), .Y(new_n630));
  INVx1_ASAP7_75t_L         g00374(.A(\a[10] ), .Y(new_n631));
  NOR2xp33_ASAP7_75t_L      g00375(.A(\a[9] ), .B(new_n631), .Y(new_n632));
  NOR2xp33_ASAP7_75t_L      g00376(.A(\a[10] ), .B(new_n550), .Y(new_n633));
  NOR2xp33_ASAP7_75t_L      g00377(.A(new_n632), .B(new_n633), .Y(new_n634));
  NOR2xp33_ASAP7_75t_L      g00378(.A(new_n630), .B(new_n634), .Y(new_n635));
  NAND2xp33_ASAP7_75t_L     g00379(.A(\a[11] ), .B(new_n631), .Y(new_n636));
  INVx1_ASAP7_75t_L         g00380(.A(\a[11] ), .Y(new_n637));
  NAND2xp33_ASAP7_75t_L     g00381(.A(\a[10] ), .B(new_n637), .Y(new_n638));
  NAND2xp33_ASAP7_75t_L     g00382(.A(new_n638), .B(new_n636), .Y(new_n639));
  NOR2xp33_ASAP7_75t_L      g00383(.A(new_n639), .B(new_n553), .Y(new_n640));
  NAND2xp33_ASAP7_75t_L     g00384(.A(new_n639), .B(new_n630), .Y(new_n641));
  NOR2xp33_ASAP7_75t_L      g00385(.A(new_n274), .B(new_n641), .Y(new_n642));
  AOI221xp5_ASAP7_75t_L     g00386(.A1(\b[1] ), .A2(new_n640), .B1(new_n635), .B2(\b[0] ), .C(new_n642), .Y(new_n643));
  NAND3xp33_ASAP7_75t_L     g00387(.A(new_n643), .B(new_n623), .C(\a[11] ), .Y(new_n644));
  INVx1_ASAP7_75t_L         g00388(.A(new_n644), .Y(new_n645));
  AOI22xp33_ASAP7_75t_L     g00389(.A1(new_n635), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n640), .Y(new_n646));
  OAI21xp33_ASAP7_75t_L     g00390(.A1(new_n641), .A2(new_n274), .B(new_n646), .Y(new_n647));
  NOR2xp33_ASAP7_75t_L      g00391(.A(new_n637), .B(new_n647), .Y(new_n648));
  O2A1O1Ixp33_ASAP7_75t_L   g00392(.A1(new_n641), .A2(new_n274), .B(new_n646), .C(\a[11] ), .Y(new_n649));
  AOI211xp5_ASAP7_75t_L     g00393(.A1(new_n623), .A2(\a[11] ), .B(new_n649), .C(new_n648), .Y(new_n650));
  OAI21xp33_ASAP7_75t_L     g00394(.A1(new_n645), .A2(new_n650), .B(new_n629), .Y(new_n651));
  A2O1A1Ixp33_ASAP7_75t_L   g00395(.A1(new_n342), .A2(new_n483), .B(new_n626), .C(new_n466), .Y(new_n652));
  INVx1_ASAP7_75t_L         g00396(.A(new_n652), .Y(new_n653));
  O2A1O1Ixp33_ASAP7_75t_L   g00397(.A1(new_n641), .A2(new_n274), .B(new_n646), .C(new_n637), .Y(new_n654));
  INVx1_ASAP7_75t_L         g00398(.A(new_n649), .Y(new_n655));
  A2O1A1Ixp33_ASAP7_75t_L   g00399(.A1(new_n554), .A2(new_n654), .B(new_n637), .C(new_n655), .Y(new_n656));
  OAI211xp5_ASAP7_75t_L     g00400(.A1(new_n628), .A2(new_n653), .B(new_n656), .C(new_n644), .Y(new_n657));
  NAND3xp33_ASAP7_75t_L     g00401(.A(new_n624), .B(new_n651), .C(new_n657), .Y(new_n658));
  NAND2xp33_ASAP7_75t_L     g00402(.A(new_n564), .B(new_n566), .Y(new_n659));
  MAJIxp5_ASAP7_75t_L       g00403(.A(new_n659), .B(new_n554), .C(new_n557), .Y(new_n660));
  AOI211xp5_ASAP7_75t_L     g00404(.A1(new_n656), .A2(new_n644), .B(new_n628), .C(new_n653), .Y(new_n661));
  INVx1_ASAP7_75t_L         g00405(.A(new_n628), .Y(new_n662));
  AOI211xp5_ASAP7_75t_L     g00406(.A1(new_n662), .A2(new_n652), .B(new_n645), .C(new_n650), .Y(new_n663));
  OAI21xp33_ASAP7_75t_L     g00407(.A1(new_n663), .A2(new_n661), .B(new_n660), .Y(new_n664));
  NOR2xp33_ASAP7_75t_L      g00408(.A(new_n384), .B(new_n375), .Y(new_n665));
  AOI221xp5_ASAP7_75t_L     g00409(.A1(\b[7] ), .A2(new_n361), .B1(new_n349), .B2(\b[6] ), .C(new_n665), .Y(new_n666));
  O2A1O1Ixp33_ASAP7_75t_L   g00410(.A1(new_n356), .A2(new_n456), .B(new_n666), .C(new_n346), .Y(new_n667));
  OAI21xp33_ASAP7_75t_L     g00411(.A1(new_n356), .A2(new_n456), .B(new_n666), .Y(new_n668));
  NAND2xp33_ASAP7_75t_L     g00412(.A(new_n346), .B(new_n668), .Y(new_n669));
  OA21x2_ASAP7_75t_L        g00413(.A1(new_n346), .A2(new_n667), .B(new_n669), .Y(new_n670));
  NAND3xp33_ASAP7_75t_L     g00414(.A(new_n658), .B(new_n664), .C(new_n670), .Y(new_n671));
  NOR3xp33_ASAP7_75t_L      g00415(.A(new_n661), .B(new_n663), .C(new_n660), .Y(new_n672));
  AOI21xp33_ASAP7_75t_L     g00416(.A1(new_n651), .A2(new_n657), .B(new_n624), .Y(new_n673));
  OAI21xp33_ASAP7_75t_L     g00417(.A1(new_n346), .A2(new_n667), .B(new_n669), .Y(new_n674));
  OAI21xp33_ASAP7_75t_L     g00418(.A1(new_n673), .A2(new_n672), .B(new_n674), .Y(new_n675));
  A2O1A1O1Ixp25_ASAP7_75t_L g00419(.A1(new_n528), .A2(new_n611), .B(new_n587), .C(new_n578), .D(new_n585), .Y(new_n676));
  NAND3xp33_ASAP7_75t_L     g00420(.A(new_n676), .B(new_n675), .C(new_n671), .Y(new_n677));
  NAND2xp33_ASAP7_75t_L     g00421(.A(new_n671), .B(new_n675), .Y(new_n678));
  A2O1A1Ixp33_ASAP7_75t_L   g00422(.A1(new_n582), .A2(new_n578), .B(new_n585), .C(new_n678), .Y(new_n679));
  INVx1_ASAP7_75t_L         g00423(.A(\b[10] ), .Y(new_n680));
  NAND2xp33_ASAP7_75t_L     g00424(.A(\b[8] ), .B(new_n286), .Y(new_n681));
  OAI221xp5_ASAP7_75t_L     g00425(.A1(new_n285), .A2(new_n590), .B1(new_n680), .B2(new_n269), .C(new_n681), .Y(new_n682));
  A2O1A1Ixp33_ASAP7_75t_L   g00426(.A1(new_n453), .A2(new_n450), .B(new_n533), .C(new_n593), .Y(new_n683));
  NOR2xp33_ASAP7_75t_L      g00427(.A(\b[9] ), .B(\b[10] ), .Y(new_n684));
  NOR2xp33_ASAP7_75t_L      g00428(.A(new_n590), .B(new_n680), .Y(new_n685));
  NOR2xp33_ASAP7_75t_L      g00429(.A(new_n684), .B(new_n685), .Y(new_n686));
  A2O1A1Ixp33_ASAP7_75t_L   g00430(.A1(new_n683), .A2(new_n596), .B(new_n595), .C(new_n686), .Y(new_n687));
  INVx1_ASAP7_75t_L         g00431(.A(new_n595), .Y(new_n688));
  OAI221xp5_ASAP7_75t_L     g00432(.A1(new_n685), .A2(new_n684), .B1(new_n594), .B2(new_n599), .C(new_n688), .Y(new_n689));
  AND2x2_ASAP7_75t_L        g00433(.A(new_n689), .B(new_n687), .Y(new_n690));
  A2O1A1Ixp33_ASAP7_75t_L   g00434(.A1(new_n690), .A2(new_n273), .B(new_n682), .C(\a[2] ), .Y(new_n691));
  NAND2xp33_ASAP7_75t_L     g00435(.A(\a[2] ), .B(new_n691), .Y(new_n692));
  A2O1A1Ixp33_ASAP7_75t_L   g00436(.A1(new_n690), .A2(new_n273), .B(new_n682), .C(new_n257), .Y(new_n693));
  NAND2xp33_ASAP7_75t_L     g00437(.A(new_n693), .B(new_n692), .Y(new_n694));
  AO21x2_ASAP7_75t_L        g00438(.A1(new_n679), .A2(new_n677), .B(new_n694), .Y(new_n695));
  NAND3xp33_ASAP7_75t_L     g00439(.A(new_n677), .B(new_n679), .C(new_n694), .Y(new_n696));
  NAND2xp33_ASAP7_75t_L     g00440(.A(new_n696), .B(new_n695), .Y(new_n697));
  XOR2x2_ASAP7_75t_L        g00441(.A(new_n697), .B(new_n622), .Y(\f[10] ));
  AOI21xp33_ASAP7_75t_L     g00442(.A1(new_n677), .A2(new_n679), .B(new_n694), .Y(new_n699));
  NAND2xp33_ASAP7_75t_L     g00443(.A(new_n664), .B(new_n658), .Y(new_n700));
  O2A1O1Ixp33_ASAP7_75t_L   g00444(.A1(new_n667), .A2(new_n346), .B(new_n669), .C(new_n700), .Y(new_n701));
  A2O1A1O1Ixp25_ASAP7_75t_L g00445(.A1(new_n578), .A2(new_n582), .B(new_n585), .C(new_n678), .D(new_n701), .Y(new_n702));
  NOR2xp33_ASAP7_75t_L      g00446(.A(new_n427), .B(new_n375), .Y(new_n703));
  AOI221xp5_ASAP7_75t_L     g00447(.A1(\b[8] ), .A2(new_n361), .B1(new_n349), .B2(\b[7] ), .C(new_n703), .Y(new_n704));
  O2A1O1Ixp33_ASAP7_75t_L   g00448(.A1(new_n356), .A2(new_n540), .B(new_n704), .C(new_n346), .Y(new_n705));
  O2A1O1Ixp33_ASAP7_75t_L   g00449(.A1(new_n356), .A2(new_n540), .B(new_n704), .C(\a[5] ), .Y(new_n706));
  INVx1_ASAP7_75t_L         g00450(.A(new_n706), .Y(new_n707));
  OAI21xp33_ASAP7_75t_L     g00451(.A1(new_n346), .A2(new_n705), .B(new_n707), .Y(new_n708));
  OAI21xp33_ASAP7_75t_L     g00452(.A1(new_n660), .A2(new_n661), .B(new_n657), .Y(new_n709));
  NAND3xp33_ASAP7_75t_L     g00453(.A(new_n630), .B(new_n636), .C(new_n638), .Y(new_n710));
  NOR2xp33_ASAP7_75t_L      g00454(.A(new_n289), .B(new_n710), .Y(new_n711));
  NAND3xp33_ASAP7_75t_L     g00455(.A(new_n553), .B(new_n634), .C(new_n639), .Y(new_n712));
  INVx1_ASAP7_75t_L         g00456(.A(new_n712), .Y(new_n713));
  AOI221xp5_ASAP7_75t_L     g00457(.A1(\b[1] ), .A2(new_n635), .B1(\b[0] ), .B2(new_n713), .C(new_n711), .Y(new_n714));
  NOR2xp33_ASAP7_75t_L      g00458(.A(new_n641), .B(new_n509), .Y(new_n715));
  INVx1_ASAP7_75t_L         g00459(.A(new_n715), .Y(new_n716));
  NAND3xp33_ASAP7_75t_L     g00460(.A(new_n714), .B(\a[11] ), .C(new_n716), .Y(new_n717));
  INVx1_ASAP7_75t_L         g00461(.A(new_n641), .Y(new_n718));
  NAND2xp33_ASAP7_75t_L     g00462(.A(\b[1] ), .B(new_n635), .Y(new_n719));
  OAI221xp5_ASAP7_75t_L     g00463(.A1(new_n710), .A2(new_n289), .B1(new_n284), .B2(new_n712), .C(new_n719), .Y(new_n720));
  A2O1A1Ixp33_ASAP7_75t_L   g00464(.A1(new_n294), .A2(new_n718), .B(new_n720), .C(new_n637), .Y(new_n721));
  NAND3xp33_ASAP7_75t_L     g00465(.A(new_n717), .B(new_n644), .C(new_n721), .Y(new_n722));
  NAND5xp2_ASAP7_75t_L      g00466(.A(\a[11] ), .B(new_n714), .C(new_n643), .D(new_n716), .E(new_n623), .Y(new_n723));
  NOR2xp33_ASAP7_75t_L      g00467(.A(new_n301), .B(new_n506), .Y(new_n724));
  AOI221xp5_ASAP7_75t_L     g00468(.A1(\b[5] ), .A2(new_n475), .B1(new_n470), .B2(\b[4] ), .C(new_n724), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g00469(.A(new_n483), .B(new_n394), .Y(new_n726));
  NAND3xp33_ASAP7_75t_L     g00470(.A(new_n726), .B(new_n725), .C(\a[8] ), .Y(new_n727));
  NAND2xp33_ASAP7_75t_L     g00471(.A(new_n391), .B(new_n393), .Y(new_n728));
  OAI21xp33_ASAP7_75t_L     g00472(.A1(new_n728), .A2(new_n477), .B(new_n725), .Y(new_n729));
  NAND2xp33_ASAP7_75t_L     g00473(.A(new_n466), .B(new_n729), .Y(new_n730));
  AND4x1_ASAP7_75t_L        g00474(.A(new_n722), .B(new_n730), .C(new_n727), .D(new_n723), .Y(new_n731));
  AOI22xp33_ASAP7_75t_L     g00475(.A1(new_n727), .A2(new_n730), .B1(new_n723), .B2(new_n722), .Y(new_n732));
  OAI21xp33_ASAP7_75t_L     g00476(.A1(new_n731), .A2(new_n732), .B(new_n709), .Y(new_n733));
  AOI21xp33_ASAP7_75t_L     g00477(.A1(new_n624), .A2(new_n651), .B(new_n663), .Y(new_n734));
  NOR2xp33_ASAP7_75t_L      g00478(.A(new_n732), .B(new_n731), .Y(new_n735));
  NAND2xp33_ASAP7_75t_L     g00479(.A(new_n735), .B(new_n734), .Y(new_n736));
  NAND3xp33_ASAP7_75t_L     g00480(.A(new_n736), .B(new_n733), .C(new_n708), .Y(new_n737));
  NOR2xp33_ASAP7_75t_L      g00481(.A(new_n346), .B(new_n705), .Y(new_n738));
  NOR2xp33_ASAP7_75t_L      g00482(.A(new_n706), .B(new_n738), .Y(new_n739));
  AND3x1_ASAP7_75t_L        g00483(.A(new_n736), .B(new_n739), .C(new_n733), .Y(new_n740));
  AOI21xp33_ASAP7_75t_L     g00484(.A1(new_n737), .A2(new_n708), .B(new_n740), .Y(new_n741));
  O2A1O1Ixp33_ASAP7_75t_L   g00485(.A1(new_n700), .A2(new_n670), .B(new_n679), .C(new_n741), .Y(new_n742));
  A2O1A1Ixp33_ASAP7_75t_L   g00486(.A1(new_n708), .A2(new_n737), .B(new_n740), .C(new_n702), .Y(new_n743));
  NOR2xp33_ASAP7_75t_L      g00487(.A(new_n590), .B(new_n287), .Y(new_n744));
  AOI221xp5_ASAP7_75t_L     g00488(.A1(\b[10] ), .A2(new_n264), .B1(\b[11] ), .B2(new_n283), .C(new_n744), .Y(new_n745));
  A2O1A1Ixp33_ASAP7_75t_L   g00489(.A1(new_n537), .A2(new_n593), .B(new_n594), .C(new_n688), .Y(new_n746));
  NOR2xp33_ASAP7_75t_L      g00490(.A(\b[10] ), .B(\b[11] ), .Y(new_n747));
  INVx1_ASAP7_75t_L         g00491(.A(\b[11] ), .Y(new_n748));
  NOR2xp33_ASAP7_75t_L      g00492(.A(new_n680), .B(new_n748), .Y(new_n749));
  NOR2xp33_ASAP7_75t_L      g00493(.A(new_n747), .B(new_n749), .Y(new_n750));
  A2O1A1Ixp33_ASAP7_75t_L   g00494(.A1(new_n746), .A2(new_n686), .B(new_n685), .C(new_n750), .Y(new_n751));
  A2O1A1O1Ixp25_ASAP7_75t_L g00495(.A1(new_n596), .A2(new_n683), .B(new_n595), .C(new_n686), .D(new_n685), .Y(new_n752));
  OAI21xp33_ASAP7_75t_L     g00496(.A1(new_n747), .A2(new_n749), .B(new_n752), .Y(new_n753));
  NAND2xp33_ASAP7_75t_L     g00497(.A(new_n751), .B(new_n753), .Y(new_n754));
  O2A1O1Ixp33_ASAP7_75t_L   g00498(.A1(new_n279), .A2(new_n754), .B(new_n745), .C(new_n257), .Y(new_n755));
  OAI21xp33_ASAP7_75t_L     g00499(.A1(new_n279), .A2(new_n754), .B(new_n745), .Y(new_n756));
  NAND2xp33_ASAP7_75t_L     g00500(.A(new_n257), .B(new_n756), .Y(new_n757));
  OAI21xp33_ASAP7_75t_L     g00501(.A1(new_n257), .A2(new_n755), .B(new_n757), .Y(new_n758));
  O2A1O1Ixp33_ASAP7_75t_L   g00502(.A1(new_n702), .A2(new_n742), .B(new_n743), .C(new_n758), .Y(new_n759));
  AO21x2_ASAP7_75t_L        g00503(.A1(new_n733), .A2(new_n736), .B(new_n739), .Y(new_n760));
  NAND3xp33_ASAP7_75t_L     g00504(.A(new_n736), .B(new_n739), .C(new_n733), .Y(new_n761));
  MAJIxp5_ASAP7_75t_L       g00505(.A(new_n588), .B(new_n584), .C(new_n575), .Y(new_n762));
  A2O1A1Ixp33_ASAP7_75t_L   g00506(.A1(new_n678), .A2(new_n762), .B(new_n701), .C(new_n741), .Y(new_n763));
  A2O1A1Ixp33_ASAP7_75t_L   g00507(.A1(new_n761), .A2(new_n760), .B(new_n742), .C(new_n763), .Y(new_n764));
  O2A1O1Ixp33_ASAP7_75t_L   g00508(.A1(new_n755), .A2(new_n257), .B(new_n757), .C(new_n764), .Y(new_n765));
  NOR2xp33_ASAP7_75t_L      g00509(.A(new_n759), .B(new_n765), .Y(new_n766));
  O2A1O1Ixp33_ASAP7_75t_L   g00510(.A1(new_n622), .A2(new_n699), .B(new_n696), .C(new_n766), .Y(new_n767));
  A2O1A1Ixp33_ASAP7_75t_L   g00511(.A1(new_n615), .A2(new_n620), .B(new_n699), .C(new_n696), .Y(new_n768));
  NOR3xp33_ASAP7_75t_L      g00512(.A(new_n765), .B(new_n759), .C(new_n768), .Y(new_n769));
  NOR2xp33_ASAP7_75t_L      g00513(.A(new_n769), .B(new_n767), .Y(\f[11] ));
  INVx1_ASAP7_75t_L         g00514(.A(new_n702), .Y(new_n771));
  INVx1_ASAP7_75t_L         g00515(.A(new_n737), .Y(new_n772));
  NAND2xp33_ASAP7_75t_L     g00516(.A(new_n761), .B(new_n760), .Y(new_n773));
  INVx1_ASAP7_75t_L         g00517(.A(\a[12] ), .Y(new_n774));
  NAND2xp33_ASAP7_75t_L     g00518(.A(\a[11] ), .B(new_n774), .Y(new_n775));
  NAND2xp33_ASAP7_75t_L     g00519(.A(\a[12] ), .B(new_n637), .Y(new_n776));
  AND2x2_ASAP7_75t_L        g00520(.A(new_n775), .B(new_n776), .Y(new_n777));
  NOR2xp33_ASAP7_75t_L      g00521(.A(new_n284), .B(new_n777), .Y(new_n778));
  A2O1A1Ixp33_ASAP7_75t_L   g00522(.A1(new_n717), .A2(new_n721), .B(new_n644), .C(new_n778), .Y(new_n779));
  NOR5xp2_ASAP7_75t_L       g00523(.A(new_n647), .B(new_n720), .C(new_n715), .D(new_n554), .E(new_n637), .Y(new_n780));
  A2O1A1Ixp33_ASAP7_75t_L   g00524(.A1(new_n775), .A2(new_n776), .B(new_n284), .C(new_n780), .Y(new_n781));
  NAND2xp33_ASAP7_75t_L     g00525(.A(\b[3] ), .B(new_n640), .Y(new_n782));
  NAND2xp33_ASAP7_75t_L     g00526(.A(\b[2] ), .B(new_n635), .Y(new_n783));
  OAI211xp5_ASAP7_75t_L     g00527(.A1(new_n712), .A2(new_n262), .B(new_n782), .C(new_n783), .Y(new_n784));
  NOR2xp33_ASAP7_75t_L      g00528(.A(new_n641), .B(new_n319), .Y(new_n785));
  A2O1A1Ixp33_ASAP7_75t_L   g00529(.A1(new_n312), .A2(new_n718), .B(new_n784), .C(\a[11] ), .Y(new_n786));
  AOI211xp5_ASAP7_75t_L     g00530(.A1(new_n312), .A2(new_n718), .B(new_n637), .C(new_n784), .Y(new_n787));
  O2A1O1Ixp33_ASAP7_75t_L   g00531(.A1(new_n784), .A2(new_n785), .B(new_n786), .C(new_n787), .Y(new_n788));
  AOI21xp33_ASAP7_75t_L     g00532(.A1(new_n781), .A2(new_n779), .B(new_n788), .Y(new_n789));
  INVx1_ASAP7_75t_L         g00533(.A(new_n789), .Y(new_n790));
  NAND3xp33_ASAP7_75t_L     g00534(.A(new_n781), .B(new_n779), .C(new_n788), .Y(new_n791));
  NOR2xp33_ASAP7_75t_L      g00535(.A(new_n332), .B(new_n506), .Y(new_n792));
  AOI221xp5_ASAP7_75t_L     g00536(.A1(\b[6] ), .A2(new_n475), .B1(new_n470), .B2(\b[5] ), .C(new_n792), .Y(new_n793));
  O2A1O1Ixp33_ASAP7_75t_L   g00537(.A1(new_n477), .A2(new_n434), .B(new_n793), .C(new_n466), .Y(new_n794));
  OAI21xp33_ASAP7_75t_L     g00538(.A1(new_n477), .A2(new_n434), .B(new_n793), .Y(new_n795));
  NAND2xp33_ASAP7_75t_L     g00539(.A(new_n466), .B(new_n795), .Y(new_n796));
  OAI21xp33_ASAP7_75t_L     g00540(.A1(new_n466), .A2(new_n794), .B(new_n796), .Y(new_n797));
  INVx1_ASAP7_75t_L         g00541(.A(new_n797), .Y(new_n798));
  NAND3xp33_ASAP7_75t_L     g00542(.A(new_n798), .B(new_n790), .C(new_n791), .Y(new_n799));
  INVx1_ASAP7_75t_L         g00543(.A(new_n791), .Y(new_n800));
  OAI21xp33_ASAP7_75t_L     g00544(.A1(new_n789), .A2(new_n800), .B(new_n797), .Y(new_n801));
  AND2x2_ASAP7_75t_L        g00545(.A(new_n723), .B(new_n722), .Y(new_n802));
  NAND2xp33_ASAP7_75t_L     g00546(.A(new_n723), .B(new_n722), .Y(new_n803));
  O2A1O1Ixp33_ASAP7_75t_L   g00547(.A1(new_n728), .A2(new_n477), .B(new_n725), .C(new_n466), .Y(new_n804));
  O2A1O1Ixp33_ASAP7_75t_L   g00548(.A1(new_n804), .A2(new_n466), .B(new_n730), .C(new_n803), .Y(new_n805));
  O2A1O1Ixp33_ASAP7_75t_L   g00549(.A1(new_n732), .A2(new_n802), .B(new_n709), .C(new_n805), .Y(new_n806));
  NAND3xp33_ASAP7_75t_L     g00550(.A(new_n806), .B(new_n801), .C(new_n799), .Y(new_n807));
  NOR3xp33_ASAP7_75t_L      g00551(.A(new_n800), .B(new_n797), .C(new_n789), .Y(new_n808));
  AOI21xp33_ASAP7_75t_L     g00552(.A1(new_n790), .A2(new_n791), .B(new_n798), .Y(new_n809));
  A2O1A1Ixp33_ASAP7_75t_L   g00553(.A1(new_n726), .A2(new_n725), .B(new_n804), .C(new_n727), .Y(new_n810));
  NAND2xp33_ASAP7_75t_L     g00554(.A(new_n810), .B(new_n802), .Y(new_n811));
  OAI21xp33_ASAP7_75t_L     g00555(.A1(new_n735), .A2(new_n734), .B(new_n811), .Y(new_n812));
  OAI21xp33_ASAP7_75t_L     g00556(.A1(new_n808), .A2(new_n809), .B(new_n812), .Y(new_n813));
  OAI22xp33_ASAP7_75t_L     g00557(.A1(new_n350), .A2(new_n534), .B1(new_n448), .B2(new_n375), .Y(new_n814));
  AOI221xp5_ASAP7_75t_L     g00558(.A1(new_n361), .A2(\b[9] ), .B1(new_n359), .B2(new_n602), .C(new_n814), .Y(new_n815));
  XNOR2x2_ASAP7_75t_L       g00559(.A(\a[5] ), .B(new_n815), .Y(new_n816));
  AOI21xp33_ASAP7_75t_L     g00560(.A1(new_n807), .A2(new_n813), .B(new_n816), .Y(new_n817));
  NOR3xp33_ASAP7_75t_L      g00561(.A(new_n812), .B(new_n809), .C(new_n808), .Y(new_n818));
  AOI21xp33_ASAP7_75t_L     g00562(.A1(new_n801), .A2(new_n799), .B(new_n806), .Y(new_n819));
  XNOR2x2_ASAP7_75t_L       g00563(.A(new_n346), .B(new_n815), .Y(new_n820));
  NOR3xp33_ASAP7_75t_L      g00564(.A(new_n820), .B(new_n818), .C(new_n819), .Y(new_n821));
  NOR2xp33_ASAP7_75t_L      g00565(.A(new_n817), .B(new_n821), .Y(new_n822));
  A2O1A1Ixp33_ASAP7_75t_L   g00566(.A1(new_n771), .A2(new_n773), .B(new_n772), .C(new_n822), .Y(new_n823));
  INVx1_ASAP7_75t_L         g00567(.A(new_n817), .Y(new_n824));
  INVx1_ASAP7_75t_L         g00568(.A(new_n821), .Y(new_n825));
  NAND2xp33_ASAP7_75t_L     g00569(.A(new_n824), .B(new_n825), .Y(new_n826));
  A2O1A1O1Ixp25_ASAP7_75t_L g00570(.A1(new_n678), .A2(new_n762), .B(new_n701), .C(new_n773), .D(new_n772), .Y(new_n827));
  NAND2xp33_ASAP7_75t_L     g00571(.A(new_n827), .B(new_n826), .Y(new_n828));
  NAND2xp33_ASAP7_75t_L     g00572(.A(new_n823), .B(new_n828), .Y(new_n829));
  NOR2xp33_ASAP7_75t_L      g00573(.A(new_n680), .B(new_n287), .Y(new_n830));
  AOI221xp5_ASAP7_75t_L     g00574(.A1(\b[11] ), .A2(new_n264), .B1(\b[12] ), .B2(new_n283), .C(new_n830), .Y(new_n831));
  NOR2xp33_ASAP7_75t_L      g00575(.A(\b[11] ), .B(\b[12] ), .Y(new_n832));
  INVx1_ASAP7_75t_L         g00576(.A(\b[12] ), .Y(new_n833));
  NOR2xp33_ASAP7_75t_L      g00577(.A(new_n748), .B(new_n833), .Y(new_n834));
  NOR2xp33_ASAP7_75t_L      g00578(.A(new_n832), .B(new_n834), .Y(new_n835));
  INVx1_ASAP7_75t_L         g00579(.A(new_n835), .Y(new_n836));
  O2A1O1Ixp33_ASAP7_75t_L   g00580(.A1(new_n680), .A2(new_n748), .B(new_n751), .C(new_n836), .Y(new_n837));
  INVx1_ASAP7_75t_L         g00581(.A(new_n837), .Y(new_n838));
  A2O1A1O1Ixp25_ASAP7_75t_L g00582(.A1(new_n686), .A2(new_n746), .B(new_n685), .C(new_n750), .D(new_n749), .Y(new_n839));
  NAND2xp33_ASAP7_75t_L     g00583(.A(new_n836), .B(new_n839), .Y(new_n840));
  NAND2xp33_ASAP7_75t_L     g00584(.A(new_n840), .B(new_n838), .Y(new_n841));
  OAI21xp33_ASAP7_75t_L     g00585(.A1(new_n279), .A2(new_n841), .B(new_n831), .Y(new_n842));
  NAND2xp33_ASAP7_75t_L     g00586(.A(\a[2] ), .B(new_n842), .Y(new_n843));
  O2A1O1Ixp33_ASAP7_75t_L   g00587(.A1(new_n279), .A2(new_n841), .B(new_n831), .C(\a[2] ), .Y(new_n844));
  AOI21xp33_ASAP7_75t_L     g00588(.A1(new_n843), .A2(\a[2] ), .B(new_n844), .Y(new_n845));
  NOR2xp33_ASAP7_75t_L      g00589(.A(new_n845), .B(new_n829), .Y(new_n846));
  A2O1A1Ixp33_ASAP7_75t_L   g00590(.A1(\a[2] ), .A2(new_n843), .B(new_n844), .C(new_n829), .Y(new_n847));
  MAJIxp5_ASAP7_75t_L       g00591(.A(new_n768), .B(new_n764), .C(new_n758), .Y(new_n848));
  O2A1O1Ixp33_ASAP7_75t_L   g00592(.A1(new_n829), .A2(new_n846), .B(new_n847), .C(new_n848), .Y(new_n849));
  OAI21xp33_ASAP7_75t_L     g00593(.A1(new_n829), .A2(new_n846), .B(new_n847), .Y(new_n850));
  INVx1_ASAP7_75t_L         g00594(.A(new_n848), .Y(new_n851));
  NOR2xp33_ASAP7_75t_L      g00595(.A(new_n851), .B(new_n850), .Y(new_n852));
  NOR2xp33_ASAP7_75t_L      g00596(.A(new_n849), .B(new_n852), .Y(\f[12] ));
  INVx1_ASAP7_75t_L         g00597(.A(new_n778), .Y(new_n854));
  MAJIxp5_ASAP7_75t_L       g00598(.A(new_n788), .B(new_n723), .C(new_n854), .Y(new_n855));
  NAND2xp33_ASAP7_75t_L     g00599(.A(\b[3] ), .B(new_n635), .Y(new_n856));
  OAI221xp5_ASAP7_75t_L     g00600(.A1(new_n710), .A2(new_n332), .B1(new_n289), .B2(new_n712), .C(new_n856), .Y(new_n857));
  A2O1A1Ixp33_ASAP7_75t_L   g00601(.A1(new_n342), .A2(new_n718), .B(new_n857), .C(\a[11] ), .Y(new_n858));
  AOI211xp5_ASAP7_75t_L     g00602(.A1(new_n342), .A2(new_n718), .B(new_n637), .C(new_n857), .Y(new_n859));
  A2O1A1O1Ixp25_ASAP7_75t_L g00603(.A1(new_n718), .A2(new_n342), .B(new_n857), .C(new_n858), .D(new_n859), .Y(new_n860));
  INVx1_ASAP7_75t_L         g00604(.A(\a[13] ), .Y(new_n861));
  NOR2xp33_ASAP7_75t_L      g00605(.A(\a[12] ), .B(new_n861), .Y(new_n862));
  NOR2xp33_ASAP7_75t_L      g00606(.A(\a[13] ), .B(new_n774), .Y(new_n863));
  OAI21xp33_ASAP7_75t_L     g00607(.A1(new_n862), .A2(new_n863), .B(new_n777), .Y(new_n864));
  NAND2xp33_ASAP7_75t_L     g00608(.A(new_n776), .B(new_n775), .Y(new_n865));
  NAND2xp33_ASAP7_75t_L     g00609(.A(\a[14] ), .B(new_n861), .Y(new_n866));
  INVx1_ASAP7_75t_L         g00610(.A(\a[14] ), .Y(new_n867));
  NAND2xp33_ASAP7_75t_L     g00611(.A(\a[13] ), .B(new_n867), .Y(new_n868));
  NAND3xp33_ASAP7_75t_L     g00612(.A(new_n865), .B(new_n866), .C(new_n868), .Y(new_n869));
  OAI22xp33_ASAP7_75t_L     g00613(.A1(new_n864), .A2(new_n284), .B1(new_n262), .B2(new_n869), .Y(new_n870));
  NAND2xp33_ASAP7_75t_L     g00614(.A(new_n868), .B(new_n866), .Y(new_n871));
  NAND2xp33_ASAP7_75t_L     g00615(.A(new_n871), .B(new_n865), .Y(new_n872));
  INVx1_ASAP7_75t_L         g00616(.A(new_n872), .Y(new_n873));
  AOI21xp33_ASAP7_75t_L     g00617(.A1(new_n275), .A2(new_n873), .B(new_n870), .Y(new_n874));
  NAND3xp33_ASAP7_75t_L     g00618(.A(new_n874), .B(new_n854), .C(\a[14] ), .Y(new_n875));
  INVx1_ASAP7_75t_L         g00619(.A(new_n875), .Y(new_n876));
  A2O1A1Ixp33_ASAP7_75t_L   g00620(.A1(new_n873), .A2(new_n275), .B(new_n870), .C(\a[14] ), .Y(new_n877));
  A2O1A1Ixp33_ASAP7_75t_L   g00621(.A1(new_n873), .A2(new_n275), .B(new_n870), .C(new_n867), .Y(new_n878));
  INVx1_ASAP7_75t_L         g00622(.A(new_n878), .Y(new_n879));
  O2A1O1Ixp33_ASAP7_75t_L   g00623(.A1(new_n854), .A2(new_n877), .B(\a[14] ), .C(new_n879), .Y(new_n880));
  OAI21xp33_ASAP7_75t_L     g00624(.A1(new_n876), .A2(new_n880), .B(new_n860), .Y(new_n881));
  A2O1A1Ixp33_ASAP7_75t_L   g00625(.A1(new_n342), .A2(new_n718), .B(new_n857), .C(new_n637), .Y(new_n882));
  INVx1_ASAP7_75t_L         g00626(.A(new_n882), .Y(new_n883));
  NOR2xp33_ASAP7_75t_L      g00627(.A(new_n862), .B(new_n863), .Y(new_n884));
  NOR2xp33_ASAP7_75t_L      g00628(.A(new_n865), .B(new_n884), .Y(new_n885));
  NOR2xp33_ASAP7_75t_L      g00629(.A(new_n871), .B(new_n777), .Y(new_n886));
  AOI22xp33_ASAP7_75t_L     g00630(.A1(new_n885), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n886), .Y(new_n887));
  O2A1O1Ixp33_ASAP7_75t_L   g00631(.A1(new_n872), .A2(new_n274), .B(new_n887), .C(new_n867), .Y(new_n888));
  A2O1A1Ixp33_ASAP7_75t_L   g00632(.A1(new_n888), .A2(new_n778), .B(new_n867), .C(new_n878), .Y(new_n889));
  OAI211xp5_ASAP7_75t_L     g00633(.A1(new_n859), .A2(new_n883), .B(new_n875), .C(new_n889), .Y(new_n890));
  NAND3xp33_ASAP7_75t_L     g00634(.A(new_n855), .B(new_n890), .C(new_n881), .Y(new_n891));
  NAND2xp33_ASAP7_75t_L     g00635(.A(\b[1] ), .B(new_n713), .Y(new_n892));
  NAND2xp33_ASAP7_75t_L     g00636(.A(new_n718), .B(new_n312), .Y(new_n893));
  NAND5xp2_ASAP7_75t_L      g00637(.A(new_n893), .B(new_n783), .C(new_n892), .D(new_n782), .E(\a[11] ), .Y(new_n894));
  A2O1A1Ixp33_ASAP7_75t_L   g00638(.A1(new_n312), .A2(new_n718), .B(new_n784), .C(new_n637), .Y(new_n895));
  NAND2xp33_ASAP7_75t_L     g00639(.A(new_n894), .B(new_n895), .Y(new_n896));
  MAJIxp5_ASAP7_75t_L       g00640(.A(new_n896), .B(new_n778), .C(new_n780), .Y(new_n897));
  AOI211xp5_ASAP7_75t_L     g00641(.A1(new_n889), .A2(new_n875), .B(new_n859), .C(new_n883), .Y(new_n898));
  NOR3xp33_ASAP7_75t_L      g00642(.A(new_n860), .B(new_n876), .C(new_n880), .Y(new_n899));
  OAI21xp33_ASAP7_75t_L     g00643(.A1(new_n898), .A2(new_n899), .B(new_n897), .Y(new_n900));
  NOR2xp33_ASAP7_75t_L      g00644(.A(new_n384), .B(new_n506), .Y(new_n901));
  AOI221xp5_ASAP7_75t_L     g00645(.A1(\b[7] ), .A2(new_n475), .B1(new_n470), .B2(\b[6] ), .C(new_n901), .Y(new_n902));
  OAI21xp33_ASAP7_75t_L     g00646(.A1(new_n477), .A2(new_n456), .B(new_n902), .Y(new_n903));
  NOR2xp33_ASAP7_75t_L      g00647(.A(new_n466), .B(new_n903), .Y(new_n904));
  O2A1O1Ixp33_ASAP7_75t_L   g00648(.A1(new_n477), .A2(new_n456), .B(new_n902), .C(\a[8] ), .Y(new_n905));
  NOR2xp33_ASAP7_75t_L      g00649(.A(new_n905), .B(new_n904), .Y(new_n906));
  NAND3xp33_ASAP7_75t_L     g00650(.A(new_n891), .B(new_n900), .C(new_n906), .Y(new_n907));
  NOR3xp33_ASAP7_75t_L      g00651(.A(new_n899), .B(new_n898), .C(new_n897), .Y(new_n908));
  AOI21xp33_ASAP7_75t_L     g00652(.A1(new_n890), .A2(new_n881), .B(new_n855), .Y(new_n909));
  O2A1O1Ixp33_ASAP7_75t_L   g00653(.A1(new_n477), .A2(new_n456), .B(new_n902), .C(new_n466), .Y(new_n910));
  INVx1_ASAP7_75t_L         g00654(.A(new_n905), .Y(new_n911));
  OAI21xp33_ASAP7_75t_L     g00655(.A1(new_n466), .A2(new_n910), .B(new_n911), .Y(new_n912));
  OAI21xp33_ASAP7_75t_L     g00656(.A1(new_n909), .A2(new_n908), .B(new_n912), .Y(new_n913));
  NAND2xp33_ASAP7_75t_L     g00657(.A(new_n907), .B(new_n913), .Y(new_n914));
  NAND3xp33_ASAP7_75t_L     g00658(.A(new_n790), .B(new_n791), .C(new_n797), .Y(new_n915));
  A2O1A1Ixp33_ASAP7_75t_L   g00659(.A1(new_n798), .A2(new_n799), .B(new_n806), .C(new_n915), .Y(new_n916));
  NOR2xp33_ASAP7_75t_L      g00660(.A(new_n914), .B(new_n916), .Y(new_n917));
  NAND3xp33_ASAP7_75t_L     g00661(.A(new_n891), .B(new_n900), .C(new_n912), .Y(new_n918));
  NOR3xp33_ASAP7_75t_L      g00662(.A(new_n908), .B(new_n909), .C(new_n912), .Y(new_n919));
  O2A1O1Ixp33_ASAP7_75t_L   g00663(.A1(new_n904), .A2(new_n905), .B(new_n918), .C(new_n919), .Y(new_n920));
  A2O1A1O1Ixp25_ASAP7_75t_L g00664(.A1(new_n799), .A2(new_n798), .B(new_n806), .C(new_n915), .D(new_n920), .Y(new_n921));
  OAI22xp33_ASAP7_75t_L     g00665(.A1(new_n350), .A2(new_n590), .B1(new_n534), .B2(new_n375), .Y(new_n922));
  AOI221xp5_ASAP7_75t_L     g00666(.A1(new_n361), .A2(\b[10] ), .B1(new_n359), .B2(new_n690), .C(new_n922), .Y(new_n923));
  XNOR2x2_ASAP7_75t_L       g00667(.A(new_n346), .B(new_n923), .Y(new_n924));
  OAI21xp33_ASAP7_75t_L     g00668(.A1(new_n917), .A2(new_n921), .B(new_n924), .Y(new_n925));
  INVx1_ASAP7_75t_L         g00669(.A(new_n701), .Y(new_n926));
  A2O1A1Ixp33_ASAP7_75t_L   g00670(.A1(new_n679), .A2(new_n926), .B(new_n741), .C(new_n737), .Y(new_n927));
  AOI21xp33_ASAP7_75t_L     g00671(.A1(new_n927), .A2(new_n824), .B(new_n821), .Y(new_n928));
  NOR3xp33_ASAP7_75t_L      g00672(.A(new_n921), .B(new_n924), .C(new_n917), .Y(new_n929));
  INVx1_ASAP7_75t_L         g00673(.A(new_n929), .Y(new_n930));
  AOI21xp33_ASAP7_75t_L     g00674(.A1(new_n925), .A2(new_n930), .B(new_n928), .Y(new_n931));
  A2O1A1O1Ixp25_ASAP7_75t_L g00675(.A1(new_n822), .A2(new_n927), .B(new_n821), .C(new_n925), .D(new_n929), .Y(new_n932));
  NOR2xp33_ASAP7_75t_L      g00676(.A(new_n748), .B(new_n287), .Y(new_n933));
  AOI221xp5_ASAP7_75t_L     g00677(.A1(\b[12] ), .A2(new_n264), .B1(\b[13] ), .B2(new_n283), .C(new_n933), .Y(new_n934));
  NOR2xp33_ASAP7_75t_L      g00678(.A(\b[12] ), .B(\b[13] ), .Y(new_n935));
  INVx1_ASAP7_75t_L         g00679(.A(\b[13] ), .Y(new_n936));
  NOR2xp33_ASAP7_75t_L      g00680(.A(new_n833), .B(new_n936), .Y(new_n937));
  NOR2xp33_ASAP7_75t_L      g00681(.A(new_n935), .B(new_n937), .Y(new_n938));
  A2O1A1Ixp33_ASAP7_75t_L   g00682(.A1(\b[12] ), .A2(\b[11] ), .B(new_n837), .C(new_n938), .Y(new_n939));
  NOR3xp33_ASAP7_75t_L      g00683(.A(new_n837), .B(new_n938), .C(new_n834), .Y(new_n940));
  INVx1_ASAP7_75t_L         g00684(.A(new_n940), .Y(new_n941));
  NAND2xp33_ASAP7_75t_L     g00685(.A(new_n939), .B(new_n941), .Y(new_n942));
  OAI21xp33_ASAP7_75t_L     g00686(.A1(new_n279), .A2(new_n942), .B(new_n934), .Y(new_n943));
  NOR2xp33_ASAP7_75t_L      g00687(.A(new_n257), .B(new_n943), .Y(new_n944));
  O2A1O1Ixp33_ASAP7_75t_L   g00688(.A1(new_n279), .A2(new_n942), .B(new_n934), .C(\a[2] ), .Y(new_n945));
  NOR2xp33_ASAP7_75t_L      g00689(.A(new_n945), .B(new_n944), .Y(new_n946));
  A2O1A1Ixp33_ASAP7_75t_L   g00690(.A1(new_n932), .A2(new_n925), .B(new_n931), .C(new_n946), .Y(new_n947));
  A2O1A1Ixp33_ASAP7_75t_L   g00691(.A1(new_n678), .A2(new_n762), .B(new_n701), .C(new_n773), .Y(new_n948));
  A2O1A1Ixp33_ASAP7_75t_L   g00692(.A1(new_n948), .A2(new_n737), .B(new_n817), .C(new_n825), .Y(new_n949));
  INVx1_ASAP7_75t_L         g00693(.A(new_n925), .Y(new_n950));
  OAI21xp33_ASAP7_75t_L     g00694(.A1(new_n929), .A2(new_n950), .B(new_n949), .Y(new_n951));
  NAND3xp33_ASAP7_75t_L     g00695(.A(new_n928), .B(new_n930), .C(new_n925), .Y(new_n952));
  OAI211xp5_ASAP7_75t_L     g00696(.A1(new_n944), .A2(new_n945), .B(new_n952), .C(new_n951), .Y(new_n953));
  NAND2xp33_ASAP7_75t_L     g00697(.A(new_n947), .B(new_n953), .Y(new_n954));
  A2O1A1Ixp33_ASAP7_75t_L   g00698(.A1(new_n850), .A2(new_n851), .B(new_n846), .C(new_n954), .Y(new_n955));
  INVx1_ASAP7_75t_L         g00699(.A(new_n955), .Y(new_n956));
  MAJIxp5_ASAP7_75t_L       g00700(.A(new_n848), .B(new_n829), .C(new_n845), .Y(new_n957));
  NOR2xp33_ASAP7_75t_L      g00701(.A(new_n954), .B(new_n957), .Y(new_n958));
  NOR2xp33_ASAP7_75t_L      g00702(.A(new_n958), .B(new_n956), .Y(\f[13] ));
  INVx1_ASAP7_75t_L         g00703(.A(\b[14] ), .Y(new_n960));
  NAND2xp33_ASAP7_75t_L     g00704(.A(\b[12] ), .B(new_n286), .Y(new_n961));
  OAI221xp5_ASAP7_75t_L     g00705(.A1(new_n285), .A2(new_n936), .B1(new_n960), .B2(new_n269), .C(new_n961), .Y(new_n962));
  NOR2xp33_ASAP7_75t_L      g00706(.A(\b[13] ), .B(\b[14] ), .Y(new_n963));
  NOR2xp33_ASAP7_75t_L      g00707(.A(new_n936), .B(new_n960), .Y(new_n964));
  NOR2xp33_ASAP7_75t_L      g00708(.A(new_n963), .B(new_n964), .Y(new_n965));
  INVx1_ASAP7_75t_L         g00709(.A(new_n965), .Y(new_n966));
  O2A1O1Ixp33_ASAP7_75t_L   g00710(.A1(new_n833), .A2(new_n936), .B(new_n939), .C(new_n966), .Y(new_n967));
  O2A1O1Ixp33_ASAP7_75t_L   g00711(.A1(new_n834), .A2(new_n837), .B(new_n938), .C(new_n937), .Y(new_n968));
  NAND2xp33_ASAP7_75t_L     g00712(.A(new_n966), .B(new_n968), .Y(new_n969));
  INVx1_ASAP7_75t_L         g00713(.A(new_n969), .Y(new_n970));
  NOR2xp33_ASAP7_75t_L      g00714(.A(new_n967), .B(new_n970), .Y(new_n971));
  A2O1A1Ixp33_ASAP7_75t_L   g00715(.A1(new_n971), .A2(new_n273), .B(new_n962), .C(\a[2] ), .Y(new_n972));
  AOI211xp5_ASAP7_75t_L     g00716(.A1(new_n971), .A2(new_n273), .B(new_n962), .C(new_n257), .Y(new_n973));
  A2O1A1O1Ixp25_ASAP7_75t_L g00717(.A1(new_n273), .A2(new_n971), .B(new_n962), .C(new_n972), .D(new_n973), .Y(new_n974));
  INVx1_ASAP7_75t_L         g00718(.A(new_n974), .Y(new_n975));
  AND2x2_ASAP7_75t_L        g00719(.A(new_n751), .B(new_n753), .Y(new_n976));
  OAI22xp33_ASAP7_75t_L     g00720(.A1(new_n350), .A2(new_n680), .B1(new_n590), .B2(new_n375), .Y(new_n977));
  AOI221xp5_ASAP7_75t_L     g00721(.A1(new_n361), .A2(\b[11] ), .B1(new_n359), .B2(new_n976), .C(new_n977), .Y(new_n978));
  XNOR2x2_ASAP7_75t_L       g00722(.A(new_n346), .B(new_n978), .Y(new_n979));
  NAND3xp33_ASAP7_75t_L     g00723(.A(new_n777), .B(new_n884), .C(new_n871), .Y(new_n980));
  NAND2xp33_ASAP7_75t_L     g00724(.A(\b[1] ), .B(new_n885), .Y(new_n981));
  OAI221xp5_ASAP7_75t_L     g00725(.A1(new_n869), .A2(new_n289), .B1(new_n284), .B2(new_n980), .C(new_n981), .Y(new_n982));
  A2O1A1Ixp33_ASAP7_75t_L   g00726(.A1(new_n294), .A2(new_n873), .B(new_n982), .C(\a[14] ), .Y(new_n983));
  NOR2xp33_ASAP7_75t_L      g00727(.A(new_n289), .B(new_n869), .Y(new_n984));
  AND3x1_ASAP7_75t_L        g00728(.A(new_n777), .B(new_n871), .C(new_n884), .Y(new_n985));
  AOI221xp5_ASAP7_75t_L     g00729(.A1(new_n885), .A2(\b[1] ), .B1(new_n985), .B2(\b[0] ), .C(new_n984), .Y(new_n986));
  O2A1O1Ixp33_ASAP7_75t_L   g00730(.A1(new_n509), .A2(new_n872), .B(new_n986), .C(\a[14] ), .Y(new_n987));
  A2O1A1O1Ixp25_ASAP7_75t_L g00731(.A1(new_n874), .A2(new_n854), .B(new_n983), .C(\a[14] ), .D(new_n987), .Y(new_n988));
  OAI21xp33_ASAP7_75t_L     g00732(.A1(new_n872), .A2(new_n274), .B(new_n887), .Y(new_n989));
  NOR2xp33_ASAP7_75t_L      g00733(.A(new_n872), .B(new_n509), .Y(new_n990));
  NOR5xp2_ASAP7_75t_L       g00734(.A(new_n989), .B(new_n982), .C(new_n990), .D(new_n778), .E(new_n867), .Y(new_n991));
  NAND2xp33_ASAP7_75t_L     g00735(.A(\b[4] ), .B(new_n635), .Y(new_n992));
  OAI221xp5_ASAP7_75t_L     g00736(.A1(new_n710), .A2(new_n384), .B1(new_n301), .B2(new_n712), .C(new_n992), .Y(new_n993));
  A2O1A1Ixp33_ASAP7_75t_L   g00737(.A1(new_n394), .A2(new_n718), .B(new_n993), .C(\a[11] ), .Y(new_n994));
  INVx1_ASAP7_75t_L         g00738(.A(new_n993), .Y(new_n995));
  O2A1O1Ixp33_ASAP7_75t_L   g00739(.A1(new_n641), .A2(new_n728), .B(new_n995), .C(\a[11] ), .Y(new_n996));
  AOI21xp33_ASAP7_75t_L     g00740(.A1(new_n994), .A2(\a[11] ), .B(new_n996), .Y(new_n997));
  NOR3xp33_ASAP7_75t_L      g00741(.A(new_n997), .B(new_n988), .C(new_n991), .Y(new_n998));
  INVx1_ASAP7_75t_L         g00742(.A(new_n990), .Y(new_n999));
  NAND3xp33_ASAP7_75t_L     g00743(.A(new_n986), .B(\a[14] ), .C(new_n999), .Y(new_n1000));
  A2O1A1Ixp33_ASAP7_75t_L   g00744(.A1(new_n294), .A2(new_n873), .B(new_n982), .C(new_n867), .Y(new_n1001));
  NAND3xp33_ASAP7_75t_L     g00745(.A(new_n875), .B(new_n1000), .C(new_n1001), .Y(new_n1002));
  NAND5xp2_ASAP7_75t_L      g00746(.A(\a[14] ), .B(new_n874), .C(new_n999), .D(new_n986), .E(new_n854), .Y(new_n1003));
  AOI221xp5_ASAP7_75t_L     g00747(.A1(new_n994), .A2(\a[11] ), .B1(new_n1003), .B2(new_n1002), .C(new_n996), .Y(new_n1004));
  OAI22xp33_ASAP7_75t_L     g00748(.A1(new_n908), .A2(new_n899), .B1(new_n1004), .B2(new_n998), .Y(new_n1005));
  AOI21xp33_ASAP7_75t_L     g00749(.A1(new_n855), .A2(new_n881), .B(new_n899), .Y(new_n1006));
  INVx1_ASAP7_75t_L         g00750(.A(new_n998), .Y(new_n1007));
  OAI21xp33_ASAP7_75t_L     g00751(.A1(new_n991), .A2(new_n988), .B(new_n997), .Y(new_n1008));
  NAND3xp33_ASAP7_75t_L     g00752(.A(new_n1006), .B(new_n1007), .C(new_n1008), .Y(new_n1009));
  NOR2xp33_ASAP7_75t_L      g00753(.A(new_n427), .B(new_n506), .Y(new_n1010));
  AOI221xp5_ASAP7_75t_L     g00754(.A1(\b[8] ), .A2(new_n475), .B1(new_n470), .B2(\b[7] ), .C(new_n1010), .Y(new_n1011));
  O2A1O1Ixp33_ASAP7_75t_L   g00755(.A1(new_n477), .A2(new_n540), .B(new_n1011), .C(new_n466), .Y(new_n1012));
  OAI21xp33_ASAP7_75t_L     g00756(.A1(new_n477), .A2(new_n540), .B(new_n1011), .Y(new_n1013));
  NAND2xp33_ASAP7_75t_L     g00757(.A(new_n466), .B(new_n1013), .Y(new_n1014));
  OA21x2_ASAP7_75t_L        g00758(.A1(new_n466), .A2(new_n1012), .B(new_n1014), .Y(new_n1015));
  NAND3xp33_ASAP7_75t_L     g00759(.A(new_n1005), .B(new_n1009), .C(new_n1015), .Y(new_n1016));
  AOI21xp33_ASAP7_75t_L     g00760(.A1(new_n1007), .A2(new_n1008), .B(new_n1006), .Y(new_n1017));
  A2O1A1O1Ixp25_ASAP7_75t_L g00761(.A1(new_n881), .A2(new_n855), .B(new_n899), .C(new_n1008), .D(new_n998), .Y(new_n1018));
  OAI21xp33_ASAP7_75t_L     g00762(.A1(new_n466), .A2(new_n1012), .B(new_n1014), .Y(new_n1019));
  A2O1A1Ixp33_ASAP7_75t_L   g00763(.A1(new_n1018), .A2(new_n1008), .B(new_n1017), .C(new_n1019), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g00764(.A(new_n1016), .B(new_n1020), .Y(new_n1021));
  A2O1A1O1Ixp25_ASAP7_75t_L g00765(.A1(new_n813), .A2(new_n915), .B(new_n920), .C(new_n918), .D(new_n1021), .Y(new_n1022));
  A2O1A1Ixp33_ASAP7_75t_L   g00766(.A1(new_n813), .A2(new_n915), .B(new_n920), .C(new_n918), .Y(new_n1023));
  AND2x2_ASAP7_75t_L        g00767(.A(new_n1016), .B(new_n1020), .Y(new_n1024));
  NOR2xp33_ASAP7_75t_L      g00768(.A(new_n1023), .B(new_n1024), .Y(new_n1025));
  OA21x2_ASAP7_75t_L        g00769(.A1(new_n1022), .A2(new_n1025), .B(new_n979), .Y(new_n1026));
  NOR3xp33_ASAP7_75t_L      g00770(.A(new_n1025), .B(new_n1022), .C(new_n979), .Y(new_n1027));
  NOR3xp33_ASAP7_75t_L      g00771(.A(new_n932), .B(new_n1026), .C(new_n1027), .Y(new_n1028));
  OAI21xp33_ASAP7_75t_L     g00772(.A1(new_n1026), .A2(new_n1027), .B(new_n932), .Y(new_n1029));
  INVx1_ASAP7_75t_L         g00773(.A(new_n1029), .Y(new_n1030));
  NOR3xp33_ASAP7_75t_L      g00774(.A(new_n1030), .B(new_n1028), .C(new_n975), .Y(new_n1031));
  NOR2xp33_ASAP7_75t_L      g00775(.A(new_n1027), .B(new_n1026), .Y(new_n1032));
  A2O1A1Ixp33_ASAP7_75t_L   g00776(.A1(new_n925), .A2(new_n949), .B(new_n929), .C(new_n1032), .Y(new_n1033));
  AOI21xp33_ASAP7_75t_L     g00777(.A1(new_n1033), .A2(new_n1029), .B(new_n974), .Y(new_n1034));
  NOR2xp33_ASAP7_75t_L      g00778(.A(new_n1031), .B(new_n1034), .Y(new_n1035));
  A2O1A1O1Ixp25_ASAP7_75t_L g00779(.A1(new_n952), .A2(new_n951), .B(new_n946), .C(new_n955), .D(new_n1035), .Y(new_n1036));
  INVx1_ASAP7_75t_L         g00780(.A(new_n932), .Y(new_n1037));
  O2A1O1Ixp33_ASAP7_75t_L   g00781(.A1(new_n950), .A2(new_n1037), .B(new_n951), .C(new_n946), .Y(new_n1038));
  AOI21xp33_ASAP7_75t_L     g00782(.A1(new_n957), .A2(new_n954), .B(new_n1038), .Y(new_n1039));
  AND2x2_ASAP7_75t_L        g00783(.A(new_n1035), .B(new_n1039), .Y(new_n1040));
  NOR2xp33_ASAP7_75t_L      g00784(.A(new_n1040), .B(new_n1036), .Y(\f[14] ));
  NOR2xp33_ASAP7_75t_L      g00785(.A(new_n1028), .B(new_n1030), .Y(new_n1042));
  INVx1_ASAP7_75t_L         g00786(.A(\b[15] ), .Y(new_n1043));
  NAND2xp33_ASAP7_75t_L     g00787(.A(\b[13] ), .B(new_n286), .Y(new_n1044));
  OAI221xp5_ASAP7_75t_L     g00788(.A1(new_n285), .A2(new_n960), .B1(new_n1043), .B2(new_n269), .C(new_n1044), .Y(new_n1045));
  NOR2xp33_ASAP7_75t_L      g00789(.A(\b[14] ), .B(\b[15] ), .Y(new_n1046));
  NOR2xp33_ASAP7_75t_L      g00790(.A(new_n960), .B(new_n1043), .Y(new_n1047));
  NOR2xp33_ASAP7_75t_L      g00791(.A(new_n1046), .B(new_n1047), .Y(new_n1048));
  A2O1A1Ixp33_ASAP7_75t_L   g00792(.A1(\b[14] ), .A2(\b[13] ), .B(new_n967), .C(new_n1048), .Y(new_n1049));
  INVx1_ASAP7_75t_L         g00793(.A(new_n1049), .Y(new_n1050));
  NOR3xp33_ASAP7_75t_L      g00794(.A(new_n967), .B(new_n1048), .C(new_n964), .Y(new_n1051));
  NOR2xp33_ASAP7_75t_L      g00795(.A(new_n1051), .B(new_n1050), .Y(new_n1052));
  A2O1A1Ixp33_ASAP7_75t_L   g00796(.A1(new_n1052), .A2(new_n273), .B(new_n1045), .C(\a[2] ), .Y(new_n1053));
  AOI211xp5_ASAP7_75t_L     g00797(.A1(new_n1052), .A2(new_n273), .B(new_n1045), .C(new_n257), .Y(new_n1054));
  A2O1A1O1Ixp25_ASAP7_75t_L g00798(.A1(new_n273), .A2(new_n1052), .B(new_n1045), .C(new_n1053), .D(new_n1054), .Y(new_n1055));
  INVx1_ASAP7_75t_L         g00799(.A(new_n1055), .Y(new_n1056));
  AND2x2_ASAP7_75t_L        g00800(.A(new_n840), .B(new_n838), .Y(new_n1057));
  NAND2xp33_ASAP7_75t_L     g00801(.A(\b[12] ), .B(new_n361), .Y(new_n1058));
  OAI221xp5_ASAP7_75t_L     g00802(.A1(new_n350), .A2(new_n748), .B1(new_n680), .B2(new_n375), .C(new_n1058), .Y(new_n1059));
  A2O1A1Ixp33_ASAP7_75t_L   g00803(.A1(new_n1057), .A2(new_n359), .B(new_n1059), .C(\a[5] ), .Y(new_n1060));
  AOI211xp5_ASAP7_75t_L     g00804(.A1(new_n1057), .A2(new_n359), .B(new_n1059), .C(new_n346), .Y(new_n1061));
  A2O1A1O1Ixp25_ASAP7_75t_L g00805(.A1(new_n1057), .A2(new_n359), .B(new_n1059), .C(new_n1060), .D(new_n1061), .Y(new_n1062));
  O2A1O1Ixp33_ASAP7_75t_L   g00806(.A1(new_n897), .A2(new_n898), .B(new_n890), .C(new_n1004), .Y(new_n1063));
  A2O1A1O1Ixp25_ASAP7_75t_L g00807(.A1(new_n1007), .A2(new_n1063), .B(new_n1006), .C(new_n1009), .D(new_n1015), .Y(new_n1064));
  INVx1_ASAP7_75t_L         g00808(.A(new_n598), .Y(new_n1065));
  NAND2xp33_ASAP7_75t_L     g00809(.A(new_n600), .B(new_n1065), .Y(new_n1066));
  NOR2xp33_ASAP7_75t_L      g00810(.A(new_n534), .B(new_n513), .Y(new_n1067));
  AOI221xp5_ASAP7_75t_L     g00811(.A1(\b[7] ), .A2(new_n560), .B1(\b[9] ), .B2(new_n475), .C(new_n1067), .Y(new_n1068));
  O2A1O1Ixp33_ASAP7_75t_L   g00812(.A1(new_n477), .A2(new_n1066), .B(new_n1068), .C(new_n466), .Y(new_n1069));
  INVx1_ASAP7_75t_L         g00813(.A(new_n1068), .Y(new_n1070));
  A2O1A1Ixp33_ASAP7_75t_L   g00814(.A1(new_n602), .A2(new_n483), .B(new_n1070), .C(new_n466), .Y(new_n1071));
  OAI21xp33_ASAP7_75t_L     g00815(.A1(new_n466), .A2(new_n1069), .B(new_n1071), .Y(new_n1072));
  INVx1_ASAP7_75t_L         g00816(.A(\a[15] ), .Y(new_n1073));
  NAND2xp33_ASAP7_75t_L     g00817(.A(\a[14] ), .B(new_n1073), .Y(new_n1074));
  NAND2xp33_ASAP7_75t_L     g00818(.A(\a[15] ), .B(new_n867), .Y(new_n1075));
  AND2x2_ASAP7_75t_L        g00819(.A(new_n1074), .B(new_n1075), .Y(new_n1076));
  NOR2xp33_ASAP7_75t_L      g00820(.A(new_n284), .B(new_n1076), .Y(new_n1077));
  INVx1_ASAP7_75t_L         g00821(.A(new_n1077), .Y(new_n1078));
  NOR2xp33_ASAP7_75t_L      g00822(.A(new_n1078), .B(new_n991), .Y(new_n1079));
  NOR2xp33_ASAP7_75t_L      g00823(.A(new_n1077), .B(new_n1003), .Y(new_n1080));
  NAND2xp33_ASAP7_75t_L     g00824(.A(\b[3] ), .B(new_n886), .Y(new_n1081));
  NAND2xp33_ASAP7_75t_L     g00825(.A(\b[1] ), .B(new_n985), .Y(new_n1082));
  NAND2xp33_ASAP7_75t_L     g00826(.A(\b[2] ), .B(new_n885), .Y(new_n1083));
  NAND2xp33_ASAP7_75t_L     g00827(.A(new_n873), .B(new_n312), .Y(new_n1084));
  NAND5xp2_ASAP7_75t_L      g00828(.A(new_n1084), .B(new_n1083), .C(new_n1082), .D(new_n1081), .E(\a[14] ), .Y(new_n1085));
  OAI211xp5_ASAP7_75t_L     g00829(.A1(new_n980), .A2(new_n262), .B(new_n1081), .C(new_n1083), .Y(new_n1086));
  A2O1A1Ixp33_ASAP7_75t_L   g00830(.A1(new_n312), .A2(new_n873), .B(new_n1086), .C(new_n867), .Y(new_n1087));
  NAND2xp33_ASAP7_75t_L     g00831(.A(new_n1085), .B(new_n1087), .Y(new_n1088));
  OAI21xp33_ASAP7_75t_L     g00832(.A1(new_n1080), .A2(new_n1079), .B(new_n1088), .Y(new_n1089));
  A2O1A1Ixp33_ASAP7_75t_L   g00833(.A1(new_n1000), .A2(new_n1001), .B(new_n875), .C(new_n1077), .Y(new_n1090));
  A2O1A1Ixp33_ASAP7_75t_L   g00834(.A1(new_n1074), .A2(new_n1075), .B(new_n284), .C(new_n991), .Y(new_n1091));
  NAND4xp25_ASAP7_75t_L     g00835(.A(new_n1084), .B(new_n1081), .C(new_n1082), .D(new_n1083), .Y(new_n1092));
  A2O1A1Ixp33_ASAP7_75t_L   g00836(.A1(new_n312), .A2(new_n873), .B(new_n1086), .C(\a[14] ), .Y(new_n1093));
  AOI211xp5_ASAP7_75t_L     g00837(.A1(new_n312), .A2(new_n873), .B(new_n867), .C(new_n1086), .Y(new_n1094));
  AOI21xp33_ASAP7_75t_L     g00838(.A1(new_n1093), .A2(new_n1092), .B(new_n1094), .Y(new_n1095));
  NAND3xp33_ASAP7_75t_L     g00839(.A(new_n1091), .B(new_n1090), .C(new_n1095), .Y(new_n1096));
  NOR2xp33_ASAP7_75t_L      g00840(.A(new_n427), .B(new_n710), .Y(new_n1097));
  AOI221xp5_ASAP7_75t_L     g00841(.A1(\b[5] ), .A2(new_n635), .B1(\b[4] ), .B2(new_n713), .C(new_n1097), .Y(new_n1098));
  O2A1O1Ixp33_ASAP7_75t_L   g00842(.A1(new_n641), .A2(new_n434), .B(new_n1098), .C(new_n637), .Y(new_n1099));
  OAI31xp33_ASAP7_75t_L     g00843(.A1(new_n433), .A2(new_n431), .A3(new_n641), .B(new_n1098), .Y(new_n1100));
  NAND2xp33_ASAP7_75t_L     g00844(.A(new_n637), .B(new_n1100), .Y(new_n1101));
  OA21x2_ASAP7_75t_L        g00845(.A1(new_n637), .A2(new_n1099), .B(new_n1101), .Y(new_n1102));
  NAND3xp33_ASAP7_75t_L     g00846(.A(new_n1096), .B(new_n1089), .C(new_n1102), .Y(new_n1103));
  AO21x2_ASAP7_75t_L        g00847(.A1(new_n1089), .A2(new_n1096), .B(new_n1102), .Y(new_n1104));
  AOI21xp33_ASAP7_75t_L     g00848(.A1(new_n1104), .A2(new_n1103), .B(new_n1018), .Y(new_n1105));
  AND3x1_ASAP7_75t_L        g00849(.A(new_n1096), .B(new_n1102), .C(new_n1089), .Y(new_n1106));
  AOI21xp33_ASAP7_75t_L     g00850(.A1(new_n1096), .A2(new_n1089), .B(new_n1102), .Y(new_n1107));
  NOR4xp25_ASAP7_75t_L      g00851(.A(new_n1106), .B(new_n998), .C(new_n1107), .D(new_n1063), .Y(new_n1108));
  OAI21xp33_ASAP7_75t_L     g00852(.A1(new_n1105), .A2(new_n1108), .B(new_n1072), .Y(new_n1109));
  A2O1A1Ixp33_ASAP7_75t_L   g00853(.A1(new_n602), .A2(new_n483), .B(new_n1070), .C(\a[8] ), .Y(new_n1110));
  NAND2xp33_ASAP7_75t_L     g00854(.A(\a[8] ), .B(new_n1110), .Y(new_n1111));
  OAI22xp33_ASAP7_75t_L     g00855(.A1(new_n1106), .A2(new_n1107), .B1(new_n998), .B2(new_n1063), .Y(new_n1112));
  NAND3xp33_ASAP7_75t_L     g00856(.A(new_n1018), .B(new_n1104), .C(new_n1103), .Y(new_n1113));
  NAND4xp25_ASAP7_75t_L     g00857(.A(new_n1112), .B(new_n1113), .C(new_n1111), .D(new_n1071), .Y(new_n1114));
  NAND2xp33_ASAP7_75t_L     g00858(.A(new_n1114), .B(new_n1109), .Y(new_n1115));
  A2O1A1Ixp33_ASAP7_75t_L   g00859(.A1(new_n1016), .A2(new_n1023), .B(new_n1064), .C(new_n1115), .Y(new_n1116));
  INVx1_ASAP7_75t_L         g00860(.A(new_n918), .Y(new_n1117));
  A2O1A1O1Ixp25_ASAP7_75t_L g00861(.A1(new_n914), .A2(new_n916), .B(new_n1117), .C(new_n1016), .D(new_n1064), .Y(new_n1118));
  NAND3xp33_ASAP7_75t_L     g00862(.A(new_n1118), .B(new_n1109), .C(new_n1114), .Y(new_n1119));
  AO21x2_ASAP7_75t_L        g00863(.A1(new_n1116), .A2(new_n1119), .B(new_n1062), .Y(new_n1120));
  A2O1A1Ixp33_ASAP7_75t_L   g00864(.A1(new_n927), .A2(new_n824), .B(new_n821), .C(new_n925), .Y(new_n1121));
  OR3x1_ASAP7_75t_L         g00865(.A(new_n1025), .B(new_n1022), .C(new_n979), .Y(new_n1122));
  A2O1A1Ixp33_ASAP7_75t_L   g00866(.A1(new_n1121), .A2(new_n930), .B(new_n1026), .C(new_n1122), .Y(new_n1123));
  INVx1_ASAP7_75t_L         g00867(.A(new_n1062), .Y(new_n1124));
  NAND3xp33_ASAP7_75t_L     g00868(.A(new_n1124), .B(new_n1116), .C(new_n1119), .Y(new_n1125));
  NAND3xp33_ASAP7_75t_L     g00869(.A(new_n1119), .B(new_n1116), .C(new_n1062), .Y(new_n1126));
  INVx1_ASAP7_75t_L         g00870(.A(new_n1126), .Y(new_n1127));
  A2O1A1Ixp33_ASAP7_75t_L   g00871(.A1(new_n1124), .A2(new_n1125), .B(new_n1127), .C(new_n1123), .Y(new_n1128));
  INVx1_ASAP7_75t_L         g00872(.A(new_n1128), .Y(new_n1129));
  NOR2xp33_ASAP7_75t_L      g00873(.A(new_n1127), .B(new_n1123), .Y(new_n1130));
  A2O1A1Ixp33_ASAP7_75t_L   g00874(.A1(new_n1130), .A2(new_n1120), .B(new_n1129), .C(new_n1056), .Y(new_n1131));
  INVx1_ASAP7_75t_L         g00875(.A(new_n1120), .Y(new_n1132));
  INVx1_ASAP7_75t_L         g00876(.A(new_n1130), .Y(new_n1133));
  OAI211xp5_ASAP7_75t_L     g00877(.A1(new_n1132), .A2(new_n1133), .B(new_n1128), .C(new_n1055), .Y(new_n1134));
  NAND2xp33_ASAP7_75t_L     g00878(.A(new_n1131), .B(new_n1134), .Y(new_n1135));
  NAND2xp33_ASAP7_75t_L     g00879(.A(new_n975), .B(new_n1042), .Y(new_n1136));
  OAI211xp5_ASAP7_75t_L     g00880(.A1(new_n1039), .A2(new_n1035), .B(new_n1134), .C(new_n1136), .Y(new_n1137));
  A2O1A1O1Ixp25_ASAP7_75t_L g00881(.A1(new_n1130), .A2(new_n1120), .B(new_n1129), .C(new_n1056), .D(new_n1137), .Y(new_n1138));
  A2O1A1O1Ixp25_ASAP7_75t_L g00882(.A1(new_n1042), .A2(new_n975), .B(new_n1036), .C(new_n1135), .D(new_n1138), .Y(\f[15] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00883(.A1(new_n1124), .A2(new_n1125), .B(new_n1133), .C(new_n1128), .Y(new_n1140));
  NOR2xp33_ASAP7_75t_L      g00884(.A(new_n1055), .B(new_n1140), .Y(new_n1141));
  A2O1A1O1Ixp25_ASAP7_75t_L g00885(.A1(new_n1042), .A2(new_n975), .B(new_n1036), .C(new_n1135), .D(new_n1141), .Y(new_n1142));
  NOR2xp33_ASAP7_75t_L      g00886(.A(new_n960), .B(new_n287), .Y(new_n1143));
  AOI221xp5_ASAP7_75t_L     g00887(.A1(\b[15] ), .A2(new_n264), .B1(\b[16] ), .B2(new_n283), .C(new_n1143), .Y(new_n1144));
  INVx1_ASAP7_75t_L         g00888(.A(new_n1144), .Y(new_n1145));
  INVx1_ASAP7_75t_L         g00889(.A(new_n939), .Y(new_n1146));
  O2A1O1Ixp33_ASAP7_75t_L   g00890(.A1(new_n937), .A2(new_n1146), .B(new_n965), .C(new_n964), .Y(new_n1147));
  INVx1_ASAP7_75t_L         g00891(.A(new_n1047), .Y(new_n1148));
  NOR2xp33_ASAP7_75t_L      g00892(.A(\b[15] ), .B(\b[16] ), .Y(new_n1149));
  INVx1_ASAP7_75t_L         g00893(.A(\b[16] ), .Y(new_n1150));
  NOR2xp33_ASAP7_75t_L      g00894(.A(new_n1043), .B(new_n1150), .Y(new_n1151));
  NOR2xp33_ASAP7_75t_L      g00895(.A(new_n1149), .B(new_n1151), .Y(new_n1152));
  INVx1_ASAP7_75t_L         g00896(.A(new_n1152), .Y(new_n1153));
  O2A1O1Ixp33_ASAP7_75t_L   g00897(.A1(new_n1046), .A2(new_n1147), .B(new_n1148), .C(new_n1153), .Y(new_n1154));
  AND3x1_ASAP7_75t_L        g00898(.A(new_n1049), .B(new_n1153), .C(new_n1148), .Y(new_n1155));
  NOR2xp33_ASAP7_75t_L      g00899(.A(new_n1154), .B(new_n1155), .Y(new_n1156));
  A2O1A1Ixp33_ASAP7_75t_L   g00900(.A1(new_n1156), .A2(new_n273), .B(new_n1145), .C(\a[2] ), .Y(new_n1157));
  INVx1_ASAP7_75t_L         g00901(.A(new_n1154), .Y(new_n1158));
  O2A1O1Ixp33_ASAP7_75t_L   g00902(.A1(new_n964), .A2(new_n967), .B(new_n1048), .C(new_n1047), .Y(new_n1159));
  NAND2xp33_ASAP7_75t_L     g00903(.A(new_n1153), .B(new_n1159), .Y(new_n1160));
  NAND2xp33_ASAP7_75t_L     g00904(.A(new_n1160), .B(new_n1158), .Y(new_n1161));
  O2A1O1Ixp33_ASAP7_75t_L   g00905(.A1(new_n279), .A2(new_n1161), .B(new_n1144), .C(\a[2] ), .Y(new_n1162));
  AOI21xp33_ASAP7_75t_L     g00906(.A1(new_n1157), .A2(\a[2] ), .B(new_n1162), .Y(new_n1163));
  INVx1_ASAP7_75t_L         g00907(.A(new_n1125), .Y(new_n1164));
  NAND2xp33_ASAP7_75t_L     g00908(.A(new_n1126), .B(new_n1120), .Y(new_n1165));
  NOR2xp33_ASAP7_75t_L      g00909(.A(new_n940), .B(new_n1146), .Y(new_n1166));
  NAND2xp33_ASAP7_75t_L     g00910(.A(\b[13] ), .B(new_n361), .Y(new_n1167));
  OAI221xp5_ASAP7_75t_L     g00911(.A1(new_n350), .A2(new_n833), .B1(new_n748), .B2(new_n375), .C(new_n1167), .Y(new_n1168));
  A2O1A1Ixp33_ASAP7_75t_L   g00912(.A1(new_n1166), .A2(new_n359), .B(new_n1168), .C(\a[5] ), .Y(new_n1169));
  AOI211xp5_ASAP7_75t_L     g00913(.A1(new_n1166), .A2(new_n359), .B(new_n1168), .C(new_n346), .Y(new_n1170));
  A2O1A1O1Ixp25_ASAP7_75t_L g00914(.A1(new_n1166), .A2(new_n359), .B(new_n1168), .C(new_n1169), .D(new_n1170), .Y(new_n1171));
  INVx1_ASAP7_75t_L         g00915(.A(new_n1171), .Y(new_n1172));
  NAND3xp33_ASAP7_75t_L     g00916(.A(new_n1112), .B(new_n1113), .C(new_n1072), .Y(new_n1173));
  A2O1A1Ixp33_ASAP7_75t_L   g00917(.A1(new_n1109), .A2(new_n1114), .B(new_n1118), .C(new_n1173), .Y(new_n1174));
  NAND2xp33_ASAP7_75t_L     g00918(.A(new_n689), .B(new_n687), .Y(new_n1175));
  NOR2xp33_ASAP7_75t_L      g00919(.A(new_n590), .B(new_n513), .Y(new_n1176));
  AOI221xp5_ASAP7_75t_L     g00920(.A1(\b[8] ), .A2(new_n560), .B1(\b[10] ), .B2(new_n475), .C(new_n1176), .Y(new_n1177));
  O2A1O1Ixp33_ASAP7_75t_L   g00921(.A1(new_n477), .A2(new_n1175), .B(new_n1177), .C(new_n466), .Y(new_n1178));
  INVx1_ASAP7_75t_L         g00922(.A(new_n1177), .Y(new_n1179));
  A2O1A1Ixp33_ASAP7_75t_L   g00923(.A1(new_n690), .A2(new_n483), .B(new_n1179), .C(new_n466), .Y(new_n1180));
  OAI21xp33_ASAP7_75t_L     g00924(.A1(new_n466), .A2(new_n1178), .B(new_n1180), .Y(new_n1181));
  NOR2xp33_ASAP7_75t_L      g00925(.A(new_n637), .B(new_n1100), .Y(new_n1182));
  O2A1O1Ixp33_ASAP7_75t_L   g00926(.A1(new_n641), .A2(new_n434), .B(new_n1098), .C(\a[11] ), .Y(new_n1183));
  OAI211xp5_ASAP7_75t_L     g00927(.A1(new_n1182), .A2(new_n1183), .B(new_n1089), .C(new_n1096), .Y(new_n1184));
  A2O1A1Ixp33_ASAP7_75t_L   g00928(.A1(new_n1103), .A2(new_n1102), .B(new_n1018), .C(new_n1184), .Y(new_n1185));
  NOR2xp33_ASAP7_75t_L      g00929(.A(new_n448), .B(new_n710), .Y(new_n1186));
  AOI221xp5_ASAP7_75t_L     g00930(.A1(\b[6] ), .A2(new_n635), .B1(\b[5] ), .B2(new_n713), .C(new_n1186), .Y(new_n1187));
  INVx1_ASAP7_75t_L         g00931(.A(new_n456), .Y(new_n1188));
  NAND2xp33_ASAP7_75t_L     g00932(.A(new_n718), .B(new_n1188), .Y(new_n1189));
  O2A1O1Ixp33_ASAP7_75t_L   g00933(.A1(new_n641), .A2(new_n456), .B(new_n1187), .C(new_n637), .Y(new_n1190));
  OAI211xp5_ASAP7_75t_L     g00934(.A1(new_n641), .A2(new_n456), .B(\a[11] ), .C(new_n1187), .Y(new_n1191));
  A2O1A1Ixp33_ASAP7_75t_L   g00935(.A1(new_n1189), .A2(new_n1187), .B(new_n1190), .C(new_n1191), .Y(new_n1192));
  MAJIxp5_ASAP7_75t_L       g00936(.A(new_n1095), .B(new_n1003), .C(new_n1078), .Y(new_n1193));
  NAND2xp33_ASAP7_75t_L     g00937(.A(\b[3] ), .B(new_n885), .Y(new_n1194));
  OAI221xp5_ASAP7_75t_L     g00938(.A1(new_n869), .A2(new_n332), .B1(new_n289), .B2(new_n980), .C(new_n1194), .Y(new_n1195));
  A2O1A1Ixp33_ASAP7_75t_L   g00939(.A1(new_n342), .A2(new_n873), .B(new_n1195), .C(\a[14] ), .Y(new_n1196));
  AOI211xp5_ASAP7_75t_L     g00940(.A1(new_n342), .A2(new_n873), .B(new_n867), .C(new_n1195), .Y(new_n1197));
  A2O1A1O1Ixp25_ASAP7_75t_L g00941(.A1(new_n873), .A2(new_n342), .B(new_n1195), .C(new_n1196), .D(new_n1197), .Y(new_n1198));
  NAND2xp33_ASAP7_75t_L     g00942(.A(new_n1075), .B(new_n1074), .Y(new_n1199));
  INVx1_ASAP7_75t_L         g00943(.A(\a[16] ), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g00944(.A(\a[15] ), .B(new_n1200), .Y(new_n1201));
  NOR2xp33_ASAP7_75t_L      g00945(.A(\a[16] ), .B(new_n1073), .Y(new_n1202));
  NOR2xp33_ASAP7_75t_L      g00946(.A(new_n1201), .B(new_n1202), .Y(new_n1203));
  NOR2xp33_ASAP7_75t_L      g00947(.A(new_n1199), .B(new_n1203), .Y(new_n1204));
  NAND2xp33_ASAP7_75t_L     g00948(.A(\a[17] ), .B(new_n1200), .Y(new_n1205));
  INVx1_ASAP7_75t_L         g00949(.A(\a[17] ), .Y(new_n1206));
  NAND2xp33_ASAP7_75t_L     g00950(.A(\a[16] ), .B(new_n1206), .Y(new_n1207));
  NAND2xp33_ASAP7_75t_L     g00951(.A(new_n1207), .B(new_n1205), .Y(new_n1208));
  NOR2xp33_ASAP7_75t_L      g00952(.A(new_n1208), .B(new_n1076), .Y(new_n1209));
  NAND2xp33_ASAP7_75t_L     g00953(.A(new_n1208), .B(new_n1199), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g00954(.A(new_n274), .B(new_n1210), .Y(new_n1211));
  AOI221xp5_ASAP7_75t_L     g00955(.A1(\b[1] ), .A2(new_n1209), .B1(new_n1204), .B2(\b[0] ), .C(new_n1211), .Y(new_n1212));
  NAND3xp33_ASAP7_75t_L     g00956(.A(new_n1212), .B(new_n1078), .C(\a[17] ), .Y(new_n1213));
  INVx1_ASAP7_75t_L         g00957(.A(new_n1213), .Y(new_n1214));
  AOI22xp33_ASAP7_75t_L     g00958(.A1(new_n1204), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n1209), .Y(new_n1215));
  AOI21xp33_ASAP7_75t_L     g00959(.A1(new_n1207), .A2(new_n1205), .B(new_n1076), .Y(new_n1216));
  NAND2xp33_ASAP7_75t_L     g00960(.A(new_n275), .B(new_n1216), .Y(new_n1217));
  NAND2xp33_ASAP7_75t_L     g00961(.A(new_n1217), .B(new_n1215), .Y(new_n1218));
  NAND2xp33_ASAP7_75t_L     g00962(.A(\a[17] ), .B(new_n1218), .Y(new_n1219));
  O2A1O1Ixp33_ASAP7_75t_L   g00963(.A1(new_n1210), .A2(new_n274), .B(new_n1215), .C(\a[17] ), .Y(new_n1220));
  O2A1O1Ixp33_ASAP7_75t_L   g00964(.A1(new_n1078), .A2(new_n1219), .B(\a[17] ), .C(new_n1220), .Y(new_n1221));
  OAI21xp33_ASAP7_75t_L     g00965(.A1(new_n1214), .A2(new_n1221), .B(new_n1198), .Y(new_n1222));
  AOI21xp33_ASAP7_75t_L     g00966(.A1(new_n342), .A2(new_n873), .B(new_n1195), .Y(new_n1223));
  NOR2xp33_ASAP7_75t_L      g00967(.A(\a[14] ), .B(new_n1223), .Y(new_n1224));
  O2A1O1Ixp33_ASAP7_75t_L   g00968(.A1(new_n1210), .A2(new_n274), .B(new_n1215), .C(new_n1206), .Y(new_n1225));
  NAND2xp33_ASAP7_75t_L     g00969(.A(new_n1206), .B(new_n1218), .Y(new_n1226));
  A2O1A1Ixp33_ASAP7_75t_L   g00970(.A1(new_n1077), .A2(new_n1225), .B(new_n1206), .C(new_n1226), .Y(new_n1227));
  OAI211xp5_ASAP7_75t_L     g00971(.A1(new_n1197), .A2(new_n1224), .B(new_n1227), .C(new_n1213), .Y(new_n1228));
  NAND3xp33_ASAP7_75t_L     g00972(.A(new_n1193), .B(new_n1222), .C(new_n1228), .Y(new_n1229));
  MAJIxp5_ASAP7_75t_L       g00973(.A(new_n1088), .B(new_n1077), .C(new_n991), .Y(new_n1230));
  AOI211xp5_ASAP7_75t_L     g00974(.A1(new_n1227), .A2(new_n1213), .B(new_n1197), .C(new_n1224), .Y(new_n1231));
  NOR3xp33_ASAP7_75t_L      g00975(.A(new_n1221), .B(new_n1198), .C(new_n1214), .Y(new_n1232));
  OAI21xp33_ASAP7_75t_L     g00976(.A1(new_n1231), .A2(new_n1232), .B(new_n1230), .Y(new_n1233));
  AO21x2_ASAP7_75t_L        g00977(.A1(new_n1229), .A2(new_n1233), .B(new_n1192), .Y(new_n1234));
  NAND3xp33_ASAP7_75t_L     g00978(.A(new_n1233), .B(new_n1229), .C(new_n1192), .Y(new_n1235));
  NAND3xp33_ASAP7_75t_L     g00979(.A(new_n1185), .B(new_n1234), .C(new_n1235), .Y(new_n1236));
  AO21x2_ASAP7_75t_L        g00980(.A1(new_n1235), .A2(new_n1234), .B(new_n1185), .Y(new_n1237));
  AO21x2_ASAP7_75t_L        g00981(.A1(new_n1236), .A2(new_n1237), .B(new_n1181), .Y(new_n1238));
  NAND3xp33_ASAP7_75t_L     g00982(.A(new_n1237), .B(new_n1236), .C(new_n1181), .Y(new_n1239));
  NAND3xp33_ASAP7_75t_L     g00983(.A(new_n1174), .B(new_n1238), .C(new_n1239), .Y(new_n1240));
  INVx1_ASAP7_75t_L         g00984(.A(new_n1173), .Y(new_n1241));
  A2O1A1O1Ixp25_ASAP7_75t_L g00985(.A1(new_n1016), .A2(new_n1023), .B(new_n1064), .C(new_n1115), .D(new_n1241), .Y(new_n1242));
  NAND2xp33_ASAP7_75t_L     g00986(.A(new_n1239), .B(new_n1238), .Y(new_n1243));
  NAND2xp33_ASAP7_75t_L     g00987(.A(new_n1242), .B(new_n1243), .Y(new_n1244));
  AOI21xp33_ASAP7_75t_L     g00988(.A1(new_n1244), .A2(new_n1240), .B(new_n1172), .Y(new_n1245));
  NOR2xp33_ASAP7_75t_L      g00989(.A(new_n1242), .B(new_n1243), .Y(new_n1246));
  AOI21xp33_ASAP7_75t_L     g00990(.A1(new_n1239), .A2(new_n1238), .B(new_n1174), .Y(new_n1247));
  NOR3xp33_ASAP7_75t_L      g00991(.A(new_n1246), .B(new_n1247), .C(new_n1171), .Y(new_n1248));
  NOR2xp33_ASAP7_75t_L      g00992(.A(new_n1245), .B(new_n1248), .Y(new_n1249));
  A2O1A1Ixp33_ASAP7_75t_L   g00993(.A1(new_n1165), .A2(new_n1123), .B(new_n1164), .C(new_n1249), .Y(new_n1250));
  O2A1O1Ixp33_ASAP7_75t_L   g00994(.A1(new_n1127), .A2(new_n1124), .B(new_n1123), .C(new_n1164), .Y(new_n1251));
  OAI21xp33_ASAP7_75t_L     g00995(.A1(new_n1247), .A2(new_n1246), .B(new_n1171), .Y(new_n1252));
  NAND3xp33_ASAP7_75t_L     g00996(.A(new_n1172), .B(new_n1244), .C(new_n1240), .Y(new_n1253));
  NAND2xp33_ASAP7_75t_L     g00997(.A(new_n1252), .B(new_n1253), .Y(new_n1254));
  NAND2xp33_ASAP7_75t_L     g00998(.A(new_n1254), .B(new_n1251), .Y(new_n1255));
  NAND3xp33_ASAP7_75t_L     g00999(.A(new_n1250), .B(new_n1255), .C(new_n1163), .Y(new_n1256));
  INVx1_ASAP7_75t_L         g01000(.A(new_n1163), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g01001(.A(new_n1254), .B(new_n1251), .Y(new_n1258));
  AOI221xp5_ASAP7_75t_L     g01002(.A1(new_n1165), .A2(new_n1123), .B1(new_n1253), .B2(new_n1252), .C(new_n1164), .Y(new_n1259));
  OAI21xp33_ASAP7_75t_L     g01003(.A1(new_n1259), .A2(new_n1258), .B(new_n1257), .Y(new_n1260));
  NAND2xp33_ASAP7_75t_L     g01004(.A(new_n1260), .B(new_n1256), .Y(new_n1261));
  XNOR2x2_ASAP7_75t_L       g01005(.A(new_n1261), .B(new_n1142), .Y(\f[16] ));
  NAND2xp33_ASAP7_75t_L     g01006(.A(new_n1255), .B(new_n1250), .Y(new_n1263));
  OAI21xp33_ASAP7_75t_L     g01007(.A1(new_n1035), .A2(new_n1039), .B(new_n1136), .Y(new_n1264));
  A2O1A1Ixp33_ASAP7_75t_L   g01008(.A1(new_n1135), .A2(new_n1264), .B(new_n1141), .C(new_n1261), .Y(new_n1265));
  A2O1A1O1Ixp25_ASAP7_75t_L g01009(.A1(new_n1123), .A2(new_n1165), .B(new_n1164), .C(new_n1252), .D(new_n1248), .Y(new_n1266));
  INVx1_ASAP7_75t_L         g01010(.A(new_n967), .Y(new_n1267));
  NAND2xp33_ASAP7_75t_L     g01011(.A(new_n969), .B(new_n1267), .Y(new_n1268));
  NOR2xp33_ASAP7_75t_L      g01012(.A(new_n833), .B(new_n375), .Y(new_n1269));
  AOI221xp5_ASAP7_75t_L     g01013(.A1(\b[14] ), .A2(new_n361), .B1(new_n349), .B2(\b[13] ), .C(new_n1269), .Y(new_n1270));
  O2A1O1Ixp33_ASAP7_75t_L   g01014(.A1(new_n356), .A2(new_n1268), .B(new_n1270), .C(new_n346), .Y(new_n1271));
  INVx1_ASAP7_75t_L         g01015(.A(new_n1271), .Y(new_n1272));
  O2A1O1Ixp33_ASAP7_75t_L   g01016(.A1(new_n356), .A2(new_n1268), .B(new_n1270), .C(\a[5] ), .Y(new_n1273));
  AOI21xp33_ASAP7_75t_L     g01017(.A1(new_n1272), .A2(\a[5] ), .B(new_n1273), .Y(new_n1274));
  NOR2xp33_ASAP7_75t_L      g01018(.A(new_n680), .B(new_n513), .Y(new_n1275));
  AOI221xp5_ASAP7_75t_L     g01019(.A1(\b[9] ), .A2(new_n560), .B1(\b[11] ), .B2(new_n475), .C(new_n1275), .Y(new_n1276));
  O2A1O1Ixp33_ASAP7_75t_L   g01020(.A1(new_n477), .A2(new_n754), .B(new_n1276), .C(new_n466), .Y(new_n1277));
  INVx1_ASAP7_75t_L         g01021(.A(new_n1277), .Y(new_n1278));
  O2A1O1Ixp33_ASAP7_75t_L   g01022(.A1(new_n477), .A2(new_n754), .B(new_n1276), .C(\a[8] ), .Y(new_n1279));
  AOI21xp33_ASAP7_75t_L     g01023(.A1(new_n1278), .A2(\a[8] ), .B(new_n1279), .Y(new_n1280));
  INVx1_ASAP7_75t_L         g01024(.A(new_n1235), .Y(new_n1281));
  AOI21xp33_ASAP7_75t_L     g01025(.A1(new_n1185), .A2(new_n1234), .B(new_n1281), .Y(new_n1282));
  OAI21xp33_ASAP7_75t_L     g01026(.A1(new_n1230), .A2(new_n1231), .B(new_n1228), .Y(new_n1283));
  NAND3xp33_ASAP7_75t_L     g01027(.A(new_n1199), .B(new_n1205), .C(new_n1207), .Y(new_n1284));
  NAND3xp33_ASAP7_75t_L     g01028(.A(new_n1076), .B(new_n1203), .C(new_n1208), .Y(new_n1285));
  NAND2xp33_ASAP7_75t_L     g01029(.A(\b[1] ), .B(new_n1204), .Y(new_n1286));
  OAI221xp5_ASAP7_75t_L     g01030(.A1(new_n1284), .A2(new_n289), .B1(new_n284), .B2(new_n1285), .C(new_n1286), .Y(new_n1287));
  A2O1A1Ixp33_ASAP7_75t_L   g01031(.A1(new_n294), .A2(new_n1216), .B(new_n1287), .C(\a[17] ), .Y(new_n1288));
  NOR2xp33_ASAP7_75t_L      g01032(.A(new_n289), .B(new_n1284), .Y(new_n1289));
  AND3x1_ASAP7_75t_L        g01033(.A(new_n1076), .B(new_n1208), .C(new_n1203), .Y(new_n1290));
  AOI221xp5_ASAP7_75t_L     g01034(.A1(new_n1204), .A2(\b[1] ), .B1(new_n1290), .B2(\b[0] ), .C(new_n1289), .Y(new_n1291));
  O2A1O1Ixp33_ASAP7_75t_L   g01035(.A1(new_n509), .A2(new_n1210), .B(new_n1291), .C(\a[17] ), .Y(new_n1292));
  A2O1A1O1Ixp25_ASAP7_75t_L g01036(.A1(new_n1212), .A2(new_n1078), .B(new_n1288), .C(\a[17] ), .D(new_n1292), .Y(new_n1293));
  NOR2xp33_ASAP7_75t_L      g01037(.A(new_n1210), .B(new_n509), .Y(new_n1294));
  NOR5xp2_ASAP7_75t_L       g01038(.A(new_n1218), .B(new_n1287), .C(new_n1294), .D(new_n1077), .E(new_n1206), .Y(new_n1295));
  NAND2xp33_ASAP7_75t_L     g01039(.A(\b[4] ), .B(new_n885), .Y(new_n1296));
  OAI221xp5_ASAP7_75t_L     g01040(.A1(new_n869), .A2(new_n384), .B1(new_n301), .B2(new_n980), .C(new_n1296), .Y(new_n1297));
  A2O1A1Ixp33_ASAP7_75t_L   g01041(.A1(new_n394), .A2(new_n873), .B(new_n1297), .C(\a[14] ), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g01042(.A(new_n384), .B(new_n869), .Y(new_n1299));
  AOI221xp5_ASAP7_75t_L     g01043(.A1(\b[3] ), .A2(new_n985), .B1(\b[4] ), .B2(new_n885), .C(new_n1299), .Y(new_n1300));
  O2A1O1Ixp33_ASAP7_75t_L   g01044(.A1(new_n872), .A2(new_n728), .B(new_n1300), .C(\a[14] ), .Y(new_n1301));
  AOI21xp33_ASAP7_75t_L     g01045(.A1(new_n1298), .A2(\a[14] ), .B(new_n1301), .Y(new_n1302));
  NOR3xp33_ASAP7_75t_L      g01046(.A(new_n1302), .B(new_n1293), .C(new_n1295), .Y(new_n1303));
  INVx1_ASAP7_75t_L         g01047(.A(new_n1294), .Y(new_n1304));
  NAND3xp33_ASAP7_75t_L     g01048(.A(new_n1291), .B(\a[17] ), .C(new_n1304), .Y(new_n1305));
  A2O1A1Ixp33_ASAP7_75t_L   g01049(.A1(new_n294), .A2(new_n1216), .B(new_n1287), .C(new_n1206), .Y(new_n1306));
  NAND3xp33_ASAP7_75t_L     g01050(.A(new_n1305), .B(new_n1306), .C(new_n1213), .Y(new_n1307));
  NAND5xp2_ASAP7_75t_L      g01051(.A(\a[17] ), .B(new_n1291), .C(new_n1212), .D(new_n1304), .E(new_n1078), .Y(new_n1308));
  AOI221xp5_ASAP7_75t_L     g01052(.A1(new_n1298), .A2(\a[14] ), .B1(new_n1308), .B2(new_n1307), .C(new_n1301), .Y(new_n1309));
  OAI21xp33_ASAP7_75t_L     g01053(.A1(new_n1303), .A2(new_n1309), .B(new_n1283), .Y(new_n1310));
  INVx1_ASAP7_75t_L         g01054(.A(new_n1303), .Y(new_n1311));
  OAI21xp33_ASAP7_75t_L     g01055(.A1(new_n1295), .A2(new_n1293), .B(new_n1302), .Y(new_n1312));
  NAND4xp25_ASAP7_75t_L     g01056(.A(new_n1229), .B(new_n1311), .C(new_n1312), .D(new_n1228), .Y(new_n1313));
  NOR2xp33_ASAP7_75t_L      g01057(.A(new_n534), .B(new_n710), .Y(new_n1314));
  AOI221xp5_ASAP7_75t_L     g01058(.A1(\b[7] ), .A2(new_n635), .B1(\b[6] ), .B2(new_n713), .C(new_n1314), .Y(new_n1315));
  OAI21xp33_ASAP7_75t_L     g01059(.A1(new_n641), .A2(new_n540), .B(new_n1315), .Y(new_n1316));
  NOR2xp33_ASAP7_75t_L      g01060(.A(new_n637), .B(new_n1316), .Y(new_n1317));
  O2A1O1Ixp33_ASAP7_75t_L   g01061(.A1(new_n641), .A2(new_n540), .B(new_n1315), .C(\a[11] ), .Y(new_n1318));
  NOR2xp33_ASAP7_75t_L      g01062(.A(new_n1318), .B(new_n1317), .Y(new_n1319));
  AND3x1_ASAP7_75t_L        g01063(.A(new_n1313), .B(new_n1319), .C(new_n1310), .Y(new_n1320));
  AOI21xp33_ASAP7_75t_L     g01064(.A1(new_n1313), .A2(new_n1310), .B(new_n1319), .Y(new_n1321));
  NOR3xp33_ASAP7_75t_L      g01065(.A(new_n1282), .B(new_n1320), .C(new_n1321), .Y(new_n1322));
  NAND3xp33_ASAP7_75t_L     g01066(.A(new_n1313), .B(new_n1310), .C(new_n1319), .Y(new_n1323));
  AO21x2_ASAP7_75t_L        g01067(.A1(new_n1310), .A2(new_n1313), .B(new_n1319), .Y(new_n1324));
  AOI221xp5_ASAP7_75t_L     g01068(.A1(new_n1185), .A2(new_n1234), .B1(new_n1323), .B2(new_n1324), .C(new_n1281), .Y(new_n1325));
  OAI21xp33_ASAP7_75t_L     g01069(.A1(new_n1325), .A2(new_n1322), .B(new_n1280), .Y(new_n1326));
  AO21x2_ASAP7_75t_L        g01070(.A1(\a[8] ), .A2(new_n1278), .B(new_n1279), .Y(new_n1327));
  AOI21xp33_ASAP7_75t_L     g01071(.A1(new_n1233), .A2(new_n1229), .B(new_n1192), .Y(new_n1328));
  A2O1A1Ixp33_ASAP7_75t_L   g01072(.A1(new_n1112), .A2(new_n1184), .B(new_n1328), .C(new_n1235), .Y(new_n1329));
  NAND3xp33_ASAP7_75t_L     g01073(.A(new_n1329), .B(new_n1323), .C(new_n1324), .Y(new_n1330));
  OAI21xp33_ASAP7_75t_L     g01074(.A1(new_n1320), .A2(new_n1321), .B(new_n1282), .Y(new_n1331));
  NAND3xp33_ASAP7_75t_L     g01075(.A(new_n1330), .B(new_n1327), .C(new_n1331), .Y(new_n1332));
  NAND2xp33_ASAP7_75t_L     g01076(.A(new_n1326), .B(new_n1332), .Y(new_n1333));
  O2A1O1Ixp33_ASAP7_75t_L   g01077(.A1(new_n1242), .A2(new_n1243), .B(new_n1239), .C(new_n1333), .Y(new_n1334));
  AOI21xp33_ASAP7_75t_L     g01078(.A1(new_n1237), .A2(new_n1236), .B(new_n1181), .Y(new_n1335));
  A2O1A1Ixp33_ASAP7_75t_L   g01079(.A1(new_n1116), .A2(new_n1173), .B(new_n1335), .C(new_n1239), .Y(new_n1336));
  AOI21xp33_ASAP7_75t_L     g01080(.A1(new_n1330), .A2(new_n1331), .B(new_n1327), .Y(new_n1337));
  NOR3xp33_ASAP7_75t_L      g01081(.A(new_n1322), .B(new_n1325), .C(new_n1280), .Y(new_n1338));
  NOR2xp33_ASAP7_75t_L      g01082(.A(new_n1338), .B(new_n1337), .Y(new_n1339));
  NOR2xp33_ASAP7_75t_L      g01083(.A(new_n1339), .B(new_n1336), .Y(new_n1340));
  OA21x2_ASAP7_75t_L        g01084(.A1(new_n1340), .A2(new_n1334), .B(new_n1274), .Y(new_n1341));
  NOR3xp33_ASAP7_75t_L      g01085(.A(new_n1274), .B(new_n1334), .C(new_n1340), .Y(new_n1342));
  NOR3xp33_ASAP7_75t_L      g01086(.A(new_n1266), .B(new_n1341), .C(new_n1342), .Y(new_n1343));
  OA21x2_ASAP7_75t_L        g01087(.A1(new_n1341), .A2(new_n1342), .B(new_n1266), .Y(new_n1344));
  NOR2xp33_ASAP7_75t_L      g01088(.A(new_n1043), .B(new_n287), .Y(new_n1345));
  AOI221xp5_ASAP7_75t_L     g01089(.A1(\b[16] ), .A2(new_n264), .B1(\b[17] ), .B2(new_n283), .C(new_n1345), .Y(new_n1346));
  INVx1_ASAP7_75t_L         g01090(.A(new_n1151), .Y(new_n1347));
  NOR2xp33_ASAP7_75t_L      g01091(.A(\b[16] ), .B(\b[17] ), .Y(new_n1348));
  INVx1_ASAP7_75t_L         g01092(.A(\b[17] ), .Y(new_n1349));
  NOR2xp33_ASAP7_75t_L      g01093(.A(new_n1150), .B(new_n1349), .Y(new_n1350));
  NOR2xp33_ASAP7_75t_L      g01094(.A(new_n1348), .B(new_n1350), .Y(new_n1351));
  INVx1_ASAP7_75t_L         g01095(.A(new_n1351), .Y(new_n1352));
  O2A1O1Ixp33_ASAP7_75t_L   g01096(.A1(new_n1153), .A2(new_n1159), .B(new_n1347), .C(new_n1352), .Y(new_n1353));
  INVx1_ASAP7_75t_L         g01097(.A(new_n1353), .Y(new_n1354));
  OAI211xp5_ASAP7_75t_L     g01098(.A1(new_n1153), .A2(new_n1159), .B(new_n1347), .C(new_n1352), .Y(new_n1355));
  NAND2xp33_ASAP7_75t_L     g01099(.A(new_n1355), .B(new_n1354), .Y(new_n1356));
  O2A1O1Ixp33_ASAP7_75t_L   g01100(.A1(new_n279), .A2(new_n1356), .B(new_n1346), .C(new_n257), .Y(new_n1357));
  INVx1_ASAP7_75t_L         g01101(.A(new_n1357), .Y(new_n1358));
  O2A1O1Ixp33_ASAP7_75t_L   g01102(.A1(new_n279), .A2(new_n1356), .B(new_n1346), .C(\a[2] ), .Y(new_n1359));
  AO21x2_ASAP7_75t_L        g01103(.A1(\a[2] ), .A2(new_n1358), .B(new_n1359), .Y(new_n1360));
  NOR3xp33_ASAP7_75t_L      g01104(.A(new_n1360), .B(new_n1344), .C(new_n1343), .Y(new_n1361));
  OA21x2_ASAP7_75t_L        g01105(.A1(new_n1343), .A2(new_n1344), .B(new_n1360), .Y(new_n1362));
  NOR2xp33_ASAP7_75t_L      g01106(.A(new_n1361), .B(new_n1362), .Y(new_n1363));
  O2A1O1Ixp33_ASAP7_75t_L   g01107(.A1(new_n1163), .A2(new_n1263), .B(new_n1265), .C(new_n1363), .Y(new_n1364));
  INVx1_ASAP7_75t_L         g01108(.A(new_n1263), .Y(new_n1365));
  A2O1A1Ixp33_ASAP7_75t_L   g01109(.A1(new_n1157), .A2(\a[2] ), .B(new_n1162), .C(new_n1365), .Y(new_n1366));
  INVx1_ASAP7_75t_L         g01110(.A(new_n1366), .Y(new_n1367));
  A2O1A1O1Ixp25_ASAP7_75t_L g01111(.A1(new_n1135), .A2(new_n1264), .B(new_n1141), .C(new_n1261), .D(new_n1367), .Y(new_n1368));
  AND2x2_ASAP7_75t_L        g01112(.A(new_n1363), .B(new_n1368), .Y(new_n1369));
  NOR2xp33_ASAP7_75t_L      g01113(.A(new_n1364), .B(new_n1369), .Y(\f[17] ));
  NOR2xp33_ASAP7_75t_L      g01114(.A(new_n1343), .B(new_n1344), .Y(new_n1371));
  INVx1_ASAP7_75t_L         g01115(.A(new_n1342), .Y(new_n1372));
  OAI21xp33_ASAP7_75t_L     g01116(.A1(new_n1341), .A2(new_n1266), .B(new_n1372), .Y(new_n1373));
  NAND2xp33_ASAP7_75t_L     g01117(.A(\b[15] ), .B(new_n361), .Y(new_n1374));
  OAI221xp5_ASAP7_75t_L     g01118(.A1(new_n350), .A2(new_n960), .B1(new_n936), .B2(new_n375), .C(new_n1374), .Y(new_n1375));
  A2O1A1Ixp33_ASAP7_75t_L   g01119(.A1(new_n1052), .A2(new_n359), .B(new_n1375), .C(\a[5] ), .Y(new_n1376));
  AOI211xp5_ASAP7_75t_L     g01120(.A1(new_n1052), .A2(new_n359), .B(new_n1375), .C(new_n346), .Y(new_n1377));
  A2O1A1O1Ixp25_ASAP7_75t_L g01121(.A1(new_n1052), .A2(new_n359), .B(new_n1375), .C(new_n1376), .D(new_n1377), .Y(new_n1378));
  INVx1_ASAP7_75t_L         g01122(.A(new_n1239), .Y(new_n1379));
  A2O1A1O1Ixp25_ASAP7_75t_L g01123(.A1(new_n1238), .A2(new_n1174), .B(new_n1379), .C(new_n1326), .D(new_n1338), .Y(new_n1380));
  OAI22xp33_ASAP7_75t_L     g01124(.A1(new_n513), .A2(new_n748), .B1(new_n680), .B2(new_n506), .Y(new_n1381));
  AOI221xp5_ASAP7_75t_L     g01125(.A1(new_n475), .A2(\b[12] ), .B1(new_n483), .B2(new_n1057), .C(new_n1381), .Y(new_n1382));
  XNOR2x2_ASAP7_75t_L       g01126(.A(new_n466), .B(new_n1382), .Y(new_n1383));
  A2O1A1O1Ixp25_ASAP7_75t_L g01127(.A1(new_n1234), .A2(new_n1185), .B(new_n1281), .C(new_n1323), .D(new_n1321), .Y(new_n1384));
  A2O1A1O1Ixp25_ASAP7_75t_L g01128(.A1(new_n1222), .A2(new_n1193), .B(new_n1232), .C(new_n1312), .D(new_n1303), .Y(new_n1385));
  INVx1_ASAP7_75t_L         g01129(.A(\a[18] ), .Y(new_n1386));
  NAND2xp33_ASAP7_75t_L     g01130(.A(\a[17] ), .B(new_n1386), .Y(new_n1387));
  NAND2xp33_ASAP7_75t_L     g01131(.A(\a[18] ), .B(new_n1206), .Y(new_n1388));
  AND2x2_ASAP7_75t_L        g01132(.A(new_n1387), .B(new_n1388), .Y(new_n1389));
  NOR2xp33_ASAP7_75t_L      g01133(.A(new_n284), .B(new_n1389), .Y(new_n1390));
  A2O1A1Ixp33_ASAP7_75t_L   g01134(.A1(new_n1305), .A2(new_n1306), .B(new_n1213), .C(new_n1390), .Y(new_n1391));
  INVx1_ASAP7_75t_L         g01135(.A(new_n1390), .Y(new_n1392));
  NAND2xp33_ASAP7_75t_L     g01136(.A(new_n1392), .B(new_n1295), .Y(new_n1393));
  NAND2xp33_ASAP7_75t_L     g01137(.A(\b[3] ), .B(new_n1209), .Y(new_n1394));
  NAND2xp33_ASAP7_75t_L     g01138(.A(\b[1] ), .B(new_n1290), .Y(new_n1395));
  NAND2xp33_ASAP7_75t_L     g01139(.A(\b[2] ), .B(new_n1204), .Y(new_n1396));
  NAND2xp33_ASAP7_75t_L     g01140(.A(new_n1216), .B(new_n312), .Y(new_n1397));
  NAND4xp25_ASAP7_75t_L     g01141(.A(new_n1397), .B(new_n1394), .C(new_n1395), .D(new_n1396), .Y(new_n1398));
  OAI211xp5_ASAP7_75t_L     g01142(.A1(new_n1285), .A2(new_n262), .B(new_n1394), .C(new_n1396), .Y(new_n1399));
  A2O1A1Ixp33_ASAP7_75t_L   g01143(.A1(new_n312), .A2(new_n1216), .B(new_n1399), .C(\a[17] ), .Y(new_n1400));
  AOI211xp5_ASAP7_75t_L     g01144(.A1(new_n312), .A2(new_n1216), .B(new_n1206), .C(new_n1399), .Y(new_n1401));
  AOI21xp33_ASAP7_75t_L     g01145(.A1(new_n1400), .A2(new_n1398), .B(new_n1401), .Y(new_n1402));
  AOI21xp33_ASAP7_75t_L     g01146(.A1(new_n1393), .A2(new_n1391), .B(new_n1402), .Y(new_n1403));
  NOR2xp33_ASAP7_75t_L      g01147(.A(new_n1392), .B(new_n1295), .Y(new_n1404));
  NOR2xp33_ASAP7_75t_L      g01148(.A(new_n1390), .B(new_n1308), .Y(new_n1405));
  NAND5xp2_ASAP7_75t_L      g01149(.A(new_n1397), .B(new_n1396), .C(new_n1395), .D(new_n1394), .E(\a[17] ), .Y(new_n1406));
  A2O1A1Ixp33_ASAP7_75t_L   g01150(.A1(new_n312), .A2(new_n1216), .B(new_n1399), .C(new_n1206), .Y(new_n1407));
  NAND2xp33_ASAP7_75t_L     g01151(.A(new_n1406), .B(new_n1407), .Y(new_n1408));
  NOR3xp33_ASAP7_75t_L      g01152(.A(new_n1404), .B(new_n1405), .C(new_n1408), .Y(new_n1409));
  NOR2xp33_ASAP7_75t_L      g01153(.A(new_n427), .B(new_n869), .Y(new_n1410));
  AOI221xp5_ASAP7_75t_L     g01154(.A1(\b[4] ), .A2(new_n985), .B1(\b[5] ), .B2(new_n885), .C(new_n1410), .Y(new_n1411));
  O2A1O1Ixp33_ASAP7_75t_L   g01155(.A1(new_n872), .A2(new_n434), .B(new_n1411), .C(new_n867), .Y(new_n1412));
  OAI31xp33_ASAP7_75t_L     g01156(.A1(new_n433), .A2(new_n431), .A3(new_n872), .B(new_n1411), .Y(new_n1413));
  NAND2xp33_ASAP7_75t_L     g01157(.A(new_n867), .B(new_n1413), .Y(new_n1414));
  OAI21xp33_ASAP7_75t_L     g01158(.A1(new_n867), .A2(new_n1412), .B(new_n1414), .Y(new_n1415));
  NOR3xp33_ASAP7_75t_L      g01159(.A(new_n1409), .B(new_n1403), .C(new_n1415), .Y(new_n1416));
  OAI21xp33_ASAP7_75t_L     g01160(.A1(new_n1405), .A2(new_n1404), .B(new_n1408), .Y(new_n1417));
  NAND3xp33_ASAP7_75t_L     g01161(.A(new_n1393), .B(new_n1391), .C(new_n1402), .Y(new_n1418));
  OA21x2_ASAP7_75t_L        g01162(.A1(new_n867), .A2(new_n1412), .B(new_n1414), .Y(new_n1419));
  AOI21xp33_ASAP7_75t_L     g01163(.A1(new_n1417), .A2(new_n1418), .B(new_n1419), .Y(new_n1420));
  OR3x1_ASAP7_75t_L         g01164(.A(new_n1385), .B(new_n1416), .C(new_n1420), .Y(new_n1421));
  NAND3xp33_ASAP7_75t_L     g01165(.A(new_n1417), .B(new_n1418), .C(new_n1415), .Y(new_n1422));
  A2O1A1Ixp33_ASAP7_75t_L   g01166(.A1(new_n1415), .A2(new_n1422), .B(new_n1416), .C(new_n1385), .Y(new_n1423));
  NAND2xp33_ASAP7_75t_L     g01167(.A(\b[8] ), .B(new_n635), .Y(new_n1424));
  OAI221xp5_ASAP7_75t_L     g01168(.A1(new_n710), .A2(new_n590), .B1(new_n448), .B2(new_n712), .C(new_n1424), .Y(new_n1425));
  A2O1A1Ixp33_ASAP7_75t_L   g01169(.A1(new_n602), .A2(new_n718), .B(new_n1425), .C(\a[11] ), .Y(new_n1426));
  NAND2xp33_ASAP7_75t_L     g01170(.A(\a[11] ), .B(new_n1426), .Y(new_n1427));
  A2O1A1Ixp33_ASAP7_75t_L   g01171(.A1(new_n602), .A2(new_n718), .B(new_n1425), .C(new_n637), .Y(new_n1428));
  AOI22xp33_ASAP7_75t_L     g01172(.A1(new_n1427), .A2(new_n1428), .B1(new_n1423), .B2(new_n1421), .Y(new_n1429));
  AND4x1_ASAP7_75t_L        g01173(.A(new_n1421), .B(new_n1428), .C(new_n1423), .D(new_n1427), .Y(new_n1430));
  NOR3xp33_ASAP7_75t_L      g01174(.A(new_n1384), .B(new_n1430), .C(new_n1429), .Y(new_n1431));
  AO22x1_ASAP7_75t_L        g01175(.A1(new_n1428), .A2(new_n1427), .B1(new_n1423), .B2(new_n1421), .Y(new_n1432));
  NAND4xp25_ASAP7_75t_L     g01176(.A(new_n1421), .B(new_n1428), .C(new_n1427), .D(new_n1423), .Y(new_n1433));
  AOI211xp5_ASAP7_75t_L     g01177(.A1(new_n1433), .A2(new_n1432), .B(new_n1321), .C(new_n1322), .Y(new_n1434));
  OA21x2_ASAP7_75t_L        g01178(.A1(new_n1431), .A2(new_n1434), .B(new_n1383), .Y(new_n1435));
  NOR3xp33_ASAP7_75t_L      g01179(.A(new_n1383), .B(new_n1431), .C(new_n1434), .Y(new_n1436));
  NOR3xp33_ASAP7_75t_L      g01180(.A(new_n1380), .B(new_n1435), .C(new_n1436), .Y(new_n1437));
  AOI21xp33_ASAP7_75t_L     g01181(.A1(new_n1174), .A2(new_n1238), .B(new_n1379), .Y(new_n1438));
  OAI21xp33_ASAP7_75t_L     g01182(.A1(new_n1337), .A2(new_n1438), .B(new_n1332), .Y(new_n1439));
  OAI21xp33_ASAP7_75t_L     g01183(.A1(new_n1431), .A2(new_n1434), .B(new_n1383), .Y(new_n1440));
  OR3x1_ASAP7_75t_L         g01184(.A(new_n1383), .B(new_n1431), .C(new_n1434), .Y(new_n1441));
  AOI21xp33_ASAP7_75t_L     g01185(.A1(new_n1441), .A2(new_n1440), .B(new_n1439), .Y(new_n1442));
  NOR3xp33_ASAP7_75t_L      g01186(.A(new_n1442), .B(new_n1437), .C(new_n1378), .Y(new_n1443));
  INVx1_ASAP7_75t_L         g01187(.A(new_n1443), .Y(new_n1444));
  OAI21xp33_ASAP7_75t_L     g01188(.A1(new_n1437), .A2(new_n1442), .B(new_n1378), .Y(new_n1445));
  NAND3xp33_ASAP7_75t_L     g01189(.A(new_n1444), .B(new_n1373), .C(new_n1445), .Y(new_n1446));
  OAI21xp33_ASAP7_75t_L     g01190(.A1(new_n1022), .A2(new_n1025), .B(new_n979), .Y(new_n1447));
  A2O1A1O1Ixp25_ASAP7_75t_L g01191(.A1(new_n925), .A2(new_n949), .B(new_n929), .C(new_n1447), .D(new_n1027), .Y(new_n1448));
  A2O1A1Ixp33_ASAP7_75t_L   g01192(.A1(new_n1126), .A2(new_n1062), .B(new_n1448), .C(new_n1125), .Y(new_n1449));
  OAI21xp33_ASAP7_75t_L     g01193(.A1(new_n1340), .A2(new_n1334), .B(new_n1274), .Y(new_n1450));
  A2O1A1O1Ixp25_ASAP7_75t_L g01194(.A1(new_n1252), .A2(new_n1449), .B(new_n1248), .C(new_n1450), .D(new_n1342), .Y(new_n1451));
  OA21x2_ASAP7_75t_L        g01195(.A1(new_n1437), .A2(new_n1442), .B(new_n1378), .Y(new_n1452));
  OAI21xp33_ASAP7_75t_L     g01196(.A1(new_n1443), .A2(new_n1452), .B(new_n1451), .Y(new_n1453));
  NOR2xp33_ASAP7_75t_L      g01197(.A(new_n1150), .B(new_n287), .Y(new_n1454));
  AOI221xp5_ASAP7_75t_L     g01198(.A1(\b[17] ), .A2(new_n264), .B1(\b[18] ), .B2(new_n283), .C(new_n1454), .Y(new_n1455));
  A2O1A1Ixp33_ASAP7_75t_L   g01199(.A1(new_n1049), .A2(new_n1148), .B(new_n1149), .C(new_n1347), .Y(new_n1456));
  NOR2xp33_ASAP7_75t_L      g01200(.A(\b[17] ), .B(\b[18] ), .Y(new_n1457));
  INVx1_ASAP7_75t_L         g01201(.A(\b[18] ), .Y(new_n1458));
  NOR2xp33_ASAP7_75t_L      g01202(.A(new_n1349), .B(new_n1458), .Y(new_n1459));
  NOR2xp33_ASAP7_75t_L      g01203(.A(new_n1457), .B(new_n1459), .Y(new_n1460));
  A2O1A1Ixp33_ASAP7_75t_L   g01204(.A1(new_n1456), .A2(new_n1351), .B(new_n1350), .C(new_n1460), .Y(new_n1461));
  NOR3xp33_ASAP7_75t_L      g01205(.A(new_n1353), .B(new_n1460), .C(new_n1350), .Y(new_n1462));
  INVx1_ASAP7_75t_L         g01206(.A(new_n1462), .Y(new_n1463));
  NAND2xp33_ASAP7_75t_L     g01207(.A(new_n1461), .B(new_n1463), .Y(new_n1464));
  O2A1O1Ixp33_ASAP7_75t_L   g01208(.A1(new_n279), .A2(new_n1464), .B(new_n1455), .C(new_n257), .Y(new_n1465));
  OAI21xp33_ASAP7_75t_L     g01209(.A1(new_n279), .A2(new_n1464), .B(new_n1455), .Y(new_n1466));
  NAND2xp33_ASAP7_75t_L     g01210(.A(new_n257), .B(new_n1466), .Y(new_n1467));
  OA21x2_ASAP7_75t_L        g01211(.A1(new_n257), .A2(new_n1465), .B(new_n1467), .Y(new_n1468));
  NAND3xp33_ASAP7_75t_L     g01212(.A(new_n1446), .B(new_n1468), .C(new_n1453), .Y(new_n1469));
  AO21x2_ASAP7_75t_L        g01213(.A1(new_n1453), .A2(new_n1446), .B(new_n1468), .Y(new_n1470));
  NAND2xp33_ASAP7_75t_L     g01214(.A(new_n1469), .B(new_n1470), .Y(new_n1471));
  A2O1A1Ixp33_ASAP7_75t_L   g01215(.A1(new_n1360), .A2(new_n1371), .B(new_n1364), .C(new_n1471), .Y(new_n1472));
  INVx1_ASAP7_75t_L         g01216(.A(new_n1472), .Y(new_n1473));
  A2O1A1Ixp33_ASAP7_75t_L   g01217(.A1(\a[2] ), .A2(new_n1358), .B(new_n1359), .C(new_n1371), .Y(new_n1474));
  A2O1A1Ixp33_ASAP7_75t_L   g01218(.A1(new_n1265), .A2(new_n1366), .B(new_n1363), .C(new_n1474), .Y(new_n1475));
  NOR2xp33_ASAP7_75t_L      g01219(.A(new_n1471), .B(new_n1475), .Y(new_n1476));
  NOR2xp33_ASAP7_75t_L      g01220(.A(new_n1476), .B(new_n1473), .Y(\f[18] ));
  NOR2xp33_ASAP7_75t_L      g01221(.A(new_n960), .B(new_n375), .Y(new_n1478));
  AOI221xp5_ASAP7_75t_L     g01222(.A1(\b[16] ), .A2(new_n361), .B1(new_n349), .B2(\b[15] ), .C(new_n1478), .Y(new_n1479));
  OAI211xp5_ASAP7_75t_L     g01223(.A1(new_n356), .A2(new_n1161), .B(\a[5] ), .C(new_n1479), .Y(new_n1480));
  INVx1_ASAP7_75t_L         g01224(.A(new_n1479), .Y(new_n1481));
  A2O1A1Ixp33_ASAP7_75t_L   g01225(.A1(new_n1156), .A2(new_n359), .B(new_n1481), .C(new_n346), .Y(new_n1482));
  NAND2xp33_ASAP7_75t_L     g01226(.A(new_n1482), .B(new_n1480), .Y(new_n1483));
  NAND3xp33_ASAP7_75t_L     g01227(.A(new_n1417), .B(new_n1419), .C(new_n1418), .Y(new_n1484));
  A2O1A1Ixp33_ASAP7_75t_L   g01228(.A1(new_n1484), .A2(new_n1419), .B(new_n1385), .C(new_n1422), .Y(new_n1485));
  NOR2xp33_ASAP7_75t_L      g01229(.A(new_n448), .B(new_n869), .Y(new_n1486));
  AOI221xp5_ASAP7_75t_L     g01230(.A1(\b[5] ), .A2(new_n985), .B1(\b[6] ), .B2(new_n885), .C(new_n1486), .Y(new_n1487));
  O2A1O1Ixp33_ASAP7_75t_L   g01231(.A1(new_n872), .A2(new_n456), .B(new_n1487), .C(new_n867), .Y(new_n1488));
  OAI21xp33_ASAP7_75t_L     g01232(.A1(new_n872), .A2(new_n456), .B(new_n1487), .Y(new_n1489));
  NAND2xp33_ASAP7_75t_L     g01233(.A(new_n867), .B(new_n1489), .Y(new_n1490));
  OAI21xp33_ASAP7_75t_L     g01234(.A1(new_n867), .A2(new_n1488), .B(new_n1490), .Y(new_n1491));
  MAJIxp5_ASAP7_75t_L       g01235(.A(new_n1402), .B(new_n1308), .C(new_n1392), .Y(new_n1492));
  NAND2xp33_ASAP7_75t_L     g01236(.A(\b[3] ), .B(new_n1204), .Y(new_n1493));
  OAI221xp5_ASAP7_75t_L     g01237(.A1(new_n1284), .A2(new_n332), .B1(new_n289), .B2(new_n1285), .C(new_n1493), .Y(new_n1494));
  AOI211xp5_ASAP7_75t_L     g01238(.A1(new_n342), .A2(new_n1216), .B(new_n1206), .C(new_n1494), .Y(new_n1495));
  INVx1_ASAP7_75t_L         g01239(.A(new_n341), .Y(new_n1496));
  NAND2xp33_ASAP7_75t_L     g01240(.A(new_n338), .B(new_n1496), .Y(new_n1497));
  NOR2xp33_ASAP7_75t_L      g01241(.A(new_n332), .B(new_n1284), .Y(new_n1498));
  AOI221xp5_ASAP7_75t_L     g01242(.A1(\b[2] ), .A2(new_n1290), .B1(\b[3] ), .B2(new_n1204), .C(new_n1498), .Y(new_n1499));
  O2A1O1Ixp33_ASAP7_75t_L   g01243(.A1(new_n1210), .A2(new_n1497), .B(new_n1499), .C(\a[17] ), .Y(new_n1500));
  INVx1_ASAP7_75t_L         g01244(.A(\a[20] ), .Y(new_n1501));
  NAND2xp33_ASAP7_75t_L     g01245(.A(new_n1388), .B(new_n1387), .Y(new_n1502));
  INVx1_ASAP7_75t_L         g01246(.A(\a[19] ), .Y(new_n1503));
  NOR2xp33_ASAP7_75t_L      g01247(.A(\a[18] ), .B(new_n1503), .Y(new_n1504));
  NOR2xp33_ASAP7_75t_L      g01248(.A(\a[19] ), .B(new_n1386), .Y(new_n1505));
  NOR2xp33_ASAP7_75t_L      g01249(.A(new_n1504), .B(new_n1505), .Y(new_n1506));
  NOR2xp33_ASAP7_75t_L      g01250(.A(new_n1502), .B(new_n1506), .Y(new_n1507));
  NAND2xp33_ASAP7_75t_L     g01251(.A(\a[20] ), .B(new_n1503), .Y(new_n1508));
  NAND2xp33_ASAP7_75t_L     g01252(.A(\a[19] ), .B(new_n1501), .Y(new_n1509));
  NAND2xp33_ASAP7_75t_L     g01253(.A(new_n1509), .B(new_n1508), .Y(new_n1510));
  NOR2xp33_ASAP7_75t_L      g01254(.A(new_n1510), .B(new_n1389), .Y(new_n1511));
  AOI22xp33_ASAP7_75t_L     g01255(.A1(new_n1507), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n1511), .Y(new_n1512));
  AOI21xp33_ASAP7_75t_L     g01256(.A1(new_n1509), .A2(new_n1508), .B(new_n1389), .Y(new_n1513));
  NAND2xp33_ASAP7_75t_L     g01257(.A(new_n275), .B(new_n1513), .Y(new_n1514));
  NAND2xp33_ASAP7_75t_L     g01258(.A(new_n1514), .B(new_n1512), .Y(new_n1515));
  NOR3xp33_ASAP7_75t_L      g01259(.A(new_n1515), .B(new_n1390), .C(new_n1501), .Y(new_n1516));
  OAI21xp33_ASAP7_75t_L     g01260(.A1(new_n1504), .A2(new_n1505), .B(new_n1389), .Y(new_n1517));
  NAND3xp33_ASAP7_75t_L     g01261(.A(new_n1502), .B(new_n1508), .C(new_n1509), .Y(new_n1518));
  OAI22xp33_ASAP7_75t_L     g01262(.A1(new_n1517), .A2(new_n284), .B1(new_n262), .B2(new_n1518), .Y(new_n1519));
  A2O1A1Ixp33_ASAP7_75t_L   g01263(.A1(new_n1513), .A2(new_n275), .B(new_n1519), .C(\a[20] ), .Y(new_n1520));
  NAND2xp33_ASAP7_75t_L     g01264(.A(new_n1510), .B(new_n1502), .Y(new_n1521));
  O2A1O1Ixp33_ASAP7_75t_L   g01265(.A1(new_n1521), .A2(new_n274), .B(new_n1512), .C(\a[20] ), .Y(new_n1522));
  O2A1O1Ixp33_ASAP7_75t_L   g01266(.A1(new_n1392), .A2(new_n1520), .B(\a[20] ), .C(new_n1522), .Y(new_n1523));
  NOR4xp25_ASAP7_75t_L      g01267(.A(new_n1523), .B(new_n1495), .C(new_n1500), .D(new_n1516), .Y(new_n1524));
  OAI211xp5_ASAP7_75t_L     g01268(.A1(new_n1497), .A2(new_n1210), .B(new_n1499), .C(\a[17] ), .Y(new_n1525));
  A2O1A1Ixp33_ASAP7_75t_L   g01269(.A1(new_n342), .A2(new_n1216), .B(new_n1494), .C(new_n1206), .Y(new_n1526));
  AOI21xp33_ASAP7_75t_L     g01270(.A1(new_n275), .A2(new_n1513), .B(new_n1519), .Y(new_n1527));
  NAND3xp33_ASAP7_75t_L     g01271(.A(new_n1527), .B(new_n1392), .C(\a[20] ), .Y(new_n1528));
  O2A1O1Ixp33_ASAP7_75t_L   g01272(.A1(new_n1521), .A2(new_n274), .B(new_n1512), .C(new_n1501), .Y(new_n1529));
  A2O1A1Ixp33_ASAP7_75t_L   g01273(.A1(new_n1513), .A2(new_n275), .B(new_n1519), .C(new_n1501), .Y(new_n1530));
  A2O1A1Ixp33_ASAP7_75t_L   g01274(.A1(new_n1529), .A2(new_n1390), .B(new_n1501), .C(new_n1530), .Y(new_n1531));
  AOI22xp33_ASAP7_75t_L     g01275(.A1(new_n1525), .A2(new_n1526), .B1(new_n1528), .B2(new_n1531), .Y(new_n1532));
  OAI21xp33_ASAP7_75t_L     g01276(.A1(new_n1524), .A2(new_n1532), .B(new_n1492), .Y(new_n1533));
  MAJIxp5_ASAP7_75t_L       g01277(.A(new_n1408), .B(new_n1390), .C(new_n1295), .Y(new_n1534));
  NAND4xp25_ASAP7_75t_L     g01278(.A(new_n1531), .B(new_n1525), .C(new_n1526), .D(new_n1528), .Y(new_n1535));
  OAI22xp33_ASAP7_75t_L     g01279(.A1(new_n1523), .A2(new_n1516), .B1(new_n1500), .B2(new_n1495), .Y(new_n1536));
  NAND3xp33_ASAP7_75t_L     g01280(.A(new_n1534), .B(new_n1535), .C(new_n1536), .Y(new_n1537));
  NAND3xp33_ASAP7_75t_L     g01281(.A(new_n1533), .B(new_n1537), .C(new_n1491), .Y(new_n1538));
  AOI21xp33_ASAP7_75t_L     g01282(.A1(new_n1533), .A2(new_n1537), .B(new_n1491), .Y(new_n1539));
  INVx1_ASAP7_75t_L         g01283(.A(new_n1539), .Y(new_n1540));
  NAND3xp33_ASAP7_75t_L     g01284(.A(new_n1485), .B(new_n1540), .C(new_n1538), .Y(new_n1541));
  O2A1O1Ixp33_ASAP7_75t_L   g01285(.A1(new_n1230), .A2(new_n1231), .B(new_n1228), .C(new_n1309), .Y(new_n1542));
  OAI22xp33_ASAP7_75t_L     g01286(.A1(new_n1542), .A2(new_n1303), .B1(new_n1420), .B2(new_n1416), .Y(new_n1543));
  OA21x2_ASAP7_75t_L        g01287(.A1(new_n867), .A2(new_n1488), .B(new_n1490), .Y(new_n1544));
  AOI21xp33_ASAP7_75t_L     g01288(.A1(new_n1536), .A2(new_n1535), .B(new_n1534), .Y(new_n1545));
  NAND2xp33_ASAP7_75t_L     g01289(.A(new_n1535), .B(new_n1536), .Y(new_n1546));
  NOR2xp33_ASAP7_75t_L      g01290(.A(new_n1492), .B(new_n1546), .Y(new_n1547));
  NOR3xp33_ASAP7_75t_L      g01291(.A(new_n1547), .B(new_n1544), .C(new_n1545), .Y(new_n1548));
  OAI211xp5_ASAP7_75t_L     g01292(.A1(new_n1548), .A2(new_n1539), .B(new_n1543), .C(new_n1422), .Y(new_n1549));
  INVx1_ASAP7_75t_L         g01293(.A(new_n635), .Y(new_n1550));
  NOR2xp33_ASAP7_75t_L      g01294(.A(new_n590), .B(new_n1550), .Y(new_n1551));
  AOI221xp5_ASAP7_75t_L     g01295(.A1(\b[8] ), .A2(new_n713), .B1(\b[10] ), .B2(new_n640), .C(new_n1551), .Y(new_n1552));
  O2A1O1Ixp33_ASAP7_75t_L   g01296(.A1(new_n641), .A2(new_n1175), .B(new_n1552), .C(new_n637), .Y(new_n1553));
  INVx1_ASAP7_75t_L         g01297(.A(new_n1553), .Y(new_n1554));
  O2A1O1Ixp33_ASAP7_75t_L   g01298(.A1(new_n641), .A2(new_n1175), .B(new_n1552), .C(\a[11] ), .Y(new_n1555));
  AOI21xp33_ASAP7_75t_L     g01299(.A1(new_n1554), .A2(\a[11] ), .B(new_n1555), .Y(new_n1556));
  AND3x1_ASAP7_75t_L        g01300(.A(new_n1541), .B(new_n1549), .C(new_n1556), .Y(new_n1557));
  AOI21xp33_ASAP7_75t_L     g01301(.A1(new_n1541), .A2(new_n1549), .B(new_n1556), .Y(new_n1558));
  OAI21xp33_ASAP7_75t_L     g01302(.A1(new_n1430), .A2(new_n1384), .B(new_n1432), .Y(new_n1559));
  NOR3xp33_ASAP7_75t_L      g01303(.A(new_n1559), .B(new_n1558), .C(new_n1557), .Y(new_n1560));
  NAND3xp33_ASAP7_75t_L     g01304(.A(new_n1541), .B(new_n1549), .C(new_n1556), .Y(new_n1561));
  AO21x2_ASAP7_75t_L        g01305(.A1(new_n1549), .A2(new_n1541), .B(new_n1556), .Y(new_n1562));
  A2O1A1O1Ixp25_ASAP7_75t_L g01306(.A1(new_n1323), .A2(new_n1329), .B(new_n1321), .C(new_n1433), .D(new_n1429), .Y(new_n1563));
  AOI21xp33_ASAP7_75t_L     g01307(.A1(new_n1562), .A2(new_n1561), .B(new_n1563), .Y(new_n1564));
  NOR2xp33_ASAP7_75t_L      g01308(.A(new_n833), .B(new_n513), .Y(new_n1565));
  AOI221xp5_ASAP7_75t_L     g01309(.A1(\b[11] ), .A2(new_n560), .B1(\b[13] ), .B2(new_n475), .C(new_n1565), .Y(new_n1566));
  INVx1_ASAP7_75t_L         g01310(.A(new_n1566), .Y(new_n1567));
  A2O1A1Ixp33_ASAP7_75t_L   g01311(.A1(new_n1166), .A2(new_n483), .B(new_n1567), .C(\a[8] ), .Y(new_n1568));
  O2A1O1Ixp33_ASAP7_75t_L   g01312(.A1(new_n477), .A2(new_n942), .B(new_n1566), .C(\a[8] ), .Y(new_n1569));
  AOI21xp33_ASAP7_75t_L     g01313(.A1(new_n1568), .A2(\a[8] ), .B(new_n1569), .Y(new_n1570));
  OAI21xp33_ASAP7_75t_L     g01314(.A1(new_n1564), .A2(new_n1560), .B(new_n1570), .Y(new_n1571));
  NAND3xp33_ASAP7_75t_L     g01315(.A(new_n1563), .B(new_n1562), .C(new_n1561), .Y(new_n1572));
  OAI21xp33_ASAP7_75t_L     g01316(.A1(new_n1557), .A2(new_n1558), .B(new_n1559), .Y(new_n1573));
  O2A1O1Ixp33_ASAP7_75t_L   g01317(.A1(new_n477), .A2(new_n942), .B(new_n1566), .C(new_n466), .Y(new_n1574));
  NOR2xp33_ASAP7_75t_L      g01318(.A(new_n466), .B(new_n1574), .Y(new_n1575));
  OAI211xp5_ASAP7_75t_L     g01319(.A1(new_n1575), .A2(new_n1569), .B(new_n1572), .C(new_n1573), .Y(new_n1576));
  OAI21xp33_ASAP7_75t_L     g01320(.A1(new_n1435), .A2(new_n1380), .B(new_n1441), .Y(new_n1577));
  NAND3xp33_ASAP7_75t_L     g01321(.A(new_n1577), .B(new_n1576), .C(new_n1571), .Y(new_n1578));
  NAND2xp33_ASAP7_75t_L     g01322(.A(new_n1576), .B(new_n1571), .Y(new_n1579));
  A2O1A1O1Ixp25_ASAP7_75t_L g01323(.A1(new_n1339), .A2(new_n1336), .B(new_n1338), .C(new_n1440), .D(new_n1436), .Y(new_n1580));
  NAND2xp33_ASAP7_75t_L     g01324(.A(new_n1579), .B(new_n1580), .Y(new_n1581));
  NAND3xp33_ASAP7_75t_L     g01325(.A(new_n1578), .B(new_n1581), .C(new_n1483), .Y(new_n1582));
  O2A1O1Ixp33_ASAP7_75t_L   g01326(.A1(new_n1380), .A2(new_n1435), .B(new_n1441), .C(new_n1579), .Y(new_n1583));
  AOI21xp33_ASAP7_75t_L     g01327(.A1(new_n1576), .A2(new_n1571), .B(new_n1577), .Y(new_n1584));
  NOR3xp33_ASAP7_75t_L      g01328(.A(new_n1584), .B(new_n1583), .C(new_n1483), .Y(new_n1585));
  AOI21xp33_ASAP7_75t_L     g01329(.A1(new_n1582), .A2(new_n1483), .B(new_n1585), .Y(new_n1586));
  OAI21xp33_ASAP7_75t_L     g01330(.A1(new_n1254), .A2(new_n1251), .B(new_n1253), .Y(new_n1587));
  A2O1A1O1Ixp25_ASAP7_75t_L g01331(.A1(new_n1450), .A2(new_n1587), .B(new_n1342), .C(new_n1445), .D(new_n1443), .Y(new_n1588));
  NAND2xp33_ASAP7_75t_L     g01332(.A(new_n1586), .B(new_n1588), .Y(new_n1589));
  NAND4xp25_ASAP7_75t_L     g01333(.A(new_n1578), .B(new_n1482), .C(new_n1581), .D(new_n1480), .Y(new_n1590));
  OAI21xp33_ASAP7_75t_L     g01334(.A1(new_n1583), .A2(new_n1584), .B(new_n1483), .Y(new_n1591));
  NAND2xp33_ASAP7_75t_L     g01335(.A(new_n1590), .B(new_n1591), .Y(new_n1592));
  A2O1A1Ixp33_ASAP7_75t_L   g01336(.A1(new_n1445), .A2(new_n1373), .B(new_n1443), .C(new_n1592), .Y(new_n1593));
  NAND2xp33_ASAP7_75t_L     g01337(.A(new_n1593), .B(new_n1589), .Y(new_n1594));
  NOR2xp33_ASAP7_75t_L      g01338(.A(new_n1349), .B(new_n287), .Y(new_n1595));
  AOI221xp5_ASAP7_75t_L     g01339(.A1(\b[18] ), .A2(new_n264), .B1(\b[19] ), .B2(new_n283), .C(new_n1595), .Y(new_n1596));
  INVx1_ASAP7_75t_L         g01340(.A(new_n1596), .Y(new_n1597));
  NOR2xp33_ASAP7_75t_L      g01341(.A(\b[18] ), .B(\b[19] ), .Y(new_n1598));
  INVx1_ASAP7_75t_L         g01342(.A(\b[19] ), .Y(new_n1599));
  NOR2xp33_ASAP7_75t_L      g01343(.A(new_n1458), .B(new_n1599), .Y(new_n1600));
  NOR2xp33_ASAP7_75t_L      g01344(.A(new_n1598), .B(new_n1600), .Y(new_n1601));
  INVx1_ASAP7_75t_L         g01345(.A(new_n1601), .Y(new_n1602));
  O2A1O1Ixp33_ASAP7_75t_L   g01346(.A1(new_n1349), .A2(new_n1458), .B(new_n1461), .C(new_n1602), .Y(new_n1603));
  A2O1A1O1Ixp25_ASAP7_75t_L g01347(.A1(new_n1351), .A2(new_n1456), .B(new_n1350), .C(new_n1460), .D(new_n1459), .Y(new_n1604));
  NAND2xp33_ASAP7_75t_L     g01348(.A(new_n1602), .B(new_n1604), .Y(new_n1605));
  INVx1_ASAP7_75t_L         g01349(.A(new_n1605), .Y(new_n1606));
  NOR2xp33_ASAP7_75t_L      g01350(.A(new_n1603), .B(new_n1606), .Y(new_n1607));
  A2O1A1Ixp33_ASAP7_75t_L   g01351(.A1(new_n1607), .A2(new_n273), .B(new_n1597), .C(\a[2] ), .Y(new_n1608));
  INVx1_ASAP7_75t_L         g01352(.A(new_n1608), .Y(new_n1609));
  A2O1A1Ixp33_ASAP7_75t_L   g01353(.A1(new_n1607), .A2(new_n273), .B(new_n1597), .C(new_n257), .Y(new_n1610));
  O2A1O1Ixp33_ASAP7_75t_L   g01354(.A1(new_n1609), .A2(new_n257), .B(new_n1610), .C(new_n1594), .Y(new_n1611));
  OAI21xp33_ASAP7_75t_L     g01355(.A1(new_n1452), .A2(new_n1451), .B(new_n1444), .Y(new_n1612));
  NOR2xp33_ASAP7_75t_L      g01356(.A(new_n1592), .B(new_n1612), .Y(new_n1613));
  NOR2xp33_ASAP7_75t_L      g01357(.A(new_n1586), .B(new_n1588), .Y(new_n1614));
  NAND2xp33_ASAP7_75t_L     g01358(.A(\a[2] ), .B(new_n1608), .Y(new_n1615));
  NAND2xp33_ASAP7_75t_L     g01359(.A(new_n1610), .B(new_n1615), .Y(new_n1616));
  OAI21xp33_ASAP7_75t_L     g01360(.A1(new_n1614), .A2(new_n1613), .B(new_n1616), .Y(new_n1617));
  NAND2xp33_ASAP7_75t_L     g01361(.A(new_n1453), .B(new_n1446), .Y(new_n1618));
  O2A1O1Ixp33_ASAP7_75t_L   g01362(.A1(new_n1465), .A2(new_n257), .B(new_n1467), .C(new_n1618), .Y(new_n1619));
  A2O1A1O1Ixp25_ASAP7_75t_L g01363(.A1(new_n1360), .A2(new_n1371), .B(new_n1364), .C(new_n1471), .D(new_n1619), .Y(new_n1620));
  O2A1O1Ixp33_ASAP7_75t_L   g01364(.A1(new_n1594), .A2(new_n1611), .B(new_n1617), .C(new_n1620), .Y(new_n1621));
  NAND4xp25_ASAP7_75t_L     g01365(.A(new_n1589), .B(new_n1593), .C(new_n1610), .D(new_n1615), .Y(new_n1622));
  NAND2xp33_ASAP7_75t_L     g01366(.A(new_n1622), .B(new_n1617), .Y(new_n1623));
  NOR3xp33_ASAP7_75t_L      g01367(.A(new_n1473), .B(new_n1623), .C(new_n1619), .Y(new_n1624));
  NOR2xp33_ASAP7_75t_L      g01368(.A(new_n1621), .B(new_n1624), .Y(\f[19] ));
  INVx1_ASAP7_75t_L         g01369(.A(new_n1594), .Y(new_n1626));
  INVx1_ASAP7_75t_L         g01370(.A(new_n1603), .Y(new_n1627));
  NAND2xp33_ASAP7_75t_L     g01371(.A(new_n1605), .B(new_n1627), .Y(new_n1628));
  O2A1O1Ixp33_ASAP7_75t_L   g01372(.A1(new_n279), .A2(new_n1628), .B(new_n1596), .C(\a[2] ), .Y(new_n1629));
  A2O1A1Ixp33_ASAP7_75t_L   g01373(.A1(\a[2] ), .A2(new_n1608), .B(new_n1629), .C(new_n1626), .Y(new_n1630));
  INVx1_ASAP7_75t_L         g01374(.A(new_n1582), .Y(new_n1631));
  INVx1_ASAP7_75t_L         g01375(.A(new_n1355), .Y(new_n1632));
  NOR2xp33_ASAP7_75t_L      g01376(.A(new_n1353), .B(new_n1632), .Y(new_n1633));
  NAND2xp33_ASAP7_75t_L     g01377(.A(\b[17] ), .B(new_n361), .Y(new_n1634));
  OAI221xp5_ASAP7_75t_L     g01378(.A1(new_n350), .A2(new_n1150), .B1(new_n1043), .B2(new_n375), .C(new_n1634), .Y(new_n1635));
  A2O1A1Ixp33_ASAP7_75t_L   g01379(.A1(new_n1633), .A2(new_n359), .B(new_n1635), .C(\a[5] ), .Y(new_n1636));
  AOI211xp5_ASAP7_75t_L     g01380(.A1(new_n1633), .A2(new_n359), .B(new_n1635), .C(new_n346), .Y(new_n1637));
  A2O1A1O1Ixp25_ASAP7_75t_L g01381(.A1(new_n1633), .A2(new_n359), .B(new_n1635), .C(new_n1636), .D(new_n1637), .Y(new_n1638));
  INVx1_ASAP7_75t_L         g01382(.A(new_n1576), .Y(new_n1639));
  NAND2xp33_ASAP7_75t_L     g01383(.A(new_n1549), .B(new_n1541), .Y(new_n1640));
  MAJIxp5_ASAP7_75t_L       g01384(.A(new_n1563), .B(new_n1640), .C(new_n1556), .Y(new_n1641));
  NOR2xp33_ASAP7_75t_L      g01385(.A(new_n680), .B(new_n1550), .Y(new_n1642));
  AOI221xp5_ASAP7_75t_L     g01386(.A1(\b[9] ), .A2(new_n713), .B1(\b[11] ), .B2(new_n640), .C(new_n1642), .Y(new_n1643));
  O2A1O1Ixp33_ASAP7_75t_L   g01387(.A1(new_n641), .A2(new_n754), .B(new_n1643), .C(new_n637), .Y(new_n1644));
  INVx1_ASAP7_75t_L         g01388(.A(new_n1643), .Y(new_n1645));
  A2O1A1Ixp33_ASAP7_75t_L   g01389(.A1(new_n976), .A2(new_n718), .B(new_n1645), .C(new_n637), .Y(new_n1646));
  OAI21xp33_ASAP7_75t_L     g01390(.A1(new_n637), .A2(new_n1644), .B(new_n1646), .Y(new_n1647));
  INVx1_ASAP7_75t_L         g01391(.A(new_n1647), .Y(new_n1648));
  AOI21xp33_ASAP7_75t_L     g01392(.A1(new_n1485), .A2(new_n1540), .B(new_n1548), .Y(new_n1649));
  A2O1A1Ixp33_ASAP7_75t_L   g01393(.A1(new_n342), .A2(new_n1216), .B(new_n1494), .C(\a[17] ), .Y(new_n1650));
  INVx1_ASAP7_75t_L         g01394(.A(new_n1650), .Y(new_n1651));
  NAND2xp33_ASAP7_75t_L     g01395(.A(new_n1528), .B(new_n1531), .Y(new_n1652));
  O2A1O1Ixp33_ASAP7_75t_L   g01396(.A1(new_n1206), .A2(new_n1651), .B(new_n1526), .C(new_n1652), .Y(new_n1653));
  NAND3xp33_ASAP7_75t_L     g01397(.A(new_n1389), .B(new_n1506), .C(new_n1510), .Y(new_n1654));
  NAND2xp33_ASAP7_75t_L     g01398(.A(\b[1] ), .B(new_n1507), .Y(new_n1655));
  OAI221xp5_ASAP7_75t_L     g01399(.A1(new_n1518), .A2(new_n289), .B1(new_n284), .B2(new_n1654), .C(new_n1655), .Y(new_n1656));
  A2O1A1Ixp33_ASAP7_75t_L   g01400(.A1(new_n294), .A2(new_n1513), .B(new_n1656), .C(\a[20] ), .Y(new_n1657));
  NOR2xp33_ASAP7_75t_L      g01401(.A(new_n289), .B(new_n1518), .Y(new_n1658));
  AND3x1_ASAP7_75t_L        g01402(.A(new_n1389), .B(new_n1510), .C(new_n1506), .Y(new_n1659));
  AOI221xp5_ASAP7_75t_L     g01403(.A1(new_n1507), .A2(\b[1] ), .B1(new_n1659), .B2(\b[0] ), .C(new_n1658), .Y(new_n1660));
  O2A1O1Ixp33_ASAP7_75t_L   g01404(.A1(new_n509), .A2(new_n1521), .B(new_n1660), .C(\a[20] ), .Y(new_n1661));
  A2O1A1O1Ixp25_ASAP7_75t_L g01405(.A1(new_n1527), .A2(new_n1392), .B(new_n1657), .C(\a[20] ), .D(new_n1661), .Y(new_n1662));
  NOR2xp33_ASAP7_75t_L      g01406(.A(new_n1521), .B(new_n509), .Y(new_n1663));
  NOR5xp2_ASAP7_75t_L       g01407(.A(new_n1515), .B(new_n1656), .C(new_n1663), .D(new_n1390), .E(new_n1501), .Y(new_n1664));
  NAND2xp33_ASAP7_75t_L     g01408(.A(\b[4] ), .B(new_n1204), .Y(new_n1665));
  OAI221xp5_ASAP7_75t_L     g01409(.A1(new_n1284), .A2(new_n384), .B1(new_n301), .B2(new_n1285), .C(new_n1665), .Y(new_n1666));
  A2O1A1Ixp33_ASAP7_75t_L   g01410(.A1(new_n394), .A2(new_n1216), .B(new_n1666), .C(\a[17] ), .Y(new_n1667));
  INVx1_ASAP7_75t_L         g01411(.A(new_n1666), .Y(new_n1668));
  O2A1O1Ixp33_ASAP7_75t_L   g01412(.A1(new_n1210), .A2(new_n728), .B(new_n1668), .C(\a[17] ), .Y(new_n1669));
  AOI21xp33_ASAP7_75t_L     g01413(.A1(new_n1667), .A2(\a[17] ), .B(new_n1669), .Y(new_n1670));
  NOR3xp33_ASAP7_75t_L      g01414(.A(new_n1670), .B(new_n1662), .C(new_n1664), .Y(new_n1671));
  INVx1_ASAP7_75t_L         g01415(.A(new_n1663), .Y(new_n1672));
  NAND3xp33_ASAP7_75t_L     g01416(.A(new_n1660), .B(\a[20] ), .C(new_n1672), .Y(new_n1673));
  A2O1A1Ixp33_ASAP7_75t_L   g01417(.A1(new_n294), .A2(new_n1513), .B(new_n1656), .C(new_n1501), .Y(new_n1674));
  NAND3xp33_ASAP7_75t_L     g01418(.A(new_n1528), .B(new_n1673), .C(new_n1674), .Y(new_n1675));
  NAND5xp2_ASAP7_75t_L      g01419(.A(\a[20] ), .B(new_n1527), .C(new_n1660), .D(new_n1672), .E(new_n1392), .Y(new_n1676));
  AOI221xp5_ASAP7_75t_L     g01420(.A1(new_n1667), .A2(\a[17] ), .B1(new_n1676), .B2(new_n1675), .C(new_n1669), .Y(new_n1677));
  OAI22xp33_ASAP7_75t_L     g01421(.A1(new_n1545), .A2(new_n1653), .B1(new_n1677), .B2(new_n1671), .Y(new_n1678));
  NOR2xp33_ASAP7_75t_L      g01422(.A(new_n1516), .B(new_n1523), .Y(new_n1679));
  A2O1A1Ixp33_ASAP7_75t_L   g01423(.A1(new_n1650), .A2(\a[17] ), .B(new_n1500), .C(new_n1679), .Y(new_n1680));
  OR3x1_ASAP7_75t_L         g01424(.A(new_n1670), .B(new_n1662), .C(new_n1664), .Y(new_n1681));
  OAI21xp33_ASAP7_75t_L     g01425(.A1(new_n1664), .A2(new_n1662), .B(new_n1670), .Y(new_n1682));
  NAND4xp25_ASAP7_75t_L     g01426(.A(new_n1533), .B(new_n1681), .C(new_n1682), .D(new_n1680), .Y(new_n1683));
  AND2x2_ASAP7_75t_L        g01427(.A(new_n537), .B(new_n539), .Y(new_n1684));
  NOR2xp33_ASAP7_75t_L      g01428(.A(new_n448), .B(new_n864), .Y(new_n1685));
  AOI221xp5_ASAP7_75t_L     g01429(.A1(\b[6] ), .A2(new_n985), .B1(\b[8] ), .B2(new_n886), .C(new_n1685), .Y(new_n1686));
  INVx1_ASAP7_75t_L         g01430(.A(new_n1686), .Y(new_n1687));
  A2O1A1Ixp33_ASAP7_75t_L   g01431(.A1(new_n1684), .A2(new_n873), .B(new_n1687), .C(\a[14] ), .Y(new_n1688));
  O2A1O1Ixp33_ASAP7_75t_L   g01432(.A1(new_n872), .A2(new_n540), .B(new_n1686), .C(\a[14] ), .Y(new_n1689));
  AOI21xp33_ASAP7_75t_L     g01433(.A1(new_n1688), .A2(\a[14] ), .B(new_n1689), .Y(new_n1690));
  AND3x1_ASAP7_75t_L        g01434(.A(new_n1678), .B(new_n1683), .C(new_n1690), .Y(new_n1691));
  AOI21xp33_ASAP7_75t_L     g01435(.A1(new_n1678), .A2(new_n1683), .B(new_n1690), .Y(new_n1692));
  NOR3xp33_ASAP7_75t_L      g01436(.A(new_n1649), .B(new_n1691), .C(new_n1692), .Y(new_n1693));
  A2O1A1Ixp33_ASAP7_75t_L   g01437(.A1(new_n1543), .A2(new_n1422), .B(new_n1539), .C(new_n1538), .Y(new_n1694));
  NOR2xp33_ASAP7_75t_L      g01438(.A(new_n1692), .B(new_n1691), .Y(new_n1695));
  NOR2xp33_ASAP7_75t_L      g01439(.A(new_n1694), .B(new_n1695), .Y(new_n1696));
  OAI21xp33_ASAP7_75t_L     g01440(.A1(new_n1693), .A2(new_n1696), .B(new_n1648), .Y(new_n1697));
  A2O1A1Ixp33_ASAP7_75t_L   g01441(.A1(new_n1540), .A2(new_n1485), .B(new_n1548), .C(new_n1695), .Y(new_n1698));
  OAI21xp33_ASAP7_75t_L     g01442(.A1(new_n1691), .A2(new_n1692), .B(new_n1649), .Y(new_n1699));
  NAND3xp33_ASAP7_75t_L     g01443(.A(new_n1698), .B(new_n1647), .C(new_n1699), .Y(new_n1700));
  NAND3xp33_ASAP7_75t_L     g01444(.A(new_n1641), .B(new_n1697), .C(new_n1700), .Y(new_n1701));
  AND2x2_ASAP7_75t_L        g01445(.A(new_n1549), .B(new_n1541), .Y(new_n1702));
  INVx1_ASAP7_75t_L         g01446(.A(new_n1556), .Y(new_n1703));
  MAJIxp5_ASAP7_75t_L       g01447(.A(new_n1559), .B(new_n1703), .C(new_n1702), .Y(new_n1704));
  AOI21xp33_ASAP7_75t_L     g01448(.A1(new_n1698), .A2(new_n1699), .B(new_n1647), .Y(new_n1705));
  NOR3xp33_ASAP7_75t_L      g01449(.A(new_n1696), .B(new_n1693), .C(new_n1648), .Y(new_n1706));
  OAI21xp33_ASAP7_75t_L     g01450(.A1(new_n1706), .A2(new_n1705), .B(new_n1704), .Y(new_n1707));
  NOR2xp33_ASAP7_75t_L      g01451(.A(new_n936), .B(new_n513), .Y(new_n1708));
  AOI221xp5_ASAP7_75t_L     g01452(.A1(\b[12] ), .A2(new_n560), .B1(\b[14] ), .B2(new_n475), .C(new_n1708), .Y(new_n1709));
  INVx1_ASAP7_75t_L         g01453(.A(new_n1709), .Y(new_n1710));
  A2O1A1Ixp33_ASAP7_75t_L   g01454(.A1(new_n971), .A2(new_n483), .B(new_n1710), .C(\a[8] ), .Y(new_n1711));
  O2A1O1Ixp33_ASAP7_75t_L   g01455(.A1(new_n477), .A2(new_n1268), .B(new_n1709), .C(\a[8] ), .Y(new_n1712));
  AOI21xp33_ASAP7_75t_L     g01456(.A1(new_n1711), .A2(\a[8] ), .B(new_n1712), .Y(new_n1713));
  NAND3xp33_ASAP7_75t_L     g01457(.A(new_n1701), .B(new_n1707), .C(new_n1713), .Y(new_n1714));
  NOR3xp33_ASAP7_75t_L      g01458(.A(new_n1704), .B(new_n1705), .C(new_n1706), .Y(new_n1715));
  AOI21xp33_ASAP7_75t_L     g01459(.A1(new_n1700), .A2(new_n1697), .B(new_n1641), .Y(new_n1716));
  O2A1O1Ixp33_ASAP7_75t_L   g01460(.A1(new_n477), .A2(new_n1268), .B(new_n1709), .C(new_n466), .Y(new_n1717));
  A2O1A1Ixp33_ASAP7_75t_L   g01461(.A1(new_n971), .A2(new_n483), .B(new_n1710), .C(new_n466), .Y(new_n1718));
  OAI21xp33_ASAP7_75t_L     g01462(.A1(new_n466), .A2(new_n1717), .B(new_n1718), .Y(new_n1719));
  OAI21xp33_ASAP7_75t_L     g01463(.A1(new_n1716), .A2(new_n1715), .B(new_n1719), .Y(new_n1720));
  NAND2xp33_ASAP7_75t_L     g01464(.A(new_n1714), .B(new_n1720), .Y(new_n1721));
  A2O1A1Ixp33_ASAP7_75t_L   g01465(.A1(new_n1577), .A2(new_n1571), .B(new_n1639), .C(new_n1721), .Y(new_n1722));
  A2O1A1O1Ixp25_ASAP7_75t_L g01466(.A1(new_n1440), .A2(new_n1439), .B(new_n1436), .C(new_n1571), .D(new_n1639), .Y(new_n1723));
  NAND3xp33_ASAP7_75t_L     g01467(.A(new_n1723), .B(new_n1720), .C(new_n1714), .Y(new_n1724));
  AOI21xp33_ASAP7_75t_L     g01468(.A1(new_n1724), .A2(new_n1722), .B(new_n1638), .Y(new_n1725));
  INVx1_ASAP7_75t_L         g01469(.A(new_n1637), .Y(new_n1726));
  A2O1A1Ixp33_ASAP7_75t_L   g01470(.A1(new_n1633), .A2(new_n359), .B(new_n1635), .C(new_n346), .Y(new_n1727));
  NAND2xp33_ASAP7_75t_L     g01471(.A(new_n1727), .B(new_n1726), .Y(new_n1728));
  AOI21xp33_ASAP7_75t_L     g01472(.A1(new_n1720), .A2(new_n1714), .B(new_n1723), .Y(new_n1729));
  OAI21xp33_ASAP7_75t_L     g01473(.A1(new_n1579), .A2(new_n1580), .B(new_n1576), .Y(new_n1730));
  NOR2xp33_ASAP7_75t_L      g01474(.A(new_n1721), .B(new_n1730), .Y(new_n1731));
  NOR3xp33_ASAP7_75t_L      g01475(.A(new_n1729), .B(new_n1731), .C(new_n1728), .Y(new_n1732));
  NOR2xp33_ASAP7_75t_L      g01476(.A(new_n1732), .B(new_n1725), .Y(new_n1733));
  A2O1A1Ixp33_ASAP7_75t_L   g01477(.A1(new_n1592), .A2(new_n1612), .B(new_n1631), .C(new_n1733), .Y(new_n1734));
  A2O1A1O1Ixp25_ASAP7_75t_L g01478(.A1(new_n1373), .A2(new_n1445), .B(new_n1443), .C(new_n1592), .D(new_n1631), .Y(new_n1735));
  OAI21xp33_ASAP7_75t_L     g01479(.A1(new_n1731), .A2(new_n1729), .B(new_n1728), .Y(new_n1736));
  NAND3xp33_ASAP7_75t_L     g01480(.A(new_n1724), .B(new_n1722), .C(new_n1638), .Y(new_n1737));
  NAND2xp33_ASAP7_75t_L     g01481(.A(new_n1737), .B(new_n1736), .Y(new_n1738));
  NAND2xp33_ASAP7_75t_L     g01482(.A(new_n1738), .B(new_n1735), .Y(new_n1739));
  NOR2xp33_ASAP7_75t_L      g01483(.A(new_n1458), .B(new_n287), .Y(new_n1740));
  AOI221xp5_ASAP7_75t_L     g01484(.A1(\b[19] ), .A2(new_n264), .B1(\b[20] ), .B2(new_n283), .C(new_n1740), .Y(new_n1741));
  INVx1_ASAP7_75t_L         g01485(.A(new_n1459), .Y(new_n1742));
  INVx1_ASAP7_75t_L         g01486(.A(new_n1600), .Y(new_n1743));
  NOR2xp33_ASAP7_75t_L      g01487(.A(\b[19] ), .B(\b[20] ), .Y(new_n1744));
  INVx1_ASAP7_75t_L         g01488(.A(\b[20] ), .Y(new_n1745));
  NOR2xp33_ASAP7_75t_L      g01489(.A(new_n1599), .B(new_n1745), .Y(new_n1746));
  NOR2xp33_ASAP7_75t_L      g01490(.A(new_n1744), .B(new_n1746), .Y(new_n1747));
  INVx1_ASAP7_75t_L         g01491(.A(new_n1747), .Y(new_n1748));
  A2O1A1O1Ixp25_ASAP7_75t_L g01492(.A1(new_n1742), .A2(new_n1461), .B(new_n1598), .C(new_n1743), .D(new_n1748), .Y(new_n1749));
  A2O1A1Ixp33_ASAP7_75t_L   g01493(.A1(new_n1461), .A2(new_n1742), .B(new_n1598), .C(new_n1743), .Y(new_n1750));
  NOR2xp33_ASAP7_75t_L      g01494(.A(new_n1747), .B(new_n1750), .Y(new_n1751));
  NOR2xp33_ASAP7_75t_L      g01495(.A(new_n1749), .B(new_n1751), .Y(new_n1752));
  NAND2xp33_ASAP7_75t_L     g01496(.A(new_n273), .B(new_n1752), .Y(new_n1753));
  OR2x4_ASAP7_75t_L         g01497(.A(new_n1749), .B(new_n1751), .Y(new_n1754));
  O2A1O1Ixp33_ASAP7_75t_L   g01498(.A1(new_n279), .A2(new_n1754), .B(new_n1741), .C(new_n257), .Y(new_n1755));
  OAI211xp5_ASAP7_75t_L     g01499(.A1(new_n279), .A2(new_n1754), .B(new_n1741), .C(\a[2] ), .Y(new_n1756));
  A2O1A1Ixp33_ASAP7_75t_L   g01500(.A1(new_n1753), .A2(new_n1741), .B(new_n1755), .C(new_n1756), .Y(new_n1757));
  AOI21xp33_ASAP7_75t_L     g01501(.A1(new_n1734), .A2(new_n1739), .B(new_n1757), .Y(new_n1758));
  O2A1O1Ixp33_ASAP7_75t_L   g01502(.A1(new_n1586), .A2(new_n1588), .B(new_n1582), .C(new_n1738), .Y(new_n1759));
  OAI21xp33_ASAP7_75t_L     g01503(.A1(new_n1586), .A2(new_n1588), .B(new_n1582), .Y(new_n1760));
  NOR2xp33_ASAP7_75t_L      g01504(.A(new_n1733), .B(new_n1760), .Y(new_n1761));
  OAI21xp33_ASAP7_75t_L     g01505(.A1(new_n279), .A2(new_n1754), .B(new_n1741), .Y(new_n1762));
  NAND2xp33_ASAP7_75t_L     g01506(.A(new_n257), .B(new_n1762), .Y(new_n1763));
  AOI211xp5_ASAP7_75t_L     g01507(.A1(new_n1763), .A2(new_n1756), .B(new_n1759), .C(new_n1761), .Y(new_n1764));
  NOR2xp33_ASAP7_75t_L      g01508(.A(new_n1758), .B(new_n1764), .Y(new_n1765));
  A2O1A1O1Ixp25_ASAP7_75t_L g01509(.A1(new_n1617), .A2(new_n1594), .B(new_n1620), .C(new_n1630), .D(new_n1765), .Y(new_n1766));
  A2O1A1O1Ixp25_ASAP7_75t_L g01510(.A1(new_n1471), .A2(new_n1475), .B(new_n1619), .C(new_n1623), .D(new_n1611), .Y(new_n1767));
  AND2x2_ASAP7_75t_L        g01511(.A(new_n1765), .B(new_n1767), .Y(new_n1768));
  NOR2xp33_ASAP7_75t_L      g01512(.A(new_n1766), .B(new_n1768), .Y(\f[20] ));
  O2A1O1Ixp33_ASAP7_75t_L   g01513(.A1(new_n1586), .A2(new_n1588), .B(new_n1582), .C(new_n1733), .Y(new_n1770));
  A2O1A1Ixp33_ASAP7_75t_L   g01514(.A1(new_n1737), .A2(new_n1736), .B(new_n1770), .C(new_n1734), .Y(new_n1771));
  NAND2xp33_ASAP7_75t_L     g01515(.A(new_n1707), .B(new_n1701), .Y(new_n1772));
  INVx1_ASAP7_75t_L         g01516(.A(new_n1051), .Y(new_n1773));
  NAND2xp33_ASAP7_75t_L     g01517(.A(new_n1049), .B(new_n1773), .Y(new_n1774));
  NOR2xp33_ASAP7_75t_L      g01518(.A(new_n960), .B(new_n513), .Y(new_n1775));
  AOI221xp5_ASAP7_75t_L     g01519(.A1(\b[13] ), .A2(new_n560), .B1(\b[15] ), .B2(new_n475), .C(new_n1775), .Y(new_n1776));
  O2A1O1Ixp33_ASAP7_75t_L   g01520(.A1(new_n477), .A2(new_n1774), .B(new_n1776), .C(new_n466), .Y(new_n1777));
  INVx1_ASAP7_75t_L         g01521(.A(new_n1776), .Y(new_n1778));
  A2O1A1Ixp33_ASAP7_75t_L   g01522(.A1(new_n1052), .A2(new_n483), .B(new_n1778), .C(new_n466), .Y(new_n1779));
  OAI21xp33_ASAP7_75t_L     g01523(.A1(new_n466), .A2(new_n1777), .B(new_n1779), .Y(new_n1780));
  NOR2xp33_ASAP7_75t_L      g01524(.A(new_n748), .B(new_n1550), .Y(new_n1781));
  AOI221xp5_ASAP7_75t_L     g01525(.A1(\b[10] ), .A2(new_n713), .B1(\b[12] ), .B2(new_n640), .C(new_n1781), .Y(new_n1782));
  INVx1_ASAP7_75t_L         g01526(.A(new_n1782), .Y(new_n1783));
  A2O1A1Ixp33_ASAP7_75t_L   g01527(.A1(new_n1057), .A2(new_n718), .B(new_n1783), .C(\a[11] ), .Y(new_n1784));
  O2A1O1Ixp33_ASAP7_75t_L   g01528(.A1(new_n641), .A2(new_n841), .B(new_n1782), .C(\a[11] ), .Y(new_n1785));
  AOI21xp33_ASAP7_75t_L     g01529(.A1(new_n1784), .A2(\a[11] ), .B(new_n1785), .Y(new_n1786));
  NAND3xp33_ASAP7_75t_L     g01530(.A(new_n1678), .B(new_n1683), .C(new_n1690), .Y(new_n1787));
  A2O1A1O1Ixp25_ASAP7_75t_L g01531(.A1(new_n1540), .A2(new_n1485), .B(new_n1548), .C(new_n1787), .D(new_n1692), .Y(new_n1788));
  A2O1A1O1Ixp25_ASAP7_75t_L g01532(.A1(new_n1535), .A2(new_n1536), .B(new_n1534), .C(new_n1680), .D(new_n1677), .Y(new_n1789));
  INVx1_ASAP7_75t_L         g01533(.A(\a[21] ), .Y(new_n1790));
  NAND2xp33_ASAP7_75t_L     g01534(.A(\a[20] ), .B(new_n1790), .Y(new_n1791));
  NAND2xp33_ASAP7_75t_L     g01535(.A(\a[21] ), .B(new_n1501), .Y(new_n1792));
  AND2x2_ASAP7_75t_L        g01536(.A(new_n1791), .B(new_n1792), .Y(new_n1793));
  NOR2xp33_ASAP7_75t_L      g01537(.A(new_n284), .B(new_n1793), .Y(new_n1794));
  INVx1_ASAP7_75t_L         g01538(.A(new_n1794), .Y(new_n1795));
  A2O1A1O1Ixp25_ASAP7_75t_L g01539(.A1(\a[20] ), .A2(new_n1657), .B(new_n1661), .C(new_n1516), .D(new_n1795), .Y(new_n1796));
  NOR2xp33_ASAP7_75t_L      g01540(.A(new_n1794), .B(new_n1676), .Y(new_n1797));
  NAND2xp33_ASAP7_75t_L     g01541(.A(\b[3] ), .B(new_n1511), .Y(new_n1798));
  NAND2xp33_ASAP7_75t_L     g01542(.A(\b[1] ), .B(new_n1659), .Y(new_n1799));
  NAND2xp33_ASAP7_75t_L     g01543(.A(\b[2] ), .B(new_n1507), .Y(new_n1800));
  NAND2xp33_ASAP7_75t_L     g01544(.A(new_n1513), .B(new_n312), .Y(new_n1801));
  NAND5xp2_ASAP7_75t_L      g01545(.A(new_n1801), .B(new_n1800), .C(new_n1799), .D(new_n1798), .E(\a[20] ), .Y(new_n1802));
  OAI211xp5_ASAP7_75t_L     g01546(.A1(new_n1654), .A2(new_n262), .B(new_n1798), .C(new_n1800), .Y(new_n1803));
  A2O1A1Ixp33_ASAP7_75t_L   g01547(.A1(new_n312), .A2(new_n1513), .B(new_n1803), .C(new_n1501), .Y(new_n1804));
  NAND2xp33_ASAP7_75t_L     g01548(.A(new_n1802), .B(new_n1804), .Y(new_n1805));
  OAI21xp33_ASAP7_75t_L     g01549(.A1(new_n1797), .A2(new_n1796), .B(new_n1805), .Y(new_n1806));
  A2O1A1Ixp33_ASAP7_75t_L   g01550(.A1(new_n1673), .A2(new_n1674), .B(new_n1528), .C(new_n1794), .Y(new_n1807));
  NAND2xp33_ASAP7_75t_L     g01551(.A(new_n1795), .B(new_n1664), .Y(new_n1808));
  AND2x2_ASAP7_75t_L        g01552(.A(new_n1802), .B(new_n1804), .Y(new_n1809));
  NAND3xp33_ASAP7_75t_L     g01553(.A(new_n1808), .B(new_n1809), .C(new_n1807), .Y(new_n1810));
  NOR2xp33_ASAP7_75t_L      g01554(.A(new_n427), .B(new_n1284), .Y(new_n1811));
  AOI221xp5_ASAP7_75t_L     g01555(.A1(\b[4] ), .A2(new_n1290), .B1(\b[5] ), .B2(new_n1204), .C(new_n1811), .Y(new_n1812));
  O2A1O1Ixp33_ASAP7_75t_L   g01556(.A1(new_n1210), .A2(new_n434), .B(new_n1812), .C(new_n1206), .Y(new_n1813));
  OAI31xp33_ASAP7_75t_L     g01557(.A1(new_n433), .A2(new_n431), .A3(new_n1210), .B(new_n1812), .Y(new_n1814));
  NAND2xp33_ASAP7_75t_L     g01558(.A(new_n1206), .B(new_n1814), .Y(new_n1815));
  OA21x2_ASAP7_75t_L        g01559(.A1(new_n1206), .A2(new_n1813), .B(new_n1815), .Y(new_n1816));
  NAND3xp33_ASAP7_75t_L     g01560(.A(new_n1806), .B(new_n1816), .C(new_n1810), .Y(new_n1817));
  AOI21xp33_ASAP7_75t_L     g01561(.A1(new_n1808), .A2(new_n1807), .B(new_n1809), .Y(new_n1818));
  NOR3xp33_ASAP7_75t_L      g01562(.A(new_n1796), .B(new_n1797), .C(new_n1805), .Y(new_n1819));
  OAI21xp33_ASAP7_75t_L     g01563(.A1(new_n1206), .A2(new_n1813), .B(new_n1815), .Y(new_n1820));
  OAI21xp33_ASAP7_75t_L     g01564(.A1(new_n1818), .A2(new_n1819), .B(new_n1820), .Y(new_n1821));
  OAI211xp5_ASAP7_75t_L     g01565(.A1(new_n1671), .A2(new_n1789), .B(new_n1817), .C(new_n1821), .Y(new_n1822));
  A2O1A1O1Ixp25_ASAP7_75t_L g01566(.A1(new_n1492), .A2(new_n1546), .B(new_n1653), .C(new_n1682), .D(new_n1671), .Y(new_n1823));
  NAND3xp33_ASAP7_75t_L     g01567(.A(new_n1806), .B(new_n1810), .C(new_n1820), .Y(new_n1824));
  NOR3xp33_ASAP7_75t_L      g01568(.A(new_n1819), .B(new_n1818), .C(new_n1820), .Y(new_n1825));
  A2O1A1Ixp33_ASAP7_75t_L   g01569(.A1(new_n1820), .A2(new_n1824), .B(new_n1825), .C(new_n1823), .Y(new_n1826));
  NOR2xp33_ASAP7_75t_L      g01570(.A(new_n534), .B(new_n864), .Y(new_n1827));
  AOI221xp5_ASAP7_75t_L     g01571(.A1(\b[7] ), .A2(new_n985), .B1(\b[9] ), .B2(new_n886), .C(new_n1827), .Y(new_n1828));
  INVx1_ASAP7_75t_L         g01572(.A(new_n1828), .Y(new_n1829));
  A2O1A1Ixp33_ASAP7_75t_L   g01573(.A1(new_n602), .A2(new_n873), .B(new_n1829), .C(\a[14] ), .Y(new_n1830));
  NAND2xp33_ASAP7_75t_L     g01574(.A(\a[14] ), .B(new_n1830), .Y(new_n1831));
  A2O1A1Ixp33_ASAP7_75t_L   g01575(.A1(new_n602), .A2(new_n873), .B(new_n1829), .C(new_n867), .Y(new_n1832));
  AOI22xp33_ASAP7_75t_L     g01576(.A1(new_n1831), .A2(new_n1832), .B1(new_n1822), .B2(new_n1826), .Y(new_n1833));
  AOI21xp33_ASAP7_75t_L     g01577(.A1(new_n1806), .A2(new_n1810), .B(new_n1816), .Y(new_n1834));
  NOR3xp33_ASAP7_75t_L      g01578(.A(new_n1823), .B(new_n1825), .C(new_n1834), .Y(new_n1835));
  AOI211xp5_ASAP7_75t_L     g01579(.A1(new_n1821), .A2(new_n1817), .B(new_n1671), .C(new_n1789), .Y(new_n1836));
  O2A1O1Ixp33_ASAP7_75t_L   g01580(.A1(new_n872), .A2(new_n1066), .B(new_n1828), .C(new_n867), .Y(new_n1837));
  OAI21xp33_ASAP7_75t_L     g01581(.A1(new_n867), .A2(new_n1837), .B(new_n1832), .Y(new_n1838));
  NOR3xp33_ASAP7_75t_L      g01582(.A(new_n1835), .B(new_n1836), .C(new_n1838), .Y(new_n1839));
  NOR3xp33_ASAP7_75t_L      g01583(.A(new_n1788), .B(new_n1833), .C(new_n1839), .Y(new_n1840));
  OAI21xp33_ASAP7_75t_L     g01584(.A1(new_n1836), .A2(new_n1835), .B(new_n1838), .Y(new_n1841));
  NAND4xp25_ASAP7_75t_L     g01585(.A(new_n1826), .B(new_n1822), .C(new_n1831), .D(new_n1832), .Y(new_n1842));
  AOI221xp5_ASAP7_75t_L     g01586(.A1(new_n1694), .A2(new_n1787), .B1(new_n1842), .B2(new_n1841), .C(new_n1692), .Y(new_n1843));
  OA21x2_ASAP7_75t_L        g01587(.A1(new_n1843), .A2(new_n1840), .B(new_n1786), .Y(new_n1844));
  NOR3xp33_ASAP7_75t_L      g01588(.A(new_n1786), .B(new_n1840), .C(new_n1843), .Y(new_n1845));
  NOR2xp33_ASAP7_75t_L      g01589(.A(new_n1845), .B(new_n1844), .Y(new_n1846));
  A2O1A1Ixp33_ASAP7_75t_L   g01590(.A1(new_n1697), .A2(new_n1641), .B(new_n1706), .C(new_n1846), .Y(new_n1847));
  INVx1_ASAP7_75t_L         g01591(.A(new_n1555), .Y(new_n1848));
  O2A1O1Ixp33_ASAP7_75t_L   g01592(.A1(new_n1553), .A2(new_n637), .B(new_n1848), .C(new_n1640), .Y(new_n1849));
  NAND2xp33_ASAP7_75t_L     g01593(.A(new_n1561), .B(new_n1562), .Y(new_n1850));
  A2O1A1O1Ixp25_ASAP7_75t_L g01594(.A1(new_n1559), .A2(new_n1850), .B(new_n1849), .C(new_n1697), .D(new_n1706), .Y(new_n1851));
  OAI21xp33_ASAP7_75t_L     g01595(.A1(new_n1844), .A2(new_n1845), .B(new_n1851), .Y(new_n1852));
  NAND3xp33_ASAP7_75t_L     g01596(.A(new_n1847), .B(new_n1780), .C(new_n1852), .Y(new_n1853));
  A2O1A1Ixp33_ASAP7_75t_L   g01597(.A1(new_n1052), .A2(new_n483), .B(new_n1778), .C(\a[8] ), .Y(new_n1854));
  O2A1O1Ixp33_ASAP7_75t_L   g01598(.A1(new_n477), .A2(new_n1774), .B(new_n1776), .C(\a[8] ), .Y(new_n1855));
  AOI21xp33_ASAP7_75t_L     g01599(.A1(new_n1854), .A2(\a[8] ), .B(new_n1855), .Y(new_n1856));
  NOR3xp33_ASAP7_75t_L      g01600(.A(new_n1851), .B(new_n1844), .C(new_n1845), .Y(new_n1857));
  A2O1A1Ixp33_ASAP7_75t_L   g01601(.A1(\a[11] ), .A2(new_n1554), .B(new_n1555), .C(new_n1702), .Y(new_n1858));
  A2O1A1Ixp33_ASAP7_75t_L   g01602(.A1(new_n1573), .A2(new_n1858), .B(new_n1705), .C(new_n1700), .Y(new_n1859));
  NOR2xp33_ASAP7_75t_L      g01603(.A(new_n1859), .B(new_n1846), .Y(new_n1860));
  OAI21xp33_ASAP7_75t_L     g01604(.A1(new_n1857), .A2(new_n1860), .B(new_n1856), .Y(new_n1861));
  NAND2xp33_ASAP7_75t_L     g01605(.A(new_n1861), .B(new_n1853), .Y(new_n1862));
  O2A1O1Ixp33_ASAP7_75t_L   g01606(.A1(new_n1772), .A2(new_n1713), .B(new_n1722), .C(new_n1862), .Y(new_n1863));
  NOR2xp33_ASAP7_75t_L      g01607(.A(new_n1716), .B(new_n1715), .Y(new_n1864));
  A2O1A1Ixp33_ASAP7_75t_L   g01608(.A1(\a[8] ), .A2(new_n1711), .B(new_n1712), .C(new_n1864), .Y(new_n1865));
  A2O1A1Ixp33_ASAP7_75t_L   g01609(.A1(new_n1713), .A2(new_n1714), .B(new_n1723), .C(new_n1865), .Y(new_n1866));
  AND2x2_ASAP7_75t_L        g01610(.A(new_n1861), .B(new_n1853), .Y(new_n1867));
  NOR2xp33_ASAP7_75t_L      g01611(.A(new_n1866), .B(new_n1867), .Y(new_n1868));
  NOR2xp33_ASAP7_75t_L      g01612(.A(new_n1150), .B(new_n375), .Y(new_n1869));
  AOI221xp5_ASAP7_75t_L     g01613(.A1(\b[18] ), .A2(new_n361), .B1(new_n349), .B2(\b[17] ), .C(new_n1869), .Y(new_n1870));
  O2A1O1Ixp33_ASAP7_75t_L   g01614(.A1(new_n356), .A2(new_n1464), .B(new_n1870), .C(new_n346), .Y(new_n1871));
  O2A1O1Ixp33_ASAP7_75t_L   g01615(.A1(new_n356), .A2(new_n1464), .B(new_n1870), .C(\a[5] ), .Y(new_n1872));
  INVx1_ASAP7_75t_L         g01616(.A(new_n1872), .Y(new_n1873));
  OAI21xp33_ASAP7_75t_L     g01617(.A1(new_n346), .A2(new_n1871), .B(new_n1873), .Y(new_n1874));
  NOR3xp33_ASAP7_75t_L      g01618(.A(new_n1868), .B(new_n1863), .C(new_n1874), .Y(new_n1875));
  NAND2xp33_ASAP7_75t_L     g01619(.A(new_n1866), .B(new_n1867), .Y(new_n1876));
  O2A1O1Ixp33_ASAP7_75t_L   g01620(.A1(new_n1717), .A2(new_n466), .B(new_n1718), .C(new_n1772), .Y(new_n1877));
  A2O1A1O1Ixp25_ASAP7_75t_L g01621(.A1(new_n1571), .A2(new_n1577), .B(new_n1639), .C(new_n1721), .D(new_n1877), .Y(new_n1878));
  NAND2xp33_ASAP7_75t_L     g01622(.A(new_n1862), .B(new_n1878), .Y(new_n1879));
  OAI21xp33_ASAP7_75t_L     g01623(.A1(new_n356), .A2(new_n1464), .B(new_n1870), .Y(new_n1880));
  NOR2xp33_ASAP7_75t_L      g01624(.A(new_n346), .B(new_n1880), .Y(new_n1881));
  NOR2xp33_ASAP7_75t_L      g01625(.A(new_n1872), .B(new_n1881), .Y(new_n1882));
  AOI21xp33_ASAP7_75t_L     g01626(.A1(new_n1876), .A2(new_n1879), .B(new_n1882), .Y(new_n1883));
  NOR2xp33_ASAP7_75t_L      g01627(.A(new_n1883), .B(new_n1875), .Y(new_n1884));
  NOR3xp33_ASAP7_75t_L      g01628(.A(new_n1729), .B(new_n1731), .C(new_n1638), .Y(new_n1885));
  A2O1A1O1Ixp25_ASAP7_75t_L g01629(.A1(new_n1592), .A2(new_n1612), .B(new_n1631), .C(new_n1738), .D(new_n1885), .Y(new_n1886));
  NAND2xp33_ASAP7_75t_L     g01630(.A(new_n1884), .B(new_n1886), .Y(new_n1887));
  NAND3xp33_ASAP7_75t_L     g01631(.A(new_n1876), .B(new_n1879), .C(new_n1882), .Y(new_n1888));
  OAI21xp33_ASAP7_75t_L     g01632(.A1(new_n1863), .A2(new_n1868), .B(new_n1874), .Y(new_n1889));
  NAND2xp33_ASAP7_75t_L     g01633(.A(new_n1888), .B(new_n1889), .Y(new_n1890));
  A2O1A1Ixp33_ASAP7_75t_L   g01634(.A1(new_n1738), .A2(new_n1760), .B(new_n1885), .C(new_n1890), .Y(new_n1891));
  NOR2xp33_ASAP7_75t_L      g01635(.A(new_n1599), .B(new_n287), .Y(new_n1892));
  AOI221xp5_ASAP7_75t_L     g01636(.A1(\b[20] ), .A2(new_n264), .B1(\b[21] ), .B2(new_n283), .C(new_n1892), .Y(new_n1893));
  NOR2xp33_ASAP7_75t_L      g01637(.A(\b[20] ), .B(\b[21] ), .Y(new_n1894));
  INVx1_ASAP7_75t_L         g01638(.A(\b[21] ), .Y(new_n1895));
  NOR2xp33_ASAP7_75t_L      g01639(.A(new_n1745), .B(new_n1895), .Y(new_n1896));
  NOR2xp33_ASAP7_75t_L      g01640(.A(new_n1894), .B(new_n1896), .Y(new_n1897));
  A2O1A1Ixp33_ASAP7_75t_L   g01641(.A1(new_n1750), .A2(new_n1747), .B(new_n1746), .C(new_n1897), .Y(new_n1898));
  O2A1O1Ixp33_ASAP7_75t_L   g01642(.A1(new_n1600), .A2(new_n1603), .B(new_n1747), .C(new_n1746), .Y(new_n1899));
  OAI21xp33_ASAP7_75t_L     g01643(.A1(new_n1894), .A2(new_n1896), .B(new_n1899), .Y(new_n1900));
  NAND2xp33_ASAP7_75t_L     g01644(.A(new_n1898), .B(new_n1900), .Y(new_n1901));
  O2A1O1Ixp33_ASAP7_75t_L   g01645(.A1(new_n279), .A2(new_n1901), .B(new_n1893), .C(new_n257), .Y(new_n1902));
  OAI21xp33_ASAP7_75t_L     g01646(.A1(new_n279), .A2(new_n1901), .B(new_n1893), .Y(new_n1903));
  NAND2xp33_ASAP7_75t_L     g01647(.A(new_n257), .B(new_n1903), .Y(new_n1904));
  OAI21xp33_ASAP7_75t_L     g01648(.A1(new_n257), .A2(new_n1902), .B(new_n1904), .Y(new_n1905));
  INVx1_ASAP7_75t_L         g01649(.A(new_n1905), .Y(new_n1906));
  NAND3xp33_ASAP7_75t_L     g01650(.A(new_n1891), .B(new_n1887), .C(new_n1906), .Y(new_n1907));
  NOR2xp33_ASAP7_75t_L      g01651(.A(new_n1731), .B(new_n1729), .Y(new_n1908));
  NAND2xp33_ASAP7_75t_L     g01652(.A(new_n1728), .B(new_n1908), .Y(new_n1909));
  A2O1A1Ixp33_ASAP7_75t_L   g01653(.A1(new_n1593), .A2(new_n1582), .B(new_n1733), .C(new_n1909), .Y(new_n1910));
  NOR2xp33_ASAP7_75t_L      g01654(.A(new_n1890), .B(new_n1910), .Y(new_n1911));
  O2A1O1Ixp33_ASAP7_75t_L   g01655(.A1(new_n1735), .A2(new_n1733), .B(new_n1909), .C(new_n1884), .Y(new_n1912));
  OAI21xp33_ASAP7_75t_L     g01656(.A1(new_n1911), .A2(new_n1912), .B(new_n1905), .Y(new_n1913));
  NAND2xp33_ASAP7_75t_L     g01657(.A(new_n1907), .B(new_n1913), .Y(new_n1914));
  A2O1A1Ixp33_ASAP7_75t_L   g01658(.A1(new_n1757), .A2(new_n1771), .B(new_n1766), .C(new_n1914), .Y(new_n1915));
  INVx1_ASAP7_75t_L         g01659(.A(new_n1915), .Y(new_n1916));
  A2O1A1Ixp33_ASAP7_75t_L   g01660(.A1(new_n1592), .A2(new_n1612), .B(new_n1631), .C(new_n1738), .Y(new_n1917));
  A2O1A1Ixp33_ASAP7_75t_L   g01661(.A1(new_n1917), .A2(new_n1760), .B(new_n1761), .C(new_n1757), .Y(new_n1918));
  OAI21xp33_ASAP7_75t_L     g01662(.A1(new_n1765), .A2(new_n1767), .B(new_n1918), .Y(new_n1919));
  NOR2xp33_ASAP7_75t_L      g01663(.A(new_n1914), .B(new_n1919), .Y(new_n1920));
  NOR2xp33_ASAP7_75t_L      g01664(.A(new_n1920), .B(new_n1916), .Y(\f[21] ));
  NAND2xp33_ASAP7_75t_L     g01665(.A(new_n1891), .B(new_n1887), .Y(new_n1922));
  NOR3xp33_ASAP7_75t_L      g01666(.A(new_n1860), .B(new_n1857), .C(new_n1856), .Y(new_n1923));
  A2O1A1O1Ixp25_ASAP7_75t_L g01667(.A1(new_n1721), .A2(new_n1730), .B(new_n1877), .C(new_n1861), .D(new_n1923), .Y(new_n1924));
  OAI22xp33_ASAP7_75t_L     g01668(.A1(new_n513), .A2(new_n1043), .B1(new_n960), .B2(new_n506), .Y(new_n1925));
  AOI221xp5_ASAP7_75t_L     g01669(.A1(new_n475), .A2(\b[16] ), .B1(new_n483), .B2(new_n1156), .C(new_n1925), .Y(new_n1926));
  XNOR2x2_ASAP7_75t_L       g01670(.A(new_n466), .B(new_n1926), .Y(new_n1927));
  OAI21xp33_ASAP7_75t_L     g01671(.A1(new_n1843), .A2(new_n1840), .B(new_n1786), .Y(new_n1928));
  A2O1A1O1Ixp25_ASAP7_75t_L g01672(.A1(new_n1697), .A2(new_n1641), .B(new_n1706), .C(new_n1928), .D(new_n1845), .Y(new_n1929));
  OAI22xp33_ASAP7_75t_L     g01673(.A1(new_n1789), .A2(new_n1671), .B1(new_n1834), .B2(new_n1825), .Y(new_n1930));
  NOR2xp33_ASAP7_75t_L      g01674(.A(new_n448), .B(new_n1284), .Y(new_n1931));
  AOI221xp5_ASAP7_75t_L     g01675(.A1(\b[5] ), .A2(new_n1290), .B1(\b[6] ), .B2(new_n1204), .C(new_n1931), .Y(new_n1932));
  O2A1O1Ixp33_ASAP7_75t_L   g01676(.A1(new_n1210), .A2(new_n456), .B(new_n1932), .C(new_n1206), .Y(new_n1933));
  OAI21xp33_ASAP7_75t_L     g01677(.A1(new_n1210), .A2(new_n456), .B(new_n1932), .Y(new_n1934));
  NAND2xp33_ASAP7_75t_L     g01678(.A(new_n1206), .B(new_n1934), .Y(new_n1935));
  OAI21xp33_ASAP7_75t_L     g01679(.A1(new_n1206), .A2(new_n1933), .B(new_n1935), .Y(new_n1936));
  INVx1_ASAP7_75t_L         g01680(.A(new_n1936), .Y(new_n1937));
  MAJIxp5_ASAP7_75t_L       g01681(.A(new_n1805), .B(new_n1794), .C(new_n1664), .Y(new_n1938));
  NOR2xp33_ASAP7_75t_L      g01682(.A(new_n332), .B(new_n1518), .Y(new_n1939));
  AOI221xp5_ASAP7_75t_L     g01683(.A1(\b[2] ), .A2(new_n1659), .B1(\b[3] ), .B2(new_n1507), .C(new_n1939), .Y(new_n1940));
  OAI211xp5_ASAP7_75t_L     g01684(.A1(new_n1497), .A2(new_n1521), .B(new_n1940), .C(\a[20] ), .Y(new_n1941));
  NAND2xp33_ASAP7_75t_L     g01685(.A(\b[3] ), .B(new_n1507), .Y(new_n1942));
  OAI221xp5_ASAP7_75t_L     g01686(.A1(new_n1518), .A2(new_n332), .B1(new_n289), .B2(new_n1654), .C(new_n1942), .Y(new_n1943));
  A2O1A1Ixp33_ASAP7_75t_L   g01687(.A1(new_n342), .A2(new_n1513), .B(new_n1943), .C(new_n1501), .Y(new_n1944));
  NAND2xp33_ASAP7_75t_L     g01688(.A(new_n1792), .B(new_n1791), .Y(new_n1945));
  INVx1_ASAP7_75t_L         g01689(.A(\a[22] ), .Y(new_n1946));
  NOR2xp33_ASAP7_75t_L      g01690(.A(\a[21] ), .B(new_n1946), .Y(new_n1947));
  NOR2xp33_ASAP7_75t_L      g01691(.A(\a[22] ), .B(new_n1790), .Y(new_n1948));
  NOR2xp33_ASAP7_75t_L      g01692(.A(new_n1947), .B(new_n1948), .Y(new_n1949));
  NOR2xp33_ASAP7_75t_L      g01693(.A(new_n1945), .B(new_n1949), .Y(new_n1950));
  NAND2xp33_ASAP7_75t_L     g01694(.A(\a[23] ), .B(new_n1946), .Y(new_n1951));
  INVx1_ASAP7_75t_L         g01695(.A(\a[23] ), .Y(new_n1952));
  NAND2xp33_ASAP7_75t_L     g01696(.A(\a[22] ), .B(new_n1952), .Y(new_n1953));
  NAND2xp33_ASAP7_75t_L     g01697(.A(new_n1953), .B(new_n1951), .Y(new_n1954));
  NOR2xp33_ASAP7_75t_L      g01698(.A(new_n1954), .B(new_n1793), .Y(new_n1955));
  NAND2xp33_ASAP7_75t_L     g01699(.A(new_n1954), .B(new_n1945), .Y(new_n1956));
  NOR2xp33_ASAP7_75t_L      g01700(.A(new_n274), .B(new_n1956), .Y(new_n1957));
  AOI221xp5_ASAP7_75t_L     g01701(.A1(\b[1] ), .A2(new_n1955), .B1(new_n1950), .B2(\b[0] ), .C(new_n1957), .Y(new_n1958));
  NAND3xp33_ASAP7_75t_L     g01702(.A(new_n1958), .B(new_n1795), .C(\a[23] ), .Y(new_n1959));
  AOI22xp33_ASAP7_75t_L     g01703(.A1(new_n1950), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n1955), .Y(new_n1960));
  O2A1O1Ixp33_ASAP7_75t_L   g01704(.A1(new_n1956), .A2(new_n274), .B(new_n1960), .C(new_n1952), .Y(new_n1961));
  OAI21xp33_ASAP7_75t_L     g01705(.A1(new_n1947), .A2(new_n1948), .B(new_n1793), .Y(new_n1962));
  OAI32xp33_ASAP7_75t_L     g01706(.A1(new_n262), .A2(new_n1954), .A3(new_n1793), .B1(new_n1962), .B2(new_n284), .Y(new_n1963));
  AOI21xp33_ASAP7_75t_L     g01707(.A1(new_n1953), .A2(new_n1951), .B(new_n1793), .Y(new_n1964));
  A2O1A1Ixp33_ASAP7_75t_L   g01708(.A1(new_n1964), .A2(new_n275), .B(new_n1963), .C(new_n1952), .Y(new_n1965));
  A2O1A1Ixp33_ASAP7_75t_L   g01709(.A1(new_n1961), .A2(new_n1794), .B(new_n1952), .C(new_n1965), .Y(new_n1966));
  NAND4xp25_ASAP7_75t_L     g01710(.A(new_n1966), .B(new_n1941), .C(new_n1944), .D(new_n1959), .Y(new_n1967));
  AOI211xp5_ASAP7_75t_L     g01711(.A1(new_n342), .A2(new_n1513), .B(new_n1501), .C(new_n1943), .Y(new_n1968));
  O2A1O1Ixp33_ASAP7_75t_L   g01712(.A1(new_n1521), .A2(new_n1497), .B(new_n1940), .C(\a[20] ), .Y(new_n1969));
  NAND2xp33_ASAP7_75t_L     g01713(.A(new_n275), .B(new_n1964), .Y(new_n1970));
  NAND2xp33_ASAP7_75t_L     g01714(.A(new_n1970), .B(new_n1960), .Y(new_n1971));
  NOR3xp33_ASAP7_75t_L      g01715(.A(new_n1971), .B(new_n1794), .C(new_n1952), .Y(new_n1972));
  NAND2xp33_ASAP7_75t_L     g01716(.A(\b[0] ), .B(new_n1950), .Y(new_n1973));
  NAND2xp33_ASAP7_75t_L     g01717(.A(\b[1] ), .B(new_n1955), .Y(new_n1974));
  AND4x1_ASAP7_75t_L        g01718(.A(new_n1970), .B(new_n1974), .C(new_n1973), .D(\a[23] ), .Y(new_n1975));
  O2A1O1Ixp33_ASAP7_75t_L   g01719(.A1(new_n1956), .A2(new_n274), .B(new_n1960), .C(\a[23] ), .Y(new_n1976));
  AOI211xp5_ASAP7_75t_L     g01720(.A1(\a[23] ), .A2(new_n1795), .B(new_n1975), .C(new_n1976), .Y(new_n1977));
  OAI22xp33_ASAP7_75t_L     g01721(.A1(new_n1977), .A2(new_n1972), .B1(new_n1969), .B2(new_n1968), .Y(new_n1978));
  AOI21xp33_ASAP7_75t_L     g01722(.A1(new_n1978), .A2(new_n1967), .B(new_n1938), .Y(new_n1979));
  NAND3xp33_ASAP7_75t_L     g01723(.A(new_n1938), .B(new_n1967), .C(new_n1978), .Y(new_n1980));
  INVx1_ASAP7_75t_L         g01724(.A(new_n1980), .Y(new_n1981));
  NOR3xp33_ASAP7_75t_L      g01725(.A(new_n1981), .B(new_n1937), .C(new_n1979), .Y(new_n1982));
  MAJIxp5_ASAP7_75t_L       g01726(.A(new_n1809), .B(new_n1676), .C(new_n1795), .Y(new_n1983));
  NAND2xp33_ASAP7_75t_L     g01727(.A(new_n1967), .B(new_n1978), .Y(new_n1984));
  NAND2xp33_ASAP7_75t_L     g01728(.A(new_n1983), .B(new_n1984), .Y(new_n1985));
  AOI21xp33_ASAP7_75t_L     g01729(.A1(new_n1985), .A2(new_n1980), .B(new_n1936), .Y(new_n1986));
  AOI211xp5_ASAP7_75t_L     g01730(.A1(new_n1930), .A2(new_n1824), .B(new_n1982), .C(new_n1986), .Y(new_n1987));
  A2O1A1Ixp33_ASAP7_75t_L   g01731(.A1(new_n1817), .A2(new_n1821), .B(new_n1823), .C(new_n1824), .Y(new_n1988));
  NAND3xp33_ASAP7_75t_L     g01732(.A(new_n1985), .B(new_n1936), .C(new_n1980), .Y(new_n1989));
  OAI21xp33_ASAP7_75t_L     g01733(.A1(new_n1979), .A2(new_n1981), .B(new_n1937), .Y(new_n1990));
  AOI21xp33_ASAP7_75t_L     g01734(.A1(new_n1990), .A2(new_n1989), .B(new_n1988), .Y(new_n1991));
  NOR2xp33_ASAP7_75t_L      g01735(.A(new_n680), .B(new_n869), .Y(new_n1992));
  AOI221xp5_ASAP7_75t_L     g01736(.A1(\b[8] ), .A2(new_n985), .B1(\b[9] ), .B2(new_n885), .C(new_n1992), .Y(new_n1993));
  O2A1O1Ixp33_ASAP7_75t_L   g01737(.A1(new_n872), .A2(new_n1175), .B(new_n1993), .C(new_n867), .Y(new_n1994));
  OAI21xp33_ASAP7_75t_L     g01738(.A1(new_n872), .A2(new_n1175), .B(new_n1993), .Y(new_n1995));
  NAND2xp33_ASAP7_75t_L     g01739(.A(new_n867), .B(new_n1995), .Y(new_n1996));
  OAI21xp33_ASAP7_75t_L     g01740(.A1(new_n867), .A2(new_n1994), .B(new_n1996), .Y(new_n1997));
  NOR3xp33_ASAP7_75t_L      g01741(.A(new_n1987), .B(new_n1991), .C(new_n1997), .Y(new_n1998));
  NAND3xp33_ASAP7_75t_L     g01742(.A(new_n1988), .B(new_n1989), .C(new_n1990), .Y(new_n1999));
  OAI211xp5_ASAP7_75t_L     g01743(.A1(new_n1986), .A2(new_n1982), .B(new_n1930), .C(new_n1824), .Y(new_n2000));
  INVx1_ASAP7_75t_L         g01744(.A(new_n1997), .Y(new_n2001));
  AOI21xp33_ASAP7_75t_L     g01745(.A1(new_n1999), .A2(new_n2000), .B(new_n2001), .Y(new_n2002));
  OAI21xp33_ASAP7_75t_L     g01746(.A1(new_n1839), .A2(new_n1788), .B(new_n1841), .Y(new_n2003));
  NOR3xp33_ASAP7_75t_L      g01747(.A(new_n2003), .B(new_n2002), .C(new_n1998), .Y(new_n2004));
  NAND3xp33_ASAP7_75t_L     g01748(.A(new_n1999), .B(new_n2001), .C(new_n2000), .Y(new_n2005));
  OAI21xp33_ASAP7_75t_L     g01749(.A1(new_n1991), .A2(new_n1987), .B(new_n1997), .Y(new_n2006));
  A2O1A1O1Ixp25_ASAP7_75t_L g01750(.A1(new_n1787), .A2(new_n1694), .B(new_n1692), .C(new_n1842), .D(new_n1833), .Y(new_n2007));
  AOI21xp33_ASAP7_75t_L     g01751(.A1(new_n2006), .A2(new_n2005), .B(new_n2007), .Y(new_n2008));
  NOR2xp33_ASAP7_75t_L      g01752(.A(new_n833), .B(new_n1550), .Y(new_n2009));
  AOI221xp5_ASAP7_75t_L     g01753(.A1(\b[11] ), .A2(new_n713), .B1(\b[13] ), .B2(new_n640), .C(new_n2009), .Y(new_n2010));
  INVx1_ASAP7_75t_L         g01754(.A(new_n2010), .Y(new_n2011));
  A2O1A1Ixp33_ASAP7_75t_L   g01755(.A1(new_n1166), .A2(new_n718), .B(new_n2011), .C(\a[11] ), .Y(new_n2012));
  O2A1O1Ixp33_ASAP7_75t_L   g01756(.A1(new_n641), .A2(new_n942), .B(new_n2010), .C(\a[11] ), .Y(new_n2013));
  AOI21xp33_ASAP7_75t_L     g01757(.A1(new_n2012), .A2(\a[11] ), .B(new_n2013), .Y(new_n2014));
  OA21x2_ASAP7_75t_L        g01758(.A1(new_n2008), .A2(new_n2004), .B(new_n2014), .Y(new_n2015));
  NOR3xp33_ASAP7_75t_L      g01759(.A(new_n2004), .B(new_n2008), .C(new_n2014), .Y(new_n2016));
  NOR3xp33_ASAP7_75t_L      g01760(.A(new_n1929), .B(new_n2015), .C(new_n2016), .Y(new_n2017));
  OAI21xp33_ASAP7_75t_L     g01761(.A1(new_n2015), .A2(new_n2016), .B(new_n1929), .Y(new_n2018));
  INVx1_ASAP7_75t_L         g01762(.A(new_n2018), .Y(new_n2019));
  NOR3xp33_ASAP7_75t_L      g01763(.A(new_n1927), .B(new_n2017), .C(new_n2019), .Y(new_n2020));
  XNOR2x2_ASAP7_75t_L       g01764(.A(\a[8] ), .B(new_n1926), .Y(new_n2021));
  INVx1_ASAP7_75t_L         g01765(.A(new_n2017), .Y(new_n2022));
  AOI21xp33_ASAP7_75t_L     g01766(.A1(new_n2022), .A2(new_n2018), .B(new_n2021), .Y(new_n2023));
  NOR3xp33_ASAP7_75t_L      g01767(.A(new_n1924), .B(new_n2020), .C(new_n2023), .Y(new_n2024));
  NAND3xp33_ASAP7_75t_L     g01768(.A(new_n2021), .B(new_n2022), .C(new_n2018), .Y(new_n2025));
  OAI21xp33_ASAP7_75t_L     g01769(.A1(new_n2017), .A2(new_n2019), .B(new_n1927), .Y(new_n2026));
  AOI221xp5_ASAP7_75t_L     g01770(.A1(new_n1861), .A2(new_n1866), .B1(new_n2026), .B2(new_n2025), .C(new_n1923), .Y(new_n2027));
  OR2x4_ASAP7_75t_L         g01771(.A(new_n2024), .B(new_n2027), .Y(new_n2028));
  NOR2xp33_ASAP7_75t_L      g01772(.A(new_n1349), .B(new_n375), .Y(new_n2029));
  AOI221xp5_ASAP7_75t_L     g01773(.A1(\b[19] ), .A2(new_n361), .B1(new_n349), .B2(\b[18] ), .C(new_n2029), .Y(new_n2030));
  INVx1_ASAP7_75t_L         g01774(.A(new_n2030), .Y(new_n2031));
  A2O1A1Ixp33_ASAP7_75t_L   g01775(.A1(new_n1607), .A2(new_n359), .B(new_n2031), .C(\a[5] ), .Y(new_n2032));
  O2A1O1Ixp33_ASAP7_75t_L   g01776(.A1(new_n356), .A2(new_n1628), .B(new_n2030), .C(\a[5] ), .Y(new_n2033));
  AOI21xp33_ASAP7_75t_L     g01777(.A1(new_n2032), .A2(\a[5] ), .B(new_n2033), .Y(new_n2034));
  NOR3xp33_ASAP7_75t_L      g01778(.A(new_n2027), .B(new_n2024), .C(new_n2034), .Y(new_n2035));
  INVx1_ASAP7_75t_L         g01779(.A(new_n2034), .Y(new_n2036));
  OAI21xp33_ASAP7_75t_L     g01780(.A1(new_n2024), .A2(new_n2027), .B(new_n2036), .Y(new_n2037));
  OAI21xp33_ASAP7_75t_L     g01781(.A1(new_n2035), .A2(new_n2028), .B(new_n2037), .Y(new_n2038));
  NAND3xp33_ASAP7_75t_L     g01782(.A(new_n1876), .B(new_n1879), .C(new_n1874), .Y(new_n2039));
  A2O1A1Ixp33_ASAP7_75t_L   g01783(.A1(new_n1909), .A2(new_n1917), .B(new_n1884), .C(new_n2039), .Y(new_n2040));
  NOR2xp33_ASAP7_75t_L      g01784(.A(new_n2038), .B(new_n2040), .Y(new_n2041));
  INVx1_ASAP7_75t_L         g01785(.A(new_n2039), .Y(new_n2042));
  A2O1A1O1Ixp25_ASAP7_75t_L g01786(.A1(new_n1760), .A2(new_n1738), .B(new_n1885), .C(new_n1890), .D(new_n2042), .Y(new_n2043));
  O2A1O1Ixp33_ASAP7_75t_L   g01787(.A1(new_n2028), .A2(new_n2035), .B(new_n2037), .C(new_n2043), .Y(new_n2044));
  INVx1_ASAP7_75t_L         g01788(.A(\b[22] ), .Y(new_n2045));
  NAND2xp33_ASAP7_75t_L     g01789(.A(\b[20] ), .B(new_n286), .Y(new_n2046));
  OAI221xp5_ASAP7_75t_L     g01790(.A1(new_n285), .A2(new_n1895), .B1(new_n2045), .B2(new_n269), .C(new_n2046), .Y(new_n2047));
  NOR2xp33_ASAP7_75t_L      g01791(.A(\b[21] ), .B(\b[22] ), .Y(new_n2048));
  NOR2xp33_ASAP7_75t_L      g01792(.A(new_n1895), .B(new_n2045), .Y(new_n2049));
  NOR2xp33_ASAP7_75t_L      g01793(.A(new_n2048), .B(new_n2049), .Y(new_n2050));
  INVx1_ASAP7_75t_L         g01794(.A(new_n2050), .Y(new_n2051));
  O2A1O1Ixp33_ASAP7_75t_L   g01795(.A1(new_n1745), .A2(new_n1895), .B(new_n1898), .C(new_n2051), .Y(new_n2052));
  INVx1_ASAP7_75t_L         g01796(.A(new_n2052), .Y(new_n2053));
  A2O1A1O1Ixp25_ASAP7_75t_L g01797(.A1(new_n1747), .A2(new_n1750), .B(new_n1746), .C(new_n1897), .D(new_n1896), .Y(new_n2054));
  NAND2xp33_ASAP7_75t_L     g01798(.A(new_n2051), .B(new_n2054), .Y(new_n2055));
  AND2x2_ASAP7_75t_L        g01799(.A(new_n2055), .B(new_n2053), .Y(new_n2056));
  A2O1A1Ixp33_ASAP7_75t_L   g01800(.A1(new_n2056), .A2(new_n273), .B(new_n2047), .C(\a[2] ), .Y(new_n2057));
  AOI211xp5_ASAP7_75t_L     g01801(.A1(new_n2056), .A2(new_n273), .B(new_n2047), .C(new_n257), .Y(new_n2058));
  A2O1A1O1Ixp25_ASAP7_75t_L g01802(.A1(new_n273), .A2(new_n2056), .B(new_n2047), .C(new_n2057), .D(new_n2058), .Y(new_n2059));
  OAI21xp33_ASAP7_75t_L     g01803(.A1(new_n2041), .A2(new_n2044), .B(new_n2059), .Y(new_n2060));
  NOR3xp33_ASAP7_75t_L      g01804(.A(new_n2044), .B(new_n2041), .C(new_n2059), .Y(new_n2061));
  INVx1_ASAP7_75t_L         g01805(.A(new_n2061), .Y(new_n2062));
  NAND2xp33_ASAP7_75t_L     g01806(.A(new_n2060), .B(new_n2062), .Y(new_n2063));
  O2A1O1Ixp33_ASAP7_75t_L   g01807(.A1(new_n1922), .A2(new_n1906), .B(new_n1915), .C(new_n2063), .Y(new_n2064));
  O2A1O1Ixp33_ASAP7_75t_L   g01808(.A1(new_n1902), .A2(new_n257), .B(new_n1904), .C(new_n1922), .Y(new_n2065));
  A2O1A1O1Ixp25_ASAP7_75t_L g01809(.A1(new_n1757), .A2(new_n1771), .B(new_n1766), .C(new_n1914), .D(new_n2065), .Y(new_n2066));
  AND2x2_ASAP7_75t_L        g01810(.A(new_n2066), .B(new_n2063), .Y(new_n2067));
  NOR2xp33_ASAP7_75t_L      g01811(.A(new_n2064), .B(new_n2067), .Y(\f[22] ));
  INVx1_ASAP7_75t_L         g01812(.A(new_n2035), .Y(new_n2069));
  A2O1A1Ixp33_ASAP7_75t_L   g01813(.A1(new_n1890), .A2(new_n1910), .B(new_n2042), .C(new_n2038), .Y(new_n2070));
  NOR2xp33_ASAP7_75t_L      g01814(.A(new_n1150), .B(new_n513), .Y(new_n2071));
  AOI221xp5_ASAP7_75t_L     g01815(.A1(\b[15] ), .A2(new_n560), .B1(\b[17] ), .B2(new_n475), .C(new_n2071), .Y(new_n2072));
  O2A1O1Ixp33_ASAP7_75t_L   g01816(.A1(new_n477), .A2(new_n1356), .B(new_n2072), .C(new_n466), .Y(new_n2073));
  INVx1_ASAP7_75t_L         g01817(.A(new_n2072), .Y(new_n2074));
  A2O1A1Ixp33_ASAP7_75t_L   g01818(.A1(new_n1633), .A2(new_n483), .B(new_n2074), .C(new_n466), .Y(new_n2075));
  OAI21xp33_ASAP7_75t_L     g01819(.A1(new_n466), .A2(new_n2073), .B(new_n2075), .Y(new_n2076));
  NAND2xp33_ASAP7_75t_L     g01820(.A(new_n2000), .B(new_n1999), .Y(new_n2077));
  MAJIxp5_ASAP7_75t_L       g01821(.A(new_n2007), .B(new_n2001), .C(new_n2077), .Y(new_n2078));
  NOR2xp33_ASAP7_75t_L      g01822(.A(new_n680), .B(new_n864), .Y(new_n2079));
  AOI221xp5_ASAP7_75t_L     g01823(.A1(\b[9] ), .A2(new_n985), .B1(\b[11] ), .B2(new_n886), .C(new_n2079), .Y(new_n2080));
  O2A1O1Ixp33_ASAP7_75t_L   g01824(.A1(new_n872), .A2(new_n754), .B(new_n2080), .C(new_n867), .Y(new_n2081));
  INVx1_ASAP7_75t_L         g01825(.A(new_n2080), .Y(new_n2082));
  A2O1A1Ixp33_ASAP7_75t_L   g01826(.A1(new_n976), .A2(new_n873), .B(new_n2082), .C(new_n867), .Y(new_n2083));
  OAI21xp33_ASAP7_75t_L     g01827(.A1(new_n867), .A2(new_n2081), .B(new_n2083), .Y(new_n2084));
  A2O1A1Ixp33_ASAP7_75t_L   g01828(.A1(new_n1930), .A2(new_n1824), .B(new_n1986), .C(new_n1989), .Y(new_n2085));
  OAI211xp5_ASAP7_75t_L     g01829(.A1(new_n1968), .A2(new_n1969), .B(new_n1966), .C(new_n1959), .Y(new_n2086));
  A2O1A1Ixp33_ASAP7_75t_L   g01830(.A1(new_n1967), .A2(new_n1978), .B(new_n1938), .C(new_n2086), .Y(new_n2087));
  NAND2xp33_ASAP7_75t_L     g01831(.A(\b[2] ), .B(new_n1955), .Y(new_n2088));
  NAND3xp33_ASAP7_75t_L     g01832(.A(new_n1793), .B(new_n1949), .C(new_n1954), .Y(new_n2089));
  NAND2xp33_ASAP7_75t_L     g01833(.A(\b[1] ), .B(new_n1950), .Y(new_n2090));
  OAI211xp5_ASAP7_75t_L     g01834(.A1(new_n284), .A2(new_n2089), .B(new_n2088), .C(new_n2090), .Y(new_n2091));
  A2O1A1Ixp33_ASAP7_75t_L   g01835(.A1(new_n294), .A2(new_n1964), .B(new_n2091), .C(\a[23] ), .Y(new_n2092));
  INVx1_ASAP7_75t_L         g01836(.A(new_n2089), .Y(new_n2093));
  NOR2xp33_ASAP7_75t_L      g01837(.A(new_n262), .B(new_n1962), .Y(new_n2094));
  AOI221xp5_ASAP7_75t_L     g01838(.A1(new_n1955), .A2(\b[2] ), .B1(new_n2093), .B2(\b[0] ), .C(new_n2094), .Y(new_n2095));
  O2A1O1Ixp33_ASAP7_75t_L   g01839(.A1(new_n509), .A2(new_n1956), .B(new_n2095), .C(\a[23] ), .Y(new_n2096));
  A2O1A1O1Ixp25_ASAP7_75t_L g01840(.A1(new_n1958), .A2(new_n1795), .B(new_n2092), .C(\a[23] ), .D(new_n2096), .Y(new_n2097));
  NOR2xp33_ASAP7_75t_L      g01841(.A(new_n1956), .B(new_n509), .Y(new_n2098));
  NOR5xp2_ASAP7_75t_L       g01842(.A(new_n1971), .B(new_n2091), .C(new_n2098), .D(new_n1794), .E(new_n1952), .Y(new_n2099));
  NAND2xp33_ASAP7_75t_L     g01843(.A(\b[4] ), .B(new_n1507), .Y(new_n2100));
  OAI221xp5_ASAP7_75t_L     g01844(.A1(new_n1518), .A2(new_n384), .B1(new_n301), .B2(new_n1654), .C(new_n2100), .Y(new_n2101));
  A2O1A1Ixp33_ASAP7_75t_L   g01845(.A1(new_n394), .A2(new_n1513), .B(new_n2101), .C(\a[20] ), .Y(new_n2102));
  INVx1_ASAP7_75t_L         g01846(.A(new_n2101), .Y(new_n2103));
  O2A1O1Ixp33_ASAP7_75t_L   g01847(.A1(new_n1521), .A2(new_n728), .B(new_n2103), .C(\a[20] ), .Y(new_n2104));
  AOI21xp33_ASAP7_75t_L     g01848(.A1(new_n2102), .A2(\a[20] ), .B(new_n2104), .Y(new_n2105));
  NOR3xp33_ASAP7_75t_L      g01849(.A(new_n2105), .B(new_n2097), .C(new_n2099), .Y(new_n2106));
  NAND2xp33_ASAP7_75t_L     g01850(.A(\b[0] ), .B(new_n2093), .Y(new_n2107));
  INVx1_ASAP7_75t_L         g01851(.A(new_n2098), .Y(new_n2108));
  NAND5xp2_ASAP7_75t_L      g01852(.A(\a[23] ), .B(new_n2107), .C(new_n2108), .D(new_n2090), .E(new_n2088), .Y(new_n2109));
  A2O1A1Ixp33_ASAP7_75t_L   g01853(.A1(new_n294), .A2(new_n1964), .B(new_n2091), .C(new_n1952), .Y(new_n2110));
  NAND3xp33_ASAP7_75t_L     g01854(.A(new_n2110), .B(new_n2109), .C(new_n1959), .Y(new_n2111));
  NAND5xp2_ASAP7_75t_L      g01855(.A(\a[23] ), .B(new_n2095), .C(new_n2108), .D(new_n1958), .E(new_n1795), .Y(new_n2112));
  AOI221xp5_ASAP7_75t_L     g01856(.A1(new_n2102), .A2(\a[20] ), .B1(new_n2112), .B2(new_n2111), .C(new_n2104), .Y(new_n2113));
  OAI21xp33_ASAP7_75t_L     g01857(.A1(new_n2106), .A2(new_n2113), .B(new_n2087), .Y(new_n2114));
  OR3x1_ASAP7_75t_L         g01858(.A(new_n2105), .B(new_n2097), .C(new_n2099), .Y(new_n2115));
  OAI21xp33_ASAP7_75t_L     g01859(.A1(new_n2099), .A2(new_n2097), .B(new_n2105), .Y(new_n2116));
  NAND4xp25_ASAP7_75t_L     g01860(.A(new_n1985), .B(new_n2116), .C(new_n2115), .D(new_n2086), .Y(new_n2117));
  OAI21xp33_ASAP7_75t_L     g01861(.A1(new_n1201), .A2(new_n1202), .B(new_n1076), .Y(new_n2118));
  NOR2xp33_ASAP7_75t_L      g01862(.A(new_n448), .B(new_n2118), .Y(new_n2119));
  AOI221xp5_ASAP7_75t_L     g01863(.A1(\b[6] ), .A2(new_n1290), .B1(\b[8] ), .B2(new_n1209), .C(new_n2119), .Y(new_n2120));
  O2A1O1Ixp33_ASAP7_75t_L   g01864(.A1(new_n1210), .A2(new_n540), .B(new_n2120), .C(new_n1206), .Y(new_n2121));
  NOR2xp33_ASAP7_75t_L      g01865(.A(new_n1206), .B(new_n2121), .Y(new_n2122));
  O2A1O1Ixp33_ASAP7_75t_L   g01866(.A1(new_n1210), .A2(new_n540), .B(new_n2120), .C(\a[17] ), .Y(new_n2123));
  NOR2xp33_ASAP7_75t_L      g01867(.A(new_n2123), .B(new_n2122), .Y(new_n2124));
  NAND3xp33_ASAP7_75t_L     g01868(.A(new_n2117), .B(new_n2124), .C(new_n2114), .Y(new_n2125));
  AO21x2_ASAP7_75t_L        g01869(.A1(new_n2114), .A2(new_n2117), .B(new_n2124), .Y(new_n2126));
  NAND3xp33_ASAP7_75t_L     g01870(.A(new_n2085), .B(new_n2125), .C(new_n2126), .Y(new_n2127));
  AO21x2_ASAP7_75t_L        g01871(.A1(new_n2126), .A2(new_n2125), .B(new_n2085), .Y(new_n2128));
  AO21x2_ASAP7_75t_L        g01872(.A1(new_n2127), .A2(new_n2128), .B(new_n2084), .Y(new_n2129));
  NAND3xp33_ASAP7_75t_L     g01873(.A(new_n2128), .B(new_n2127), .C(new_n2084), .Y(new_n2130));
  NAND3xp33_ASAP7_75t_L     g01874(.A(new_n2078), .B(new_n2129), .C(new_n2130), .Y(new_n2131));
  NOR2xp33_ASAP7_75t_L      g01875(.A(new_n1991), .B(new_n1987), .Y(new_n2132));
  MAJIxp5_ASAP7_75t_L       g01876(.A(new_n2003), .B(new_n1997), .C(new_n2132), .Y(new_n2133));
  AOI21xp33_ASAP7_75t_L     g01877(.A1(new_n2128), .A2(new_n2127), .B(new_n2084), .Y(new_n2134));
  AND3x1_ASAP7_75t_L        g01878(.A(new_n2128), .B(new_n2127), .C(new_n2084), .Y(new_n2135));
  OAI21xp33_ASAP7_75t_L     g01879(.A1(new_n2134), .A2(new_n2135), .B(new_n2133), .Y(new_n2136));
  NOR2xp33_ASAP7_75t_L      g01880(.A(new_n936), .B(new_n1550), .Y(new_n2137));
  AOI221xp5_ASAP7_75t_L     g01881(.A1(\b[12] ), .A2(new_n713), .B1(\b[14] ), .B2(new_n640), .C(new_n2137), .Y(new_n2138));
  INVx1_ASAP7_75t_L         g01882(.A(new_n2138), .Y(new_n2139));
  A2O1A1Ixp33_ASAP7_75t_L   g01883(.A1(new_n971), .A2(new_n718), .B(new_n2139), .C(\a[11] ), .Y(new_n2140));
  O2A1O1Ixp33_ASAP7_75t_L   g01884(.A1(new_n641), .A2(new_n1268), .B(new_n2138), .C(\a[11] ), .Y(new_n2141));
  AOI21xp33_ASAP7_75t_L     g01885(.A1(new_n2140), .A2(\a[11] ), .B(new_n2141), .Y(new_n2142));
  NAND3xp33_ASAP7_75t_L     g01886(.A(new_n2131), .B(new_n2136), .C(new_n2142), .Y(new_n2143));
  NOR3xp33_ASAP7_75t_L      g01887(.A(new_n2133), .B(new_n2135), .C(new_n2134), .Y(new_n2144));
  AOI21xp33_ASAP7_75t_L     g01888(.A1(new_n2129), .A2(new_n2130), .B(new_n2078), .Y(new_n2145));
  INVx1_ASAP7_75t_L         g01889(.A(new_n2142), .Y(new_n2146));
  OAI21xp33_ASAP7_75t_L     g01890(.A1(new_n2144), .A2(new_n2145), .B(new_n2146), .Y(new_n2147));
  OAI21xp33_ASAP7_75t_L     g01891(.A1(new_n2008), .A2(new_n2004), .B(new_n2014), .Y(new_n2148));
  A2O1A1O1Ixp25_ASAP7_75t_L g01892(.A1(new_n1928), .A2(new_n1859), .B(new_n1845), .C(new_n2148), .D(new_n2016), .Y(new_n2149));
  AOI21xp33_ASAP7_75t_L     g01893(.A1(new_n2147), .A2(new_n2143), .B(new_n2149), .Y(new_n2150));
  NOR3xp33_ASAP7_75t_L      g01894(.A(new_n2146), .B(new_n2145), .C(new_n2144), .Y(new_n2151));
  AOI21xp33_ASAP7_75t_L     g01895(.A1(new_n2131), .A2(new_n2136), .B(new_n2142), .Y(new_n2152));
  INVx1_ASAP7_75t_L         g01896(.A(new_n2016), .Y(new_n2153));
  OAI21xp33_ASAP7_75t_L     g01897(.A1(new_n2015), .A2(new_n1929), .B(new_n2153), .Y(new_n2154));
  NOR3xp33_ASAP7_75t_L      g01898(.A(new_n2154), .B(new_n2151), .C(new_n2152), .Y(new_n2155));
  OAI21xp33_ASAP7_75t_L     g01899(.A1(new_n2150), .A2(new_n2155), .B(new_n2076), .Y(new_n2156));
  A2O1A1Ixp33_ASAP7_75t_L   g01900(.A1(new_n1633), .A2(new_n483), .B(new_n2074), .C(\a[8] ), .Y(new_n2157));
  O2A1O1Ixp33_ASAP7_75t_L   g01901(.A1(new_n477), .A2(new_n1356), .B(new_n2072), .C(\a[8] ), .Y(new_n2158));
  AOI21xp33_ASAP7_75t_L     g01902(.A1(new_n2157), .A2(\a[8] ), .B(new_n2158), .Y(new_n2159));
  OAI21xp33_ASAP7_75t_L     g01903(.A1(new_n2152), .A2(new_n2151), .B(new_n2154), .Y(new_n2160));
  NAND3xp33_ASAP7_75t_L     g01904(.A(new_n2149), .B(new_n2147), .C(new_n2143), .Y(new_n2161));
  NAND3xp33_ASAP7_75t_L     g01905(.A(new_n2161), .B(new_n2160), .C(new_n2159), .Y(new_n2162));
  NAND2xp33_ASAP7_75t_L     g01906(.A(new_n2162), .B(new_n2156), .Y(new_n2163));
  O2A1O1Ixp33_ASAP7_75t_L   g01907(.A1(new_n1924), .A2(new_n2023), .B(new_n2025), .C(new_n2163), .Y(new_n2164));
  OAI21xp33_ASAP7_75t_L     g01908(.A1(new_n2023), .A2(new_n1924), .B(new_n2025), .Y(new_n2165));
  NOR3xp33_ASAP7_75t_L      g01909(.A(new_n2155), .B(new_n2150), .C(new_n2159), .Y(new_n2166));
  O2A1O1Ixp33_ASAP7_75t_L   g01910(.A1(new_n2159), .A2(new_n2166), .B(new_n2162), .C(new_n2165), .Y(new_n2167));
  NOR2xp33_ASAP7_75t_L      g01911(.A(new_n1458), .B(new_n375), .Y(new_n2168));
  AOI221xp5_ASAP7_75t_L     g01912(.A1(\b[20] ), .A2(new_n361), .B1(new_n349), .B2(\b[19] ), .C(new_n2168), .Y(new_n2169));
  INVx1_ASAP7_75t_L         g01913(.A(new_n2169), .Y(new_n2170));
  A2O1A1Ixp33_ASAP7_75t_L   g01914(.A1(new_n1752), .A2(new_n359), .B(new_n2170), .C(\a[5] ), .Y(new_n2171));
  NAND2xp33_ASAP7_75t_L     g01915(.A(\a[5] ), .B(new_n2171), .Y(new_n2172));
  A2O1A1Ixp33_ASAP7_75t_L   g01916(.A1(new_n1752), .A2(new_n359), .B(new_n2170), .C(new_n346), .Y(new_n2173));
  AND2x2_ASAP7_75t_L        g01917(.A(new_n2173), .B(new_n2172), .Y(new_n2174));
  OAI21xp33_ASAP7_75t_L     g01918(.A1(new_n2167), .A2(new_n2164), .B(new_n2174), .Y(new_n2175));
  NAND3xp33_ASAP7_75t_L     g01919(.A(new_n2165), .B(new_n2156), .C(new_n2162), .Y(new_n2176));
  A2O1A1O1Ixp25_ASAP7_75t_L g01920(.A1(new_n1861), .A2(new_n1866), .B(new_n1923), .C(new_n2026), .D(new_n2020), .Y(new_n2177));
  NAND2xp33_ASAP7_75t_L     g01921(.A(new_n2163), .B(new_n2177), .Y(new_n2178));
  NAND2xp33_ASAP7_75t_L     g01922(.A(new_n2173), .B(new_n2172), .Y(new_n2179));
  NAND3xp33_ASAP7_75t_L     g01923(.A(new_n2178), .B(new_n2176), .C(new_n2179), .Y(new_n2180));
  NAND4xp25_ASAP7_75t_L     g01924(.A(new_n2070), .B(new_n2175), .C(new_n2180), .D(new_n2069), .Y(new_n2181));
  NAND2xp33_ASAP7_75t_L     g01925(.A(new_n2180), .B(new_n2175), .Y(new_n2182));
  A2O1A1Ixp33_ASAP7_75t_L   g01926(.A1(new_n2038), .A2(new_n2040), .B(new_n2035), .C(new_n2182), .Y(new_n2183));
  NAND2xp33_ASAP7_75t_L     g01927(.A(new_n2183), .B(new_n2181), .Y(new_n2184));
  NOR2xp33_ASAP7_75t_L      g01928(.A(new_n1895), .B(new_n287), .Y(new_n2185));
  AOI221xp5_ASAP7_75t_L     g01929(.A1(\b[22] ), .A2(new_n264), .B1(\b[23] ), .B2(new_n283), .C(new_n2185), .Y(new_n2186));
  NOR2xp33_ASAP7_75t_L      g01930(.A(\b[22] ), .B(\b[23] ), .Y(new_n2187));
  INVx1_ASAP7_75t_L         g01931(.A(\b[23] ), .Y(new_n2188));
  NOR2xp33_ASAP7_75t_L      g01932(.A(new_n2045), .B(new_n2188), .Y(new_n2189));
  NOR2xp33_ASAP7_75t_L      g01933(.A(new_n2187), .B(new_n2189), .Y(new_n2190));
  A2O1A1Ixp33_ASAP7_75t_L   g01934(.A1(\b[22] ), .A2(\b[21] ), .B(new_n2052), .C(new_n2190), .Y(new_n2191));
  INVx1_ASAP7_75t_L         g01935(.A(new_n2049), .Y(new_n2192));
  OAI211xp5_ASAP7_75t_L     g01936(.A1(new_n2187), .A2(new_n2189), .B(new_n2053), .C(new_n2192), .Y(new_n2193));
  NAND2xp33_ASAP7_75t_L     g01937(.A(new_n2191), .B(new_n2193), .Y(new_n2194));
  O2A1O1Ixp33_ASAP7_75t_L   g01938(.A1(new_n279), .A2(new_n2194), .B(new_n2186), .C(new_n257), .Y(new_n2195));
  O2A1O1Ixp33_ASAP7_75t_L   g01939(.A1(new_n279), .A2(new_n2194), .B(new_n2186), .C(\a[2] ), .Y(new_n2196));
  INVx1_ASAP7_75t_L         g01940(.A(new_n2196), .Y(new_n2197));
  O2A1O1Ixp33_ASAP7_75t_L   g01941(.A1(new_n2195), .A2(new_n257), .B(new_n2197), .C(new_n2184), .Y(new_n2198));
  INVx1_ASAP7_75t_L         g01942(.A(new_n2195), .Y(new_n2199));
  A2O1A1Ixp33_ASAP7_75t_L   g01943(.A1(\a[2] ), .A2(new_n2199), .B(new_n2196), .C(new_n2184), .Y(new_n2200));
  A2O1A1O1Ixp25_ASAP7_75t_L g01944(.A1(new_n1914), .A2(new_n1919), .B(new_n2065), .C(new_n2060), .D(new_n2061), .Y(new_n2201));
  O2A1O1Ixp33_ASAP7_75t_L   g01945(.A1(new_n2184), .A2(new_n2198), .B(new_n2200), .C(new_n2201), .Y(new_n2202));
  OA211x2_ASAP7_75t_L       g01946(.A1(new_n2184), .A2(new_n2198), .B(new_n2200), .C(new_n2201), .Y(new_n2203));
  NOR2xp33_ASAP7_75t_L      g01947(.A(new_n2202), .B(new_n2203), .Y(\f[23] ));
  INVx1_ASAP7_75t_L         g01948(.A(\b[24] ), .Y(new_n2205));
  NAND2xp33_ASAP7_75t_L     g01949(.A(\b[22] ), .B(new_n286), .Y(new_n2206));
  OAI221xp5_ASAP7_75t_L     g01950(.A1(new_n285), .A2(new_n2188), .B1(new_n2205), .B2(new_n269), .C(new_n2206), .Y(new_n2207));
  INVx1_ASAP7_75t_L         g01951(.A(new_n1896), .Y(new_n2208));
  A2O1A1Ixp33_ASAP7_75t_L   g01952(.A1(new_n1898), .A2(new_n2208), .B(new_n2048), .C(new_n2192), .Y(new_n2209));
  NOR2xp33_ASAP7_75t_L      g01953(.A(\b[23] ), .B(\b[24] ), .Y(new_n2210));
  NOR2xp33_ASAP7_75t_L      g01954(.A(new_n2188), .B(new_n2205), .Y(new_n2211));
  NOR2xp33_ASAP7_75t_L      g01955(.A(new_n2210), .B(new_n2211), .Y(new_n2212));
  A2O1A1Ixp33_ASAP7_75t_L   g01956(.A1(new_n2209), .A2(new_n2190), .B(new_n2189), .C(new_n2212), .Y(new_n2213));
  O2A1O1Ixp33_ASAP7_75t_L   g01957(.A1(new_n2049), .A2(new_n2052), .B(new_n2190), .C(new_n2189), .Y(new_n2214));
  OAI21xp33_ASAP7_75t_L     g01958(.A1(new_n2210), .A2(new_n2211), .B(new_n2214), .Y(new_n2215));
  AND2x2_ASAP7_75t_L        g01959(.A(new_n2213), .B(new_n2215), .Y(new_n2216));
  A2O1A1Ixp33_ASAP7_75t_L   g01960(.A1(new_n2216), .A2(new_n273), .B(new_n2207), .C(\a[2] ), .Y(new_n2217));
  AOI211xp5_ASAP7_75t_L     g01961(.A1(new_n2216), .A2(new_n273), .B(new_n2207), .C(new_n257), .Y(new_n2218));
  A2O1A1O1Ixp25_ASAP7_75t_L g01962(.A1(new_n273), .A2(new_n2216), .B(new_n2207), .C(new_n2217), .D(new_n2218), .Y(new_n2219));
  INVx1_ASAP7_75t_L         g01963(.A(new_n1924), .Y(new_n2220));
  A2O1A1Ixp33_ASAP7_75t_L   g01964(.A1(new_n2026), .A2(new_n2220), .B(new_n2020), .C(new_n2163), .Y(new_n2221));
  INVx1_ASAP7_75t_L         g01965(.A(new_n2221), .Y(new_n2222));
  O2A1O1Ixp33_ASAP7_75t_L   g01966(.A1(new_n2177), .A2(new_n2222), .B(new_n2178), .C(new_n2174), .Y(new_n2223));
  A2O1A1O1Ixp25_ASAP7_75t_L g01967(.A1(new_n2038), .A2(new_n2040), .B(new_n2035), .C(new_n2182), .D(new_n2223), .Y(new_n2224));
  NOR2xp33_ASAP7_75t_L      g01968(.A(new_n1599), .B(new_n375), .Y(new_n2225));
  AOI221xp5_ASAP7_75t_L     g01969(.A1(\b[21] ), .A2(new_n361), .B1(new_n349), .B2(\b[20] ), .C(new_n2225), .Y(new_n2226));
  O2A1O1Ixp33_ASAP7_75t_L   g01970(.A1(new_n356), .A2(new_n1901), .B(new_n2226), .C(new_n346), .Y(new_n2227));
  NOR2xp33_ASAP7_75t_L      g01971(.A(new_n346), .B(new_n2227), .Y(new_n2228));
  O2A1O1Ixp33_ASAP7_75t_L   g01972(.A1(new_n356), .A2(new_n1901), .B(new_n2226), .C(\a[5] ), .Y(new_n2229));
  NOR2xp33_ASAP7_75t_L      g01973(.A(new_n2229), .B(new_n2228), .Y(new_n2230));
  INVx1_ASAP7_75t_L         g01974(.A(new_n2229), .Y(new_n2231));
  OAI21xp33_ASAP7_75t_L     g01975(.A1(new_n346), .A2(new_n2227), .B(new_n2231), .Y(new_n2232));
  INVx1_ASAP7_75t_L         g01976(.A(new_n2166), .Y(new_n2233));
  A2O1A1Ixp33_ASAP7_75t_L   g01977(.A1(new_n2162), .A2(new_n2159), .B(new_n2177), .C(new_n2233), .Y(new_n2234));
  NAND2xp33_ASAP7_75t_L     g01978(.A(new_n1997), .B(new_n2132), .Y(new_n2235));
  OAI21xp33_ASAP7_75t_L     g01979(.A1(new_n1998), .A2(new_n2002), .B(new_n2003), .Y(new_n2236));
  A2O1A1Ixp33_ASAP7_75t_L   g01980(.A1(new_n2236), .A2(new_n2235), .B(new_n2134), .C(new_n2130), .Y(new_n2237));
  NOR2xp33_ASAP7_75t_L      g01981(.A(new_n748), .B(new_n864), .Y(new_n2238));
  AOI221xp5_ASAP7_75t_L     g01982(.A1(\b[10] ), .A2(new_n985), .B1(\b[12] ), .B2(new_n886), .C(new_n2238), .Y(new_n2239));
  INVx1_ASAP7_75t_L         g01983(.A(new_n2239), .Y(new_n2240));
  A2O1A1Ixp33_ASAP7_75t_L   g01984(.A1(new_n1057), .A2(new_n873), .B(new_n2240), .C(\a[14] ), .Y(new_n2241));
  O2A1O1Ixp33_ASAP7_75t_L   g01985(.A1(new_n872), .A2(new_n841), .B(new_n2239), .C(\a[14] ), .Y(new_n2242));
  AOI21xp33_ASAP7_75t_L     g01986(.A1(new_n2241), .A2(\a[14] ), .B(new_n2242), .Y(new_n2243));
  AOI21xp33_ASAP7_75t_L     g01987(.A1(new_n2117), .A2(new_n2114), .B(new_n2124), .Y(new_n2244));
  A2O1A1O1Ixp25_ASAP7_75t_L g01988(.A1(new_n1990), .A2(new_n1988), .B(new_n1982), .C(new_n2125), .D(new_n2244), .Y(new_n2245));
  A2O1A1O1Ixp25_ASAP7_75t_L g01989(.A1(new_n1967), .A2(new_n1978), .B(new_n1938), .C(new_n2086), .D(new_n2113), .Y(new_n2246));
  INVx1_ASAP7_75t_L         g01990(.A(\a[24] ), .Y(new_n2247));
  NAND2xp33_ASAP7_75t_L     g01991(.A(\a[23] ), .B(new_n2247), .Y(new_n2248));
  NAND2xp33_ASAP7_75t_L     g01992(.A(\a[24] ), .B(new_n1952), .Y(new_n2249));
  AND2x2_ASAP7_75t_L        g01993(.A(new_n2248), .B(new_n2249), .Y(new_n2250));
  NOR2xp33_ASAP7_75t_L      g01994(.A(new_n284), .B(new_n2250), .Y(new_n2251));
  INVx1_ASAP7_75t_L         g01995(.A(new_n2251), .Y(new_n2252));
  NOR2xp33_ASAP7_75t_L      g01996(.A(new_n2252), .B(new_n2099), .Y(new_n2253));
  NOR2xp33_ASAP7_75t_L      g01997(.A(new_n2251), .B(new_n2112), .Y(new_n2254));
  NAND2xp33_ASAP7_75t_L     g01998(.A(\b[3] ), .B(new_n1955), .Y(new_n2255));
  NAND2xp33_ASAP7_75t_L     g01999(.A(\b[1] ), .B(new_n2093), .Y(new_n2256));
  NAND2xp33_ASAP7_75t_L     g02000(.A(\b[2] ), .B(new_n1950), .Y(new_n2257));
  NAND2xp33_ASAP7_75t_L     g02001(.A(new_n1964), .B(new_n312), .Y(new_n2258));
  NAND5xp2_ASAP7_75t_L      g02002(.A(new_n2258), .B(new_n2257), .C(new_n2256), .D(new_n2255), .E(\a[23] ), .Y(new_n2259));
  OAI211xp5_ASAP7_75t_L     g02003(.A1(new_n2089), .A2(new_n262), .B(new_n2255), .C(new_n2257), .Y(new_n2260));
  A2O1A1Ixp33_ASAP7_75t_L   g02004(.A1(new_n312), .A2(new_n1964), .B(new_n2260), .C(new_n1952), .Y(new_n2261));
  NAND2xp33_ASAP7_75t_L     g02005(.A(new_n2259), .B(new_n2261), .Y(new_n2262));
  OAI21xp33_ASAP7_75t_L     g02006(.A1(new_n2254), .A2(new_n2253), .B(new_n2262), .Y(new_n2263));
  A2O1A1Ixp33_ASAP7_75t_L   g02007(.A1(new_n2110), .A2(new_n2109), .B(new_n1959), .C(new_n2251), .Y(new_n2264));
  NAND2xp33_ASAP7_75t_L     g02008(.A(new_n2252), .B(new_n2099), .Y(new_n2265));
  AND2x2_ASAP7_75t_L        g02009(.A(new_n2259), .B(new_n2261), .Y(new_n2266));
  NAND3xp33_ASAP7_75t_L     g02010(.A(new_n2265), .B(new_n2264), .C(new_n2266), .Y(new_n2267));
  NOR2xp33_ASAP7_75t_L      g02011(.A(new_n427), .B(new_n1518), .Y(new_n2268));
  AOI221xp5_ASAP7_75t_L     g02012(.A1(\b[4] ), .A2(new_n1659), .B1(\b[5] ), .B2(new_n1507), .C(new_n2268), .Y(new_n2269));
  OAI21xp33_ASAP7_75t_L     g02013(.A1(new_n1521), .A2(new_n434), .B(new_n2269), .Y(new_n2270));
  NOR2xp33_ASAP7_75t_L      g02014(.A(new_n1501), .B(new_n2270), .Y(new_n2271));
  O2A1O1Ixp33_ASAP7_75t_L   g02015(.A1(new_n1521), .A2(new_n434), .B(new_n2269), .C(\a[20] ), .Y(new_n2272));
  NOR2xp33_ASAP7_75t_L      g02016(.A(new_n2272), .B(new_n2271), .Y(new_n2273));
  NAND3xp33_ASAP7_75t_L     g02017(.A(new_n2273), .B(new_n2267), .C(new_n2263), .Y(new_n2274));
  AOI21xp33_ASAP7_75t_L     g02018(.A1(new_n2265), .A2(new_n2264), .B(new_n2266), .Y(new_n2275));
  NOR3xp33_ASAP7_75t_L      g02019(.A(new_n2253), .B(new_n2254), .C(new_n2262), .Y(new_n2276));
  O2A1O1Ixp33_ASAP7_75t_L   g02020(.A1(new_n1521), .A2(new_n434), .B(new_n2269), .C(new_n1501), .Y(new_n2277));
  INVx1_ASAP7_75t_L         g02021(.A(new_n2272), .Y(new_n2278));
  OAI21xp33_ASAP7_75t_L     g02022(.A1(new_n1501), .A2(new_n2277), .B(new_n2278), .Y(new_n2279));
  OAI21xp33_ASAP7_75t_L     g02023(.A1(new_n2275), .A2(new_n2276), .B(new_n2279), .Y(new_n2280));
  OAI211xp5_ASAP7_75t_L     g02024(.A1(new_n2106), .A2(new_n2246), .B(new_n2274), .C(new_n2280), .Y(new_n2281));
  INVx1_ASAP7_75t_L         g02025(.A(new_n2086), .Y(new_n2282));
  A2O1A1O1Ixp25_ASAP7_75t_L g02026(.A1(new_n1983), .A2(new_n1984), .B(new_n2282), .C(new_n2116), .D(new_n2106), .Y(new_n2283));
  NAND3xp33_ASAP7_75t_L     g02027(.A(new_n2279), .B(new_n2263), .C(new_n2267), .Y(new_n2284));
  NOR3xp33_ASAP7_75t_L      g02028(.A(new_n2279), .B(new_n2276), .C(new_n2275), .Y(new_n2285));
  A2O1A1Ixp33_ASAP7_75t_L   g02029(.A1(new_n2279), .A2(new_n2284), .B(new_n2285), .C(new_n2283), .Y(new_n2286));
  NOR2xp33_ASAP7_75t_L      g02030(.A(new_n590), .B(new_n1284), .Y(new_n2287));
  AOI221xp5_ASAP7_75t_L     g02031(.A1(\b[7] ), .A2(new_n1290), .B1(\b[8] ), .B2(new_n1204), .C(new_n2287), .Y(new_n2288));
  INVx1_ASAP7_75t_L         g02032(.A(new_n2288), .Y(new_n2289));
  A2O1A1Ixp33_ASAP7_75t_L   g02033(.A1(new_n602), .A2(new_n1216), .B(new_n2289), .C(\a[17] ), .Y(new_n2290));
  NAND2xp33_ASAP7_75t_L     g02034(.A(\a[17] ), .B(new_n2290), .Y(new_n2291));
  A2O1A1Ixp33_ASAP7_75t_L   g02035(.A1(new_n602), .A2(new_n1216), .B(new_n2289), .C(new_n1206), .Y(new_n2292));
  AOI22xp33_ASAP7_75t_L     g02036(.A1(new_n2291), .A2(new_n2292), .B1(new_n2281), .B2(new_n2286), .Y(new_n2293));
  AOI21xp33_ASAP7_75t_L     g02037(.A1(new_n2263), .A2(new_n2267), .B(new_n2273), .Y(new_n2294));
  NOR3xp33_ASAP7_75t_L      g02038(.A(new_n2283), .B(new_n2285), .C(new_n2294), .Y(new_n2295));
  AOI211xp5_ASAP7_75t_L     g02039(.A1(new_n2274), .A2(new_n2280), .B(new_n2246), .C(new_n2106), .Y(new_n2296));
  NAND2xp33_ASAP7_75t_L     g02040(.A(new_n2292), .B(new_n2291), .Y(new_n2297));
  NOR3xp33_ASAP7_75t_L      g02041(.A(new_n2297), .B(new_n2296), .C(new_n2295), .Y(new_n2298));
  NOR3xp33_ASAP7_75t_L      g02042(.A(new_n2245), .B(new_n2293), .C(new_n2298), .Y(new_n2299));
  OAI21xp33_ASAP7_75t_L     g02043(.A1(new_n2295), .A2(new_n2296), .B(new_n2297), .Y(new_n2300));
  NAND4xp25_ASAP7_75t_L     g02044(.A(new_n2286), .B(new_n2281), .C(new_n2291), .D(new_n2292), .Y(new_n2301));
  AOI221xp5_ASAP7_75t_L     g02045(.A1(new_n2085), .A2(new_n2125), .B1(new_n2301), .B2(new_n2300), .C(new_n2244), .Y(new_n2302));
  OAI21xp33_ASAP7_75t_L     g02046(.A1(new_n2302), .A2(new_n2299), .B(new_n2243), .Y(new_n2303));
  NOR3xp33_ASAP7_75t_L      g02047(.A(new_n2299), .B(new_n2302), .C(new_n2243), .Y(new_n2304));
  INVx1_ASAP7_75t_L         g02048(.A(new_n2304), .Y(new_n2305));
  NAND3xp33_ASAP7_75t_L     g02049(.A(new_n2237), .B(new_n2305), .C(new_n2303), .Y(new_n2306));
  AOI21xp33_ASAP7_75t_L     g02050(.A1(new_n2078), .A2(new_n2129), .B(new_n2135), .Y(new_n2307));
  INVx1_ASAP7_75t_L         g02051(.A(new_n2303), .Y(new_n2308));
  OAI21xp33_ASAP7_75t_L     g02052(.A1(new_n2304), .A2(new_n2308), .B(new_n2307), .Y(new_n2309));
  NAND2xp33_ASAP7_75t_L     g02053(.A(new_n2309), .B(new_n2306), .Y(new_n2310));
  NOR2xp33_ASAP7_75t_L      g02054(.A(new_n960), .B(new_n1550), .Y(new_n2311));
  AOI221xp5_ASAP7_75t_L     g02055(.A1(\b[13] ), .A2(new_n713), .B1(\b[15] ), .B2(new_n640), .C(new_n2311), .Y(new_n2312));
  O2A1O1Ixp33_ASAP7_75t_L   g02056(.A1(new_n641), .A2(new_n1774), .B(new_n2312), .C(new_n637), .Y(new_n2313));
  INVx1_ASAP7_75t_L         g02057(.A(new_n2313), .Y(new_n2314));
  O2A1O1Ixp33_ASAP7_75t_L   g02058(.A1(new_n641), .A2(new_n1774), .B(new_n2312), .C(\a[11] ), .Y(new_n2315));
  AO21x2_ASAP7_75t_L        g02059(.A1(\a[11] ), .A2(new_n2314), .B(new_n2315), .Y(new_n2316));
  NOR2xp33_ASAP7_75t_L      g02060(.A(new_n2316), .B(new_n2310), .Y(new_n2317));
  AOI21xp33_ASAP7_75t_L     g02061(.A1(new_n2314), .A2(\a[11] ), .B(new_n2315), .Y(new_n2318));
  AOI21xp33_ASAP7_75t_L     g02062(.A1(new_n2306), .A2(new_n2309), .B(new_n2318), .Y(new_n2319));
  NAND2xp33_ASAP7_75t_L     g02063(.A(new_n2136), .B(new_n2131), .Y(new_n2320));
  MAJIxp5_ASAP7_75t_L       g02064(.A(new_n2149), .B(new_n2320), .C(new_n2142), .Y(new_n2321));
  NOR3xp33_ASAP7_75t_L      g02065(.A(new_n2317), .B(new_n2321), .C(new_n2319), .Y(new_n2322));
  NAND3xp33_ASAP7_75t_L     g02066(.A(new_n2318), .B(new_n2306), .C(new_n2309), .Y(new_n2323));
  NAND2xp33_ASAP7_75t_L     g02067(.A(new_n2316), .B(new_n2310), .Y(new_n2324));
  NOR2xp33_ASAP7_75t_L      g02068(.A(new_n2145), .B(new_n2144), .Y(new_n2325));
  MAJIxp5_ASAP7_75t_L       g02069(.A(new_n2154), .B(new_n2325), .C(new_n2146), .Y(new_n2326));
  AOI21xp33_ASAP7_75t_L     g02070(.A1(new_n2324), .A2(new_n2323), .B(new_n2326), .Y(new_n2327));
  INVx1_ASAP7_75t_L         g02071(.A(new_n1461), .Y(new_n2328));
  NOR2xp33_ASAP7_75t_L      g02072(.A(new_n1462), .B(new_n2328), .Y(new_n2329));
  NOR2xp33_ASAP7_75t_L      g02073(.A(new_n1349), .B(new_n513), .Y(new_n2330));
  AOI221xp5_ASAP7_75t_L     g02074(.A1(\b[16] ), .A2(new_n560), .B1(\b[18] ), .B2(new_n475), .C(new_n2330), .Y(new_n2331));
  INVx1_ASAP7_75t_L         g02075(.A(new_n2331), .Y(new_n2332));
  A2O1A1Ixp33_ASAP7_75t_L   g02076(.A1(new_n2329), .A2(new_n483), .B(new_n2332), .C(\a[8] ), .Y(new_n2333));
  O2A1O1Ixp33_ASAP7_75t_L   g02077(.A1(new_n477), .A2(new_n1464), .B(new_n2331), .C(\a[8] ), .Y(new_n2334));
  AOI21xp33_ASAP7_75t_L     g02078(.A1(new_n2333), .A2(\a[8] ), .B(new_n2334), .Y(new_n2335));
  OAI21xp33_ASAP7_75t_L     g02079(.A1(new_n2327), .A2(new_n2322), .B(new_n2335), .Y(new_n2336));
  NAND3xp33_ASAP7_75t_L     g02080(.A(new_n2326), .B(new_n2324), .C(new_n2323), .Y(new_n2337));
  OAI21xp33_ASAP7_75t_L     g02081(.A1(new_n2319), .A2(new_n2317), .B(new_n2321), .Y(new_n2338));
  O2A1O1Ixp33_ASAP7_75t_L   g02082(.A1(new_n477), .A2(new_n1464), .B(new_n2331), .C(new_n466), .Y(new_n2339));
  NOR2xp33_ASAP7_75t_L      g02083(.A(new_n466), .B(new_n2339), .Y(new_n2340));
  OAI211xp5_ASAP7_75t_L     g02084(.A1(new_n2340), .A2(new_n2334), .B(new_n2337), .C(new_n2338), .Y(new_n2341));
  NAND3xp33_ASAP7_75t_L     g02085(.A(new_n2234), .B(new_n2336), .C(new_n2341), .Y(new_n2342));
  A2O1A1O1Ixp25_ASAP7_75t_L g02086(.A1(new_n2026), .A2(new_n2220), .B(new_n2020), .C(new_n2163), .D(new_n2166), .Y(new_n2343));
  NAND2xp33_ASAP7_75t_L     g02087(.A(new_n2336), .B(new_n2341), .Y(new_n2344));
  NAND2xp33_ASAP7_75t_L     g02088(.A(new_n2344), .B(new_n2343), .Y(new_n2345));
  NAND3xp33_ASAP7_75t_L     g02089(.A(new_n2342), .B(new_n2232), .C(new_n2345), .Y(new_n2346));
  INVx1_ASAP7_75t_L         g02090(.A(new_n2346), .Y(new_n2347));
  NAND3xp33_ASAP7_75t_L     g02091(.A(new_n2342), .B(new_n2230), .C(new_n2345), .Y(new_n2348));
  O2A1O1Ixp33_ASAP7_75t_L   g02092(.A1(new_n2230), .A2(new_n2347), .B(new_n2348), .C(new_n2224), .Y(new_n2349));
  NOR2xp33_ASAP7_75t_L      g02093(.A(new_n2344), .B(new_n2343), .Y(new_n2350));
  AOI21xp33_ASAP7_75t_L     g02094(.A1(new_n2341), .A2(new_n2336), .B(new_n2234), .Y(new_n2351));
  NOR3xp33_ASAP7_75t_L      g02095(.A(new_n2351), .B(new_n2350), .C(new_n2232), .Y(new_n2352));
  A2O1A1Ixp33_ASAP7_75t_L   g02096(.A1(new_n2232), .A2(new_n2346), .B(new_n2352), .C(new_n2224), .Y(new_n2353));
  O2A1O1Ixp33_ASAP7_75t_L   g02097(.A1(new_n2224), .A2(new_n2349), .B(new_n2353), .C(new_n2219), .Y(new_n2354));
  O2A1O1Ixp33_ASAP7_75t_L   g02098(.A1(new_n2020), .A2(new_n2024), .B(new_n2221), .C(new_n2167), .Y(new_n2355));
  OAI21xp33_ASAP7_75t_L     g02099(.A1(new_n2350), .A2(new_n2351), .B(new_n2232), .Y(new_n2356));
  NAND2xp33_ASAP7_75t_L     g02100(.A(new_n2356), .B(new_n2348), .Y(new_n2357));
  O2A1O1Ixp33_ASAP7_75t_L   g02101(.A1(new_n2355), .A2(new_n2174), .B(new_n2183), .C(new_n2357), .Y(new_n2358));
  A2O1A1Ixp33_ASAP7_75t_L   g02102(.A1(new_n2028), .A2(new_n2037), .B(new_n2043), .C(new_n2069), .Y(new_n2359));
  AOI221xp5_ASAP7_75t_L     g02103(.A1(new_n2348), .A2(new_n2356), .B1(new_n2182), .B2(new_n2359), .C(new_n2223), .Y(new_n2360));
  OAI21xp33_ASAP7_75t_L     g02104(.A1(new_n2360), .A2(new_n2358), .B(new_n2219), .Y(new_n2361));
  AOI21xp33_ASAP7_75t_L     g02105(.A1(new_n2199), .A2(\a[2] ), .B(new_n2196), .Y(new_n2362));
  MAJIxp5_ASAP7_75t_L       g02106(.A(new_n2201), .B(new_n2184), .C(new_n2362), .Y(new_n2363));
  INVx1_ASAP7_75t_L         g02107(.A(new_n2363), .Y(new_n2364));
  O2A1O1Ixp33_ASAP7_75t_L   g02108(.A1(new_n2219), .A2(new_n2354), .B(new_n2361), .C(new_n2364), .Y(new_n2365));
  O2A1O1Ixp33_ASAP7_75t_L   g02109(.A1(new_n2228), .A2(new_n2229), .B(new_n2346), .C(new_n2352), .Y(new_n2366));
  A2O1A1Ixp33_ASAP7_75t_L   g02110(.A1(new_n2182), .A2(new_n2359), .B(new_n2223), .C(new_n2366), .Y(new_n2367));
  INVx1_ASAP7_75t_L         g02111(.A(new_n2219), .Y(new_n2368));
  NAND3xp33_ASAP7_75t_L     g02112(.A(new_n2367), .B(new_n2353), .C(new_n2368), .Y(new_n2369));
  NAND2xp33_ASAP7_75t_L     g02113(.A(new_n2361), .B(new_n2369), .Y(new_n2370));
  NOR2xp33_ASAP7_75t_L      g02114(.A(new_n2370), .B(new_n2363), .Y(new_n2371));
  NOR2xp33_ASAP7_75t_L      g02115(.A(new_n2371), .B(new_n2365), .Y(\f[24] ));
  O2A1O1Ixp33_ASAP7_75t_L   g02116(.A1(new_n2198), .A2(new_n2202), .B(new_n2370), .C(new_n2354), .Y(new_n2373));
  NOR2xp33_ASAP7_75t_L      g02117(.A(new_n2188), .B(new_n287), .Y(new_n2374));
  AOI221xp5_ASAP7_75t_L     g02118(.A1(\b[24] ), .A2(new_n264), .B1(\b[25] ), .B2(new_n283), .C(new_n2374), .Y(new_n2375));
  NOR2xp33_ASAP7_75t_L      g02119(.A(\b[24] ), .B(\b[25] ), .Y(new_n2376));
  INVx1_ASAP7_75t_L         g02120(.A(\b[25] ), .Y(new_n2377));
  NOR2xp33_ASAP7_75t_L      g02121(.A(new_n2205), .B(new_n2377), .Y(new_n2378));
  NOR2xp33_ASAP7_75t_L      g02122(.A(new_n2376), .B(new_n2378), .Y(new_n2379));
  INVx1_ASAP7_75t_L         g02123(.A(new_n2379), .Y(new_n2380));
  O2A1O1Ixp33_ASAP7_75t_L   g02124(.A1(new_n2188), .A2(new_n2205), .B(new_n2213), .C(new_n2380), .Y(new_n2381));
  INVx1_ASAP7_75t_L         g02125(.A(new_n2381), .Y(new_n2382));
  A2O1A1O1Ixp25_ASAP7_75t_L g02126(.A1(new_n2190), .A2(new_n2209), .B(new_n2189), .C(new_n2212), .D(new_n2211), .Y(new_n2383));
  NAND2xp33_ASAP7_75t_L     g02127(.A(new_n2380), .B(new_n2383), .Y(new_n2384));
  NAND2xp33_ASAP7_75t_L     g02128(.A(new_n2384), .B(new_n2382), .Y(new_n2385));
  O2A1O1Ixp33_ASAP7_75t_L   g02129(.A1(new_n279), .A2(new_n2385), .B(new_n2375), .C(new_n257), .Y(new_n2386));
  NOR2xp33_ASAP7_75t_L      g02130(.A(new_n257), .B(new_n2386), .Y(new_n2387));
  O2A1O1Ixp33_ASAP7_75t_L   g02131(.A1(new_n279), .A2(new_n2385), .B(new_n2375), .C(\a[2] ), .Y(new_n2388));
  NOR2xp33_ASAP7_75t_L      g02132(.A(new_n2388), .B(new_n2387), .Y(new_n2389));
  NOR3xp33_ASAP7_75t_L      g02133(.A(new_n2322), .B(new_n2327), .C(new_n2335), .Y(new_n2390));
  A2O1A1O1Ixp25_ASAP7_75t_L g02134(.A1(new_n2163), .A2(new_n2165), .B(new_n2166), .C(new_n2336), .D(new_n2390), .Y(new_n2391));
  NAND2xp33_ASAP7_75t_L     g02135(.A(new_n2267), .B(new_n2263), .Y(new_n2392));
  MAJIxp5_ASAP7_75t_L       g02136(.A(new_n2283), .B(new_n2273), .C(new_n2392), .Y(new_n2393));
  NOR2xp33_ASAP7_75t_L      g02137(.A(new_n448), .B(new_n1518), .Y(new_n2394));
  AOI221xp5_ASAP7_75t_L     g02138(.A1(\b[5] ), .A2(new_n1659), .B1(\b[6] ), .B2(new_n1507), .C(new_n2394), .Y(new_n2395));
  O2A1O1Ixp33_ASAP7_75t_L   g02139(.A1(new_n1521), .A2(new_n456), .B(new_n2395), .C(new_n1501), .Y(new_n2396));
  OAI21xp33_ASAP7_75t_L     g02140(.A1(new_n1521), .A2(new_n456), .B(new_n2395), .Y(new_n2397));
  NAND2xp33_ASAP7_75t_L     g02141(.A(new_n1501), .B(new_n2397), .Y(new_n2398));
  OAI21xp33_ASAP7_75t_L     g02142(.A1(new_n1501), .A2(new_n2396), .B(new_n2398), .Y(new_n2399));
  MAJIxp5_ASAP7_75t_L       g02143(.A(new_n2266), .B(new_n2112), .C(new_n2252), .Y(new_n2400));
  NOR2xp33_ASAP7_75t_L      g02144(.A(new_n301), .B(new_n1962), .Y(new_n2401));
  AOI221xp5_ASAP7_75t_L     g02145(.A1(new_n1955), .A2(\b[4] ), .B1(new_n2093), .B2(\b[2] ), .C(new_n2401), .Y(new_n2402));
  OAI211xp5_ASAP7_75t_L     g02146(.A1(new_n1497), .A2(new_n1956), .B(new_n2402), .C(\a[23] ), .Y(new_n2403));
  NAND2xp33_ASAP7_75t_L     g02147(.A(\b[4] ), .B(new_n1955), .Y(new_n2404));
  OAI221xp5_ASAP7_75t_L     g02148(.A1(new_n1962), .A2(new_n301), .B1(new_n289), .B2(new_n2089), .C(new_n2404), .Y(new_n2405));
  A2O1A1Ixp33_ASAP7_75t_L   g02149(.A1(new_n342), .A2(new_n1964), .B(new_n2405), .C(new_n1952), .Y(new_n2406));
  INVx1_ASAP7_75t_L         g02150(.A(\a[25] ), .Y(new_n2407));
  NOR2xp33_ASAP7_75t_L      g02151(.A(\a[24] ), .B(new_n2407), .Y(new_n2408));
  NOR2xp33_ASAP7_75t_L      g02152(.A(\a[25] ), .B(new_n2247), .Y(new_n2409));
  OAI21xp33_ASAP7_75t_L     g02153(.A1(new_n2408), .A2(new_n2409), .B(new_n2250), .Y(new_n2410));
  NAND2xp33_ASAP7_75t_L     g02154(.A(new_n2249), .B(new_n2248), .Y(new_n2411));
  NAND2xp33_ASAP7_75t_L     g02155(.A(\a[26] ), .B(new_n2407), .Y(new_n2412));
  INVx1_ASAP7_75t_L         g02156(.A(\a[26] ), .Y(new_n2413));
  NAND2xp33_ASAP7_75t_L     g02157(.A(\a[25] ), .B(new_n2413), .Y(new_n2414));
  NAND3xp33_ASAP7_75t_L     g02158(.A(new_n2411), .B(new_n2412), .C(new_n2414), .Y(new_n2415));
  OAI22xp33_ASAP7_75t_L     g02159(.A1(new_n2410), .A2(new_n284), .B1(new_n262), .B2(new_n2415), .Y(new_n2416));
  AOI21xp33_ASAP7_75t_L     g02160(.A1(new_n2414), .A2(new_n2412), .B(new_n2250), .Y(new_n2417));
  AOI21xp33_ASAP7_75t_L     g02161(.A1(new_n275), .A2(new_n2417), .B(new_n2416), .Y(new_n2418));
  NAND3xp33_ASAP7_75t_L     g02162(.A(new_n2418), .B(new_n2252), .C(\a[26] ), .Y(new_n2419));
  NOR2xp33_ASAP7_75t_L      g02163(.A(new_n2408), .B(new_n2409), .Y(new_n2420));
  NOR2xp33_ASAP7_75t_L      g02164(.A(new_n2411), .B(new_n2420), .Y(new_n2421));
  NAND2xp33_ASAP7_75t_L     g02165(.A(new_n2414), .B(new_n2412), .Y(new_n2422));
  NOR2xp33_ASAP7_75t_L      g02166(.A(new_n2422), .B(new_n2250), .Y(new_n2423));
  AOI22xp33_ASAP7_75t_L     g02167(.A1(new_n2421), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n2423), .Y(new_n2424));
  INVx1_ASAP7_75t_L         g02168(.A(new_n2417), .Y(new_n2425));
  O2A1O1Ixp33_ASAP7_75t_L   g02169(.A1(new_n2425), .A2(new_n274), .B(new_n2424), .C(new_n2413), .Y(new_n2426));
  A2O1A1Ixp33_ASAP7_75t_L   g02170(.A1(new_n2417), .A2(new_n275), .B(new_n2416), .C(new_n2413), .Y(new_n2427));
  A2O1A1Ixp33_ASAP7_75t_L   g02171(.A1(new_n2426), .A2(new_n2251), .B(new_n2413), .C(new_n2427), .Y(new_n2428));
  NAND4xp25_ASAP7_75t_L     g02172(.A(new_n2428), .B(new_n2403), .C(new_n2406), .D(new_n2419), .Y(new_n2429));
  INVx1_ASAP7_75t_L         g02173(.A(new_n2429), .Y(new_n2430));
  AOI22xp33_ASAP7_75t_L     g02174(.A1(new_n2403), .A2(new_n2406), .B1(new_n2419), .B2(new_n2428), .Y(new_n2431));
  OAI21xp33_ASAP7_75t_L     g02175(.A1(new_n2431), .A2(new_n2430), .B(new_n2400), .Y(new_n2432));
  MAJIxp5_ASAP7_75t_L       g02176(.A(new_n2262), .B(new_n2251), .C(new_n2099), .Y(new_n2433));
  AOI211xp5_ASAP7_75t_L     g02177(.A1(new_n342), .A2(new_n1964), .B(new_n1952), .C(new_n2405), .Y(new_n2434));
  O2A1O1Ixp33_ASAP7_75t_L   g02178(.A1(new_n1956), .A2(new_n1497), .B(new_n2402), .C(\a[23] ), .Y(new_n2435));
  OAI21xp33_ASAP7_75t_L     g02179(.A1(new_n2425), .A2(new_n274), .B(new_n2424), .Y(new_n2436));
  NOR3xp33_ASAP7_75t_L      g02180(.A(new_n2436), .B(new_n2251), .C(new_n2413), .Y(new_n2437));
  A2O1A1Ixp33_ASAP7_75t_L   g02181(.A1(new_n2417), .A2(new_n275), .B(new_n2416), .C(\a[26] ), .Y(new_n2438));
  O2A1O1Ixp33_ASAP7_75t_L   g02182(.A1(new_n2425), .A2(new_n274), .B(new_n2424), .C(\a[26] ), .Y(new_n2439));
  O2A1O1Ixp33_ASAP7_75t_L   g02183(.A1(new_n2252), .A2(new_n2438), .B(\a[26] ), .C(new_n2439), .Y(new_n2440));
  OAI22xp33_ASAP7_75t_L     g02184(.A1(new_n2440), .A2(new_n2437), .B1(new_n2435), .B2(new_n2434), .Y(new_n2441));
  NAND3xp33_ASAP7_75t_L     g02185(.A(new_n2433), .B(new_n2429), .C(new_n2441), .Y(new_n2442));
  NAND3xp33_ASAP7_75t_L     g02186(.A(new_n2432), .B(new_n2399), .C(new_n2442), .Y(new_n2443));
  INVx1_ASAP7_75t_L         g02187(.A(new_n2399), .Y(new_n2444));
  AOI21xp33_ASAP7_75t_L     g02188(.A1(new_n2441), .A2(new_n2429), .B(new_n2433), .Y(new_n2445));
  NAND2xp33_ASAP7_75t_L     g02189(.A(new_n2429), .B(new_n2441), .Y(new_n2446));
  NOR2xp33_ASAP7_75t_L      g02190(.A(new_n2400), .B(new_n2446), .Y(new_n2447));
  OAI21xp33_ASAP7_75t_L     g02191(.A1(new_n2445), .A2(new_n2447), .B(new_n2444), .Y(new_n2448));
  NAND3xp33_ASAP7_75t_L     g02192(.A(new_n2393), .B(new_n2443), .C(new_n2448), .Y(new_n2449));
  OAI22xp33_ASAP7_75t_L     g02193(.A1(new_n2285), .A2(new_n2294), .B1(new_n2106), .B2(new_n2246), .Y(new_n2450));
  NOR3xp33_ASAP7_75t_L      g02194(.A(new_n2444), .B(new_n2445), .C(new_n2447), .Y(new_n2451));
  AOI21xp33_ASAP7_75t_L     g02195(.A1(new_n2432), .A2(new_n2442), .B(new_n2399), .Y(new_n2452));
  OAI211xp5_ASAP7_75t_L     g02196(.A1(new_n2452), .A2(new_n2451), .B(new_n2450), .C(new_n2284), .Y(new_n2453));
  NOR2xp33_ASAP7_75t_L      g02197(.A(new_n680), .B(new_n1284), .Y(new_n2454));
  AOI221xp5_ASAP7_75t_L     g02198(.A1(\b[8] ), .A2(new_n1290), .B1(\b[9] ), .B2(new_n1204), .C(new_n2454), .Y(new_n2455));
  O2A1O1Ixp33_ASAP7_75t_L   g02199(.A1(new_n1210), .A2(new_n1175), .B(new_n2455), .C(new_n1206), .Y(new_n2456));
  OAI21xp33_ASAP7_75t_L     g02200(.A1(new_n1210), .A2(new_n1175), .B(new_n2455), .Y(new_n2457));
  NAND2xp33_ASAP7_75t_L     g02201(.A(new_n1206), .B(new_n2457), .Y(new_n2458));
  OAI21xp33_ASAP7_75t_L     g02202(.A1(new_n1206), .A2(new_n2456), .B(new_n2458), .Y(new_n2459));
  INVx1_ASAP7_75t_L         g02203(.A(new_n2459), .Y(new_n2460));
  NAND3xp33_ASAP7_75t_L     g02204(.A(new_n2460), .B(new_n2449), .C(new_n2453), .Y(new_n2461));
  O2A1O1Ixp33_ASAP7_75t_L   g02205(.A1(new_n2271), .A2(new_n2272), .B(new_n2284), .C(new_n2285), .Y(new_n2462));
  NAND2xp33_ASAP7_75t_L     g02206(.A(new_n2443), .B(new_n2448), .Y(new_n2463));
  O2A1O1Ixp33_ASAP7_75t_L   g02207(.A1(new_n2283), .A2(new_n2462), .B(new_n2284), .C(new_n2463), .Y(new_n2464));
  AOI21xp33_ASAP7_75t_L     g02208(.A1(new_n2448), .A2(new_n2443), .B(new_n2393), .Y(new_n2465));
  OAI21xp33_ASAP7_75t_L     g02209(.A1(new_n2465), .A2(new_n2464), .B(new_n2459), .Y(new_n2466));
  A2O1A1O1Ixp25_ASAP7_75t_L g02210(.A1(new_n2125), .A2(new_n2085), .B(new_n2244), .C(new_n2301), .D(new_n2293), .Y(new_n2467));
  NAND3xp33_ASAP7_75t_L     g02211(.A(new_n2467), .B(new_n2466), .C(new_n2461), .Y(new_n2468));
  NOR3xp33_ASAP7_75t_L      g02212(.A(new_n2464), .B(new_n2465), .C(new_n2459), .Y(new_n2469));
  AOI21xp33_ASAP7_75t_L     g02213(.A1(new_n2449), .A2(new_n2453), .B(new_n2460), .Y(new_n2470));
  OAI21xp33_ASAP7_75t_L     g02214(.A1(new_n2298), .A2(new_n2245), .B(new_n2300), .Y(new_n2471));
  OAI21xp33_ASAP7_75t_L     g02215(.A1(new_n2470), .A2(new_n2469), .B(new_n2471), .Y(new_n2472));
  NOR2xp33_ASAP7_75t_L      g02216(.A(new_n833), .B(new_n864), .Y(new_n2473));
  AOI221xp5_ASAP7_75t_L     g02217(.A1(\b[11] ), .A2(new_n985), .B1(\b[13] ), .B2(new_n886), .C(new_n2473), .Y(new_n2474));
  INVx1_ASAP7_75t_L         g02218(.A(new_n2474), .Y(new_n2475));
  A2O1A1Ixp33_ASAP7_75t_L   g02219(.A1(new_n1166), .A2(new_n873), .B(new_n2475), .C(\a[14] ), .Y(new_n2476));
  O2A1O1Ixp33_ASAP7_75t_L   g02220(.A1(new_n872), .A2(new_n942), .B(new_n2474), .C(\a[14] ), .Y(new_n2477));
  AO21x2_ASAP7_75t_L        g02221(.A1(\a[14] ), .A2(new_n2476), .B(new_n2477), .Y(new_n2478));
  AOI21xp33_ASAP7_75t_L     g02222(.A1(new_n2472), .A2(new_n2468), .B(new_n2478), .Y(new_n2479));
  NOR3xp33_ASAP7_75t_L      g02223(.A(new_n2471), .B(new_n2470), .C(new_n2469), .Y(new_n2480));
  AOI21xp33_ASAP7_75t_L     g02224(.A1(new_n2466), .A2(new_n2461), .B(new_n2467), .Y(new_n2481));
  AOI21xp33_ASAP7_75t_L     g02225(.A1(new_n2476), .A2(\a[14] ), .B(new_n2477), .Y(new_n2482));
  NOR3xp33_ASAP7_75t_L      g02226(.A(new_n2480), .B(new_n2481), .C(new_n2482), .Y(new_n2483));
  A2O1A1O1Ixp25_ASAP7_75t_L g02227(.A1(new_n2129), .A2(new_n2078), .B(new_n2135), .C(new_n2303), .D(new_n2304), .Y(new_n2484));
  OR3x1_ASAP7_75t_L         g02228(.A(new_n2484), .B(new_n2479), .C(new_n2483), .Y(new_n2485));
  OAI21xp33_ASAP7_75t_L     g02229(.A1(new_n2479), .A2(new_n2483), .B(new_n2484), .Y(new_n2486));
  NOR2xp33_ASAP7_75t_L      g02230(.A(new_n1043), .B(new_n1550), .Y(new_n2487));
  AOI221xp5_ASAP7_75t_L     g02231(.A1(\b[14] ), .A2(new_n713), .B1(\b[16] ), .B2(new_n640), .C(new_n2487), .Y(new_n2488));
  INVx1_ASAP7_75t_L         g02232(.A(new_n2488), .Y(new_n2489));
  A2O1A1Ixp33_ASAP7_75t_L   g02233(.A1(new_n1156), .A2(new_n718), .B(new_n2489), .C(\a[11] ), .Y(new_n2490));
  AOI211xp5_ASAP7_75t_L     g02234(.A1(new_n1156), .A2(new_n718), .B(new_n2489), .C(new_n637), .Y(new_n2491));
  A2O1A1O1Ixp25_ASAP7_75t_L g02235(.A1(new_n1156), .A2(new_n718), .B(new_n2489), .C(new_n2490), .D(new_n2491), .Y(new_n2492));
  NAND3xp33_ASAP7_75t_L     g02236(.A(new_n2485), .B(new_n2486), .C(new_n2492), .Y(new_n2493));
  NOR3xp33_ASAP7_75t_L      g02237(.A(new_n2484), .B(new_n2483), .C(new_n2479), .Y(new_n2494));
  OAI21xp33_ASAP7_75t_L     g02238(.A1(new_n2481), .A2(new_n2480), .B(new_n2482), .Y(new_n2495));
  NAND3xp33_ASAP7_75t_L     g02239(.A(new_n2468), .B(new_n2472), .C(new_n2478), .Y(new_n2496));
  AOI221xp5_ASAP7_75t_L     g02240(.A1(new_n2237), .A2(new_n2303), .B1(new_n2496), .B2(new_n2495), .C(new_n2304), .Y(new_n2497));
  O2A1O1Ixp33_ASAP7_75t_L   g02241(.A1(new_n641), .A2(new_n1161), .B(new_n2488), .C(\a[11] ), .Y(new_n2498));
  OAI22xp33_ASAP7_75t_L     g02242(.A1(new_n2494), .A2(new_n2497), .B1(new_n2498), .B2(new_n2491), .Y(new_n2499));
  AND2x2_ASAP7_75t_L        g02243(.A(new_n2499), .B(new_n2493), .Y(new_n2500));
  INVx1_ASAP7_75t_L         g02244(.A(new_n2315), .Y(new_n2501));
  O2A1O1Ixp33_ASAP7_75t_L   g02245(.A1(new_n2313), .A2(new_n637), .B(new_n2501), .C(new_n2310), .Y(new_n2502));
  O2A1O1Ixp33_ASAP7_75t_L   g02246(.A1(new_n2316), .A2(new_n2317), .B(new_n2321), .C(new_n2502), .Y(new_n2503));
  NAND2xp33_ASAP7_75t_L     g02247(.A(new_n2503), .B(new_n2500), .Y(new_n2504));
  NOR2xp33_ASAP7_75t_L      g02248(.A(new_n2497), .B(new_n2494), .Y(new_n2505));
  A2O1A1Ixp33_ASAP7_75t_L   g02249(.A1(\a[11] ), .A2(new_n2490), .B(new_n2498), .C(new_n2505), .Y(new_n2506));
  INVx1_ASAP7_75t_L         g02250(.A(new_n2499), .Y(new_n2507));
  NAND3xp33_ASAP7_75t_L     g02251(.A(new_n2306), .B(new_n2316), .C(new_n2309), .Y(new_n2508));
  A2O1A1Ixp33_ASAP7_75t_L   g02252(.A1(new_n2318), .A2(new_n2323), .B(new_n2326), .C(new_n2508), .Y(new_n2509));
  A2O1A1Ixp33_ASAP7_75t_L   g02253(.A1(new_n2506), .A2(new_n2505), .B(new_n2507), .C(new_n2509), .Y(new_n2510));
  NOR2xp33_ASAP7_75t_L      g02254(.A(new_n1458), .B(new_n513), .Y(new_n2511));
  AOI221xp5_ASAP7_75t_L     g02255(.A1(\b[17] ), .A2(new_n560), .B1(\b[19] ), .B2(new_n475), .C(new_n2511), .Y(new_n2512));
  INVx1_ASAP7_75t_L         g02256(.A(new_n2512), .Y(new_n2513));
  A2O1A1Ixp33_ASAP7_75t_L   g02257(.A1(new_n1607), .A2(new_n483), .B(new_n2513), .C(\a[8] ), .Y(new_n2514));
  O2A1O1Ixp33_ASAP7_75t_L   g02258(.A1(new_n477), .A2(new_n1628), .B(new_n2512), .C(\a[8] ), .Y(new_n2515));
  AOI21xp33_ASAP7_75t_L     g02259(.A1(new_n2514), .A2(\a[8] ), .B(new_n2515), .Y(new_n2516));
  NAND3xp33_ASAP7_75t_L     g02260(.A(new_n2504), .B(new_n2510), .C(new_n2516), .Y(new_n2517));
  AO21x2_ASAP7_75t_L        g02261(.A1(new_n2510), .A2(new_n2504), .B(new_n2516), .Y(new_n2518));
  AOI21xp33_ASAP7_75t_L     g02262(.A1(new_n2518), .A2(new_n2517), .B(new_n2391), .Y(new_n2519));
  NAND2xp33_ASAP7_75t_L     g02263(.A(new_n2517), .B(new_n2518), .Y(new_n2520));
  NAND2xp33_ASAP7_75t_L     g02264(.A(new_n2391), .B(new_n2520), .Y(new_n2521));
  NAND2xp33_ASAP7_75t_L     g02265(.A(new_n2055), .B(new_n2053), .Y(new_n2522));
  NOR2xp33_ASAP7_75t_L      g02266(.A(new_n1745), .B(new_n375), .Y(new_n2523));
  AOI221xp5_ASAP7_75t_L     g02267(.A1(\b[22] ), .A2(new_n361), .B1(new_n349), .B2(\b[21] ), .C(new_n2523), .Y(new_n2524));
  O2A1O1Ixp33_ASAP7_75t_L   g02268(.A1(new_n356), .A2(new_n2522), .B(new_n2524), .C(new_n346), .Y(new_n2525));
  INVx1_ASAP7_75t_L         g02269(.A(new_n2525), .Y(new_n2526));
  O2A1O1Ixp33_ASAP7_75t_L   g02270(.A1(new_n356), .A2(new_n2522), .B(new_n2524), .C(\a[5] ), .Y(new_n2527));
  AO21x2_ASAP7_75t_L        g02271(.A1(\a[5] ), .A2(new_n2526), .B(new_n2527), .Y(new_n2528));
  O2A1O1Ixp33_ASAP7_75t_L   g02272(.A1(new_n2391), .A2(new_n2519), .B(new_n2521), .C(new_n2528), .Y(new_n2529));
  NAND2xp33_ASAP7_75t_L     g02273(.A(new_n2499), .B(new_n2493), .Y(new_n2530));
  XNOR2x2_ASAP7_75t_L       g02274(.A(new_n2530), .B(new_n2509), .Y(new_n2531));
  NOR2xp33_ASAP7_75t_L      g02275(.A(new_n2516), .B(new_n2531), .Y(new_n2532));
  INVx1_ASAP7_75t_L         g02276(.A(new_n2391), .Y(new_n2533));
  O2A1O1Ixp33_ASAP7_75t_L   g02277(.A1(new_n2516), .A2(new_n2532), .B(new_n2517), .C(new_n2533), .Y(new_n2534));
  NOR2xp33_ASAP7_75t_L      g02278(.A(new_n2391), .B(new_n2520), .Y(new_n2535));
  AOI21xp33_ASAP7_75t_L     g02279(.A1(new_n2526), .A2(\a[5] ), .B(new_n2527), .Y(new_n2536));
  NOR3xp33_ASAP7_75t_L      g02280(.A(new_n2535), .B(new_n2536), .C(new_n2534), .Y(new_n2537));
  NOR2xp33_ASAP7_75t_L      g02281(.A(new_n2537), .B(new_n2529), .Y(new_n2538));
  O2A1O1Ixp33_ASAP7_75t_L   g02282(.A1(new_n2224), .A2(new_n2366), .B(new_n2346), .C(new_n2538), .Y(new_n2539));
  A2O1A1Ixp33_ASAP7_75t_L   g02283(.A1(new_n2356), .A2(new_n2348), .B(new_n2224), .C(new_n2346), .Y(new_n2540));
  INVx1_ASAP7_75t_L         g02284(.A(new_n2519), .Y(new_n2541));
  A2O1A1Ixp33_ASAP7_75t_L   g02285(.A1(new_n2541), .A2(new_n2520), .B(new_n2535), .C(new_n2536), .Y(new_n2542));
  OAI211xp5_ASAP7_75t_L     g02286(.A1(new_n2519), .A2(new_n2391), .B(new_n2521), .C(new_n2528), .Y(new_n2543));
  NAND2xp33_ASAP7_75t_L     g02287(.A(new_n2543), .B(new_n2542), .Y(new_n2544));
  NOR2xp33_ASAP7_75t_L      g02288(.A(new_n2540), .B(new_n2544), .Y(new_n2545));
  NOR3xp33_ASAP7_75t_L      g02289(.A(new_n2539), .B(new_n2545), .C(new_n2389), .Y(new_n2546));
  INVx1_ASAP7_75t_L         g02290(.A(new_n2546), .Y(new_n2547));
  OAI21xp33_ASAP7_75t_L     g02291(.A1(new_n2545), .A2(new_n2539), .B(new_n2389), .Y(new_n2548));
  NAND2xp33_ASAP7_75t_L     g02292(.A(new_n2548), .B(new_n2547), .Y(new_n2549));
  XOR2x2_ASAP7_75t_L        g02293(.A(new_n2549), .B(new_n2373), .Y(\f[25] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02294(.A1(new_n2182), .A2(new_n2359), .B(new_n2223), .C(new_n2357), .D(new_n2347), .Y(new_n2551));
  O2A1O1Ixp33_ASAP7_75t_L   g02295(.A1(new_n2391), .A2(new_n2519), .B(new_n2521), .C(new_n2536), .Y(new_n2552));
  INVx1_ASAP7_75t_L         g02296(.A(new_n2552), .Y(new_n2553));
  NAND2xp33_ASAP7_75t_L     g02297(.A(new_n2486), .B(new_n2485), .Y(new_n2554));
  INVx1_ASAP7_75t_L         g02298(.A(new_n2490), .Y(new_n2555));
  INVx1_ASAP7_75t_L         g02299(.A(new_n2498), .Y(new_n2556));
  O2A1O1Ixp33_ASAP7_75t_L   g02300(.A1(new_n2555), .A2(new_n637), .B(new_n2556), .C(new_n2554), .Y(new_n2557));
  A2O1A1O1Ixp25_ASAP7_75t_L g02301(.A1(new_n2303), .A2(new_n2237), .B(new_n2304), .C(new_n2495), .D(new_n2483), .Y(new_n2558));
  XNOR2x2_ASAP7_75t_L       g02302(.A(new_n2393), .B(new_n2463), .Y(new_n2559));
  MAJIxp5_ASAP7_75t_L       g02303(.A(new_n2471), .B(new_n2459), .C(new_n2559), .Y(new_n2560));
  NOR2xp33_ASAP7_75t_L      g02304(.A(new_n680), .B(new_n2118), .Y(new_n2561));
  AOI221xp5_ASAP7_75t_L     g02305(.A1(\b[9] ), .A2(new_n1290), .B1(\b[11] ), .B2(new_n1209), .C(new_n2561), .Y(new_n2562));
  O2A1O1Ixp33_ASAP7_75t_L   g02306(.A1(new_n1210), .A2(new_n754), .B(new_n2562), .C(new_n1206), .Y(new_n2563));
  INVx1_ASAP7_75t_L         g02307(.A(new_n2562), .Y(new_n2564));
  A2O1A1Ixp33_ASAP7_75t_L   g02308(.A1(new_n976), .A2(new_n1216), .B(new_n2564), .C(new_n1206), .Y(new_n2565));
  OAI21xp33_ASAP7_75t_L     g02309(.A1(new_n1206), .A2(new_n2563), .B(new_n2565), .Y(new_n2566));
  A2O1A1Ixp33_ASAP7_75t_L   g02310(.A1(new_n2450), .A2(new_n2284), .B(new_n2452), .C(new_n2443), .Y(new_n2567));
  A2O1A1Ixp33_ASAP7_75t_L   g02311(.A1(new_n342), .A2(new_n1964), .B(new_n2405), .C(\a[23] ), .Y(new_n2568));
  INVx1_ASAP7_75t_L         g02312(.A(new_n2568), .Y(new_n2569));
  NAND2xp33_ASAP7_75t_L     g02313(.A(new_n2419), .B(new_n2428), .Y(new_n2570));
  O2A1O1Ixp33_ASAP7_75t_L   g02314(.A1(new_n1952), .A2(new_n2569), .B(new_n2406), .C(new_n2570), .Y(new_n2571));
  NAND3xp33_ASAP7_75t_L     g02315(.A(new_n2250), .B(new_n2420), .C(new_n2422), .Y(new_n2572));
  NAND2xp33_ASAP7_75t_L     g02316(.A(\b[1] ), .B(new_n2421), .Y(new_n2573));
  OAI221xp5_ASAP7_75t_L     g02317(.A1(new_n2415), .A2(new_n289), .B1(new_n284), .B2(new_n2572), .C(new_n2573), .Y(new_n2574));
  A2O1A1Ixp33_ASAP7_75t_L   g02318(.A1(new_n294), .A2(new_n2417), .B(new_n2574), .C(\a[26] ), .Y(new_n2575));
  NOR2xp33_ASAP7_75t_L      g02319(.A(new_n289), .B(new_n2415), .Y(new_n2576));
  AND3x1_ASAP7_75t_L        g02320(.A(new_n2250), .B(new_n2422), .C(new_n2420), .Y(new_n2577));
  AOI221xp5_ASAP7_75t_L     g02321(.A1(new_n2421), .A2(\b[1] ), .B1(new_n2577), .B2(\b[0] ), .C(new_n2576), .Y(new_n2578));
  O2A1O1Ixp33_ASAP7_75t_L   g02322(.A1(new_n509), .A2(new_n2425), .B(new_n2578), .C(\a[26] ), .Y(new_n2579));
  A2O1A1O1Ixp25_ASAP7_75t_L g02323(.A1(new_n2418), .A2(new_n2252), .B(new_n2575), .C(\a[26] ), .D(new_n2579), .Y(new_n2580));
  NAND2xp33_ASAP7_75t_L     g02324(.A(new_n2417), .B(new_n294), .Y(new_n2581));
  INVx1_ASAP7_75t_L         g02325(.A(new_n2581), .Y(new_n2582));
  NOR5xp2_ASAP7_75t_L       g02326(.A(new_n2436), .B(new_n2574), .C(new_n2582), .D(new_n2251), .E(new_n2413), .Y(new_n2583));
  NAND2xp33_ASAP7_75t_L     g02327(.A(\b[5] ), .B(new_n1955), .Y(new_n2584));
  OAI221xp5_ASAP7_75t_L     g02328(.A1(new_n1962), .A2(new_n332), .B1(new_n301), .B2(new_n2089), .C(new_n2584), .Y(new_n2585));
  A2O1A1Ixp33_ASAP7_75t_L   g02329(.A1(new_n394), .A2(new_n1964), .B(new_n2585), .C(\a[23] ), .Y(new_n2586));
  NOR2xp33_ASAP7_75t_L      g02330(.A(new_n332), .B(new_n1962), .Y(new_n2587));
  AOI221xp5_ASAP7_75t_L     g02331(.A1(new_n1955), .A2(\b[5] ), .B1(new_n2093), .B2(\b[3] ), .C(new_n2587), .Y(new_n2588));
  O2A1O1Ixp33_ASAP7_75t_L   g02332(.A1(new_n728), .A2(new_n1956), .B(new_n2588), .C(\a[23] ), .Y(new_n2589));
  AOI21xp33_ASAP7_75t_L     g02333(.A1(new_n2586), .A2(\a[23] ), .B(new_n2589), .Y(new_n2590));
  NOR3xp33_ASAP7_75t_L      g02334(.A(new_n2590), .B(new_n2580), .C(new_n2583), .Y(new_n2591));
  NAND3xp33_ASAP7_75t_L     g02335(.A(new_n2578), .B(\a[26] ), .C(new_n2581), .Y(new_n2592));
  A2O1A1Ixp33_ASAP7_75t_L   g02336(.A1(new_n294), .A2(new_n2417), .B(new_n2574), .C(new_n2413), .Y(new_n2593));
  NAND3xp33_ASAP7_75t_L     g02337(.A(new_n2419), .B(new_n2592), .C(new_n2593), .Y(new_n2594));
  NAND5xp2_ASAP7_75t_L      g02338(.A(\a[26] ), .B(new_n2418), .C(new_n2581), .D(new_n2578), .E(new_n2252), .Y(new_n2595));
  AOI221xp5_ASAP7_75t_L     g02339(.A1(new_n2586), .A2(\a[23] ), .B1(new_n2595), .B2(new_n2594), .C(new_n2589), .Y(new_n2596));
  OAI22xp33_ASAP7_75t_L     g02340(.A1(new_n2445), .A2(new_n2571), .B1(new_n2596), .B2(new_n2591), .Y(new_n2597));
  NOR2xp33_ASAP7_75t_L      g02341(.A(new_n2437), .B(new_n2440), .Y(new_n2598));
  A2O1A1Ixp33_ASAP7_75t_L   g02342(.A1(new_n2568), .A2(\a[23] ), .B(new_n2435), .C(new_n2598), .Y(new_n2599));
  OR3x1_ASAP7_75t_L         g02343(.A(new_n2590), .B(new_n2580), .C(new_n2583), .Y(new_n2600));
  OAI21xp33_ASAP7_75t_L     g02344(.A1(new_n2583), .A2(new_n2580), .B(new_n2590), .Y(new_n2601));
  NAND4xp25_ASAP7_75t_L     g02345(.A(new_n2432), .B(new_n2601), .C(new_n2600), .D(new_n2599), .Y(new_n2602));
  NOR2xp33_ASAP7_75t_L      g02346(.A(new_n448), .B(new_n1517), .Y(new_n2603));
  AOI221xp5_ASAP7_75t_L     g02347(.A1(\b[6] ), .A2(new_n1659), .B1(\b[8] ), .B2(new_n1511), .C(new_n2603), .Y(new_n2604));
  O2A1O1Ixp33_ASAP7_75t_L   g02348(.A1(new_n1521), .A2(new_n540), .B(new_n2604), .C(new_n1501), .Y(new_n2605));
  NOR2xp33_ASAP7_75t_L      g02349(.A(new_n1501), .B(new_n2605), .Y(new_n2606));
  O2A1O1Ixp33_ASAP7_75t_L   g02350(.A1(new_n1521), .A2(new_n540), .B(new_n2604), .C(\a[20] ), .Y(new_n2607));
  NOR2xp33_ASAP7_75t_L      g02351(.A(new_n2607), .B(new_n2606), .Y(new_n2608));
  NAND3xp33_ASAP7_75t_L     g02352(.A(new_n2602), .B(new_n2608), .C(new_n2597), .Y(new_n2609));
  AOI21xp33_ASAP7_75t_L     g02353(.A1(new_n2602), .A2(new_n2597), .B(new_n2608), .Y(new_n2610));
  INVx1_ASAP7_75t_L         g02354(.A(new_n2610), .Y(new_n2611));
  NAND3xp33_ASAP7_75t_L     g02355(.A(new_n2567), .B(new_n2611), .C(new_n2609), .Y(new_n2612));
  AO21x2_ASAP7_75t_L        g02356(.A1(new_n2609), .A2(new_n2611), .B(new_n2567), .Y(new_n2613));
  AOI21xp33_ASAP7_75t_L     g02357(.A1(new_n2613), .A2(new_n2612), .B(new_n2566), .Y(new_n2614));
  AND3x1_ASAP7_75t_L        g02358(.A(new_n2613), .B(new_n2612), .C(new_n2566), .Y(new_n2615));
  NOR3xp33_ASAP7_75t_L      g02359(.A(new_n2560), .B(new_n2614), .C(new_n2615), .Y(new_n2616));
  NAND2xp33_ASAP7_75t_L     g02360(.A(new_n2453), .B(new_n2449), .Y(new_n2617));
  MAJIxp5_ASAP7_75t_L       g02361(.A(new_n2467), .B(new_n2617), .C(new_n2460), .Y(new_n2618));
  AO21x2_ASAP7_75t_L        g02362(.A1(new_n2612), .A2(new_n2613), .B(new_n2566), .Y(new_n2619));
  NAND3xp33_ASAP7_75t_L     g02363(.A(new_n2613), .B(new_n2612), .C(new_n2566), .Y(new_n2620));
  AOI21xp33_ASAP7_75t_L     g02364(.A1(new_n2619), .A2(new_n2620), .B(new_n2618), .Y(new_n2621));
  NOR2xp33_ASAP7_75t_L      g02365(.A(new_n936), .B(new_n864), .Y(new_n2622));
  AOI221xp5_ASAP7_75t_L     g02366(.A1(\b[12] ), .A2(new_n985), .B1(\b[14] ), .B2(new_n886), .C(new_n2622), .Y(new_n2623));
  O2A1O1Ixp33_ASAP7_75t_L   g02367(.A1(new_n872), .A2(new_n1268), .B(new_n2623), .C(new_n867), .Y(new_n2624));
  INVx1_ASAP7_75t_L         g02368(.A(new_n2623), .Y(new_n2625));
  A2O1A1Ixp33_ASAP7_75t_L   g02369(.A1(new_n971), .A2(new_n873), .B(new_n2625), .C(new_n867), .Y(new_n2626));
  OAI21xp33_ASAP7_75t_L     g02370(.A1(new_n867), .A2(new_n2624), .B(new_n2626), .Y(new_n2627));
  NOR3xp33_ASAP7_75t_L      g02371(.A(new_n2616), .B(new_n2621), .C(new_n2627), .Y(new_n2628));
  NAND3xp33_ASAP7_75t_L     g02372(.A(new_n2618), .B(new_n2619), .C(new_n2620), .Y(new_n2629));
  OAI21xp33_ASAP7_75t_L     g02373(.A1(new_n2614), .A2(new_n2615), .B(new_n2560), .Y(new_n2630));
  A2O1A1Ixp33_ASAP7_75t_L   g02374(.A1(new_n971), .A2(new_n873), .B(new_n2625), .C(\a[14] ), .Y(new_n2631));
  O2A1O1Ixp33_ASAP7_75t_L   g02375(.A1(new_n872), .A2(new_n1268), .B(new_n2623), .C(\a[14] ), .Y(new_n2632));
  AOI21xp33_ASAP7_75t_L     g02376(.A1(new_n2631), .A2(\a[14] ), .B(new_n2632), .Y(new_n2633));
  AOI21xp33_ASAP7_75t_L     g02377(.A1(new_n2629), .A2(new_n2630), .B(new_n2633), .Y(new_n2634));
  NOR3xp33_ASAP7_75t_L      g02378(.A(new_n2558), .B(new_n2628), .C(new_n2634), .Y(new_n2635));
  OAI21xp33_ASAP7_75t_L     g02379(.A1(new_n2479), .A2(new_n2484), .B(new_n2496), .Y(new_n2636));
  NAND3xp33_ASAP7_75t_L     g02380(.A(new_n2629), .B(new_n2630), .C(new_n2633), .Y(new_n2637));
  OAI21xp33_ASAP7_75t_L     g02381(.A1(new_n2621), .A2(new_n2616), .B(new_n2627), .Y(new_n2638));
  AOI21xp33_ASAP7_75t_L     g02382(.A1(new_n2638), .A2(new_n2637), .B(new_n2636), .Y(new_n2639));
  NOR2xp33_ASAP7_75t_L      g02383(.A(new_n1150), .B(new_n1550), .Y(new_n2640));
  AOI221xp5_ASAP7_75t_L     g02384(.A1(\b[15] ), .A2(new_n713), .B1(\b[17] ), .B2(new_n640), .C(new_n2640), .Y(new_n2641));
  O2A1O1Ixp33_ASAP7_75t_L   g02385(.A1(new_n641), .A2(new_n1356), .B(new_n2641), .C(new_n637), .Y(new_n2642));
  INVx1_ASAP7_75t_L         g02386(.A(new_n2641), .Y(new_n2643));
  A2O1A1Ixp33_ASAP7_75t_L   g02387(.A1(new_n1633), .A2(new_n718), .B(new_n2643), .C(new_n637), .Y(new_n2644));
  OAI21xp33_ASAP7_75t_L     g02388(.A1(new_n637), .A2(new_n2642), .B(new_n2644), .Y(new_n2645));
  OAI21xp33_ASAP7_75t_L     g02389(.A1(new_n2639), .A2(new_n2635), .B(new_n2645), .Y(new_n2646));
  NAND3xp33_ASAP7_75t_L     g02390(.A(new_n2636), .B(new_n2637), .C(new_n2638), .Y(new_n2647));
  OAI21xp33_ASAP7_75t_L     g02391(.A1(new_n2634), .A2(new_n2628), .B(new_n2558), .Y(new_n2648));
  A2O1A1Ixp33_ASAP7_75t_L   g02392(.A1(new_n1633), .A2(new_n718), .B(new_n2643), .C(\a[11] ), .Y(new_n2649));
  O2A1O1Ixp33_ASAP7_75t_L   g02393(.A1(new_n641), .A2(new_n1356), .B(new_n2641), .C(\a[11] ), .Y(new_n2650));
  AOI21xp33_ASAP7_75t_L     g02394(.A1(new_n2649), .A2(\a[11] ), .B(new_n2650), .Y(new_n2651));
  NAND3xp33_ASAP7_75t_L     g02395(.A(new_n2647), .B(new_n2651), .C(new_n2648), .Y(new_n2652));
  AOI221xp5_ASAP7_75t_L     g02396(.A1(new_n2652), .A2(new_n2646), .B1(new_n2530), .B2(new_n2509), .C(new_n2557), .Y(new_n2653));
  NAND2xp33_ASAP7_75t_L     g02397(.A(new_n2652), .B(new_n2646), .Y(new_n2654));
  O2A1O1Ixp33_ASAP7_75t_L   g02398(.A1(new_n2503), .A2(new_n2500), .B(new_n2506), .C(new_n2654), .Y(new_n2655));
  NOR2xp33_ASAP7_75t_L      g02399(.A(new_n1599), .B(new_n513), .Y(new_n2656));
  AOI221xp5_ASAP7_75t_L     g02400(.A1(\b[18] ), .A2(new_n560), .B1(\b[20] ), .B2(new_n475), .C(new_n2656), .Y(new_n2657));
  INVx1_ASAP7_75t_L         g02401(.A(new_n2657), .Y(new_n2658));
  A2O1A1Ixp33_ASAP7_75t_L   g02402(.A1(new_n1752), .A2(new_n483), .B(new_n2658), .C(\a[8] ), .Y(new_n2659));
  INVx1_ASAP7_75t_L         g02403(.A(new_n2659), .Y(new_n2660));
  A2O1A1Ixp33_ASAP7_75t_L   g02404(.A1(new_n1752), .A2(new_n483), .B(new_n2658), .C(new_n466), .Y(new_n2661));
  OAI21xp33_ASAP7_75t_L     g02405(.A1(new_n466), .A2(new_n2660), .B(new_n2661), .Y(new_n2662));
  NOR3xp33_ASAP7_75t_L      g02406(.A(new_n2662), .B(new_n2655), .C(new_n2653), .Y(new_n2663));
  OAI211xp5_ASAP7_75t_L     g02407(.A1(new_n2500), .A2(new_n2503), .B(new_n2654), .C(new_n2506), .Y(new_n2664));
  AOI21xp33_ASAP7_75t_L     g02408(.A1(new_n2647), .A2(new_n2648), .B(new_n2651), .Y(new_n2665));
  NOR3xp33_ASAP7_75t_L      g02409(.A(new_n2635), .B(new_n2639), .C(new_n2645), .Y(new_n2666));
  NOR2xp33_ASAP7_75t_L      g02410(.A(new_n2665), .B(new_n2666), .Y(new_n2667));
  A2O1A1Ixp33_ASAP7_75t_L   g02411(.A1(new_n2530), .A2(new_n2509), .B(new_n2557), .C(new_n2667), .Y(new_n2668));
  INVx1_ASAP7_75t_L         g02412(.A(new_n2661), .Y(new_n2669));
  AOI21xp33_ASAP7_75t_L     g02413(.A1(new_n2659), .A2(\a[8] ), .B(new_n2669), .Y(new_n2670));
  AOI21xp33_ASAP7_75t_L     g02414(.A1(new_n2668), .A2(new_n2664), .B(new_n2670), .Y(new_n2671));
  NOR2xp33_ASAP7_75t_L      g02415(.A(new_n2671), .B(new_n2663), .Y(new_n2672));
  MAJx2_ASAP7_75t_L         g02416(.A(new_n2391), .B(new_n2516), .C(new_n2531), .Y(new_n2673));
  NAND2xp33_ASAP7_75t_L     g02417(.A(new_n2672), .B(new_n2673), .Y(new_n2674));
  NAND3xp33_ASAP7_75t_L     g02418(.A(new_n2668), .B(new_n2664), .C(new_n2670), .Y(new_n2675));
  OAI21xp33_ASAP7_75t_L     g02419(.A1(new_n2653), .A2(new_n2655), .B(new_n2662), .Y(new_n2676));
  NAND2xp33_ASAP7_75t_L     g02420(.A(new_n2676), .B(new_n2675), .Y(new_n2677));
  A2O1A1Ixp33_ASAP7_75t_L   g02421(.A1(new_n2520), .A2(new_n2533), .B(new_n2532), .C(new_n2677), .Y(new_n2678));
  AND2x2_ASAP7_75t_L        g02422(.A(new_n2191), .B(new_n2193), .Y(new_n2679));
  NOR2xp33_ASAP7_75t_L      g02423(.A(new_n1895), .B(new_n375), .Y(new_n2680));
  AOI221xp5_ASAP7_75t_L     g02424(.A1(\b[23] ), .A2(new_n361), .B1(new_n349), .B2(\b[22] ), .C(new_n2680), .Y(new_n2681));
  INVx1_ASAP7_75t_L         g02425(.A(new_n2681), .Y(new_n2682));
  A2O1A1Ixp33_ASAP7_75t_L   g02426(.A1(new_n2679), .A2(new_n359), .B(new_n2682), .C(\a[5] ), .Y(new_n2683));
  NAND2xp33_ASAP7_75t_L     g02427(.A(\a[5] ), .B(new_n2683), .Y(new_n2684));
  O2A1O1Ixp33_ASAP7_75t_L   g02428(.A1(new_n356), .A2(new_n2194), .B(new_n2681), .C(\a[5] ), .Y(new_n2685));
  INVx1_ASAP7_75t_L         g02429(.A(new_n2685), .Y(new_n2686));
  NAND4xp25_ASAP7_75t_L     g02430(.A(new_n2674), .B(new_n2678), .C(new_n2686), .D(new_n2684), .Y(new_n2687));
  MAJIxp5_ASAP7_75t_L       g02431(.A(new_n2391), .B(new_n2516), .C(new_n2531), .Y(new_n2688));
  NOR2xp33_ASAP7_75t_L      g02432(.A(new_n2688), .B(new_n2677), .Y(new_n2689));
  NOR2xp33_ASAP7_75t_L      g02433(.A(new_n2672), .B(new_n2673), .Y(new_n2690));
  O2A1O1Ixp33_ASAP7_75t_L   g02434(.A1(new_n356), .A2(new_n2194), .B(new_n2681), .C(new_n346), .Y(new_n2691));
  OAI21xp33_ASAP7_75t_L     g02435(.A1(new_n346), .A2(new_n2691), .B(new_n2686), .Y(new_n2692));
  OAI21xp33_ASAP7_75t_L     g02436(.A1(new_n2689), .A2(new_n2690), .B(new_n2692), .Y(new_n2693));
  NAND2xp33_ASAP7_75t_L     g02437(.A(new_n2687), .B(new_n2693), .Y(new_n2694));
  O2A1O1Ixp33_ASAP7_75t_L   g02438(.A1(new_n2551), .A2(new_n2538), .B(new_n2553), .C(new_n2694), .Y(new_n2695));
  A2O1A1Ixp33_ASAP7_75t_L   g02439(.A1(new_n2542), .A2(new_n2543), .B(new_n2551), .C(new_n2553), .Y(new_n2696));
  NAND2xp33_ASAP7_75t_L     g02440(.A(new_n2678), .B(new_n2674), .Y(new_n2697));
  O2A1O1Ixp33_ASAP7_75t_L   g02441(.A1(new_n2691), .A2(new_n346), .B(new_n2686), .C(new_n2697), .Y(new_n2698));
  O2A1O1Ixp33_ASAP7_75t_L   g02442(.A1(new_n2697), .A2(new_n2698), .B(new_n2693), .C(new_n2696), .Y(new_n2699));
  NOR2xp33_ASAP7_75t_L      g02443(.A(new_n2205), .B(new_n287), .Y(new_n2700));
  AOI221xp5_ASAP7_75t_L     g02444(.A1(\b[25] ), .A2(new_n264), .B1(\b[26] ), .B2(new_n283), .C(new_n2700), .Y(new_n2701));
  NOR2xp33_ASAP7_75t_L      g02445(.A(\b[25] ), .B(\b[26] ), .Y(new_n2702));
  INVx1_ASAP7_75t_L         g02446(.A(\b[26] ), .Y(new_n2703));
  NOR2xp33_ASAP7_75t_L      g02447(.A(new_n2377), .B(new_n2703), .Y(new_n2704));
  NOR2xp33_ASAP7_75t_L      g02448(.A(new_n2702), .B(new_n2704), .Y(new_n2705));
  A2O1A1Ixp33_ASAP7_75t_L   g02449(.A1(\b[25] ), .A2(\b[24] ), .B(new_n2381), .C(new_n2705), .Y(new_n2706));
  OR3x1_ASAP7_75t_L         g02450(.A(new_n2381), .B(new_n2378), .C(new_n2705), .Y(new_n2707));
  NAND2xp33_ASAP7_75t_L     g02451(.A(new_n2706), .B(new_n2707), .Y(new_n2708));
  INVx1_ASAP7_75t_L         g02452(.A(new_n2708), .Y(new_n2709));
  NAND2xp33_ASAP7_75t_L     g02453(.A(new_n273), .B(new_n2709), .Y(new_n2710));
  O2A1O1Ixp33_ASAP7_75t_L   g02454(.A1(new_n279), .A2(new_n2708), .B(new_n2701), .C(new_n257), .Y(new_n2711));
  OAI211xp5_ASAP7_75t_L     g02455(.A1(new_n279), .A2(new_n2708), .B(new_n2701), .C(\a[2] ), .Y(new_n2712));
  A2O1A1Ixp33_ASAP7_75t_L   g02456(.A1(new_n2710), .A2(new_n2701), .B(new_n2711), .C(new_n2712), .Y(new_n2713));
  OAI21xp33_ASAP7_75t_L     g02457(.A1(new_n2695), .A2(new_n2699), .B(new_n2713), .Y(new_n2714));
  INVx1_ASAP7_75t_L         g02458(.A(new_n2714), .Y(new_n2715));
  NOR3xp33_ASAP7_75t_L      g02459(.A(new_n2699), .B(new_n2695), .C(new_n2713), .Y(new_n2716));
  NOR2xp33_ASAP7_75t_L      g02460(.A(new_n2716), .B(new_n2715), .Y(new_n2717));
  INVx1_ASAP7_75t_L         g02461(.A(new_n2717), .Y(new_n2718));
  O2A1O1Ixp33_ASAP7_75t_L   g02462(.A1(new_n2373), .A2(new_n2549), .B(new_n2547), .C(new_n2718), .Y(new_n2719));
  A2O1A1O1Ixp25_ASAP7_75t_L g02463(.A1(new_n2370), .A2(new_n2363), .B(new_n2354), .C(new_n2548), .D(new_n2546), .Y(new_n2720));
  INVx1_ASAP7_75t_L         g02464(.A(new_n2720), .Y(new_n2721));
  NOR2xp33_ASAP7_75t_L      g02465(.A(new_n2721), .B(new_n2717), .Y(new_n2722));
  NOR2xp33_ASAP7_75t_L      g02466(.A(new_n2722), .B(new_n2719), .Y(\f[26] ));
  NAND2xp33_ASAP7_75t_L     g02467(.A(new_n2664), .B(new_n2668), .Y(new_n2724));
  O2A1O1Ixp33_ASAP7_75t_L   g02468(.A1(new_n2660), .A2(new_n466), .B(new_n2661), .C(new_n2724), .Y(new_n2725));
  NAND2xp33_ASAP7_75t_L     g02469(.A(new_n2459), .B(new_n2559), .Y(new_n2726));
  A2O1A1Ixp33_ASAP7_75t_L   g02470(.A1(new_n2472), .A2(new_n2726), .B(new_n2614), .C(new_n2620), .Y(new_n2727));
  NOR2xp33_ASAP7_75t_L      g02471(.A(new_n748), .B(new_n2118), .Y(new_n2728));
  AOI221xp5_ASAP7_75t_L     g02472(.A1(\b[10] ), .A2(new_n1290), .B1(\b[12] ), .B2(new_n1209), .C(new_n2728), .Y(new_n2729));
  INVx1_ASAP7_75t_L         g02473(.A(new_n2729), .Y(new_n2730));
  A2O1A1Ixp33_ASAP7_75t_L   g02474(.A1(new_n1057), .A2(new_n1216), .B(new_n2730), .C(\a[17] ), .Y(new_n2731));
  O2A1O1Ixp33_ASAP7_75t_L   g02475(.A1(new_n1210), .A2(new_n841), .B(new_n2729), .C(\a[17] ), .Y(new_n2732));
  AOI21xp33_ASAP7_75t_L     g02476(.A1(new_n2731), .A2(\a[17] ), .B(new_n2732), .Y(new_n2733));
  A2O1A1O1Ixp25_ASAP7_75t_L g02477(.A1(new_n2448), .A2(new_n2393), .B(new_n2451), .C(new_n2609), .D(new_n2610), .Y(new_n2734));
  A2O1A1O1Ixp25_ASAP7_75t_L g02478(.A1(new_n2429), .A2(new_n2441), .B(new_n2433), .C(new_n2599), .D(new_n2596), .Y(new_n2735));
  INVx1_ASAP7_75t_L         g02479(.A(\a[27] ), .Y(new_n2736));
  NAND2xp33_ASAP7_75t_L     g02480(.A(\a[26] ), .B(new_n2736), .Y(new_n2737));
  NAND2xp33_ASAP7_75t_L     g02481(.A(\a[27] ), .B(new_n2413), .Y(new_n2738));
  AND2x2_ASAP7_75t_L        g02482(.A(new_n2737), .B(new_n2738), .Y(new_n2739));
  NOR2xp33_ASAP7_75t_L      g02483(.A(new_n284), .B(new_n2739), .Y(new_n2740));
  INVx1_ASAP7_75t_L         g02484(.A(new_n2740), .Y(new_n2741));
  A2O1A1O1Ixp25_ASAP7_75t_L g02485(.A1(\a[26] ), .A2(new_n2575), .B(new_n2579), .C(new_n2437), .D(new_n2741), .Y(new_n2742));
  NOR2xp33_ASAP7_75t_L      g02486(.A(new_n2740), .B(new_n2595), .Y(new_n2743));
  NAND2xp33_ASAP7_75t_L     g02487(.A(\b[3] ), .B(new_n2423), .Y(new_n2744));
  NAND2xp33_ASAP7_75t_L     g02488(.A(\b[1] ), .B(new_n2577), .Y(new_n2745));
  NAND2xp33_ASAP7_75t_L     g02489(.A(\b[2] ), .B(new_n2421), .Y(new_n2746));
  NAND2xp33_ASAP7_75t_L     g02490(.A(new_n2417), .B(new_n312), .Y(new_n2747));
  NAND5xp2_ASAP7_75t_L      g02491(.A(new_n2747), .B(new_n2746), .C(new_n2745), .D(new_n2744), .E(\a[26] ), .Y(new_n2748));
  OAI211xp5_ASAP7_75t_L     g02492(.A1(new_n2572), .A2(new_n262), .B(new_n2744), .C(new_n2746), .Y(new_n2749));
  A2O1A1Ixp33_ASAP7_75t_L   g02493(.A1(new_n312), .A2(new_n2417), .B(new_n2749), .C(new_n2413), .Y(new_n2750));
  NAND2xp33_ASAP7_75t_L     g02494(.A(new_n2748), .B(new_n2750), .Y(new_n2751));
  OAI21xp33_ASAP7_75t_L     g02495(.A1(new_n2743), .A2(new_n2742), .B(new_n2751), .Y(new_n2752));
  A2O1A1Ixp33_ASAP7_75t_L   g02496(.A1(new_n2592), .A2(new_n2593), .B(new_n2419), .C(new_n2740), .Y(new_n2753));
  NAND2xp33_ASAP7_75t_L     g02497(.A(new_n2741), .B(new_n2583), .Y(new_n2754));
  AND2x2_ASAP7_75t_L        g02498(.A(new_n2748), .B(new_n2750), .Y(new_n2755));
  NAND3xp33_ASAP7_75t_L     g02499(.A(new_n2754), .B(new_n2755), .C(new_n2753), .Y(new_n2756));
  NOR2xp33_ASAP7_75t_L      g02500(.A(new_n384), .B(new_n1962), .Y(new_n2757));
  AOI221xp5_ASAP7_75t_L     g02501(.A1(new_n1955), .A2(\b[6] ), .B1(new_n2093), .B2(\b[4] ), .C(new_n2757), .Y(new_n2758));
  O2A1O1Ixp33_ASAP7_75t_L   g02502(.A1(new_n1956), .A2(new_n434), .B(new_n2758), .C(new_n1952), .Y(new_n2759));
  OAI31xp33_ASAP7_75t_L     g02503(.A1(new_n433), .A2(new_n431), .A3(new_n1956), .B(new_n2758), .Y(new_n2760));
  NAND2xp33_ASAP7_75t_L     g02504(.A(new_n1952), .B(new_n2760), .Y(new_n2761));
  OA21x2_ASAP7_75t_L        g02505(.A1(new_n1952), .A2(new_n2759), .B(new_n2761), .Y(new_n2762));
  NAND3xp33_ASAP7_75t_L     g02506(.A(new_n2752), .B(new_n2762), .C(new_n2756), .Y(new_n2763));
  AOI21xp33_ASAP7_75t_L     g02507(.A1(new_n2752), .A2(new_n2756), .B(new_n2762), .Y(new_n2764));
  INVx1_ASAP7_75t_L         g02508(.A(new_n2764), .Y(new_n2765));
  OAI211xp5_ASAP7_75t_L     g02509(.A1(new_n2591), .A2(new_n2735), .B(new_n2765), .C(new_n2763), .Y(new_n2766));
  A2O1A1O1Ixp25_ASAP7_75t_L g02510(.A1(new_n2400), .A2(new_n2446), .B(new_n2571), .C(new_n2601), .D(new_n2591), .Y(new_n2767));
  OAI21xp33_ASAP7_75t_L     g02511(.A1(new_n1952), .A2(new_n2759), .B(new_n2761), .Y(new_n2768));
  NAND3xp33_ASAP7_75t_L     g02512(.A(new_n2752), .B(new_n2756), .C(new_n2768), .Y(new_n2769));
  AOI21xp33_ASAP7_75t_L     g02513(.A1(new_n2754), .A2(new_n2753), .B(new_n2755), .Y(new_n2770));
  NOR3xp33_ASAP7_75t_L      g02514(.A(new_n2742), .B(new_n2743), .C(new_n2751), .Y(new_n2771));
  NOR3xp33_ASAP7_75t_L      g02515(.A(new_n2771), .B(new_n2770), .C(new_n2768), .Y(new_n2772));
  A2O1A1Ixp33_ASAP7_75t_L   g02516(.A1(new_n2768), .A2(new_n2769), .B(new_n2772), .C(new_n2767), .Y(new_n2773));
  NOR2xp33_ASAP7_75t_L      g02517(.A(new_n534), .B(new_n1517), .Y(new_n2774));
  AOI221xp5_ASAP7_75t_L     g02518(.A1(\b[7] ), .A2(new_n1659), .B1(\b[9] ), .B2(new_n1511), .C(new_n2774), .Y(new_n2775));
  INVx1_ASAP7_75t_L         g02519(.A(new_n2775), .Y(new_n2776));
  A2O1A1Ixp33_ASAP7_75t_L   g02520(.A1(new_n602), .A2(new_n1513), .B(new_n2776), .C(\a[20] ), .Y(new_n2777));
  NAND2xp33_ASAP7_75t_L     g02521(.A(\a[20] ), .B(new_n2777), .Y(new_n2778));
  A2O1A1Ixp33_ASAP7_75t_L   g02522(.A1(new_n602), .A2(new_n1513), .B(new_n2776), .C(new_n1501), .Y(new_n2779));
  AOI22xp33_ASAP7_75t_L     g02523(.A1(new_n2778), .A2(new_n2779), .B1(new_n2773), .B2(new_n2766), .Y(new_n2780));
  NOR3xp33_ASAP7_75t_L      g02524(.A(new_n2767), .B(new_n2772), .C(new_n2764), .Y(new_n2781));
  OA21x2_ASAP7_75t_L        g02525(.A1(new_n2772), .A2(new_n2764), .B(new_n2767), .Y(new_n2782));
  O2A1O1Ixp33_ASAP7_75t_L   g02526(.A1(new_n1521), .A2(new_n1066), .B(new_n2775), .C(new_n1501), .Y(new_n2783));
  OAI21xp33_ASAP7_75t_L     g02527(.A1(new_n1501), .A2(new_n2783), .B(new_n2779), .Y(new_n2784));
  NOR3xp33_ASAP7_75t_L      g02528(.A(new_n2782), .B(new_n2784), .C(new_n2781), .Y(new_n2785));
  NOR3xp33_ASAP7_75t_L      g02529(.A(new_n2734), .B(new_n2780), .C(new_n2785), .Y(new_n2786));
  OAI21xp33_ASAP7_75t_L     g02530(.A1(new_n2781), .A2(new_n2782), .B(new_n2784), .Y(new_n2787));
  NAND4xp25_ASAP7_75t_L     g02531(.A(new_n2766), .B(new_n2773), .C(new_n2779), .D(new_n2778), .Y(new_n2788));
  AOI221xp5_ASAP7_75t_L     g02532(.A1(new_n2567), .A2(new_n2609), .B1(new_n2787), .B2(new_n2788), .C(new_n2610), .Y(new_n2789));
  OAI21xp33_ASAP7_75t_L     g02533(.A1(new_n2786), .A2(new_n2789), .B(new_n2733), .Y(new_n2790));
  NOR3xp33_ASAP7_75t_L      g02534(.A(new_n2789), .B(new_n2786), .C(new_n2733), .Y(new_n2791));
  INVx1_ASAP7_75t_L         g02535(.A(new_n2791), .Y(new_n2792));
  NAND3xp33_ASAP7_75t_L     g02536(.A(new_n2727), .B(new_n2790), .C(new_n2792), .Y(new_n2793));
  AOI21xp33_ASAP7_75t_L     g02537(.A1(new_n2618), .A2(new_n2619), .B(new_n2615), .Y(new_n2794));
  INVx1_ASAP7_75t_L         g02538(.A(new_n2790), .Y(new_n2795));
  OAI21xp33_ASAP7_75t_L     g02539(.A1(new_n2795), .A2(new_n2791), .B(new_n2794), .Y(new_n2796));
  NOR2xp33_ASAP7_75t_L      g02540(.A(new_n960), .B(new_n864), .Y(new_n2797));
  AOI221xp5_ASAP7_75t_L     g02541(.A1(\b[13] ), .A2(new_n985), .B1(\b[15] ), .B2(new_n886), .C(new_n2797), .Y(new_n2798));
  INVx1_ASAP7_75t_L         g02542(.A(new_n2798), .Y(new_n2799));
  A2O1A1Ixp33_ASAP7_75t_L   g02543(.A1(new_n1052), .A2(new_n873), .B(new_n2799), .C(\a[14] ), .Y(new_n2800));
  O2A1O1Ixp33_ASAP7_75t_L   g02544(.A1(new_n872), .A2(new_n1774), .B(new_n2798), .C(\a[14] ), .Y(new_n2801));
  AOI21xp33_ASAP7_75t_L     g02545(.A1(new_n2800), .A2(\a[14] ), .B(new_n2801), .Y(new_n2802));
  NAND3xp33_ASAP7_75t_L     g02546(.A(new_n2793), .B(new_n2802), .C(new_n2796), .Y(new_n2803));
  NOR3xp33_ASAP7_75t_L      g02547(.A(new_n2794), .B(new_n2795), .C(new_n2791), .Y(new_n2804));
  AOI21xp33_ASAP7_75t_L     g02548(.A1(new_n2792), .A2(new_n2790), .B(new_n2727), .Y(new_n2805));
  O2A1O1Ixp33_ASAP7_75t_L   g02549(.A1(new_n872), .A2(new_n1774), .B(new_n2798), .C(new_n867), .Y(new_n2806));
  A2O1A1Ixp33_ASAP7_75t_L   g02550(.A1(new_n1052), .A2(new_n873), .B(new_n2799), .C(new_n867), .Y(new_n2807));
  OAI21xp33_ASAP7_75t_L     g02551(.A1(new_n867), .A2(new_n2806), .B(new_n2807), .Y(new_n2808));
  OAI21xp33_ASAP7_75t_L     g02552(.A1(new_n2805), .A2(new_n2804), .B(new_n2808), .Y(new_n2809));
  NOR2xp33_ASAP7_75t_L      g02553(.A(new_n2621), .B(new_n2616), .Y(new_n2810));
  MAJIxp5_ASAP7_75t_L       g02554(.A(new_n2636), .B(new_n2627), .C(new_n2810), .Y(new_n2811));
  NAND3xp33_ASAP7_75t_L     g02555(.A(new_n2811), .B(new_n2809), .C(new_n2803), .Y(new_n2812));
  NOR3xp33_ASAP7_75t_L      g02556(.A(new_n2804), .B(new_n2805), .C(new_n2808), .Y(new_n2813));
  AOI21xp33_ASAP7_75t_L     g02557(.A1(new_n2793), .A2(new_n2796), .B(new_n2802), .Y(new_n2814));
  NAND2xp33_ASAP7_75t_L     g02558(.A(new_n2630), .B(new_n2629), .Y(new_n2815));
  MAJIxp5_ASAP7_75t_L       g02559(.A(new_n2558), .B(new_n2633), .C(new_n2815), .Y(new_n2816));
  OAI21xp33_ASAP7_75t_L     g02560(.A1(new_n2814), .A2(new_n2813), .B(new_n2816), .Y(new_n2817));
  NOR2xp33_ASAP7_75t_L      g02561(.A(new_n1349), .B(new_n1550), .Y(new_n2818));
  AOI221xp5_ASAP7_75t_L     g02562(.A1(\b[16] ), .A2(new_n713), .B1(\b[18] ), .B2(new_n640), .C(new_n2818), .Y(new_n2819));
  INVx1_ASAP7_75t_L         g02563(.A(new_n2819), .Y(new_n2820));
  A2O1A1Ixp33_ASAP7_75t_L   g02564(.A1(new_n2329), .A2(new_n718), .B(new_n2820), .C(\a[11] ), .Y(new_n2821));
  O2A1O1Ixp33_ASAP7_75t_L   g02565(.A1(new_n641), .A2(new_n1464), .B(new_n2819), .C(\a[11] ), .Y(new_n2822));
  AOI21xp33_ASAP7_75t_L     g02566(.A1(new_n2821), .A2(\a[11] ), .B(new_n2822), .Y(new_n2823));
  NAND3xp33_ASAP7_75t_L     g02567(.A(new_n2812), .B(new_n2817), .C(new_n2823), .Y(new_n2824));
  NOR3xp33_ASAP7_75t_L      g02568(.A(new_n2816), .B(new_n2814), .C(new_n2813), .Y(new_n2825));
  AOI21xp33_ASAP7_75t_L     g02569(.A1(new_n2809), .A2(new_n2803), .B(new_n2811), .Y(new_n2826));
  O2A1O1Ixp33_ASAP7_75t_L   g02570(.A1(new_n641), .A2(new_n1464), .B(new_n2819), .C(new_n637), .Y(new_n2827));
  A2O1A1Ixp33_ASAP7_75t_L   g02571(.A1(new_n2329), .A2(new_n718), .B(new_n2820), .C(new_n637), .Y(new_n2828));
  OAI21xp33_ASAP7_75t_L     g02572(.A1(new_n637), .A2(new_n2827), .B(new_n2828), .Y(new_n2829));
  OAI21xp33_ASAP7_75t_L     g02573(.A1(new_n2826), .A2(new_n2825), .B(new_n2829), .Y(new_n2830));
  A2O1A1O1Ixp25_ASAP7_75t_L g02574(.A1(new_n2530), .A2(new_n2509), .B(new_n2557), .C(new_n2652), .D(new_n2665), .Y(new_n2831));
  NAND3xp33_ASAP7_75t_L     g02575(.A(new_n2831), .B(new_n2830), .C(new_n2824), .Y(new_n2832));
  A2O1A1Ixp33_ASAP7_75t_L   g02576(.A1(new_n2492), .A2(new_n2493), .B(new_n2503), .C(new_n2506), .Y(new_n2833));
  NAND2xp33_ASAP7_75t_L     g02577(.A(new_n2824), .B(new_n2830), .Y(new_n2834));
  A2O1A1Ixp33_ASAP7_75t_L   g02578(.A1(new_n2667), .A2(new_n2833), .B(new_n2665), .C(new_n2834), .Y(new_n2835));
  AND2x2_ASAP7_75t_L        g02579(.A(new_n1898), .B(new_n1900), .Y(new_n2836));
  NOR2xp33_ASAP7_75t_L      g02580(.A(new_n1745), .B(new_n513), .Y(new_n2837));
  AOI221xp5_ASAP7_75t_L     g02581(.A1(\b[19] ), .A2(new_n560), .B1(\b[21] ), .B2(new_n475), .C(new_n2837), .Y(new_n2838));
  INVx1_ASAP7_75t_L         g02582(.A(new_n2838), .Y(new_n2839));
  A2O1A1Ixp33_ASAP7_75t_L   g02583(.A1(new_n2836), .A2(new_n483), .B(new_n2839), .C(\a[8] ), .Y(new_n2840));
  O2A1O1Ixp33_ASAP7_75t_L   g02584(.A1(new_n477), .A2(new_n1901), .B(new_n2838), .C(\a[8] ), .Y(new_n2841));
  AO21x2_ASAP7_75t_L        g02585(.A1(\a[8] ), .A2(new_n2840), .B(new_n2841), .Y(new_n2842));
  AOI21xp33_ASAP7_75t_L     g02586(.A1(new_n2835), .A2(new_n2832), .B(new_n2842), .Y(new_n2843));
  NOR3xp33_ASAP7_75t_L      g02587(.A(new_n2834), .B(new_n2655), .C(new_n2665), .Y(new_n2844));
  AOI21xp33_ASAP7_75t_L     g02588(.A1(new_n2830), .A2(new_n2824), .B(new_n2831), .Y(new_n2845));
  AOI21xp33_ASAP7_75t_L     g02589(.A1(new_n2840), .A2(\a[8] ), .B(new_n2841), .Y(new_n2846));
  NOR3xp33_ASAP7_75t_L      g02590(.A(new_n2844), .B(new_n2845), .C(new_n2846), .Y(new_n2847));
  NOR2xp33_ASAP7_75t_L      g02591(.A(new_n2843), .B(new_n2847), .Y(new_n2848));
  A2O1A1Ixp33_ASAP7_75t_L   g02592(.A1(new_n2677), .A2(new_n2688), .B(new_n2725), .C(new_n2848), .Y(new_n2849));
  NOR2xp33_ASAP7_75t_L      g02593(.A(new_n2653), .B(new_n2655), .Y(new_n2850));
  MAJIxp5_ASAP7_75t_L       g02594(.A(new_n2688), .B(new_n2662), .C(new_n2850), .Y(new_n2851));
  OAI21xp33_ASAP7_75t_L     g02595(.A1(new_n2843), .A2(new_n2847), .B(new_n2851), .Y(new_n2852));
  NAND2xp33_ASAP7_75t_L     g02596(.A(new_n2213), .B(new_n2215), .Y(new_n2853));
  NOR2xp33_ASAP7_75t_L      g02597(.A(new_n2045), .B(new_n375), .Y(new_n2854));
  AOI221xp5_ASAP7_75t_L     g02598(.A1(\b[24] ), .A2(new_n361), .B1(new_n349), .B2(\b[23] ), .C(new_n2854), .Y(new_n2855));
  O2A1O1Ixp33_ASAP7_75t_L   g02599(.A1(new_n356), .A2(new_n2853), .B(new_n2855), .C(new_n346), .Y(new_n2856));
  OAI21xp33_ASAP7_75t_L     g02600(.A1(new_n356), .A2(new_n2853), .B(new_n2855), .Y(new_n2857));
  NAND2xp33_ASAP7_75t_L     g02601(.A(new_n346), .B(new_n2857), .Y(new_n2858));
  OA21x2_ASAP7_75t_L        g02602(.A1(new_n346), .A2(new_n2856), .B(new_n2858), .Y(new_n2859));
  NAND3xp33_ASAP7_75t_L     g02603(.A(new_n2849), .B(new_n2852), .C(new_n2859), .Y(new_n2860));
  NOR3xp33_ASAP7_75t_L      g02604(.A(new_n2851), .B(new_n2847), .C(new_n2843), .Y(new_n2861));
  OAI21xp33_ASAP7_75t_L     g02605(.A1(new_n2845), .A2(new_n2844), .B(new_n2846), .Y(new_n2862));
  NAND3xp33_ASAP7_75t_L     g02606(.A(new_n2835), .B(new_n2842), .C(new_n2832), .Y(new_n2863));
  AOI221xp5_ASAP7_75t_L     g02607(.A1(new_n2677), .A2(new_n2688), .B1(new_n2863), .B2(new_n2862), .C(new_n2725), .Y(new_n2864));
  NOR2xp33_ASAP7_75t_L      g02608(.A(new_n346), .B(new_n2857), .Y(new_n2865));
  O2A1O1Ixp33_ASAP7_75t_L   g02609(.A1(new_n356), .A2(new_n2853), .B(new_n2855), .C(\a[5] ), .Y(new_n2866));
  OAI22xp33_ASAP7_75t_L     g02610(.A1(new_n2861), .A2(new_n2864), .B1(new_n2866), .B2(new_n2865), .Y(new_n2867));
  NAND2xp33_ASAP7_75t_L     g02611(.A(new_n2867), .B(new_n2860), .Y(new_n2868));
  O2A1O1Ixp33_ASAP7_75t_L   g02612(.A1(new_n2529), .A2(new_n2537), .B(new_n2540), .C(new_n2552), .Y(new_n2869));
  INVx1_ASAP7_75t_L         g02613(.A(new_n2698), .Y(new_n2870));
  A2O1A1Ixp33_ASAP7_75t_L   g02614(.A1(new_n2687), .A2(new_n2693), .B(new_n2869), .C(new_n2870), .Y(new_n2871));
  NOR2xp33_ASAP7_75t_L      g02615(.A(new_n2868), .B(new_n2871), .Y(new_n2872));
  A2O1A1Ixp33_ASAP7_75t_L   g02616(.A1(new_n2694), .A2(new_n2696), .B(new_n2698), .C(new_n2868), .Y(new_n2873));
  INVx1_ASAP7_75t_L         g02617(.A(new_n2873), .Y(new_n2874));
  NOR2xp33_ASAP7_75t_L      g02618(.A(new_n2377), .B(new_n287), .Y(new_n2875));
  AOI221xp5_ASAP7_75t_L     g02619(.A1(\b[26] ), .A2(new_n264), .B1(\b[27] ), .B2(new_n283), .C(new_n2875), .Y(new_n2876));
  INVx1_ASAP7_75t_L         g02620(.A(new_n2876), .Y(new_n2877));
  NOR2xp33_ASAP7_75t_L      g02621(.A(\b[26] ), .B(\b[27] ), .Y(new_n2878));
  INVx1_ASAP7_75t_L         g02622(.A(\b[27] ), .Y(new_n2879));
  NOR2xp33_ASAP7_75t_L      g02623(.A(new_n2703), .B(new_n2879), .Y(new_n2880));
  NOR2xp33_ASAP7_75t_L      g02624(.A(new_n2878), .B(new_n2880), .Y(new_n2881));
  INVx1_ASAP7_75t_L         g02625(.A(new_n2881), .Y(new_n2882));
  O2A1O1Ixp33_ASAP7_75t_L   g02626(.A1(new_n2377), .A2(new_n2703), .B(new_n2706), .C(new_n2882), .Y(new_n2883));
  INVx1_ASAP7_75t_L         g02627(.A(new_n2883), .Y(new_n2884));
  O2A1O1Ixp33_ASAP7_75t_L   g02628(.A1(new_n2378), .A2(new_n2381), .B(new_n2705), .C(new_n2704), .Y(new_n2885));
  NAND2xp33_ASAP7_75t_L     g02629(.A(new_n2882), .B(new_n2885), .Y(new_n2886));
  AND2x2_ASAP7_75t_L        g02630(.A(new_n2886), .B(new_n2884), .Y(new_n2887));
  A2O1A1Ixp33_ASAP7_75t_L   g02631(.A1(new_n2887), .A2(new_n273), .B(new_n2877), .C(\a[2] ), .Y(new_n2888));
  NAND2xp33_ASAP7_75t_L     g02632(.A(new_n2886), .B(new_n2884), .Y(new_n2889));
  O2A1O1Ixp33_ASAP7_75t_L   g02633(.A1(new_n279), .A2(new_n2889), .B(new_n2876), .C(new_n257), .Y(new_n2890));
  NOR2xp33_ASAP7_75t_L      g02634(.A(new_n257), .B(new_n2890), .Y(new_n2891));
  A2O1A1O1Ixp25_ASAP7_75t_L g02635(.A1(new_n273), .A2(new_n2887), .B(new_n2877), .C(new_n2888), .D(new_n2891), .Y(new_n2892));
  OAI21xp33_ASAP7_75t_L     g02636(.A1(new_n2872), .A2(new_n2874), .B(new_n2892), .Y(new_n2893));
  NOR3xp33_ASAP7_75t_L      g02637(.A(new_n2874), .B(new_n2872), .C(new_n2892), .Y(new_n2894));
  INVx1_ASAP7_75t_L         g02638(.A(new_n2894), .Y(new_n2895));
  NAND2xp33_ASAP7_75t_L     g02639(.A(new_n2893), .B(new_n2895), .Y(new_n2896));
  O2A1O1Ixp33_ASAP7_75t_L   g02640(.A1(new_n2720), .A2(new_n2718), .B(new_n2714), .C(new_n2896), .Y(new_n2897));
  OAI21xp33_ASAP7_75t_L     g02641(.A1(new_n2716), .A2(new_n2720), .B(new_n2714), .Y(new_n2898));
  AOI21xp33_ASAP7_75t_L     g02642(.A1(new_n2895), .A2(new_n2893), .B(new_n2898), .Y(new_n2899));
  NOR2xp33_ASAP7_75t_L      g02643(.A(new_n2899), .B(new_n2897), .Y(\f[27] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02644(.A1(new_n2721), .A2(new_n2717), .B(new_n2715), .C(new_n2893), .D(new_n2894), .Y(new_n2901));
  NOR2xp33_ASAP7_75t_L      g02645(.A(new_n2188), .B(new_n375), .Y(new_n2902));
  AOI221xp5_ASAP7_75t_L     g02646(.A1(\b[25] ), .A2(new_n361), .B1(new_n349), .B2(\b[24] ), .C(new_n2902), .Y(new_n2903));
  O2A1O1Ixp33_ASAP7_75t_L   g02647(.A1(new_n356), .A2(new_n2385), .B(new_n2903), .C(new_n346), .Y(new_n2904));
  NOR2xp33_ASAP7_75t_L      g02648(.A(new_n346), .B(new_n2904), .Y(new_n2905));
  O2A1O1Ixp33_ASAP7_75t_L   g02649(.A1(new_n356), .A2(new_n2385), .B(new_n2903), .C(\a[5] ), .Y(new_n2906));
  NOR2xp33_ASAP7_75t_L      g02650(.A(new_n2906), .B(new_n2905), .Y(new_n2907));
  A2O1A1Ixp33_ASAP7_75t_L   g02651(.A1(new_n2763), .A2(new_n2762), .B(new_n2767), .C(new_n2769), .Y(new_n2908));
  NOR2xp33_ASAP7_75t_L      g02652(.A(new_n427), .B(new_n1962), .Y(new_n2909));
  AOI221xp5_ASAP7_75t_L     g02653(.A1(new_n1955), .A2(\b[7] ), .B1(new_n2093), .B2(\b[5] ), .C(new_n2909), .Y(new_n2910));
  O2A1O1Ixp33_ASAP7_75t_L   g02654(.A1(new_n1956), .A2(new_n456), .B(new_n2910), .C(new_n1952), .Y(new_n2911));
  OAI21xp33_ASAP7_75t_L     g02655(.A1(new_n1956), .A2(new_n456), .B(new_n2910), .Y(new_n2912));
  NAND2xp33_ASAP7_75t_L     g02656(.A(new_n1952), .B(new_n2912), .Y(new_n2913));
  OAI21xp33_ASAP7_75t_L     g02657(.A1(new_n1952), .A2(new_n2911), .B(new_n2913), .Y(new_n2914));
  MAJIxp5_ASAP7_75t_L       g02658(.A(new_n2755), .B(new_n2595), .C(new_n2741), .Y(new_n2915));
  NOR2xp33_ASAP7_75t_L      g02659(.A(new_n332), .B(new_n2415), .Y(new_n2916));
  AOI221xp5_ASAP7_75t_L     g02660(.A1(\b[2] ), .A2(new_n2577), .B1(\b[3] ), .B2(new_n2421), .C(new_n2916), .Y(new_n2917));
  OAI211xp5_ASAP7_75t_L     g02661(.A1(new_n1497), .A2(new_n2425), .B(new_n2917), .C(\a[26] ), .Y(new_n2918));
  NAND2xp33_ASAP7_75t_L     g02662(.A(\b[3] ), .B(new_n2421), .Y(new_n2919));
  OAI221xp5_ASAP7_75t_L     g02663(.A1(new_n2415), .A2(new_n332), .B1(new_n289), .B2(new_n2572), .C(new_n2919), .Y(new_n2920));
  A2O1A1Ixp33_ASAP7_75t_L   g02664(.A1(new_n342), .A2(new_n2417), .B(new_n2920), .C(new_n2413), .Y(new_n2921));
  INVx1_ASAP7_75t_L         g02665(.A(\a[28] ), .Y(new_n2922));
  NOR2xp33_ASAP7_75t_L      g02666(.A(\a[27] ), .B(new_n2922), .Y(new_n2923));
  NOR2xp33_ASAP7_75t_L      g02667(.A(\a[28] ), .B(new_n2736), .Y(new_n2924));
  OAI21xp33_ASAP7_75t_L     g02668(.A1(new_n2923), .A2(new_n2924), .B(new_n2739), .Y(new_n2925));
  NAND2xp33_ASAP7_75t_L     g02669(.A(new_n2738), .B(new_n2737), .Y(new_n2926));
  NAND2xp33_ASAP7_75t_L     g02670(.A(\a[29] ), .B(new_n2922), .Y(new_n2927));
  INVx1_ASAP7_75t_L         g02671(.A(\a[29] ), .Y(new_n2928));
  NAND2xp33_ASAP7_75t_L     g02672(.A(\a[28] ), .B(new_n2928), .Y(new_n2929));
  NAND3xp33_ASAP7_75t_L     g02673(.A(new_n2926), .B(new_n2927), .C(new_n2929), .Y(new_n2930));
  OAI22xp33_ASAP7_75t_L     g02674(.A1(new_n2925), .A2(new_n284), .B1(new_n262), .B2(new_n2930), .Y(new_n2931));
  AOI21xp33_ASAP7_75t_L     g02675(.A1(new_n2929), .A2(new_n2927), .B(new_n2739), .Y(new_n2932));
  AOI21xp33_ASAP7_75t_L     g02676(.A1(new_n275), .A2(new_n2932), .B(new_n2931), .Y(new_n2933));
  NAND3xp33_ASAP7_75t_L     g02677(.A(new_n2933), .B(new_n2741), .C(\a[29] ), .Y(new_n2934));
  NOR2xp33_ASAP7_75t_L      g02678(.A(new_n2923), .B(new_n2924), .Y(new_n2935));
  NOR2xp33_ASAP7_75t_L      g02679(.A(new_n2926), .B(new_n2935), .Y(new_n2936));
  NAND2xp33_ASAP7_75t_L     g02680(.A(new_n2929), .B(new_n2927), .Y(new_n2937));
  NOR2xp33_ASAP7_75t_L      g02681(.A(new_n2937), .B(new_n2739), .Y(new_n2938));
  AOI22xp33_ASAP7_75t_L     g02682(.A1(new_n2936), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n2938), .Y(new_n2939));
  INVx1_ASAP7_75t_L         g02683(.A(new_n2932), .Y(new_n2940));
  O2A1O1Ixp33_ASAP7_75t_L   g02684(.A1(new_n2940), .A2(new_n274), .B(new_n2939), .C(new_n2928), .Y(new_n2941));
  A2O1A1Ixp33_ASAP7_75t_L   g02685(.A1(new_n2932), .A2(new_n275), .B(new_n2931), .C(new_n2928), .Y(new_n2942));
  A2O1A1Ixp33_ASAP7_75t_L   g02686(.A1(new_n2941), .A2(new_n2740), .B(new_n2928), .C(new_n2942), .Y(new_n2943));
  NAND4xp25_ASAP7_75t_L     g02687(.A(new_n2943), .B(new_n2918), .C(new_n2921), .D(new_n2934), .Y(new_n2944));
  AOI211xp5_ASAP7_75t_L     g02688(.A1(new_n342), .A2(new_n2417), .B(new_n2413), .C(new_n2920), .Y(new_n2945));
  O2A1O1Ixp33_ASAP7_75t_L   g02689(.A1(new_n2425), .A2(new_n1497), .B(new_n2917), .C(\a[26] ), .Y(new_n2946));
  NAND2xp33_ASAP7_75t_L     g02690(.A(new_n275), .B(new_n2932), .Y(new_n2947));
  NAND2xp33_ASAP7_75t_L     g02691(.A(new_n2947), .B(new_n2939), .Y(new_n2948));
  NOR3xp33_ASAP7_75t_L      g02692(.A(new_n2948), .B(new_n2740), .C(new_n2928), .Y(new_n2949));
  A2O1A1Ixp33_ASAP7_75t_L   g02693(.A1(new_n2932), .A2(new_n275), .B(new_n2931), .C(\a[29] ), .Y(new_n2950));
  O2A1O1Ixp33_ASAP7_75t_L   g02694(.A1(new_n2940), .A2(new_n274), .B(new_n2939), .C(\a[29] ), .Y(new_n2951));
  O2A1O1Ixp33_ASAP7_75t_L   g02695(.A1(new_n2741), .A2(new_n2950), .B(\a[29] ), .C(new_n2951), .Y(new_n2952));
  OAI22xp33_ASAP7_75t_L     g02696(.A1(new_n2952), .A2(new_n2949), .B1(new_n2946), .B2(new_n2945), .Y(new_n2953));
  NAND2xp33_ASAP7_75t_L     g02697(.A(new_n2944), .B(new_n2953), .Y(new_n2954));
  NAND2xp33_ASAP7_75t_L     g02698(.A(new_n2915), .B(new_n2954), .Y(new_n2955));
  MAJIxp5_ASAP7_75t_L       g02699(.A(new_n2751), .B(new_n2740), .C(new_n2583), .Y(new_n2956));
  NAND3xp33_ASAP7_75t_L     g02700(.A(new_n2956), .B(new_n2944), .C(new_n2953), .Y(new_n2957));
  NAND3xp33_ASAP7_75t_L     g02701(.A(new_n2955), .B(new_n2914), .C(new_n2957), .Y(new_n2958));
  INVx1_ASAP7_75t_L         g02702(.A(new_n2914), .Y(new_n2959));
  AOI21xp33_ASAP7_75t_L     g02703(.A1(new_n2953), .A2(new_n2944), .B(new_n2956), .Y(new_n2960));
  INVx1_ASAP7_75t_L         g02704(.A(new_n2957), .Y(new_n2961));
  OAI21xp33_ASAP7_75t_L     g02705(.A1(new_n2960), .A2(new_n2961), .B(new_n2959), .Y(new_n2962));
  NAND3xp33_ASAP7_75t_L     g02706(.A(new_n2908), .B(new_n2958), .C(new_n2962), .Y(new_n2963));
  OAI22xp33_ASAP7_75t_L     g02707(.A1(new_n2735), .A2(new_n2591), .B1(new_n2764), .B2(new_n2772), .Y(new_n2964));
  NOR3xp33_ASAP7_75t_L      g02708(.A(new_n2961), .B(new_n2959), .C(new_n2960), .Y(new_n2965));
  AOI21xp33_ASAP7_75t_L     g02709(.A1(new_n2955), .A2(new_n2957), .B(new_n2914), .Y(new_n2966));
  OAI211xp5_ASAP7_75t_L     g02710(.A1(new_n2966), .A2(new_n2965), .B(new_n2964), .C(new_n2769), .Y(new_n2967));
  NOR2xp33_ASAP7_75t_L      g02711(.A(new_n680), .B(new_n1518), .Y(new_n2968));
  AOI221xp5_ASAP7_75t_L     g02712(.A1(\b[8] ), .A2(new_n1659), .B1(\b[9] ), .B2(new_n1507), .C(new_n2968), .Y(new_n2969));
  O2A1O1Ixp33_ASAP7_75t_L   g02713(.A1(new_n1521), .A2(new_n1175), .B(new_n2969), .C(new_n1501), .Y(new_n2970));
  OAI21xp33_ASAP7_75t_L     g02714(.A1(new_n1521), .A2(new_n1175), .B(new_n2969), .Y(new_n2971));
  NAND2xp33_ASAP7_75t_L     g02715(.A(new_n1501), .B(new_n2971), .Y(new_n2972));
  OAI21xp33_ASAP7_75t_L     g02716(.A1(new_n1501), .A2(new_n2970), .B(new_n2972), .Y(new_n2973));
  INVx1_ASAP7_75t_L         g02717(.A(new_n2973), .Y(new_n2974));
  NAND3xp33_ASAP7_75t_L     g02718(.A(new_n2963), .B(new_n2974), .C(new_n2967), .Y(new_n2975));
  AOI211xp5_ASAP7_75t_L     g02719(.A1(new_n2964), .A2(new_n2769), .B(new_n2965), .C(new_n2966), .Y(new_n2976));
  AOI21xp33_ASAP7_75t_L     g02720(.A1(new_n2962), .A2(new_n2958), .B(new_n2908), .Y(new_n2977));
  OAI21xp33_ASAP7_75t_L     g02721(.A1(new_n2977), .A2(new_n2976), .B(new_n2973), .Y(new_n2978));
  A2O1A1O1Ixp25_ASAP7_75t_L g02722(.A1(new_n2609), .A2(new_n2567), .B(new_n2610), .C(new_n2788), .D(new_n2780), .Y(new_n2979));
  NAND3xp33_ASAP7_75t_L     g02723(.A(new_n2979), .B(new_n2978), .C(new_n2975), .Y(new_n2980));
  NOR3xp33_ASAP7_75t_L      g02724(.A(new_n2976), .B(new_n2977), .C(new_n2973), .Y(new_n2981));
  AOI21xp33_ASAP7_75t_L     g02725(.A1(new_n2963), .A2(new_n2967), .B(new_n2974), .Y(new_n2982));
  OAI21xp33_ASAP7_75t_L     g02726(.A1(new_n2785), .A2(new_n2734), .B(new_n2787), .Y(new_n2983));
  OAI21xp33_ASAP7_75t_L     g02727(.A1(new_n2981), .A2(new_n2982), .B(new_n2983), .Y(new_n2984));
  NOR2xp33_ASAP7_75t_L      g02728(.A(new_n833), .B(new_n2118), .Y(new_n2985));
  AOI221xp5_ASAP7_75t_L     g02729(.A1(\b[11] ), .A2(new_n1290), .B1(\b[13] ), .B2(new_n1209), .C(new_n2985), .Y(new_n2986));
  INVx1_ASAP7_75t_L         g02730(.A(new_n2986), .Y(new_n2987));
  A2O1A1Ixp33_ASAP7_75t_L   g02731(.A1(new_n1166), .A2(new_n1216), .B(new_n2987), .C(\a[17] ), .Y(new_n2988));
  O2A1O1Ixp33_ASAP7_75t_L   g02732(.A1(new_n1210), .A2(new_n942), .B(new_n2986), .C(\a[17] ), .Y(new_n2989));
  AOI21xp33_ASAP7_75t_L     g02733(.A1(new_n2988), .A2(\a[17] ), .B(new_n2989), .Y(new_n2990));
  NAND3xp33_ASAP7_75t_L     g02734(.A(new_n2980), .B(new_n2984), .C(new_n2990), .Y(new_n2991));
  NOR3xp33_ASAP7_75t_L      g02735(.A(new_n2983), .B(new_n2982), .C(new_n2981), .Y(new_n2992));
  AOI21xp33_ASAP7_75t_L     g02736(.A1(new_n2978), .A2(new_n2975), .B(new_n2979), .Y(new_n2993));
  AO21x2_ASAP7_75t_L        g02737(.A1(\a[17] ), .A2(new_n2988), .B(new_n2989), .Y(new_n2994));
  OAI21xp33_ASAP7_75t_L     g02738(.A1(new_n2993), .A2(new_n2992), .B(new_n2994), .Y(new_n2995));
  AOI221xp5_ASAP7_75t_L     g02739(.A1(new_n2995), .A2(new_n2991), .B1(new_n2727), .B2(new_n2790), .C(new_n2791), .Y(new_n2996));
  NOR3xp33_ASAP7_75t_L      g02740(.A(new_n2992), .B(new_n2993), .C(new_n2994), .Y(new_n2997));
  AOI21xp33_ASAP7_75t_L     g02741(.A1(new_n2980), .A2(new_n2984), .B(new_n2990), .Y(new_n2998));
  A2O1A1O1Ixp25_ASAP7_75t_L g02742(.A1(new_n2619), .A2(new_n2618), .B(new_n2615), .C(new_n2790), .D(new_n2791), .Y(new_n2999));
  NOR3xp33_ASAP7_75t_L      g02743(.A(new_n2999), .B(new_n2998), .C(new_n2997), .Y(new_n3000));
  NOR2xp33_ASAP7_75t_L      g02744(.A(new_n1043), .B(new_n864), .Y(new_n3001));
  AOI221xp5_ASAP7_75t_L     g02745(.A1(\b[14] ), .A2(new_n985), .B1(\b[16] ), .B2(new_n886), .C(new_n3001), .Y(new_n3002));
  OAI311xp33_ASAP7_75t_L    g02746(.A1(new_n1155), .A2(new_n872), .A3(new_n1154), .B1(\a[14] ), .C1(new_n3002), .Y(new_n3003));
  INVx1_ASAP7_75t_L         g02747(.A(new_n3002), .Y(new_n3004));
  A2O1A1Ixp33_ASAP7_75t_L   g02748(.A1(new_n1156), .A2(new_n873), .B(new_n3004), .C(new_n867), .Y(new_n3005));
  AND2x2_ASAP7_75t_L        g02749(.A(new_n3003), .B(new_n3005), .Y(new_n3006));
  OAI21xp33_ASAP7_75t_L     g02750(.A1(new_n2996), .A2(new_n3000), .B(new_n3006), .Y(new_n3007));
  AOI21xp33_ASAP7_75t_L     g02751(.A1(new_n2995), .A2(new_n2991), .B(new_n2999), .Y(new_n3008));
  OAI21xp33_ASAP7_75t_L     g02752(.A1(new_n2997), .A2(new_n2998), .B(new_n2999), .Y(new_n3009));
  NAND2xp33_ASAP7_75t_L     g02753(.A(new_n3003), .B(new_n3005), .Y(new_n3010));
  OAI211xp5_ASAP7_75t_L     g02754(.A1(new_n2999), .A2(new_n3008), .B(new_n3009), .C(new_n3010), .Y(new_n3011));
  NAND2xp33_ASAP7_75t_L     g02755(.A(new_n3007), .B(new_n3011), .Y(new_n3012));
  NAND2xp33_ASAP7_75t_L     g02756(.A(new_n2796), .B(new_n2793), .Y(new_n3013));
  MAJIxp5_ASAP7_75t_L       g02757(.A(new_n2811), .B(new_n3013), .C(new_n2802), .Y(new_n3014));
  NOR2xp33_ASAP7_75t_L      g02758(.A(new_n3012), .B(new_n3014), .Y(new_n3015));
  NOR2xp33_ASAP7_75t_L      g02759(.A(new_n2805), .B(new_n2804), .Y(new_n3016));
  MAJIxp5_ASAP7_75t_L       g02760(.A(new_n2816), .B(new_n2808), .C(new_n3016), .Y(new_n3017));
  AOI21xp33_ASAP7_75t_L     g02761(.A1(new_n3011), .A2(new_n3007), .B(new_n3017), .Y(new_n3018));
  NOR2xp33_ASAP7_75t_L      g02762(.A(new_n1458), .B(new_n1550), .Y(new_n3019));
  AOI221xp5_ASAP7_75t_L     g02763(.A1(\b[17] ), .A2(new_n713), .B1(\b[19] ), .B2(new_n640), .C(new_n3019), .Y(new_n3020));
  O2A1O1Ixp33_ASAP7_75t_L   g02764(.A1(new_n641), .A2(new_n1628), .B(new_n3020), .C(new_n637), .Y(new_n3021));
  INVx1_ASAP7_75t_L         g02765(.A(new_n3020), .Y(new_n3022));
  A2O1A1Ixp33_ASAP7_75t_L   g02766(.A1(new_n1607), .A2(new_n718), .B(new_n3022), .C(new_n637), .Y(new_n3023));
  OAI21xp33_ASAP7_75t_L     g02767(.A1(new_n637), .A2(new_n3021), .B(new_n3023), .Y(new_n3024));
  NOR3xp33_ASAP7_75t_L      g02768(.A(new_n3015), .B(new_n3018), .C(new_n3024), .Y(new_n3025));
  NAND3xp33_ASAP7_75t_L     g02769(.A(new_n3017), .B(new_n3011), .C(new_n3007), .Y(new_n3026));
  NAND2xp33_ASAP7_75t_L     g02770(.A(new_n3012), .B(new_n3014), .Y(new_n3027));
  A2O1A1Ixp33_ASAP7_75t_L   g02771(.A1(new_n1607), .A2(new_n718), .B(new_n3022), .C(\a[11] ), .Y(new_n3028));
  O2A1O1Ixp33_ASAP7_75t_L   g02772(.A1(new_n641), .A2(new_n1628), .B(new_n3020), .C(\a[11] ), .Y(new_n3029));
  AOI21xp33_ASAP7_75t_L     g02773(.A1(new_n3028), .A2(\a[11] ), .B(new_n3029), .Y(new_n3030));
  AOI21xp33_ASAP7_75t_L     g02774(.A1(new_n3026), .A2(new_n3027), .B(new_n3030), .Y(new_n3031));
  NOR2xp33_ASAP7_75t_L      g02775(.A(new_n3031), .B(new_n3025), .Y(new_n3032));
  NAND2xp33_ASAP7_75t_L     g02776(.A(new_n2817), .B(new_n2812), .Y(new_n3033));
  O2A1O1Ixp33_ASAP7_75t_L   g02777(.A1(new_n2827), .A2(new_n637), .B(new_n2828), .C(new_n3033), .Y(new_n3034));
  A2O1A1O1Ixp25_ASAP7_75t_L g02778(.A1(new_n2833), .A2(new_n2667), .B(new_n2665), .C(new_n2834), .D(new_n3034), .Y(new_n3035));
  NAND2xp33_ASAP7_75t_L     g02779(.A(new_n3032), .B(new_n3035), .Y(new_n3036));
  NAND3xp33_ASAP7_75t_L     g02780(.A(new_n3026), .B(new_n3027), .C(new_n3030), .Y(new_n3037));
  OAI21xp33_ASAP7_75t_L     g02781(.A1(new_n3018), .A2(new_n3015), .B(new_n3024), .Y(new_n3038));
  NAND2xp33_ASAP7_75t_L     g02782(.A(new_n3037), .B(new_n3038), .Y(new_n3039));
  MAJIxp5_ASAP7_75t_L       g02783(.A(new_n2831), .B(new_n3033), .C(new_n2823), .Y(new_n3040));
  NAND2xp33_ASAP7_75t_L     g02784(.A(new_n3040), .B(new_n3039), .Y(new_n3041));
  NOR2xp33_ASAP7_75t_L      g02785(.A(new_n1895), .B(new_n513), .Y(new_n3042));
  AOI221xp5_ASAP7_75t_L     g02786(.A1(\b[20] ), .A2(new_n560), .B1(\b[22] ), .B2(new_n475), .C(new_n3042), .Y(new_n3043));
  O2A1O1Ixp33_ASAP7_75t_L   g02787(.A1(new_n477), .A2(new_n2522), .B(new_n3043), .C(new_n466), .Y(new_n3044));
  O2A1O1Ixp33_ASAP7_75t_L   g02788(.A1(new_n477), .A2(new_n2522), .B(new_n3043), .C(\a[8] ), .Y(new_n3045));
  INVx1_ASAP7_75t_L         g02789(.A(new_n3045), .Y(new_n3046));
  OAI21xp33_ASAP7_75t_L     g02790(.A1(new_n466), .A2(new_n3044), .B(new_n3046), .Y(new_n3047));
  AOI21xp33_ASAP7_75t_L     g02791(.A1(new_n3036), .A2(new_n3041), .B(new_n3047), .Y(new_n3048));
  NOR2xp33_ASAP7_75t_L      g02792(.A(new_n3040), .B(new_n3039), .Y(new_n3049));
  O2A1O1Ixp33_ASAP7_75t_L   g02793(.A1(new_n3033), .A2(new_n2823), .B(new_n2835), .C(new_n3032), .Y(new_n3050));
  INVx1_ASAP7_75t_L         g02794(.A(new_n3044), .Y(new_n3051));
  AOI21xp33_ASAP7_75t_L     g02795(.A1(new_n3051), .A2(\a[8] ), .B(new_n3045), .Y(new_n3052));
  NOR3xp33_ASAP7_75t_L      g02796(.A(new_n3050), .B(new_n3052), .C(new_n3049), .Y(new_n3053));
  A2O1A1O1Ixp25_ASAP7_75t_L g02797(.A1(new_n2688), .A2(new_n2677), .B(new_n2725), .C(new_n2862), .D(new_n2847), .Y(new_n3054));
  NOR3xp33_ASAP7_75t_L      g02798(.A(new_n3054), .B(new_n3053), .C(new_n3048), .Y(new_n3055));
  OAI21xp33_ASAP7_75t_L     g02799(.A1(new_n3049), .A2(new_n3050), .B(new_n3052), .Y(new_n3056));
  NAND3xp33_ASAP7_75t_L     g02800(.A(new_n3036), .B(new_n3047), .C(new_n3041), .Y(new_n3057));
  OAI21xp33_ASAP7_75t_L     g02801(.A1(new_n2843), .A2(new_n2851), .B(new_n2863), .Y(new_n3058));
  AOI21xp33_ASAP7_75t_L     g02802(.A1(new_n3057), .A2(new_n3056), .B(new_n3058), .Y(new_n3059));
  NOR3xp33_ASAP7_75t_L      g02803(.A(new_n3059), .B(new_n2907), .C(new_n3055), .Y(new_n3060));
  NAND3xp33_ASAP7_75t_L     g02804(.A(new_n3058), .B(new_n3057), .C(new_n3056), .Y(new_n3061));
  OAI21xp33_ASAP7_75t_L     g02805(.A1(new_n3048), .A2(new_n3053), .B(new_n3054), .Y(new_n3062));
  NAND3xp33_ASAP7_75t_L     g02806(.A(new_n3061), .B(new_n2907), .C(new_n3062), .Y(new_n3063));
  OAI21xp33_ASAP7_75t_L     g02807(.A1(new_n2907), .A2(new_n3060), .B(new_n3063), .Y(new_n3064));
  NOR3xp33_ASAP7_75t_L      g02808(.A(new_n2861), .B(new_n2859), .C(new_n2864), .Y(new_n3065));
  INVx1_ASAP7_75t_L         g02809(.A(new_n3065), .Y(new_n3066));
  A2O1A1O1Ixp25_ASAP7_75t_L g02810(.A1(new_n2544), .A2(new_n2540), .B(new_n2552), .C(new_n2694), .D(new_n2698), .Y(new_n3067));
  A2O1A1Ixp33_ASAP7_75t_L   g02811(.A1(new_n2860), .A2(new_n2867), .B(new_n3067), .C(new_n3066), .Y(new_n3068));
  NOR2xp33_ASAP7_75t_L      g02812(.A(new_n3064), .B(new_n3068), .Y(new_n3069));
  NOR4xp25_ASAP7_75t_L      g02813(.A(new_n3059), .B(new_n2906), .C(new_n3055), .D(new_n2905), .Y(new_n3070));
  AOI21xp33_ASAP7_75t_L     g02814(.A1(new_n3061), .A2(new_n3062), .B(new_n2907), .Y(new_n3071));
  NOR2xp33_ASAP7_75t_L      g02815(.A(new_n3071), .B(new_n3070), .Y(new_n3072));
  A2O1A1O1Ixp25_ASAP7_75t_L g02816(.A1(new_n2867), .A2(new_n2860), .B(new_n3067), .C(new_n3066), .D(new_n3072), .Y(new_n3073));
  NOR2xp33_ASAP7_75t_L      g02817(.A(new_n2703), .B(new_n287), .Y(new_n3074));
  AOI221xp5_ASAP7_75t_L     g02818(.A1(\b[27] ), .A2(new_n264), .B1(\b[28] ), .B2(new_n283), .C(new_n3074), .Y(new_n3075));
  INVx1_ASAP7_75t_L         g02819(.A(new_n3075), .Y(new_n3076));
  INVx1_ASAP7_75t_L         g02820(.A(new_n2880), .Y(new_n3077));
  NOR2xp33_ASAP7_75t_L      g02821(.A(\b[27] ), .B(\b[28] ), .Y(new_n3078));
  INVx1_ASAP7_75t_L         g02822(.A(\b[28] ), .Y(new_n3079));
  NOR2xp33_ASAP7_75t_L      g02823(.A(new_n2879), .B(new_n3079), .Y(new_n3080));
  NOR2xp33_ASAP7_75t_L      g02824(.A(new_n3078), .B(new_n3080), .Y(new_n3081));
  INVx1_ASAP7_75t_L         g02825(.A(new_n3081), .Y(new_n3082));
  O2A1O1Ixp33_ASAP7_75t_L   g02826(.A1(new_n2882), .A2(new_n2885), .B(new_n3077), .C(new_n3082), .Y(new_n3083));
  NOR3xp33_ASAP7_75t_L      g02827(.A(new_n2883), .B(new_n3081), .C(new_n2880), .Y(new_n3084));
  NOR2xp33_ASAP7_75t_L      g02828(.A(new_n3083), .B(new_n3084), .Y(new_n3085));
  A2O1A1Ixp33_ASAP7_75t_L   g02829(.A1(new_n3085), .A2(new_n273), .B(new_n3076), .C(\a[2] ), .Y(new_n3086));
  INVx1_ASAP7_75t_L         g02830(.A(new_n3085), .Y(new_n3087));
  O2A1O1Ixp33_ASAP7_75t_L   g02831(.A1(new_n279), .A2(new_n3087), .B(new_n3075), .C(\a[2] ), .Y(new_n3088));
  AOI21xp33_ASAP7_75t_L     g02832(.A1(new_n3086), .A2(\a[2] ), .B(new_n3088), .Y(new_n3089));
  OAI21xp33_ASAP7_75t_L     g02833(.A1(new_n3073), .A2(new_n3069), .B(new_n3089), .Y(new_n3090));
  NOR3xp33_ASAP7_75t_L      g02834(.A(new_n3069), .B(new_n3073), .C(new_n3089), .Y(new_n3091));
  INVx1_ASAP7_75t_L         g02835(.A(new_n3091), .Y(new_n3092));
  NAND2xp33_ASAP7_75t_L     g02836(.A(new_n3090), .B(new_n3092), .Y(new_n3093));
  XOR2x2_ASAP7_75t_L        g02837(.A(new_n2901), .B(new_n3093), .Y(\f[28] ));
  NOR2xp33_ASAP7_75t_L      g02838(.A(new_n2879), .B(new_n287), .Y(new_n3095));
  AOI221xp5_ASAP7_75t_L     g02839(.A1(\b[28] ), .A2(new_n264), .B1(\b[29] ), .B2(new_n283), .C(new_n3095), .Y(new_n3096));
  NOR2xp33_ASAP7_75t_L      g02840(.A(\b[28] ), .B(\b[29] ), .Y(new_n3097));
  INVx1_ASAP7_75t_L         g02841(.A(\b[29] ), .Y(new_n3098));
  NOR2xp33_ASAP7_75t_L      g02842(.A(new_n3079), .B(new_n3098), .Y(new_n3099));
  NOR2xp33_ASAP7_75t_L      g02843(.A(new_n3097), .B(new_n3099), .Y(new_n3100));
  A2O1A1Ixp33_ASAP7_75t_L   g02844(.A1(\b[28] ), .A2(\b[27] ), .B(new_n3083), .C(new_n3100), .Y(new_n3101));
  O2A1O1Ixp33_ASAP7_75t_L   g02845(.A1(new_n2880), .A2(new_n2883), .B(new_n3081), .C(new_n3080), .Y(new_n3102));
  OAI21xp33_ASAP7_75t_L     g02846(.A1(new_n3097), .A2(new_n3099), .B(new_n3102), .Y(new_n3103));
  NAND2xp33_ASAP7_75t_L     g02847(.A(new_n3101), .B(new_n3103), .Y(new_n3104));
  O2A1O1Ixp33_ASAP7_75t_L   g02848(.A1(new_n279), .A2(new_n3104), .B(new_n3096), .C(new_n257), .Y(new_n3105));
  OAI21xp33_ASAP7_75t_L     g02849(.A1(new_n279), .A2(new_n3104), .B(new_n3096), .Y(new_n3106));
  NAND2xp33_ASAP7_75t_L     g02850(.A(new_n257), .B(new_n3106), .Y(new_n3107));
  OA21x2_ASAP7_75t_L        g02851(.A1(new_n257), .A2(new_n3105), .B(new_n3107), .Y(new_n3108));
  NOR2xp33_ASAP7_75t_L      g02852(.A(new_n2205), .B(new_n375), .Y(new_n3109));
  AOI221xp5_ASAP7_75t_L     g02853(.A1(\b[26] ), .A2(new_n361), .B1(new_n349), .B2(\b[25] ), .C(new_n3109), .Y(new_n3110));
  O2A1O1Ixp33_ASAP7_75t_L   g02854(.A1(new_n356), .A2(new_n2708), .B(new_n3110), .C(new_n346), .Y(new_n3111));
  INVx1_ASAP7_75t_L         g02855(.A(new_n3111), .Y(new_n3112));
  O2A1O1Ixp33_ASAP7_75t_L   g02856(.A1(new_n356), .A2(new_n2708), .B(new_n3110), .C(\a[5] ), .Y(new_n3113));
  INVx1_ASAP7_75t_L         g02857(.A(new_n3113), .Y(new_n3114));
  NAND2xp33_ASAP7_75t_L     g02858(.A(new_n3027), .B(new_n3026), .Y(new_n3115));
  O2A1O1Ixp33_ASAP7_75t_L   g02859(.A1(new_n3021), .A2(new_n637), .B(new_n3023), .C(new_n3115), .Y(new_n3116));
  O2A1O1Ixp33_ASAP7_75t_L   g02860(.A1(new_n3025), .A2(new_n3024), .B(new_n3040), .C(new_n3116), .Y(new_n3117));
  NAND3xp33_ASAP7_75t_L     g02861(.A(new_n2963), .B(new_n2967), .C(new_n2973), .Y(new_n3118));
  NOR2xp33_ASAP7_75t_L      g02862(.A(new_n680), .B(new_n1517), .Y(new_n3119));
  AOI221xp5_ASAP7_75t_L     g02863(.A1(\b[9] ), .A2(new_n1659), .B1(\b[11] ), .B2(new_n1511), .C(new_n3119), .Y(new_n3120));
  O2A1O1Ixp33_ASAP7_75t_L   g02864(.A1(new_n1521), .A2(new_n754), .B(new_n3120), .C(new_n1501), .Y(new_n3121));
  INVx1_ASAP7_75t_L         g02865(.A(new_n3120), .Y(new_n3122));
  A2O1A1Ixp33_ASAP7_75t_L   g02866(.A1(new_n976), .A2(new_n1513), .B(new_n3122), .C(new_n1501), .Y(new_n3123));
  OAI21xp33_ASAP7_75t_L     g02867(.A1(new_n1501), .A2(new_n3121), .B(new_n3123), .Y(new_n3124));
  A2O1A1Ixp33_ASAP7_75t_L   g02868(.A1(new_n2964), .A2(new_n2769), .B(new_n2966), .C(new_n2958), .Y(new_n3125));
  OAI211xp5_ASAP7_75t_L     g02869(.A1(new_n2945), .A2(new_n2946), .B(new_n2943), .C(new_n2934), .Y(new_n3126));
  A2O1A1Ixp33_ASAP7_75t_L   g02870(.A1(new_n2944), .A2(new_n2953), .B(new_n2956), .C(new_n3126), .Y(new_n3127));
  NOR2xp33_ASAP7_75t_L      g02871(.A(new_n289), .B(new_n2930), .Y(new_n3128));
  AND3x1_ASAP7_75t_L        g02872(.A(new_n2739), .B(new_n2937), .C(new_n2935), .Y(new_n3129));
  AOI221xp5_ASAP7_75t_L     g02873(.A1(new_n2936), .A2(\b[1] ), .B1(new_n3129), .B2(\b[0] ), .C(new_n3128), .Y(new_n3130));
  NAND2xp33_ASAP7_75t_L     g02874(.A(new_n2932), .B(new_n294), .Y(new_n3131));
  NAND3xp33_ASAP7_75t_L     g02875(.A(new_n3130), .B(\a[29] ), .C(new_n3131), .Y(new_n3132));
  NAND3xp33_ASAP7_75t_L     g02876(.A(new_n2739), .B(new_n2935), .C(new_n2937), .Y(new_n3133));
  NAND2xp33_ASAP7_75t_L     g02877(.A(\b[1] ), .B(new_n2936), .Y(new_n3134));
  OAI221xp5_ASAP7_75t_L     g02878(.A1(new_n2930), .A2(new_n289), .B1(new_n284), .B2(new_n3133), .C(new_n3134), .Y(new_n3135));
  A2O1A1Ixp33_ASAP7_75t_L   g02879(.A1(new_n294), .A2(new_n2932), .B(new_n3135), .C(new_n2928), .Y(new_n3136));
  NAND3xp33_ASAP7_75t_L     g02880(.A(new_n2934), .B(new_n3132), .C(new_n3136), .Y(new_n3137));
  INVx1_ASAP7_75t_L         g02881(.A(new_n3137), .Y(new_n3138));
  INVx1_ASAP7_75t_L         g02882(.A(new_n3131), .Y(new_n3139));
  NOR5xp2_ASAP7_75t_L       g02883(.A(new_n2948), .B(new_n3135), .C(new_n3139), .D(new_n2740), .E(new_n2928), .Y(new_n3140));
  NAND2xp33_ASAP7_75t_L     g02884(.A(\b[4] ), .B(new_n2421), .Y(new_n3141));
  OAI221xp5_ASAP7_75t_L     g02885(.A1(new_n2415), .A2(new_n384), .B1(new_n301), .B2(new_n2572), .C(new_n3141), .Y(new_n3142));
  A2O1A1Ixp33_ASAP7_75t_L   g02886(.A1(new_n394), .A2(new_n2417), .B(new_n3142), .C(\a[26] ), .Y(new_n3143));
  INVx1_ASAP7_75t_L         g02887(.A(new_n3142), .Y(new_n3144));
  O2A1O1Ixp33_ASAP7_75t_L   g02888(.A1(new_n2425), .A2(new_n728), .B(new_n3144), .C(\a[26] ), .Y(new_n3145));
  AOI21xp33_ASAP7_75t_L     g02889(.A1(new_n3143), .A2(\a[26] ), .B(new_n3145), .Y(new_n3146));
  NOR3xp33_ASAP7_75t_L      g02890(.A(new_n3138), .B(new_n3140), .C(new_n3146), .Y(new_n3147));
  NAND5xp2_ASAP7_75t_L      g02891(.A(\a[29] ), .B(new_n2933), .C(new_n3131), .D(new_n3130), .E(new_n2741), .Y(new_n3148));
  AOI221xp5_ASAP7_75t_L     g02892(.A1(new_n3143), .A2(\a[26] ), .B1(new_n3148), .B2(new_n3137), .C(new_n3145), .Y(new_n3149));
  OAI21xp33_ASAP7_75t_L     g02893(.A1(new_n3147), .A2(new_n3149), .B(new_n3127), .Y(new_n3150));
  OR3x1_ASAP7_75t_L         g02894(.A(new_n3138), .B(new_n3140), .C(new_n3146), .Y(new_n3151));
  OAI21xp33_ASAP7_75t_L     g02895(.A1(new_n3140), .A2(new_n3138), .B(new_n3146), .Y(new_n3152));
  NAND4xp25_ASAP7_75t_L     g02896(.A(new_n2955), .B(new_n3152), .C(new_n3151), .D(new_n3126), .Y(new_n3153));
  NOR2xp33_ASAP7_75t_L      g02897(.A(new_n448), .B(new_n1962), .Y(new_n3154));
  AOI221xp5_ASAP7_75t_L     g02898(.A1(new_n1955), .A2(\b[8] ), .B1(new_n2093), .B2(\b[6] ), .C(new_n3154), .Y(new_n3155));
  O2A1O1Ixp33_ASAP7_75t_L   g02899(.A1(new_n1956), .A2(new_n540), .B(new_n3155), .C(new_n1952), .Y(new_n3156));
  NOR2xp33_ASAP7_75t_L      g02900(.A(new_n1952), .B(new_n3156), .Y(new_n3157));
  O2A1O1Ixp33_ASAP7_75t_L   g02901(.A1(new_n1956), .A2(new_n540), .B(new_n3155), .C(\a[23] ), .Y(new_n3158));
  NOR2xp33_ASAP7_75t_L      g02902(.A(new_n3158), .B(new_n3157), .Y(new_n3159));
  NAND3xp33_ASAP7_75t_L     g02903(.A(new_n3153), .B(new_n3150), .C(new_n3159), .Y(new_n3160));
  AO21x2_ASAP7_75t_L        g02904(.A1(new_n3150), .A2(new_n3153), .B(new_n3159), .Y(new_n3161));
  NAND3xp33_ASAP7_75t_L     g02905(.A(new_n3125), .B(new_n3160), .C(new_n3161), .Y(new_n3162));
  A2O1A1Ixp33_ASAP7_75t_L   g02906(.A1(new_n2432), .A2(new_n2599), .B(new_n2596), .C(new_n2600), .Y(new_n3163));
  INVx1_ASAP7_75t_L         g02907(.A(new_n2769), .Y(new_n3164));
  O2A1O1Ixp33_ASAP7_75t_L   g02908(.A1(new_n2772), .A2(new_n2764), .B(new_n3163), .C(new_n3164), .Y(new_n3165));
  AND3x1_ASAP7_75t_L        g02909(.A(new_n3153), .B(new_n3150), .C(new_n3159), .Y(new_n3166));
  AOI21xp33_ASAP7_75t_L     g02910(.A1(new_n3153), .A2(new_n3150), .B(new_n3159), .Y(new_n3167));
  OAI221xp5_ASAP7_75t_L     g02911(.A1(new_n3165), .A2(new_n2966), .B1(new_n3166), .B2(new_n3167), .C(new_n2958), .Y(new_n3168));
  AOI21xp33_ASAP7_75t_L     g02912(.A1(new_n3168), .A2(new_n3162), .B(new_n3124), .Y(new_n3169));
  AND3x1_ASAP7_75t_L        g02913(.A(new_n3168), .B(new_n3162), .C(new_n3124), .Y(new_n3170));
  AOI211xp5_ASAP7_75t_L     g02914(.A1(new_n2984), .A2(new_n3118), .B(new_n3169), .C(new_n3170), .Y(new_n3171));
  A2O1A1Ixp33_ASAP7_75t_L   g02915(.A1(new_n2974), .A2(new_n2975), .B(new_n2979), .C(new_n3118), .Y(new_n3172));
  AO21x2_ASAP7_75t_L        g02916(.A1(new_n3162), .A2(new_n3168), .B(new_n3124), .Y(new_n3173));
  NAND3xp33_ASAP7_75t_L     g02917(.A(new_n3168), .B(new_n3162), .C(new_n3124), .Y(new_n3174));
  AOI21xp33_ASAP7_75t_L     g02918(.A1(new_n3174), .A2(new_n3173), .B(new_n3172), .Y(new_n3175));
  NOR2xp33_ASAP7_75t_L      g02919(.A(new_n936), .B(new_n2118), .Y(new_n3176));
  AOI221xp5_ASAP7_75t_L     g02920(.A1(\b[12] ), .A2(new_n1290), .B1(\b[14] ), .B2(new_n1209), .C(new_n3176), .Y(new_n3177));
  O2A1O1Ixp33_ASAP7_75t_L   g02921(.A1(new_n1210), .A2(new_n1268), .B(new_n3177), .C(new_n1206), .Y(new_n3178));
  INVx1_ASAP7_75t_L         g02922(.A(new_n3177), .Y(new_n3179));
  A2O1A1Ixp33_ASAP7_75t_L   g02923(.A1(new_n971), .A2(new_n1216), .B(new_n3179), .C(new_n1206), .Y(new_n3180));
  OAI21xp33_ASAP7_75t_L     g02924(.A1(new_n1206), .A2(new_n3178), .B(new_n3180), .Y(new_n3181));
  NOR3xp33_ASAP7_75t_L      g02925(.A(new_n3171), .B(new_n3175), .C(new_n3181), .Y(new_n3182));
  OA21x2_ASAP7_75t_L        g02926(.A1(new_n3175), .A2(new_n3171), .B(new_n3181), .Y(new_n3183));
  NAND2xp33_ASAP7_75t_L     g02927(.A(new_n2984), .B(new_n2980), .Y(new_n3184));
  MAJIxp5_ASAP7_75t_L       g02928(.A(new_n2999), .B(new_n3184), .C(new_n2990), .Y(new_n3185));
  NOR3xp33_ASAP7_75t_L      g02929(.A(new_n3185), .B(new_n3183), .C(new_n3182), .Y(new_n3186));
  OA21x2_ASAP7_75t_L        g02930(.A1(new_n3182), .A2(new_n3183), .B(new_n3185), .Y(new_n3187));
  NOR2xp33_ASAP7_75t_L      g02931(.A(new_n1150), .B(new_n864), .Y(new_n3188));
  AOI221xp5_ASAP7_75t_L     g02932(.A1(\b[15] ), .A2(new_n985), .B1(\b[17] ), .B2(new_n886), .C(new_n3188), .Y(new_n3189));
  O2A1O1Ixp33_ASAP7_75t_L   g02933(.A1(new_n872), .A2(new_n1356), .B(new_n3189), .C(new_n867), .Y(new_n3190));
  INVx1_ASAP7_75t_L         g02934(.A(new_n3189), .Y(new_n3191));
  A2O1A1Ixp33_ASAP7_75t_L   g02935(.A1(new_n1633), .A2(new_n873), .B(new_n3191), .C(new_n867), .Y(new_n3192));
  OAI21xp33_ASAP7_75t_L     g02936(.A1(new_n867), .A2(new_n3190), .B(new_n3192), .Y(new_n3193));
  NOR3xp33_ASAP7_75t_L      g02937(.A(new_n3187), .B(new_n3193), .C(new_n3186), .Y(new_n3194));
  INVx1_ASAP7_75t_L         g02938(.A(new_n3184), .Y(new_n3195));
  A2O1A1Ixp33_ASAP7_75t_L   g02939(.A1(\a[17] ), .A2(new_n2988), .B(new_n2989), .C(new_n3195), .Y(new_n3196));
  AO21x2_ASAP7_75t_L        g02940(.A1(new_n2991), .A2(new_n2995), .B(new_n2999), .Y(new_n3197));
  OR3x1_ASAP7_75t_L         g02941(.A(new_n3171), .B(new_n3175), .C(new_n3181), .Y(new_n3198));
  OAI21xp33_ASAP7_75t_L     g02942(.A1(new_n3175), .A2(new_n3171), .B(new_n3181), .Y(new_n3199));
  NAND4xp25_ASAP7_75t_L     g02943(.A(new_n3197), .B(new_n3198), .C(new_n3199), .D(new_n3196), .Y(new_n3200));
  OAI21xp33_ASAP7_75t_L     g02944(.A1(new_n3182), .A2(new_n3183), .B(new_n3185), .Y(new_n3201));
  A2O1A1Ixp33_ASAP7_75t_L   g02945(.A1(new_n1633), .A2(new_n873), .B(new_n3191), .C(\a[14] ), .Y(new_n3202));
  O2A1O1Ixp33_ASAP7_75t_L   g02946(.A1(new_n872), .A2(new_n1356), .B(new_n3189), .C(\a[14] ), .Y(new_n3203));
  AOI21xp33_ASAP7_75t_L     g02947(.A1(new_n3202), .A2(\a[14] ), .B(new_n3203), .Y(new_n3204));
  AOI21xp33_ASAP7_75t_L     g02948(.A1(new_n3200), .A2(new_n3201), .B(new_n3204), .Y(new_n3205));
  NOR2xp33_ASAP7_75t_L      g02949(.A(new_n3205), .B(new_n3194), .Y(new_n3206));
  O2A1O1Ixp33_ASAP7_75t_L   g02950(.A1(new_n2806), .A2(new_n867), .B(new_n2807), .C(new_n3013), .Y(new_n3207));
  O2A1O1Ixp33_ASAP7_75t_L   g02951(.A1(new_n2999), .A2(new_n3008), .B(new_n3009), .C(new_n3006), .Y(new_n3208));
  O2A1O1Ixp33_ASAP7_75t_L   g02952(.A1(new_n3207), .A2(new_n2826), .B(new_n3012), .C(new_n3208), .Y(new_n3209));
  NAND2xp33_ASAP7_75t_L     g02953(.A(new_n3206), .B(new_n3209), .Y(new_n3210));
  A2O1A1Ixp33_ASAP7_75t_L   g02954(.A1(new_n2793), .A2(new_n2792), .B(new_n3008), .C(new_n3009), .Y(new_n3211));
  NAND3xp33_ASAP7_75t_L     g02955(.A(new_n3200), .B(new_n3201), .C(new_n3204), .Y(new_n3212));
  OAI21xp33_ASAP7_75t_L     g02956(.A1(new_n3186), .A2(new_n3187), .B(new_n3193), .Y(new_n3213));
  NAND2xp33_ASAP7_75t_L     g02957(.A(new_n3212), .B(new_n3213), .Y(new_n3214));
  A2O1A1Ixp33_ASAP7_75t_L   g02958(.A1(new_n3010), .A2(new_n3211), .B(new_n3018), .C(new_n3214), .Y(new_n3215));
  NOR2xp33_ASAP7_75t_L      g02959(.A(new_n1599), .B(new_n1550), .Y(new_n3216));
  AOI221xp5_ASAP7_75t_L     g02960(.A1(\b[18] ), .A2(new_n713), .B1(\b[20] ), .B2(new_n640), .C(new_n3216), .Y(new_n3217));
  INVx1_ASAP7_75t_L         g02961(.A(new_n3217), .Y(new_n3218));
  A2O1A1Ixp33_ASAP7_75t_L   g02962(.A1(new_n1752), .A2(new_n718), .B(new_n3218), .C(\a[11] ), .Y(new_n3219));
  O2A1O1Ixp33_ASAP7_75t_L   g02963(.A1(new_n641), .A2(new_n1754), .B(new_n3217), .C(\a[11] ), .Y(new_n3220));
  AOI21xp33_ASAP7_75t_L     g02964(.A1(new_n3219), .A2(\a[11] ), .B(new_n3220), .Y(new_n3221));
  INVx1_ASAP7_75t_L         g02965(.A(new_n3221), .Y(new_n3222));
  NAND3xp33_ASAP7_75t_L     g02966(.A(new_n3222), .B(new_n3215), .C(new_n3210), .Y(new_n3223));
  NOR2xp33_ASAP7_75t_L      g02967(.A(new_n3018), .B(new_n3015), .Y(new_n3224));
  A2O1A1Ixp33_ASAP7_75t_L   g02968(.A1(\a[11] ), .A2(new_n3028), .B(new_n3029), .C(new_n3224), .Y(new_n3225));
  AOI21xp33_ASAP7_75t_L     g02969(.A1(new_n3215), .A2(new_n3210), .B(new_n3222), .Y(new_n3226));
  O2A1O1Ixp33_ASAP7_75t_L   g02970(.A1(new_n3032), .A2(new_n3035), .B(new_n3225), .C(new_n3226), .Y(new_n3227));
  INVx1_ASAP7_75t_L         g02971(.A(new_n3208), .Y(new_n3228));
  A2O1A1Ixp33_ASAP7_75t_L   g02972(.A1(new_n3006), .A2(new_n3007), .B(new_n3017), .C(new_n3228), .Y(new_n3229));
  NOR2xp33_ASAP7_75t_L      g02973(.A(new_n3214), .B(new_n3229), .Y(new_n3230));
  NOR2xp33_ASAP7_75t_L      g02974(.A(new_n3206), .B(new_n3209), .Y(new_n3231));
  OAI21xp33_ASAP7_75t_L     g02975(.A1(new_n3230), .A2(new_n3231), .B(new_n3221), .Y(new_n3232));
  NAND4xp25_ASAP7_75t_L     g02976(.A(new_n3041), .B(new_n3223), .C(new_n3232), .D(new_n3225), .Y(new_n3233));
  A2O1A1Ixp33_ASAP7_75t_L   g02977(.A1(new_n3223), .A2(new_n3227), .B(new_n3117), .C(new_n3233), .Y(new_n3234));
  AOI21xp33_ASAP7_75t_L     g02978(.A1(new_n3232), .A2(new_n3223), .B(new_n3117), .Y(new_n3235));
  NOR3xp33_ASAP7_75t_L      g02979(.A(new_n3231), .B(new_n3230), .C(new_n3221), .Y(new_n3236));
  A2O1A1O1Ixp25_ASAP7_75t_L g02980(.A1(new_n3040), .A2(new_n3039), .B(new_n3116), .C(new_n3232), .D(new_n3236), .Y(new_n3237));
  NOR2xp33_ASAP7_75t_L      g02981(.A(new_n2045), .B(new_n513), .Y(new_n3238));
  AOI221xp5_ASAP7_75t_L     g02982(.A1(\b[21] ), .A2(new_n560), .B1(\b[23] ), .B2(new_n475), .C(new_n3238), .Y(new_n3239));
  O2A1O1Ixp33_ASAP7_75t_L   g02983(.A1(new_n477), .A2(new_n2194), .B(new_n3239), .C(new_n466), .Y(new_n3240));
  INVx1_ASAP7_75t_L         g02984(.A(new_n3239), .Y(new_n3241));
  A2O1A1Ixp33_ASAP7_75t_L   g02985(.A1(new_n2679), .A2(new_n483), .B(new_n3241), .C(new_n466), .Y(new_n3242));
  OAI21xp33_ASAP7_75t_L     g02986(.A1(new_n466), .A2(new_n3240), .B(new_n3242), .Y(new_n3243));
  A2O1A1Ixp33_ASAP7_75t_L   g02987(.A1(new_n3237), .A2(new_n3232), .B(new_n3235), .C(new_n3243), .Y(new_n3244));
  A2O1A1Ixp33_ASAP7_75t_L   g02988(.A1(new_n2679), .A2(new_n483), .B(new_n3241), .C(\a[8] ), .Y(new_n3245));
  O2A1O1Ixp33_ASAP7_75t_L   g02989(.A1(new_n477), .A2(new_n2194), .B(new_n3239), .C(\a[8] ), .Y(new_n3246));
  AOI21xp33_ASAP7_75t_L     g02990(.A1(new_n3245), .A2(\a[8] ), .B(new_n3246), .Y(new_n3247));
  AOI211xp5_ASAP7_75t_L     g02991(.A1(new_n3237), .A2(new_n3232), .B(new_n3247), .C(new_n3235), .Y(new_n3248));
  OAI21xp33_ASAP7_75t_L     g02992(.A1(new_n3048), .A2(new_n3054), .B(new_n3057), .Y(new_n3249));
  A2O1A1Ixp33_ASAP7_75t_L   g02993(.A1(new_n3244), .A2(new_n3234), .B(new_n3248), .C(new_n3249), .Y(new_n3250));
  A2O1A1Ixp33_ASAP7_75t_L   g02994(.A1(new_n3237), .A2(new_n3232), .B(new_n3235), .C(new_n3247), .Y(new_n3251));
  A2O1A1Ixp33_ASAP7_75t_L   g02995(.A1(new_n3030), .A2(new_n3037), .B(new_n3035), .C(new_n3225), .Y(new_n3252));
  OAI21xp33_ASAP7_75t_L     g02996(.A1(new_n3236), .A2(new_n3226), .B(new_n3252), .Y(new_n3253));
  NAND3xp33_ASAP7_75t_L     g02997(.A(new_n3253), .B(new_n3233), .C(new_n3243), .Y(new_n3254));
  A2O1A1Ixp33_ASAP7_75t_L   g02998(.A1(\a[8] ), .A2(new_n2659), .B(new_n2669), .C(new_n2850), .Y(new_n3255));
  OAI21xp33_ASAP7_75t_L     g02999(.A1(new_n2672), .A2(new_n2673), .B(new_n3255), .Y(new_n3256));
  A2O1A1O1Ixp25_ASAP7_75t_L g03000(.A1(new_n2848), .A2(new_n3256), .B(new_n2847), .C(new_n3056), .D(new_n3053), .Y(new_n3257));
  NAND3xp33_ASAP7_75t_L     g03001(.A(new_n3257), .B(new_n3254), .C(new_n3251), .Y(new_n3258));
  NAND2xp33_ASAP7_75t_L     g03002(.A(new_n3250), .B(new_n3258), .Y(new_n3259));
  O2A1O1Ixp33_ASAP7_75t_L   g03003(.A1(new_n346), .A2(new_n3111), .B(new_n3114), .C(new_n3259), .Y(new_n3260));
  INVx1_ASAP7_75t_L         g03004(.A(new_n3260), .Y(new_n3261));
  AO21x2_ASAP7_75t_L        g03005(.A1(\a[5] ), .A2(new_n3112), .B(new_n3113), .Y(new_n3262));
  NOR2xp33_ASAP7_75t_L      g03006(.A(new_n3262), .B(new_n3259), .Y(new_n3263));
  A2O1A1O1Ixp25_ASAP7_75t_L g03007(.A1(new_n3112), .A2(\a[5] ), .B(new_n3113), .C(new_n3261), .D(new_n3263), .Y(new_n3264));
  A2O1A1O1Ixp25_ASAP7_75t_L g03008(.A1(new_n2868), .A2(new_n2871), .B(new_n3065), .C(new_n3064), .D(new_n3060), .Y(new_n3265));
  AOI21xp33_ASAP7_75t_L     g03009(.A1(new_n3254), .A2(new_n3251), .B(new_n3257), .Y(new_n3266));
  A2O1A1O1Ixp25_ASAP7_75t_L g03010(.A1(new_n3223), .A2(new_n3227), .B(new_n3117), .C(new_n3233), .D(new_n3243), .Y(new_n3267));
  NOR3xp33_ASAP7_75t_L      g03011(.A(new_n3249), .B(new_n3248), .C(new_n3267), .Y(new_n3268));
  OAI21xp33_ASAP7_75t_L     g03012(.A1(new_n3268), .A2(new_n3266), .B(new_n3262), .Y(new_n3269));
  O2A1O1Ixp33_ASAP7_75t_L   g03013(.A1(new_n3259), .A2(new_n3260), .B(new_n3269), .C(new_n3265), .Y(new_n3270));
  AOI21xp33_ASAP7_75t_L     g03014(.A1(new_n3112), .A2(\a[5] ), .B(new_n3113), .Y(new_n3271));
  NAND3xp33_ASAP7_75t_L     g03015(.A(new_n3258), .B(new_n3250), .C(new_n3271), .Y(new_n3272));
  NAND2xp33_ASAP7_75t_L     g03016(.A(new_n3272), .B(new_n3269), .Y(new_n3273));
  A2O1A1Ixp33_ASAP7_75t_L   g03017(.A1(new_n3064), .A2(new_n3068), .B(new_n3060), .C(new_n3273), .Y(new_n3274));
  A2O1A1Ixp33_ASAP7_75t_L   g03018(.A1(new_n3064), .A2(new_n3068), .B(new_n3060), .C(new_n3274), .Y(new_n3275));
  O2A1O1Ixp33_ASAP7_75t_L   g03019(.A1(new_n3270), .A2(new_n3264), .B(new_n3275), .C(new_n3108), .Y(new_n3276));
  INVx1_ASAP7_75t_L         g03020(.A(new_n3060), .Y(new_n3277));
  A2O1A1O1Ixp25_ASAP7_75t_L g03021(.A1(new_n2696), .A2(new_n2694), .B(new_n2698), .C(new_n2868), .D(new_n3065), .Y(new_n3278));
  O2A1O1Ixp33_ASAP7_75t_L   g03022(.A1(new_n3072), .A2(new_n3278), .B(new_n3277), .C(new_n3273), .Y(new_n3279));
  A2O1A1Ixp33_ASAP7_75t_L   g03023(.A1(new_n3274), .A2(new_n3273), .B(new_n3279), .C(new_n3108), .Y(new_n3280));
  A2O1A1O1Ixp25_ASAP7_75t_L g03024(.A1(new_n2893), .A2(new_n2898), .B(new_n2894), .C(new_n3090), .D(new_n3091), .Y(new_n3281));
  O2A1O1Ixp33_ASAP7_75t_L   g03025(.A1(new_n3108), .A2(new_n3276), .B(new_n3280), .C(new_n3281), .Y(new_n3282));
  OA211x2_ASAP7_75t_L       g03026(.A1(new_n3108), .A2(new_n3276), .B(new_n3280), .C(new_n3281), .Y(new_n3283));
  NOR2xp33_ASAP7_75t_L      g03027(.A(new_n3282), .B(new_n3283), .Y(\f[29] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03028(.A1(new_n3223), .A2(new_n3227), .B(new_n3117), .C(new_n3233), .D(new_n3247), .Y(new_n3285));
  O2A1O1Ixp33_ASAP7_75t_L   g03029(.A1(new_n3267), .A2(new_n3243), .B(new_n3249), .C(new_n3285), .Y(new_n3286));
  A2O1A1Ixp33_ASAP7_75t_L   g03030(.A1(new_n2984), .A2(new_n3118), .B(new_n3169), .C(new_n3174), .Y(new_n3287));
  NOR2xp33_ASAP7_75t_L      g03031(.A(new_n748), .B(new_n1517), .Y(new_n3288));
  AOI221xp5_ASAP7_75t_L     g03032(.A1(\b[10] ), .A2(new_n1659), .B1(\b[12] ), .B2(new_n1511), .C(new_n3288), .Y(new_n3289));
  INVx1_ASAP7_75t_L         g03033(.A(new_n3289), .Y(new_n3290));
  A2O1A1Ixp33_ASAP7_75t_L   g03034(.A1(new_n1057), .A2(new_n1513), .B(new_n3290), .C(\a[20] ), .Y(new_n3291));
  O2A1O1Ixp33_ASAP7_75t_L   g03035(.A1(new_n1521), .A2(new_n841), .B(new_n3289), .C(\a[20] ), .Y(new_n3292));
  AOI21xp33_ASAP7_75t_L     g03036(.A1(new_n3291), .A2(\a[20] ), .B(new_n3292), .Y(new_n3293));
  A2O1A1O1Ixp25_ASAP7_75t_L g03037(.A1(new_n2962), .A2(new_n2908), .B(new_n2965), .C(new_n3160), .D(new_n3167), .Y(new_n3294));
  INVx1_ASAP7_75t_L         g03038(.A(new_n3126), .Y(new_n3295));
  A2O1A1Ixp33_ASAP7_75t_L   g03039(.A1(new_n2954), .A2(new_n2915), .B(new_n3295), .C(new_n3152), .Y(new_n3296));
  A2O1A1Ixp33_ASAP7_75t_L   g03040(.A1(new_n294), .A2(new_n2932), .B(new_n3135), .C(\a[29] ), .Y(new_n3297));
  O2A1O1Ixp33_ASAP7_75t_L   g03041(.A1(new_n509), .A2(new_n2940), .B(new_n3130), .C(\a[29] ), .Y(new_n3298));
  INVx1_ASAP7_75t_L         g03042(.A(\a[30] ), .Y(new_n3299));
  NAND2xp33_ASAP7_75t_L     g03043(.A(\a[29] ), .B(new_n3299), .Y(new_n3300));
  NAND2xp33_ASAP7_75t_L     g03044(.A(\a[30] ), .B(new_n2928), .Y(new_n3301));
  AND2x2_ASAP7_75t_L        g03045(.A(new_n3300), .B(new_n3301), .Y(new_n3302));
  NOR2xp33_ASAP7_75t_L      g03046(.A(new_n284), .B(new_n3302), .Y(new_n3303));
  INVx1_ASAP7_75t_L         g03047(.A(new_n3303), .Y(new_n3304));
  A2O1A1O1Ixp25_ASAP7_75t_L g03048(.A1(\a[29] ), .A2(new_n3297), .B(new_n3298), .C(new_n2949), .D(new_n3304), .Y(new_n3305));
  NOR2xp33_ASAP7_75t_L      g03049(.A(new_n3303), .B(new_n3148), .Y(new_n3306));
  NAND2xp33_ASAP7_75t_L     g03050(.A(\b[3] ), .B(new_n2938), .Y(new_n3307));
  NAND2xp33_ASAP7_75t_L     g03051(.A(\b[1] ), .B(new_n3129), .Y(new_n3308));
  NAND2xp33_ASAP7_75t_L     g03052(.A(\b[2] ), .B(new_n2936), .Y(new_n3309));
  NAND2xp33_ASAP7_75t_L     g03053(.A(new_n2932), .B(new_n312), .Y(new_n3310));
  NAND5xp2_ASAP7_75t_L      g03054(.A(new_n3310), .B(new_n3309), .C(new_n3308), .D(new_n3307), .E(\a[29] ), .Y(new_n3311));
  OAI211xp5_ASAP7_75t_L     g03055(.A1(new_n3133), .A2(new_n262), .B(new_n3307), .C(new_n3309), .Y(new_n3312));
  A2O1A1Ixp33_ASAP7_75t_L   g03056(.A1(new_n312), .A2(new_n2932), .B(new_n3312), .C(new_n2928), .Y(new_n3313));
  NAND2xp33_ASAP7_75t_L     g03057(.A(new_n3311), .B(new_n3313), .Y(new_n3314));
  OAI21xp33_ASAP7_75t_L     g03058(.A1(new_n3306), .A2(new_n3305), .B(new_n3314), .Y(new_n3315));
  A2O1A1Ixp33_ASAP7_75t_L   g03059(.A1(new_n3132), .A2(new_n3136), .B(new_n2934), .C(new_n3303), .Y(new_n3316));
  A2O1A1Ixp33_ASAP7_75t_L   g03060(.A1(new_n3300), .A2(new_n3301), .B(new_n284), .C(new_n3140), .Y(new_n3317));
  NAND4xp25_ASAP7_75t_L     g03061(.A(new_n3310), .B(new_n3307), .C(new_n3308), .D(new_n3309), .Y(new_n3318));
  A2O1A1Ixp33_ASAP7_75t_L   g03062(.A1(new_n312), .A2(new_n2932), .B(new_n3312), .C(\a[29] ), .Y(new_n3319));
  AOI211xp5_ASAP7_75t_L     g03063(.A1(new_n312), .A2(new_n2932), .B(new_n2928), .C(new_n3312), .Y(new_n3320));
  AOI21xp33_ASAP7_75t_L     g03064(.A1(new_n3319), .A2(new_n3318), .B(new_n3320), .Y(new_n3321));
  NAND3xp33_ASAP7_75t_L     g03065(.A(new_n3317), .B(new_n3316), .C(new_n3321), .Y(new_n3322));
  NOR2xp33_ASAP7_75t_L      g03066(.A(new_n427), .B(new_n2415), .Y(new_n3323));
  AOI221xp5_ASAP7_75t_L     g03067(.A1(\b[4] ), .A2(new_n2577), .B1(\b[5] ), .B2(new_n2421), .C(new_n3323), .Y(new_n3324));
  OA211x2_ASAP7_75t_L       g03068(.A1(new_n2425), .A2(new_n434), .B(\a[26] ), .C(new_n3324), .Y(new_n3325));
  O2A1O1Ixp33_ASAP7_75t_L   g03069(.A1(new_n2425), .A2(new_n434), .B(new_n3324), .C(\a[26] ), .Y(new_n3326));
  NOR2xp33_ASAP7_75t_L      g03070(.A(new_n3326), .B(new_n3325), .Y(new_n3327));
  AND3x1_ASAP7_75t_L        g03071(.A(new_n3322), .B(new_n3315), .C(new_n3327), .Y(new_n3328));
  AOI21xp33_ASAP7_75t_L     g03072(.A1(new_n3322), .A2(new_n3315), .B(new_n3327), .Y(new_n3329));
  AO211x2_ASAP7_75t_L       g03073(.A1(new_n3296), .A2(new_n3151), .B(new_n3329), .C(new_n3328), .Y(new_n3330));
  A2O1A1O1Ixp25_ASAP7_75t_L g03074(.A1(new_n2915), .A2(new_n2954), .B(new_n3295), .C(new_n3152), .D(new_n3147), .Y(new_n3331));
  OAI21xp33_ASAP7_75t_L     g03075(.A1(new_n3328), .A2(new_n3329), .B(new_n3331), .Y(new_n3332));
  NOR2xp33_ASAP7_75t_L      g03076(.A(new_n534), .B(new_n1962), .Y(new_n3333));
  AOI221xp5_ASAP7_75t_L     g03077(.A1(new_n1955), .A2(\b[9] ), .B1(new_n2093), .B2(\b[7] ), .C(new_n3333), .Y(new_n3334));
  INVx1_ASAP7_75t_L         g03078(.A(new_n3334), .Y(new_n3335));
  A2O1A1Ixp33_ASAP7_75t_L   g03079(.A1(new_n602), .A2(new_n1964), .B(new_n3335), .C(\a[23] ), .Y(new_n3336));
  NAND2xp33_ASAP7_75t_L     g03080(.A(\a[23] ), .B(new_n3336), .Y(new_n3337));
  A2O1A1Ixp33_ASAP7_75t_L   g03081(.A1(new_n602), .A2(new_n1964), .B(new_n3335), .C(new_n1952), .Y(new_n3338));
  AOI22xp33_ASAP7_75t_L     g03082(.A1(new_n3337), .A2(new_n3338), .B1(new_n3332), .B2(new_n3330), .Y(new_n3339));
  NOR3xp33_ASAP7_75t_L      g03083(.A(new_n3331), .B(new_n3328), .C(new_n3329), .Y(new_n3340));
  OA21x2_ASAP7_75t_L        g03084(.A1(new_n3328), .A2(new_n3329), .B(new_n3331), .Y(new_n3341));
  NAND2xp33_ASAP7_75t_L     g03085(.A(new_n3338), .B(new_n3337), .Y(new_n3342));
  NOR3xp33_ASAP7_75t_L      g03086(.A(new_n3342), .B(new_n3341), .C(new_n3340), .Y(new_n3343));
  NOR3xp33_ASAP7_75t_L      g03087(.A(new_n3294), .B(new_n3339), .C(new_n3343), .Y(new_n3344));
  OAI21xp33_ASAP7_75t_L     g03088(.A1(new_n3340), .A2(new_n3341), .B(new_n3342), .Y(new_n3345));
  NAND4xp25_ASAP7_75t_L     g03089(.A(new_n3330), .B(new_n3332), .C(new_n3338), .D(new_n3337), .Y(new_n3346));
  AOI221xp5_ASAP7_75t_L     g03090(.A1(new_n3125), .A2(new_n3160), .B1(new_n3345), .B2(new_n3346), .C(new_n3167), .Y(new_n3347));
  OAI21xp33_ASAP7_75t_L     g03091(.A1(new_n3347), .A2(new_n3344), .B(new_n3293), .Y(new_n3348));
  NOR3xp33_ASAP7_75t_L      g03092(.A(new_n3344), .B(new_n3347), .C(new_n3293), .Y(new_n3349));
  INVx1_ASAP7_75t_L         g03093(.A(new_n3349), .Y(new_n3350));
  NAND3xp33_ASAP7_75t_L     g03094(.A(new_n3287), .B(new_n3348), .C(new_n3350), .Y(new_n3351));
  INVx1_ASAP7_75t_L         g03095(.A(new_n3118), .Y(new_n3352));
  NAND2xp33_ASAP7_75t_L     g03096(.A(new_n2978), .B(new_n2975), .Y(new_n3353));
  A2O1A1O1Ixp25_ASAP7_75t_L g03097(.A1(new_n2983), .A2(new_n3353), .B(new_n3352), .C(new_n3173), .D(new_n3170), .Y(new_n3354));
  INVx1_ASAP7_75t_L         g03098(.A(new_n3348), .Y(new_n3355));
  OAI21xp33_ASAP7_75t_L     g03099(.A1(new_n3349), .A2(new_n3355), .B(new_n3354), .Y(new_n3356));
  NOR2xp33_ASAP7_75t_L      g03100(.A(new_n960), .B(new_n2118), .Y(new_n3357));
  AOI221xp5_ASAP7_75t_L     g03101(.A1(\b[13] ), .A2(new_n1290), .B1(\b[15] ), .B2(new_n1209), .C(new_n3357), .Y(new_n3358));
  INVx1_ASAP7_75t_L         g03102(.A(new_n3358), .Y(new_n3359));
  A2O1A1Ixp33_ASAP7_75t_L   g03103(.A1(new_n1052), .A2(new_n1216), .B(new_n3359), .C(\a[17] ), .Y(new_n3360));
  O2A1O1Ixp33_ASAP7_75t_L   g03104(.A1(new_n1210), .A2(new_n1774), .B(new_n3358), .C(\a[17] ), .Y(new_n3361));
  AOI21xp33_ASAP7_75t_L     g03105(.A1(new_n3360), .A2(\a[17] ), .B(new_n3361), .Y(new_n3362));
  NAND3xp33_ASAP7_75t_L     g03106(.A(new_n3351), .B(new_n3362), .C(new_n3356), .Y(new_n3363));
  NOR3xp33_ASAP7_75t_L      g03107(.A(new_n3354), .B(new_n3355), .C(new_n3349), .Y(new_n3364));
  AOI21xp33_ASAP7_75t_L     g03108(.A1(new_n3350), .A2(new_n3348), .B(new_n3287), .Y(new_n3365));
  O2A1O1Ixp33_ASAP7_75t_L   g03109(.A1(new_n1210), .A2(new_n1774), .B(new_n3358), .C(new_n1206), .Y(new_n3366));
  A2O1A1Ixp33_ASAP7_75t_L   g03110(.A1(new_n1052), .A2(new_n1216), .B(new_n3359), .C(new_n1206), .Y(new_n3367));
  OAI21xp33_ASAP7_75t_L     g03111(.A1(new_n1206), .A2(new_n3366), .B(new_n3367), .Y(new_n3368));
  OAI21xp33_ASAP7_75t_L     g03112(.A1(new_n3364), .A2(new_n3365), .B(new_n3368), .Y(new_n3369));
  NOR2xp33_ASAP7_75t_L      g03113(.A(new_n3175), .B(new_n3171), .Y(new_n3370));
  MAJIxp5_ASAP7_75t_L       g03114(.A(new_n3185), .B(new_n3181), .C(new_n3370), .Y(new_n3371));
  NAND3xp33_ASAP7_75t_L     g03115(.A(new_n3371), .B(new_n3369), .C(new_n3363), .Y(new_n3372));
  NAND2xp33_ASAP7_75t_L     g03116(.A(new_n3181), .B(new_n3370), .Y(new_n3373));
  INVx1_ASAP7_75t_L         g03117(.A(new_n3373), .Y(new_n3374));
  NAND2xp33_ASAP7_75t_L     g03118(.A(new_n3363), .B(new_n3369), .Y(new_n3375));
  OAI21xp33_ASAP7_75t_L     g03119(.A1(new_n3374), .A2(new_n3187), .B(new_n3375), .Y(new_n3376));
  NOR2xp33_ASAP7_75t_L      g03120(.A(new_n1349), .B(new_n864), .Y(new_n3377));
  AOI221xp5_ASAP7_75t_L     g03121(.A1(\b[16] ), .A2(new_n985), .B1(\b[18] ), .B2(new_n886), .C(new_n3377), .Y(new_n3378));
  INVx1_ASAP7_75t_L         g03122(.A(new_n3378), .Y(new_n3379));
  A2O1A1Ixp33_ASAP7_75t_L   g03123(.A1(new_n2329), .A2(new_n873), .B(new_n3379), .C(\a[14] ), .Y(new_n3380));
  O2A1O1Ixp33_ASAP7_75t_L   g03124(.A1(new_n872), .A2(new_n1464), .B(new_n3378), .C(\a[14] ), .Y(new_n3381));
  AOI21xp33_ASAP7_75t_L     g03125(.A1(new_n3380), .A2(\a[14] ), .B(new_n3381), .Y(new_n3382));
  NAND3xp33_ASAP7_75t_L     g03126(.A(new_n3376), .B(new_n3372), .C(new_n3382), .Y(new_n3383));
  AND4x1_ASAP7_75t_L        g03127(.A(new_n3201), .B(new_n3373), .C(new_n3369), .D(new_n3363), .Y(new_n3384));
  AOI21xp33_ASAP7_75t_L     g03128(.A1(new_n3369), .A2(new_n3363), .B(new_n3371), .Y(new_n3385));
  O2A1O1Ixp33_ASAP7_75t_L   g03129(.A1(new_n872), .A2(new_n1464), .B(new_n3378), .C(new_n867), .Y(new_n3386));
  A2O1A1Ixp33_ASAP7_75t_L   g03130(.A1(new_n2329), .A2(new_n873), .B(new_n3379), .C(new_n867), .Y(new_n3387));
  OAI21xp33_ASAP7_75t_L     g03131(.A1(new_n867), .A2(new_n3386), .B(new_n3387), .Y(new_n3388));
  OAI21xp33_ASAP7_75t_L     g03132(.A1(new_n3385), .A2(new_n3384), .B(new_n3388), .Y(new_n3389));
  NAND2xp33_ASAP7_75t_L     g03133(.A(new_n3389), .B(new_n3383), .Y(new_n3390));
  NOR2xp33_ASAP7_75t_L      g03134(.A(new_n3186), .B(new_n3187), .Y(new_n3391));
  A2O1A1Ixp33_ASAP7_75t_L   g03135(.A1(\a[14] ), .A2(new_n3202), .B(new_n3203), .C(new_n3391), .Y(new_n3392));
  A2O1A1Ixp33_ASAP7_75t_L   g03136(.A1(new_n3228), .A2(new_n3027), .B(new_n3206), .C(new_n3392), .Y(new_n3393));
  NOR2xp33_ASAP7_75t_L      g03137(.A(new_n3390), .B(new_n3393), .Y(new_n3394));
  NOR3xp33_ASAP7_75t_L      g03138(.A(new_n3384), .B(new_n3385), .C(new_n3388), .Y(new_n3395));
  AOI21xp33_ASAP7_75t_L     g03139(.A1(new_n3376), .A2(new_n3372), .B(new_n3382), .Y(new_n3396));
  NOR2xp33_ASAP7_75t_L      g03140(.A(new_n3395), .B(new_n3396), .Y(new_n3397));
  MAJIxp5_ASAP7_75t_L       g03141(.A(new_n3229), .B(new_n3391), .C(new_n3193), .Y(new_n3398));
  NOR2xp33_ASAP7_75t_L      g03142(.A(new_n3398), .B(new_n3397), .Y(new_n3399));
  NOR2xp33_ASAP7_75t_L      g03143(.A(new_n1895), .B(new_n710), .Y(new_n3400));
  AOI221xp5_ASAP7_75t_L     g03144(.A1(\b[20] ), .A2(new_n635), .B1(\b[19] ), .B2(new_n713), .C(new_n3400), .Y(new_n3401));
  O2A1O1Ixp33_ASAP7_75t_L   g03145(.A1(new_n641), .A2(new_n1901), .B(new_n3401), .C(new_n637), .Y(new_n3402));
  OAI21xp33_ASAP7_75t_L     g03146(.A1(new_n641), .A2(new_n1901), .B(new_n3401), .Y(new_n3403));
  NAND2xp33_ASAP7_75t_L     g03147(.A(new_n637), .B(new_n3403), .Y(new_n3404));
  OAI21xp33_ASAP7_75t_L     g03148(.A1(new_n637), .A2(new_n3402), .B(new_n3404), .Y(new_n3405));
  NOR3xp33_ASAP7_75t_L      g03149(.A(new_n3394), .B(new_n3399), .C(new_n3405), .Y(new_n3406));
  NAND2xp33_ASAP7_75t_L     g03150(.A(new_n3398), .B(new_n3397), .Y(new_n3407));
  INVx1_ASAP7_75t_L         g03151(.A(new_n3392), .Y(new_n3408));
  A2O1A1Ixp33_ASAP7_75t_L   g03152(.A1(new_n3214), .A2(new_n3229), .B(new_n3408), .C(new_n3390), .Y(new_n3409));
  OA21x2_ASAP7_75t_L        g03153(.A1(new_n637), .A2(new_n3402), .B(new_n3404), .Y(new_n3410));
  AOI21xp33_ASAP7_75t_L     g03154(.A1(new_n3409), .A2(new_n3407), .B(new_n3410), .Y(new_n3411));
  NOR3xp33_ASAP7_75t_L      g03155(.A(new_n3237), .B(new_n3406), .C(new_n3411), .Y(new_n3412));
  NAND3xp33_ASAP7_75t_L     g03156(.A(new_n3410), .B(new_n3409), .C(new_n3407), .Y(new_n3413));
  OAI21xp33_ASAP7_75t_L     g03157(.A1(new_n3399), .A2(new_n3394), .B(new_n3405), .Y(new_n3414));
  AOI211xp5_ASAP7_75t_L     g03158(.A1(new_n3414), .A2(new_n3413), .B(new_n3236), .C(new_n3227), .Y(new_n3415));
  NOR2xp33_ASAP7_75t_L      g03159(.A(new_n2188), .B(new_n513), .Y(new_n3416));
  AOI221xp5_ASAP7_75t_L     g03160(.A1(\b[22] ), .A2(new_n560), .B1(\b[24] ), .B2(new_n475), .C(new_n3416), .Y(new_n3417));
  O2A1O1Ixp33_ASAP7_75t_L   g03161(.A1(new_n477), .A2(new_n2853), .B(new_n3417), .C(new_n466), .Y(new_n3418));
  O2A1O1Ixp33_ASAP7_75t_L   g03162(.A1(new_n477), .A2(new_n2853), .B(new_n3417), .C(\a[8] ), .Y(new_n3419));
  INVx1_ASAP7_75t_L         g03163(.A(new_n3419), .Y(new_n3420));
  OAI21xp33_ASAP7_75t_L     g03164(.A1(new_n466), .A2(new_n3418), .B(new_n3420), .Y(new_n3421));
  OAI21xp33_ASAP7_75t_L     g03165(.A1(new_n3412), .A2(new_n3415), .B(new_n3421), .Y(new_n3422));
  OAI211xp5_ASAP7_75t_L     g03166(.A1(new_n3236), .A2(new_n3227), .B(new_n3413), .C(new_n3414), .Y(new_n3423));
  NAND3xp33_ASAP7_75t_L     g03167(.A(new_n3409), .B(new_n3407), .C(new_n3405), .Y(new_n3424));
  A2O1A1Ixp33_ASAP7_75t_L   g03168(.A1(new_n3405), .A2(new_n3424), .B(new_n3406), .C(new_n3237), .Y(new_n3425));
  INVx1_ASAP7_75t_L         g03169(.A(new_n3418), .Y(new_n3426));
  AOI21xp33_ASAP7_75t_L     g03170(.A1(new_n3426), .A2(\a[8] ), .B(new_n3419), .Y(new_n3427));
  NAND3xp33_ASAP7_75t_L     g03171(.A(new_n3423), .B(new_n3425), .C(new_n3427), .Y(new_n3428));
  NAND2xp33_ASAP7_75t_L     g03172(.A(new_n3422), .B(new_n3428), .Y(new_n3429));
  NAND2xp33_ASAP7_75t_L     g03173(.A(new_n3286), .B(new_n3429), .Y(new_n3430));
  A2O1A1Ixp33_ASAP7_75t_L   g03174(.A1(new_n3247), .A2(new_n3251), .B(new_n3257), .C(new_n3244), .Y(new_n3431));
  AOI21xp33_ASAP7_75t_L     g03175(.A1(new_n3423), .A2(new_n3425), .B(new_n3427), .Y(new_n3432));
  NOR3xp33_ASAP7_75t_L      g03176(.A(new_n3415), .B(new_n3412), .C(new_n3421), .Y(new_n3433));
  NOR2xp33_ASAP7_75t_L      g03177(.A(new_n3433), .B(new_n3432), .Y(new_n3434));
  NAND2xp33_ASAP7_75t_L     g03178(.A(new_n3434), .B(new_n3431), .Y(new_n3435));
  NOR2xp33_ASAP7_75t_L      g03179(.A(new_n2377), .B(new_n375), .Y(new_n3436));
  AOI221xp5_ASAP7_75t_L     g03180(.A1(\b[27] ), .A2(new_n361), .B1(new_n349), .B2(\b[26] ), .C(new_n3436), .Y(new_n3437));
  INVx1_ASAP7_75t_L         g03181(.A(new_n3437), .Y(new_n3438));
  A2O1A1Ixp33_ASAP7_75t_L   g03182(.A1(new_n2887), .A2(new_n359), .B(new_n3438), .C(\a[5] ), .Y(new_n3439));
  O2A1O1Ixp33_ASAP7_75t_L   g03183(.A1(new_n356), .A2(new_n2889), .B(new_n3437), .C(\a[5] ), .Y(new_n3440));
  AOI21xp33_ASAP7_75t_L     g03184(.A1(new_n3439), .A2(\a[5] ), .B(new_n3440), .Y(new_n3441));
  NAND3xp33_ASAP7_75t_L     g03185(.A(new_n3435), .B(new_n3430), .C(new_n3441), .Y(new_n3442));
  NAND2xp33_ASAP7_75t_L     g03186(.A(new_n3251), .B(new_n3254), .Y(new_n3443));
  AOI221xp5_ASAP7_75t_L     g03187(.A1(new_n3428), .A2(new_n3422), .B1(new_n3249), .B2(new_n3443), .C(new_n3285), .Y(new_n3444));
  NOR2xp33_ASAP7_75t_L      g03188(.A(new_n3286), .B(new_n3429), .Y(new_n3445));
  O2A1O1Ixp33_ASAP7_75t_L   g03189(.A1(new_n356), .A2(new_n2889), .B(new_n3437), .C(new_n346), .Y(new_n3446));
  A2O1A1Ixp33_ASAP7_75t_L   g03190(.A1(new_n2887), .A2(new_n359), .B(new_n3438), .C(new_n346), .Y(new_n3447));
  OAI21xp33_ASAP7_75t_L     g03191(.A1(new_n346), .A2(new_n3446), .B(new_n3447), .Y(new_n3448));
  OAI21xp33_ASAP7_75t_L     g03192(.A1(new_n3444), .A2(new_n3445), .B(new_n3448), .Y(new_n3449));
  NAND2xp33_ASAP7_75t_L     g03193(.A(new_n3449), .B(new_n3442), .Y(new_n3450));
  A2O1A1O1Ixp25_ASAP7_75t_L g03194(.A1(new_n3064), .A2(new_n3068), .B(new_n3060), .C(new_n3273), .D(new_n3260), .Y(new_n3451));
  XNOR2x2_ASAP7_75t_L       g03195(.A(new_n3450), .B(new_n3451), .Y(new_n3452));
  NOR2xp33_ASAP7_75t_L      g03196(.A(new_n3079), .B(new_n287), .Y(new_n3453));
  AOI221xp5_ASAP7_75t_L     g03197(.A1(\b[29] ), .A2(new_n264), .B1(\b[30] ), .B2(new_n283), .C(new_n3453), .Y(new_n3454));
  NOR2xp33_ASAP7_75t_L      g03198(.A(\b[29] ), .B(\b[30] ), .Y(new_n3455));
  INVx1_ASAP7_75t_L         g03199(.A(\b[30] ), .Y(new_n3456));
  NOR2xp33_ASAP7_75t_L      g03200(.A(new_n3098), .B(new_n3456), .Y(new_n3457));
  NOR2xp33_ASAP7_75t_L      g03201(.A(new_n3455), .B(new_n3457), .Y(new_n3458));
  INVx1_ASAP7_75t_L         g03202(.A(new_n3458), .Y(new_n3459));
  O2A1O1Ixp33_ASAP7_75t_L   g03203(.A1(new_n3079), .A2(new_n3098), .B(new_n3101), .C(new_n3459), .Y(new_n3460));
  INVx1_ASAP7_75t_L         g03204(.A(new_n3460), .Y(new_n3461));
  O2A1O1Ixp33_ASAP7_75t_L   g03205(.A1(new_n3080), .A2(new_n3083), .B(new_n3100), .C(new_n3099), .Y(new_n3462));
  NAND2xp33_ASAP7_75t_L     g03206(.A(new_n3459), .B(new_n3462), .Y(new_n3463));
  NAND2xp33_ASAP7_75t_L     g03207(.A(new_n3463), .B(new_n3461), .Y(new_n3464));
  O2A1O1Ixp33_ASAP7_75t_L   g03208(.A1(new_n279), .A2(new_n3464), .B(new_n3454), .C(new_n257), .Y(new_n3465));
  OAI21xp33_ASAP7_75t_L     g03209(.A1(new_n279), .A2(new_n3464), .B(new_n3454), .Y(new_n3466));
  NAND2xp33_ASAP7_75t_L     g03210(.A(new_n257), .B(new_n3466), .Y(new_n3467));
  OAI21xp33_ASAP7_75t_L     g03211(.A1(new_n257), .A2(new_n3465), .B(new_n3467), .Y(new_n3468));
  NAND2xp33_ASAP7_75t_L     g03212(.A(new_n3468), .B(new_n3452), .Y(new_n3469));
  O2A1O1Ixp33_ASAP7_75t_L   g03213(.A1(new_n3465), .A2(new_n257), .B(new_n3467), .C(new_n3452), .Y(new_n3470));
  AOI21xp33_ASAP7_75t_L     g03214(.A1(new_n3469), .A2(new_n3452), .B(new_n3470), .Y(new_n3471));
  A2O1A1O1Ixp25_ASAP7_75t_L g03215(.A1(new_n3261), .A2(new_n3262), .B(new_n3263), .C(new_n3274), .D(new_n3279), .Y(new_n3472));
  MAJIxp5_ASAP7_75t_L       g03216(.A(new_n3281), .B(new_n3472), .C(new_n3108), .Y(new_n3473));
  XNOR2x2_ASAP7_75t_L       g03217(.A(new_n3473), .B(new_n3471), .Y(\f[30] ));
  NOR2xp33_ASAP7_75t_L      g03218(.A(new_n3385), .B(new_n3384), .Y(new_n3475));
  A2O1A1Ixp33_ASAP7_75t_L   g03219(.A1(\a[14] ), .A2(new_n3380), .B(new_n3381), .C(new_n3475), .Y(new_n3476));
  OAI211xp5_ASAP7_75t_L     g03220(.A1(new_n3325), .A2(new_n3326), .B(new_n3322), .C(new_n3315), .Y(new_n3477));
  A2O1A1O1Ixp25_ASAP7_75t_L g03221(.A1(new_n2944), .A2(new_n2953), .B(new_n2956), .C(new_n3126), .D(new_n3149), .Y(new_n3478));
  OAI22xp33_ASAP7_75t_L     g03222(.A1(new_n3328), .A2(new_n3329), .B1(new_n3147), .B2(new_n3478), .Y(new_n3479));
  NOR2xp33_ASAP7_75t_L      g03223(.A(new_n448), .B(new_n2415), .Y(new_n3480));
  AOI221xp5_ASAP7_75t_L     g03224(.A1(\b[5] ), .A2(new_n2577), .B1(\b[6] ), .B2(new_n2421), .C(new_n3480), .Y(new_n3481));
  O2A1O1Ixp33_ASAP7_75t_L   g03225(.A1(new_n2425), .A2(new_n456), .B(new_n3481), .C(new_n2413), .Y(new_n3482));
  OAI21xp33_ASAP7_75t_L     g03226(.A1(new_n2425), .A2(new_n456), .B(new_n3481), .Y(new_n3483));
  NAND2xp33_ASAP7_75t_L     g03227(.A(new_n2413), .B(new_n3483), .Y(new_n3484));
  OAI21xp33_ASAP7_75t_L     g03228(.A1(new_n2413), .A2(new_n3482), .B(new_n3484), .Y(new_n3485));
  MAJIxp5_ASAP7_75t_L       g03229(.A(new_n3321), .B(new_n3148), .C(new_n3304), .Y(new_n3486));
  NAND2xp33_ASAP7_75t_L     g03230(.A(\b[3] ), .B(new_n2936), .Y(new_n3487));
  OAI221xp5_ASAP7_75t_L     g03231(.A1(new_n2930), .A2(new_n332), .B1(new_n289), .B2(new_n3133), .C(new_n3487), .Y(new_n3488));
  AOI211xp5_ASAP7_75t_L     g03232(.A1(new_n342), .A2(new_n2932), .B(new_n2928), .C(new_n3488), .Y(new_n3489));
  NOR2xp33_ASAP7_75t_L      g03233(.A(new_n332), .B(new_n2930), .Y(new_n3490));
  AOI221xp5_ASAP7_75t_L     g03234(.A1(\b[2] ), .A2(new_n3129), .B1(\b[3] ), .B2(new_n2936), .C(new_n3490), .Y(new_n3491));
  O2A1O1Ixp33_ASAP7_75t_L   g03235(.A1(new_n2940), .A2(new_n1497), .B(new_n3491), .C(\a[29] ), .Y(new_n3492));
  INVx1_ASAP7_75t_L         g03236(.A(\a[32] ), .Y(new_n3493));
  NAND2xp33_ASAP7_75t_L     g03237(.A(new_n3301), .B(new_n3300), .Y(new_n3494));
  INVx1_ASAP7_75t_L         g03238(.A(\a[31] ), .Y(new_n3495));
  NOR2xp33_ASAP7_75t_L      g03239(.A(\a[30] ), .B(new_n3495), .Y(new_n3496));
  NOR2xp33_ASAP7_75t_L      g03240(.A(\a[31] ), .B(new_n3299), .Y(new_n3497));
  NOR2xp33_ASAP7_75t_L      g03241(.A(new_n3496), .B(new_n3497), .Y(new_n3498));
  NOR2xp33_ASAP7_75t_L      g03242(.A(new_n3494), .B(new_n3498), .Y(new_n3499));
  NAND2xp33_ASAP7_75t_L     g03243(.A(\a[32] ), .B(new_n3495), .Y(new_n3500));
  NAND2xp33_ASAP7_75t_L     g03244(.A(\a[31] ), .B(new_n3493), .Y(new_n3501));
  NAND2xp33_ASAP7_75t_L     g03245(.A(new_n3501), .B(new_n3500), .Y(new_n3502));
  NOR2xp33_ASAP7_75t_L      g03246(.A(new_n3502), .B(new_n3302), .Y(new_n3503));
  AOI22xp33_ASAP7_75t_L     g03247(.A1(new_n3499), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n3503), .Y(new_n3504));
  AOI21xp33_ASAP7_75t_L     g03248(.A1(new_n3501), .A2(new_n3500), .B(new_n3302), .Y(new_n3505));
  NAND2xp33_ASAP7_75t_L     g03249(.A(new_n275), .B(new_n3505), .Y(new_n3506));
  NAND2xp33_ASAP7_75t_L     g03250(.A(new_n3506), .B(new_n3504), .Y(new_n3507));
  NOR3xp33_ASAP7_75t_L      g03251(.A(new_n3507), .B(new_n3303), .C(new_n3493), .Y(new_n3508));
  OAI21xp33_ASAP7_75t_L     g03252(.A1(new_n3496), .A2(new_n3497), .B(new_n3302), .Y(new_n3509));
  NAND3xp33_ASAP7_75t_L     g03253(.A(new_n3494), .B(new_n3500), .C(new_n3501), .Y(new_n3510));
  OAI22xp33_ASAP7_75t_L     g03254(.A1(new_n3509), .A2(new_n284), .B1(new_n262), .B2(new_n3510), .Y(new_n3511));
  A2O1A1Ixp33_ASAP7_75t_L   g03255(.A1(new_n3505), .A2(new_n275), .B(new_n3511), .C(\a[32] ), .Y(new_n3512));
  INVx1_ASAP7_75t_L         g03256(.A(new_n3505), .Y(new_n3513));
  O2A1O1Ixp33_ASAP7_75t_L   g03257(.A1(new_n3513), .A2(new_n274), .B(new_n3504), .C(\a[32] ), .Y(new_n3514));
  O2A1O1Ixp33_ASAP7_75t_L   g03258(.A1(new_n3304), .A2(new_n3512), .B(\a[32] ), .C(new_n3514), .Y(new_n3515));
  NOR4xp25_ASAP7_75t_L      g03259(.A(new_n3515), .B(new_n3489), .C(new_n3492), .D(new_n3508), .Y(new_n3516));
  A2O1A1Ixp33_ASAP7_75t_L   g03260(.A1(new_n342), .A2(new_n2932), .B(new_n3488), .C(\a[29] ), .Y(new_n3517));
  A2O1A1O1Ixp25_ASAP7_75t_L g03261(.A1(new_n2932), .A2(new_n342), .B(new_n3488), .C(new_n3517), .D(new_n3489), .Y(new_n3518));
  AOI21xp33_ASAP7_75t_L     g03262(.A1(new_n275), .A2(new_n3505), .B(new_n3511), .Y(new_n3519));
  NAND3xp33_ASAP7_75t_L     g03263(.A(new_n3519), .B(new_n3304), .C(\a[32] ), .Y(new_n3520));
  O2A1O1Ixp33_ASAP7_75t_L   g03264(.A1(new_n3513), .A2(new_n274), .B(new_n3504), .C(new_n3493), .Y(new_n3521));
  A2O1A1Ixp33_ASAP7_75t_L   g03265(.A1(new_n3505), .A2(new_n275), .B(new_n3511), .C(new_n3493), .Y(new_n3522));
  A2O1A1Ixp33_ASAP7_75t_L   g03266(.A1(new_n3521), .A2(new_n3303), .B(new_n3493), .C(new_n3522), .Y(new_n3523));
  AOI21xp33_ASAP7_75t_L     g03267(.A1(new_n3523), .A2(new_n3520), .B(new_n3518), .Y(new_n3524));
  OAI21xp33_ASAP7_75t_L     g03268(.A1(new_n3516), .A2(new_n3524), .B(new_n3486), .Y(new_n3525));
  MAJIxp5_ASAP7_75t_L       g03269(.A(new_n3314), .B(new_n3303), .C(new_n3140), .Y(new_n3526));
  OAI211xp5_ASAP7_75t_L     g03270(.A1(new_n1497), .A2(new_n2940), .B(new_n3491), .C(\a[29] ), .Y(new_n3527));
  A2O1A1Ixp33_ASAP7_75t_L   g03271(.A1(new_n342), .A2(new_n2932), .B(new_n3488), .C(new_n2928), .Y(new_n3528));
  NAND4xp25_ASAP7_75t_L     g03272(.A(new_n3523), .B(new_n3527), .C(new_n3528), .D(new_n3520), .Y(new_n3529));
  OAI22xp33_ASAP7_75t_L     g03273(.A1(new_n3515), .A2(new_n3508), .B1(new_n3492), .B2(new_n3489), .Y(new_n3530));
  NAND3xp33_ASAP7_75t_L     g03274(.A(new_n3526), .B(new_n3529), .C(new_n3530), .Y(new_n3531));
  NAND3xp33_ASAP7_75t_L     g03275(.A(new_n3525), .B(new_n3531), .C(new_n3485), .Y(new_n3532));
  INVx1_ASAP7_75t_L         g03276(.A(new_n3532), .Y(new_n3533));
  AOI21xp33_ASAP7_75t_L     g03277(.A1(new_n3525), .A2(new_n3531), .B(new_n3485), .Y(new_n3534));
  AOI211xp5_ASAP7_75t_L     g03278(.A1(new_n3479), .A2(new_n3477), .B(new_n3533), .C(new_n3534), .Y(new_n3535));
  NAND3xp33_ASAP7_75t_L     g03279(.A(new_n3322), .B(new_n3315), .C(new_n3327), .Y(new_n3536));
  A2O1A1Ixp33_ASAP7_75t_L   g03280(.A1(new_n3536), .A2(new_n3327), .B(new_n3331), .C(new_n3477), .Y(new_n3537));
  INVx1_ASAP7_75t_L         g03281(.A(new_n3534), .Y(new_n3538));
  AOI21xp33_ASAP7_75t_L     g03282(.A1(new_n3538), .A2(new_n3532), .B(new_n3537), .Y(new_n3539));
  NOR2xp33_ASAP7_75t_L      g03283(.A(new_n590), .B(new_n1962), .Y(new_n3540));
  AOI221xp5_ASAP7_75t_L     g03284(.A1(new_n1955), .A2(\b[10] ), .B1(new_n2093), .B2(\b[8] ), .C(new_n3540), .Y(new_n3541));
  O2A1O1Ixp33_ASAP7_75t_L   g03285(.A1(new_n1956), .A2(new_n1175), .B(new_n3541), .C(new_n1952), .Y(new_n3542));
  OAI21xp33_ASAP7_75t_L     g03286(.A1(new_n1956), .A2(new_n1175), .B(new_n3541), .Y(new_n3543));
  NAND2xp33_ASAP7_75t_L     g03287(.A(new_n1952), .B(new_n3543), .Y(new_n3544));
  OAI21xp33_ASAP7_75t_L     g03288(.A1(new_n1952), .A2(new_n3542), .B(new_n3544), .Y(new_n3545));
  NOR3xp33_ASAP7_75t_L      g03289(.A(new_n3535), .B(new_n3539), .C(new_n3545), .Y(new_n3546));
  NAND3xp33_ASAP7_75t_L     g03290(.A(new_n3537), .B(new_n3532), .C(new_n3538), .Y(new_n3547));
  OAI211xp5_ASAP7_75t_L     g03291(.A1(new_n3534), .A2(new_n3533), .B(new_n3479), .C(new_n3477), .Y(new_n3548));
  INVx1_ASAP7_75t_L         g03292(.A(new_n3545), .Y(new_n3549));
  AOI21xp33_ASAP7_75t_L     g03293(.A1(new_n3547), .A2(new_n3548), .B(new_n3549), .Y(new_n3550));
  OAI21xp33_ASAP7_75t_L     g03294(.A1(new_n3343), .A2(new_n3294), .B(new_n3345), .Y(new_n3551));
  NOR3xp33_ASAP7_75t_L      g03295(.A(new_n3551), .B(new_n3550), .C(new_n3546), .Y(new_n3552));
  NAND3xp33_ASAP7_75t_L     g03296(.A(new_n3547), .B(new_n3549), .C(new_n3548), .Y(new_n3553));
  OAI21xp33_ASAP7_75t_L     g03297(.A1(new_n3539), .A2(new_n3535), .B(new_n3545), .Y(new_n3554));
  A2O1A1O1Ixp25_ASAP7_75t_L g03298(.A1(new_n3160), .A2(new_n3125), .B(new_n3167), .C(new_n3346), .D(new_n3339), .Y(new_n3555));
  AOI21xp33_ASAP7_75t_L     g03299(.A1(new_n3554), .A2(new_n3553), .B(new_n3555), .Y(new_n3556));
  NOR2xp33_ASAP7_75t_L      g03300(.A(new_n833), .B(new_n1517), .Y(new_n3557));
  AOI221xp5_ASAP7_75t_L     g03301(.A1(\b[11] ), .A2(new_n1659), .B1(\b[13] ), .B2(new_n1511), .C(new_n3557), .Y(new_n3558));
  INVx1_ASAP7_75t_L         g03302(.A(new_n3558), .Y(new_n3559));
  A2O1A1Ixp33_ASAP7_75t_L   g03303(.A1(new_n1166), .A2(new_n1513), .B(new_n3559), .C(\a[20] ), .Y(new_n3560));
  O2A1O1Ixp33_ASAP7_75t_L   g03304(.A1(new_n1521), .A2(new_n942), .B(new_n3558), .C(\a[20] ), .Y(new_n3561));
  AOI21xp33_ASAP7_75t_L     g03305(.A1(new_n3560), .A2(\a[20] ), .B(new_n3561), .Y(new_n3562));
  OAI21xp33_ASAP7_75t_L     g03306(.A1(new_n3556), .A2(new_n3552), .B(new_n3562), .Y(new_n3563));
  NAND3xp33_ASAP7_75t_L     g03307(.A(new_n3555), .B(new_n3554), .C(new_n3553), .Y(new_n3564));
  OAI21xp33_ASAP7_75t_L     g03308(.A1(new_n3546), .A2(new_n3550), .B(new_n3551), .Y(new_n3565));
  AO21x2_ASAP7_75t_L        g03309(.A1(\a[20] ), .A2(new_n3560), .B(new_n3561), .Y(new_n3566));
  NAND3xp33_ASAP7_75t_L     g03310(.A(new_n3564), .B(new_n3565), .C(new_n3566), .Y(new_n3567));
  OAI21xp33_ASAP7_75t_L     g03311(.A1(new_n3355), .A2(new_n3354), .B(new_n3350), .Y(new_n3568));
  NAND3xp33_ASAP7_75t_L     g03312(.A(new_n3568), .B(new_n3567), .C(new_n3563), .Y(new_n3569));
  AOI21xp33_ASAP7_75t_L     g03313(.A1(new_n3564), .A2(new_n3565), .B(new_n3566), .Y(new_n3570));
  NOR3xp33_ASAP7_75t_L      g03314(.A(new_n3552), .B(new_n3556), .C(new_n3562), .Y(new_n3571));
  A2O1A1O1Ixp25_ASAP7_75t_L g03315(.A1(new_n3173), .A2(new_n3172), .B(new_n3170), .C(new_n3348), .D(new_n3349), .Y(new_n3572));
  OAI21xp33_ASAP7_75t_L     g03316(.A1(new_n3570), .A2(new_n3571), .B(new_n3572), .Y(new_n3573));
  NOR2xp33_ASAP7_75t_L      g03317(.A(new_n1043), .B(new_n2118), .Y(new_n3574));
  AOI221xp5_ASAP7_75t_L     g03318(.A1(\b[14] ), .A2(new_n1290), .B1(\b[16] ), .B2(new_n1209), .C(new_n3574), .Y(new_n3575));
  OAI311xp33_ASAP7_75t_L    g03319(.A1(new_n1155), .A2(new_n1210), .A3(new_n1154), .B1(\a[17] ), .C1(new_n3575), .Y(new_n3576));
  INVx1_ASAP7_75t_L         g03320(.A(new_n3575), .Y(new_n3577));
  A2O1A1Ixp33_ASAP7_75t_L   g03321(.A1(new_n1156), .A2(new_n1216), .B(new_n3577), .C(new_n1206), .Y(new_n3578));
  NAND4xp25_ASAP7_75t_L     g03322(.A(new_n3569), .B(new_n3578), .C(new_n3576), .D(new_n3573), .Y(new_n3579));
  NOR3xp33_ASAP7_75t_L      g03323(.A(new_n3572), .B(new_n3571), .C(new_n3570), .Y(new_n3580));
  AOI221xp5_ASAP7_75t_L     g03324(.A1(new_n3287), .A2(new_n3348), .B1(new_n3563), .B2(new_n3567), .C(new_n3349), .Y(new_n3581));
  NAND2xp33_ASAP7_75t_L     g03325(.A(new_n3576), .B(new_n3578), .Y(new_n3582));
  OAI21xp33_ASAP7_75t_L     g03326(.A1(new_n3581), .A2(new_n3580), .B(new_n3582), .Y(new_n3583));
  NAND2xp33_ASAP7_75t_L     g03327(.A(new_n3583), .B(new_n3579), .Y(new_n3584));
  NAND2xp33_ASAP7_75t_L     g03328(.A(new_n3356), .B(new_n3351), .Y(new_n3585));
  MAJIxp5_ASAP7_75t_L       g03329(.A(new_n3371), .B(new_n3585), .C(new_n3362), .Y(new_n3586));
  NOR2xp33_ASAP7_75t_L      g03330(.A(new_n3586), .B(new_n3584), .Y(new_n3587));
  NOR3xp33_ASAP7_75t_L      g03331(.A(new_n3580), .B(new_n3581), .C(new_n3582), .Y(new_n3588));
  OA21x2_ASAP7_75t_L        g03332(.A1(new_n3581), .A2(new_n3580), .B(new_n3582), .Y(new_n3589));
  NOR2xp33_ASAP7_75t_L      g03333(.A(new_n3588), .B(new_n3589), .Y(new_n3590));
  O2A1O1Ixp33_ASAP7_75t_L   g03334(.A1(new_n3585), .A2(new_n3362), .B(new_n3376), .C(new_n3590), .Y(new_n3591));
  NOR2xp33_ASAP7_75t_L      g03335(.A(new_n1458), .B(new_n864), .Y(new_n3592));
  AOI221xp5_ASAP7_75t_L     g03336(.A1(\b[17] ), .A2(new_n985), .B1(\b[19] ), .B2(new_n886), .C(new_n3592), .Y(new_n3593));
  O2A1O1Ixp33_ASAP7_75t_L   g03337(.A1(new_n872), .A2(new_n1628), .B(new_n3593), .C(new_n867), .Y(new_n3594));
  INVx1_ASAP7_75t_L         g03338(.A(new_n3593), .Y(new_n3595));
  A2O1A1Ixp33_ASAP7_75t_L   g03339(.A1(new_n1607), .A2(new_n873), .B(new_n3595), .C(new_n867), .Y(new_n3596));
  OAI21xp33_ASAP7_75t_L     g03340(.A1(new_n867), .A2(new_n3594), .B(new_n3596), .Y(new_n3597));
  NOR3xp33_ASAP7_75t_L      g03341(.A(new_n3591), .B(new_n3597), .C(new_n3587), .Y(new_n3598));
  O2A1O1Ixp33_ASAP7_75t_L   g03342(.A1(new_n3366), .A2(new_n1206), .B(new_n3367), .C(new_n3585), .Y(new_n3599));
  INVx1_ASAP7_75t_L         g03343(.A(new_n3599), .Y(new_n3600));
  NAND3xp33_ASAP7_75t_L     g03344(.A(new_n3590), .B(new_n3376), .C(new_n3600), .Y(new_n3601));
  NOR2xp33_ASAP7_75t_L      g03345(.A(new_n3581), .B(new_n3580), .Y(new_n3602));
  NAND2xp33_ASAP7_75t_L     g03346(.A(new_n3582), .B(new_n3602), .Y(new_n3603));
  A2O1A1Ixp33_ASAP7_75t_L   g03347(.A1(new_n3603), .A2(new_n3602), .B(new_n3589), .C(new_n3586), .Y(new_n3604));
  A2O1A1Ixp33_ASAP7_75t_L   g03348(.A1(new_n1607), .A2(new_n873), .B(new_n3595), .C(\a[14] ), .Y(new_n3605));
  O2A1O1Ixp33_ASAP7_75t_L   g03349(.A1(new_n872), .A2(new_n1628), .B(new_n3593), .C(\a[14] ), .Y(new_n3606));
  AOI21xp33_ASAP7_75t_L     g03350(.A1(new_n3605), .A2(\a[14] ), .B(new_n3606), .Y(new_n3607));
  AOI21xp33_ASAP7_75t_L     g03351(.A1(new_n3601), .A2(new_n3604), .B(new_n3607), .Y(new_n3608));
  NOR2xp33_ASAP7_75t_L      g03352(.A(new_n3608), .B(new_n3598), .Y(new_n3609));
  NAND3xp33_ASAP7_75t_L     g03353(.A(new_n3609), .B(new_n3409), .C(new_n3476), .Y(new_n3610));
  NAND3xp33_ASAP7_75t_L     g03354(.A(new_n3601), .B(new_n3604), .C(new_n3607), .Y(new_n3611));
  OAI21xp33_ASAP7_75t_L     g03355(.A1(new_n3587), .A2(new_n3591), .B(new_n3597), .Y(new_n3612));
  NAND2xp33_ASAP7_75t_L     g03356(.A(new_n3611), .B(new_n3612), .Y(new_n3613));
  A2O1A1Ixp33_ASAP7_75t_L   g03357(.A1(new_n3382), .A2(new_n3383), .B(new_n3398), .C(new_n3476), .Y(new_n3614));
  NAND2xp33_ASAP7_75t_L     g03358(.A(new_n3613), .B(new_n3614), .Y(new_n3615));
  NOR2xp33_ASAP7_75t_L      g03359(.A(new_n1895), .B(new_n1550), .Y(new_n3616));
  AOI221xp5_ASAP7_75t_L     g03360(.A1(\b[20] ), .A2(new_n713), .B1(\b[22] ), .B2(new_n640), .C(new_n3616), .Y(new_n3617));
  O2A1O1Ixp33_ASAP7_75t_L   g03361(.A1(new_n641), .A2(new_n2522), .B(new_n3617), .C(new_n637), .Y(new_n3618));
  O2A1O1Ixp33_ASAP7_75t_L   g03362(.A1(new_n641), .A2(new_n2522), .B(new_n3617), .C(\a[11] ), .Y(new_n3619));
  INVx1_ASAP7_75t_L         g03363(.A(new_n3619), .Y(new_n3620));
  OA21x2_ASAP7_75t_L        g03364(.A1(new_n637), .A2(new_n3618), .B(new_n3620), .Y(new_n3621));
  NAND3xp33_ASAP7_75t_L     g03365(.A(new_n3610), .B(new_n3621), .C(new_n3615), .Y(new_n3622));
  NOR2xp33_ASAP7_75t_L      g03366(.A(new_n3613), .B(new_n3614), .Y(new_n3623));
  AOI21xp33_ASAP7_75t_L     g03367(.A1(new_n3409), .A2(new_n3476), .B(new_n3609), .Y(new_n3624));
  OAI21xp33_ASAP7_75t_L     g03368(.A1(new_n637), .A2(new_n3618), .B(new_n3620), .Y(new_n3625));
  OAI21xp33_ASAP7_75t_L     g03369(.A1(new_n3623), .A2(new_n3624), .B(new_n3625), .Y(new_n3626));
  OAI22xp33_ASAP7_75t_L     g03370(.A1(new_n3227), .A2(new_n3236), .B1(new_n3411), .B2(new_n3406), .Y(new_n3627));
  NAND4xp25_ASAP7_75t_L     g03371(.A(new_n3627), .B(new_n3424), .C(new_n3622), .D(new_n3626), .Y(new_n3628));
  NOR3xp33_ASAP7_75t_L      g03372(.A(new_n3624), .B(new_n3623), .C(new_n3625), .Y(new_n3629));
  AOI21xp33_ASAP7_75t_L     g03373(.A1(new_n3610), .A2(new_n3615), .B(new_n3621), .Y(new_n3630));
  A2O1A1Ixp33_ASAP7_75t_L   g03374(.A1(new_n3413), .A2(new_n3410), .B(new_n3237), .C(new_n3424), .Y(new_n3631));
  OAI21xp33_ASAP7_75t_L     g03375(.A1(new_n3630), .A2(new_n3629), .B(new_n3631), .Y(new_n3632));
  NOR2xp33_ASAP7_75t_L      g03376(.A(new_n2205), .B(new_n513), .Y(new_n3633));
  AOI221xp5_ASAP7_75t_L     g03377(.A1(\b[23] ), .A2(new_n560), .B1(\b[25] ), .B2(new_n475), .C(new_n3633), .Y(new_n3634));
  O2A1O1Ixp33_ASAP7_75t_L   g03378(.A1(new_n477), .A2(new_n2385), .B(new_n3634), .C(new_n466), .Y(new_n3635));
  INVx1_ASAP7_75t_L         g03379(.A(new_n3635), .Y(new_n3636));
  O2A1O1Ixp33_ASAP7_75t_L   g03380(.A1(new_n477), .A2(new_n2385), .B(new_n3634), .C(\a[8] ), .Y(new_n3637));
  AOI21xp33_ASAP7_75t_L     g03381(.A1(new_n3636), .A2(\a[8] ), .B(new_n3637), .Y(new_n3638));
  NAND3xp33_ASAP7_75t_L     g03382(.A(new_n3628), .B(new_n3638), .C(new_n3632), .Y(new_n3639));
  NOR3xp33_ASAP7_75t_L      g03383(.A(new_n3631), .B(new_n3630), .C(new_n3629), .Y(new_n3640));
  AOI22xp33_ASAP7_75t_L     g03384(.A1(new_n3626), .A2(new_n3622), .B1(new_n3424), .B2(new_n3627), .Y(new_n3641));
  INVx1_ASAP7_75t_L         g03385(.A(new_n3637), .Y(new_n3642));
  OAI21xp33_ASAP7_75t_L     g03386(.A1(new_n466), .A2(new_n3635), .B(new_n3642), .Y(new_n3643));
  OAI21xp33_ASAP7_75t_L     g03387(.A1(new_n3640), .A2(new_n3641), .B(new_n3643), .Y(new_n3644));
  NAND2xp33_ASAP7_75t_L     g03388(.A(new_n3639), .B(new_n3644), .Y(new_n3645));
  OAI21xp33_ASAP7_75t_L     g03389(.A1(new_n3433), .A2(new_n3286), .B(new_n3422), .Y(new_n3646));
  NOR2xp33_ASAP7_75t_L      g03390(.A(new_n3646), .B(new_n3645), .Y(new_n3647));
  A2O1A1O1Ixp25_ASAP7_75t_L g03391(.A1(new_n3249), .A2(new_n3443), .B(new_n3285), .C(new_n3428), .D(new_n3432), .Y(new_n3648));
  AOI21xp33_ASAP7_75t_L     g03392(.A1(new_n3644), .A2(new_n3639), .B(new_n3648), .Y(new_n3649));
  OAI22xp33_ASAP7_75t_L     g03393(.A1(new_n350), .A2(new_n2879), .B1(new_n2703), .B2(new_n375), .Y(new_n3650));
  AOI221xp5_ASAP7_75t_L     g03394(.A1(new_n361), .A2(\b[28] ), .B1(new_n359), .B2(new_n3085), .C(new_n3650), .Y(new_n3651));
  XNOR2x2_ASAP7_75t_L       g03395(.A(\a[5] ), .B(new_n3651), .Y(new_n3652));
  NOR3xp33_ASAP7_75t_L      g03396(.A(new_n3647), .B(new_n3649), .C(new_n3652), .Y(new_n3653));
  NAND3xp33_ASAP7_75t_L     g03397(.A(new_n3648), .B(new_n3644), .C(new_n3639), .Y(new_n3654));
  NAND2xp33_ASAP7_75t_L     g03398(.A(new_n3646), .B(new_n3645), .Y(new_n3655));
  XNOR2x2_ASAP7_75t_L       g03399(.A(new_n346), .B(new_n3651), .Y(new_n3656));
  AOI21xp33_ASAP7_75t_L     g03400(.A1(new_n3654), .A2(new_n3655), .B(new_n3656), .Y(new_n3657));
  NOR2xp33_ASAP7_75t_L      g03401(.A(new_n3657), .B(new_n3653), .Y(new_n3658));
  A2O1A1Ixp33_ASAP7_75t_L   g03402(.A1(new_n2873), .A2(new_n3066), .B(new_n3072), .C(new_n3277), .Y(new_n3659));
  NAND3xp33_ASAP7_75t_L     g03403(.A(new_n3435), .B(new_n3448), .C(new_n3430), .Y(new_n3660));
  INVx1_ASAP7_75t_L         g03404(.A(new_n3660), .Y(new_n3661));
  A2O1A1O1Ixp25_ASAP7_75t_L g03405(.A1(new_n3273), .A2(new_n3659), .B(new_n3260), .C(new_n3450), .D(new_n3661), .Y(new_n3662));
  NAND2xp33_ASAP7_75t_L     g03406(.A(new_n3658), .B(new_n3662), .Y(new_n3663));
  A2O1A1Ixp33_ASAP7_75t_L   g03407(.A1(new_n3272), .A2(new_n3271), .B(new_n3265), .C(new_n3261), .Y(new_n3664));
  NAND3xp33_ASAP7_75t_L     g03408(.A(new_n3654), .B(new_n3655), .C(new_n3656), .Y(new_n3665));
  OAI21xp33_ASAP7_75t_L     g03409(.A1(new_n3649), .A2(new_n3647), .B(new_n3652), .Y(new_n3666));
  NAND2xp33_ASAP7_75t_L     g03410(.A(new_n3665), .B(new_n3666), .Y(new_n3667));
  A2O1A1Ixp33_ASAP7_75t_L   g03411(.A1(new_n3664), .A2(new_n3450), .B(new_n3661), .C(new_n3667), .Y(new_n3668));
  NAND2xp33_ASAP7_75t_L     g03412(.A(new_n3668), .B(new_n3663), .Y(new_n3669));
  NOR2xp33_ASAP7_75t_L      g03413(.A(new_n3098), .B(new_n287), .Y(new_n3670));
  AOI221xp5_ASAP7_75t_L     g03414(.A1(\b[30] ), .A2(new_n264), .B1(\b[31] ), .B2(new_n283), .C(new_n3670), .Y(new_n3671));
  INVx1_ASAP7_75t_L         g03415(.A(new_n3457), .Y(new_n3672));
  NOR2xp33_ASAP7_75t_L      g03416(.A(\b[30] ), .B(\b[31] ), .Y(new_n3673));
  INVx1_ASAP7_75t_L         g03417(.A(\b[31] ), .Y(new_n3674));
  NOR2xp33_ASAP7_75t_L      g03418(.A(new_n3456), .B(new_n3674), .Y(new_n3675));
  NOR2xp33_ASAP7_75t_L      g03419(.A(new_n3673), .B(new_n3675), .Y(new_n3676));
  INVx1_ASAP7_75t_L         g03420(.A(new_n3676), .Y(new_n3677));
  O2A1O1Ixp33_ASAP7_75t_L   g03421(.A1(new_n3459), .A2(new_n3462), .B(new_n3672), .C(new_n3677), .Y(new_n3678));
  INVx1_ASAP7_75t_L         g03422(.A(new_n3678), .Y(new_n3679));
  NAND3xp33_ASAP7_75t_L     g03423(.A(new_n3461), .B(new_n3672), .C(new_n3677), .Y(new_n3680));
  NAND2xp33_ASAP7_75t_L     g03424(.A(new_n3679), .B(new_n3680), .Y(new_n3681));
  O2A1O1Ixp33_ASAP7_75t_L   g03425(.A1(new_n279), .A2(new_n3681), .B(new_n3671), .C(new_n257), .Y(new_n3682));
  O2A1O1Ixp33_ASAP7_75t_L   g03426(.A1(new_n279), .A2(new_n3681), .B(new_n3671), .C(\a[2] ), .Y(new_n3683));
  INVx1_ASAP7_75t_L         g03427(.A(new_n3683), .Y(new_n3684));
  O2A1O1Ixp33_ASAP7_75t_L   g03428(.A1(new_n3682), .A2(new_n257), .B(new_n3684), .C(new_n3669), .Y(new_n3685));
  INVx1_ASAP7_75t_L         g03429(.A(new_n3682), .Y(new_n3686));
  A2O1A1Ixp33_ASAP7_75t_L   g03430(.A1(\a[2] ), .A2(new_n3686), .B(new_n3683), .C(new_n3669), .Y(new_n3687));
  MAJIxp5_ASAP7_75t_L       g03431(.A(new_n3473), .B(new_n3452), .C(new_n3468), .Y(new_n3688));
  O2A1O1Ixp33_ASAP7_75t_L   g03432(.A1(new_n3669), .A2(new_n3685), .B(new_n3687), .C(new_n3688), .Y(new_n3689));
  OAI21xp33_ASAP7_75t_L     g03433(.A1(new_n3669), .A2(new_n3685), .B(new_n3687), .Y(new_n3690));
  INVx1_ASAP7_75t_L         g03434(.A(new_n3688), .Y(new_n3691));
  NOR2xp33_ASAP7_75t_L      g03435(.A(new_n3691), .B(new_n3690), .Y(new_n3692));
  NOR2xp33_ASAP7_75t_L      g03436(.A(new_n3689), .B(new_n3692), .Y(\f[31] ));
  AOI21xp33_ASAP7_75t_L     g03437(.A1(new_n3686), .A2(\a[2] ), .B(new_n3683), .Y(new_n3694));
  MAJIxp5_ASAP7_75t_L       g03438(.A(new_n3688), .B(new_n3669), .C(new_n3694), .Y(new_n3695));
  XOR2x2_ASAP7_75t_L        g03439(.A(new_n3613), .B(new_n3614), .Y(new_n3696));
  MAJIxp5_ASAP7_75t_L       g03440(.A(new_n3631), .B(new_n3625), .C(new_n3696), .Y(new_n3697));
  OAI21xp33_ASAP7_75t_L     g03441(.A1(new_n3570), .A2(new_n3572), .B(new_n3567), .Y(new_n3698));
  NAND2xp33_ASAP7_75t_L     g03442(.A(new_n3548), .B(new_n3547), .Y(new_n3699));
  MAJIxp5_ASAP7_75t_L       g03443(.A(new_n3555), .B(new_n3699), .C(new_n3549), .Y(new_n3700));
  NOR2xp33_ASAP7_75t_L      g03444(.A(new_n3508), .B(new_n3515), .Y(new_n3701));
  A2O1A1Ixp33_ASAP7_75t_L   g03445(.A1(new_n3517), .A2(\a[29] ), .B(new_n3492), .C(new_n3701), .Y(new_n3702));
  NAND3xp33_ASAP7_75t_L     g03446(.A(new_n3302), .B(new_n3498), .C(new_n3502), .Y(new_n3703));
  NAND2xp33_ASAP7_75t_L     g03447(.A(\b[1] ), .B(new_n3499), .Y(new_n3704));
  OAI221xp5_ASAP7_75t_L     g03448(.A1(new_n3510), .A2(new_n289), .B1(new_n284), .B2(new_n3703), .C(new_n3704), .Y(new_n3705));
  A2O1A1Ixp33_ASAP7_75t_L   g03449(.A1(new_n294), .A2(new_n3505), .B(new_n3705), .C(\a[32] ), .Y(new_n3706));
  NOR2xp33_ASAP7_75t_L      g03450(.A(new_n289), .B(new_n3510), .Y(new_n3707));
  AND3x1_ASAP7_75t_L        g03451(.A(new_n3302), .B(new_n3502), .C(new_n3498), .Y(new_n3708));
  AOI221xp5_ASAP7_75t_L     g03452(.A1(new_n3499), .A2(\b[1] ), .B1(new_n3708), .B2(\b[0] ), .C(new_n3707), .Y(new_n3709));
  O2A1O1Ixp33_ASAP7_75t_L   g03453(.A1(new_n509), .A2(new_n3513), .B(new_n3709), .C(\a[32] ), .Y(new_n3710));
  A2O1A1O1Ixp25_ASAP7_75t_L g03454(.A1(new_n3519), .A2(new_n3304), .B(new_n3706), .C(\a[32] ), .D(new_n3710), .Y(new_n3711));
  NAND2xp33_ASAP7_75t_L     g03455(.A(new_n3505), .B(new_n294), .Y(new_n3712));
  INVx1_ASAP7_75t_L         g03456(.A(new_n3712), .Y(new_n3713));
  NOR5xp2_ASAP7_75t_L       g03457(.A(new_n3507), .B(new_n3705), .C(new_n3713), .D(new_n3303), .E(new_n3493), .Y(new_n3714));
  NAND2xp33_ASAP7_75t_L     g03458(.A(\b[4] ), .B(new_n2936), .Y(new_n3715));
  OAI221xp5_ASAP7_75t_L     g03459(.A1(new_n2930), .A2(new_n384), .B1(new_n301), .B2(new_n3133), .C(new_n3715), .Y(new_n3716));
  A2O1A1Ixp33_ASAP7_75t_L   g03460(.A1(new_n394), .A2(new_n2932), .B(new_n3716), .C(\a[29] ), .Y(new_n3717));
  INVx1_ASAP7_75t_L         g03461(.A(new_n3716), .Y(new_n3718));
  O2A1O1Ixp33_ASAP7_75t_L   g03462(.A1(new_n2940), .A2(new_n728), .B(new_n3718), .C(\a[29] ), .Y(new_n3719));
  AOI21xp33_ASAP7_75t_L     g03463(.A1(new_n3717), .A2(\a[29] ), .B(new_n3719), .Y(new_n3720));
  OR3x1_ASAP7_75t_L         g03464(.A(new_n3720), .B(new_n3711), .C(new_n3714), .Y(new_n3721));
  OAI21xp33_ASAP7_75t_L     g03465(.A1(new_n3714), .A2(new_n3711), .B(new_n3720), .Y(new_n3722));
  AOI22xp33_ASAP7_75t_L     g03466(.A1(new_n3721), .A2(new_n3722), .B1(new_n3702), .B2(new_n3525), .Y(new_n3723));
  NAND2xp33_ASAP7_75t_L     g03467(.A(new_n3520), .B(new_n3523), .Y(new_n3724));
  MAJIxp5_ASAP7_75t_L       g03468(.A(new_n3526), .B(new_n3724), .C(new_n3518), .Y(new_n3725));
  NOR3xp33_ASAP7_75t_L      g03469(.A(new_n3720), .B(new_n3711), .C(new_n3714), .Y(new_n3726));
  NAND3xp33_ASAP7_75t_L     g03470(.A(new_n3709), .B(\a[32] ), .C(new_n3712), .Y(new_n3727));
  A2O1A1Ixp33_ASAP7_75t_L   g03471(.A1(new_n294), .A2(new_n3505), .B(new_n3705), .C(new_n3493), .Y(new_n3728));
  NAND3xp33_ASAP7_75t_L     g03472(.A(new_n3520), .B(new_n3727), .C(new_n3728), .Y(new_n3729));
  NAND5xp2_ASAP7_75t_L      g03473(.A(\a[32] ), .B(new_n3519), .C(new_n3712), .D(new_n3709), .E(new_n3304), .Y(new_n3730));
  AOI221xp5_ASAP7_75t_L     g03474(.A1(new_n3717), .A2(\a[29] ), .B1(new_n3730), .B2(new_n3729), .C(new_n3719), .Y(new_n3731));
  NOR3xp33_ASAP7_75t_L      g03475(.A(new_n3725), .B(new_n3726), .C(new_n3731), .Y(new_n3732));
  NOR2xp33_ASAP7_75t_L      g03476(.A(new_n534), .B(new_n2415), .Y(new_n3733));
  AOI221xp5_ASAP7_75t_L     g03477(.A1(\b[6] ), .A2(new_n2577), .B1(\b[7] ), .B2(new_n2421), .C(new_n3733), .Y(new_n3734));
  OAI21xp33_ASAP7_75t_L     g03478(.A1(new_n2425), .A2(new_n540), .B(new_n3734), .Y(new_n3735));
  NOR2xp33_ASAP7_75t_L      g03479(.A(new_n2413), .B(new_n3735), .Y(new_n3736));
  O2A1O1Ixp33_ASAP7_75t_L   g03480(.A1(new_n2425), .A2(new_n540), .B(new_n3734), .C(\a[26] ), .Y(new_n3737));
  NOR2xp33_ASAP7_75t_L      g03481(.A(new_n3737), .B(new_n3736), .Y(new_n3738));
  OAI21xp33_ASAP7_75t_L     g03482(.A1(new_n3732), .A2(new_n3723), .B(new_n3738), .Y(new_n3739));
  OAI21xp33_ASAP7_75t_L     g03483(.A1(new_n3726), .A2(new_n3731), .B(new_n3725), .Y(new_n3740));
  NAND4xp25_ASAP7_75t_L     g03484(.A(new_n3525), .B(new_n3721), .C(new_n3722), .D(new_n3702), .Y(new_n3741));
  O2A1O1Ixp33_ASAP7_75t_L   g03485(.A1(new_n2425), .A2(new_n540), .B(new_n3734), .C(new_n2413), .Y(new_n3742));
  INVx1_ASAP7_75t_L         g03486(.A(new_n3737), .Y(new_n3743));
  OAI21xp33_ASAP7_75t_L     g03487(.A1(new_n2413), .A2(new_n3742), .B(new_n3743), .Y(new_n3744));
  NAND3xp33_ASAP7_75t_L     g03488(.A(new_n3741), .B(new_n3744), .C(new_n3740), .Y(new_n3745));
  NAND2xp33_ASAP7_75t_L     g03489(.A(new_n3745), .B(new_n3739), .Y(new_n3746));
  A2O1A1Ixp33_ASAP7_75t_L   g03490(.A1(new_n3479), .A2(new_n3477), .B(new_n3534), .C(new_n3532), .Y(new_n3747));
  NOR2xp33_ASAP7_75t_L      g03491(.A(new_n3747), .B(new_n3746), .Y(new_n3748));
  INVx1_ASAP7_75t_L         g03492(.A(new_n3725), .Y(new_n3749));
  A2O1A1O1Ixp25_ASAP7_75t_L g03493(.A1(new_n3529), .A2(new_n3530), .B(new_n3526), .C(new_n3702), .D(new_n3731), .Y(new_n3750));
  A2O1A1O1Ixp25_ASAP7_75t_L g03494(.A1(new_n3721), .A2(new_n3750), .B(new_n3749), .C(new_n3741), .D(new_n3738), .Y(new_n3751));
  AOI21xp33_ASAP7_75t_L     g03495(.A1(new_n3537), .A2(new_n3538), .B(new_n3533), .Y(new_n3752));
  O2A1O1Ixp33_ASAP7_75t_L   g03496(.A1(new_n3738), .A2(new_n3751), .B(new_n3739), .C(new_n3752), .Y(new_n3753));
  NOR2xp33_ASAP7_75t_L      g03497(.A(new_n680), .B(new_n1962), .Y(new_n3754));
  AOI221xp5_ASAP7_75t_L     g03498(.A1(new_n1955), .A2(\b[11] ), .B1(new_n2093), .B2(\b[9] ), .C(new_n3754), .Y(new_n3755));
  O2A1O1Ixp33_ASAP7_75t_L   g03499(.A1(new_n1956), .A2(new_n754), .B(new_n3755), .C(new_n1952), .Y(new_n3756));
  INVx1_ASAP7_75t_L         g03500(.A(new_n3755), .Y(new_n3757));
  A2O1A1Ixp33_ASAP7_75t_L   g03501(.A1(new_n976), .A2(new_n1964), .B(new_n3757), .C(new_n1952), .Y(new_n3758));
  OAI21xp33_ASAP7_75t_L     g03502(.A1(new_n1952), .A2(new_n3756), .B(new_n3758), .Y(new_n3759));
  INVx1_ASAP7_75t_L         g03503(.A(new_n3759), .Y(new_n3760));
  NOR3xp33_ASAP7_75t_L      g03504(.A(new_n3753), .B(new_n3760), .C(new_n3748), .Y(new_n3761));
  NAND3xp33_ASAP7_75t_L     g03505(.A(new_n3752), .B(new_n3745), .C(new_n3739), .Y(new_n3762));
  NAND2xp33_ASAP7_75t_L     g03506(.A(new_n3529), .B(new_n3530), .Y(new_n3763));
  INVx1_ASAP7_75t_L         g03507(.A(new_n3517), .Y(new_n3764));
  O2A1O1Ixp33_ASAP7_75t_L   g03508(.A1(new_n2928), .A2(new_n3764), .B(new_n3528), .C(new_n3724), .Y(new_n3765));
  A2O1A1O1Ixp25_ASAP7_75t_L g03509(.A1(new_n3486), .A2(new_n3763), .B(new_n3765), .C(new_n3722), .D(new_n3726), .Y(new_n3766));
  A2O1A1Ixp33_ASAP7_75t_L   g03510(.A1(new_n3766), .A2(new_n3722), .B(new_n3723), .C(new_n3744), .Y(new_n3767));
  A2O1A1O1Ixp25_ASAP7_75t_L g03511(.A1(new_n3721), .A2(new_n3750), .B(new_n3749), .C(new_n3741), .D(new_n3744), .Y(new_n3768));
  A2O1A1Ixp33_ASAP7_75t_L   g03512(.A1(new_n3767), .A2(new_n3744), .B(new_n3768), .C(new_n3747), .Y(new_n3769));
  AOI21xp33_ASAP7_75t_L     g03513(.A1(new_n3762), .A2(new_n3769), .B(new_n3759), .Y(new_n3770));
  OAI21xp33_ASAP7_75t_L     g03514(.A1(new_n3761), .A2(new_n3770), .B(new_n3700), .Y(new_n3771));
  NOR2xp33_ASAP7_75t_L      g03515(.A(new_n3539), .B(new_n3535), .Y(new_n3772));
  MAJIxp5_ASAP7_75t_L       g03516(.A(new_n3551), .B(new_n3545), .C(new_n3772), .Y(new_n3773));
  NAND3xp33_ASAP7_75t_L     g03517(.A(new_n3762), .B(new_n3769), .C(new_n3759), .Y(new_n3774));
  OAI21xp33_ASAP7_75t_L     g03518(.A1(new_n3748), .A2(new_n3753), .B(new_n3760), .Y(new_n3775));
  NAND3xp33_ASAP7_75t_L     g03519(.A(new_n3773), .B(new_n3774), .C(new_n3775), .Y(new_n3776));
  NOR2xp33_ASAP7_75t_L      g03520(.A(new_n936), .B(new_n1517), .Y(new_n3777));
  AOI221xp5_ASAP7_75t_L     g03521(.A1(\b[12] ), .A2(new_n1659), .B1(\b[14] ), .B2(new_n1511), .C(new_n3777), .Y(new_n3778));
  INVx1_ASAP7_75t_L         g03522(.A(new_n3778), .Y(new_n3779));
  A2O1A1Ixp33_ASAP7_75t_L   g03523(.A1(new_n971), .A2(new_n1513), .B(new_n3779), .C(\a[20] ), .Y(new_n3780));
  O2A1O1Ixp33_ASAP7_75t_L   g03524(.A1(new_n1521), .A2(new_n1268), .B(new_n3778), .C(\a[20] ), .Y(new_n3781));
  AOI21xp33_ASAP7_75t_L     g03525(.A1(new_n3780), .A2(\a[20] ), .B(new_n3781), .Y(new_n3782));
  NAND3xp33_ASAP7_75t_L     g03526(.A(new_n3776), .B(new_n3782), .C(new_n3771), .Y(new_n3783));
  AOI21xp33_ASAP7_75t_L     g03527(.A1(new_n3775), .A2(new_n3774), .B(new_n3773), .Y(new_n3784));
  O2A1O1Ixp33_ASAP7_75t_L   g03528(.A1(new_n3542), .A2(new_n1952), .B(new_n3544), .C(new_n3699), .Y(new_n3785));
  NAND2xp33_ASAP7_75t_L     g03529(.A(new_n3553), .B(new_n3554), .Y(new_n3786));
  A2O1A1O1Ixp25_ASAP7_75t_L g03530(.A1(new_n3551), .A2(new_n3786), .B(new_n3785), .C(new_n3775), .D(new_n3761), .Y(new_n3787));
  AO21x2_ASAP7_75t_L        g03531(.A1(\a[20] ), .A2(new_n3780), .B(new_n3781), .Y(new_n3788));
  A2O1A1Ixp33_ASAP7_75t_L   g03532(.A1(new_n3787), .A2(new_n3775), .B(new_n3784), .C(new_n3788), .Y(new_n3789));
  NAND3xp33_ASAP7_75t_L     g03533(.A(new_n3698), .B(new_n3783), .C(new_n3789), .Y(new_n3790));
  A2O1A1O1Ixp25_ASAP7_75t_L g03534(.A1(new_n3348), .A2(new_n3287), .B(new_n3349), .C(new_n3563), .D(new_n3571), .Y(new_n3791));
  AOI211xp5_ASAP7_75t_L     g03535(.A1(new_n3787), .A2(new_n3775), .B(new_n3788), .C(new_n3784), .Y(new_n3792));
  NAND2xp33_ASAP7_75t_L     g03536(.A(new_n3545), .B(new_n3772), .Y(new_n3793));
  A2O1A1O1Ixp25_ASAP7_75t_L g03537(.A1(new_n3553), .A2(new_n3549), .B(new_n3555), .C(new_n3793), .D(new_n3770), .Y(new_n3794));
  A2O1A1O1Ixp25_ASAP7_75t_L g03538(.A1(new_n3774), .A2(new_n3794), .B(new_n3773), .C(new_n3776), .D(new_n3782), .Y(new_n3795));
  OAI21xp33_ASAP7_75t_L     g03539(.A1(new_n3792), .A2(new_n3795), .B(new_n3791), .Y(new_n3796));
  NOR2xp33_ASAP7_75t_L      g03540(.A(new_n1150), .B(new_n2118), .Y(new_n3797));
  AOI221xp5_ASAP7_75t_L     g03541(.A1(\b[15] ), .A2(new_n1290), .B1(\b[17] ), .B2(new_n1209), .C(new_n3797), .Y(new_n3798));
  INVx1_ASAP7_75t_L         g03542(.A(new_n3798), .Y(new_n3799));
  A2O1A1Ixp33_ASAP7_75t_L   g03543(.A1(new_n1633), .A2(new_n1216), .B(new_n3799), .C(\a[17] ), .Y(new_n3800));
  NAND2xp33_ASAP7_75t_L     g03544(.A(\a[17] ), .B(new_n3800), .Y(new_n3801));
  A2O1A1Ixp33_ASAP7_75t_L   g03545(.A1(new_n1633), .A2(new_n1216), .B(new_n3799), .C(new_n1206), .Y(new_n3802));
  NAND4xp25_ASAP7_75t_L     g03546(.A(new_n3790), .B(new_n3802), .C(new_n3796), .D(new_n3801), .Y(new_n3803));
  NOR3xp33_ASAP7_75t_L      g03547(.A(new_n3791), .B(new_n3792), .C(new_n3795), .Y(new_n3804));
  AOI21xp33_ASAP7_75t_L     g03548(.A1(new_n3789), .A2(new_n3783), .B(new_n3698), .Y(new_n3805));
  O2A1O1Ixp33_ASAP7_75t_L   g03549(.A1(new_n1210), .A2(new_n1356), .B(new_n3798), .C(new_n1206), .Y(new_n3806));
  OAI21xp33_ASAP7_75t_L     g03550(.A1(new_n1206), .A2(new_n3806), .B(new_n3802), .Y(new_n3807));
  OAI21xp33_ASAP7_75t_L     g03551(.A1(new_n3805), .A2(new_n3804), .B(new_n3807), .Y(new_n3808));
  NAND2xp33_ASAP7_75t_L     g03552(.A(new_n3803), .B(new_n3808), .Y(new_n3809));
  A2O1A1Ixp33_ASAP7_75t_L   g03553(.A1(new_n3376), .A2(new_n3600), .B(new_n3590), .C(new_n3603), .Y(new_n3810));
  NOR2xp33_ASAP7_75t_L      g03554(.A(new_n3809), .B(new_n3810), .Y(new_n3811));
  INVx1_ASAP7_75t_L         g03555(.A(new_n3586), .Y(new_n3812));
  AND2x2_ASAP7_75t_L        g03556(.A(new_n3803), .B(new_n3808), .Y(new_n3813));
  O2A1O1Ixp33_ASAP7_75t_L   g03557(.A1(new_n3590), .A2(new_n3812), .B(new_n3603), .C(new_n3813), .Y(new_n3814));
  NOR2xp33_ASAP7_75t_L      g03558(.A(new_n1599), .B(new_n864), .Y(new_n3815));
  AOI221xp5_ASAP7_75t_L     g03559(.A1(\b[18] ), .A2(new_n985), .B1(\b[20] ), .B2(new_n886), .C(new_n3815), .Y(new_n3816));
  INVx1_ASAP7_75t_L         g03560(.A(new_n3816), .Y(new_n3817));
  A2O1A1Ixp33_ASAP7_75t_L   g03561(.A1(new_n1752), .A2(new_n873), .B(new_n3817), .C(\a[14] ), .Y(new_n3818));
  O2A1O1Ixp33_ASAP7_75t_L   g03562(.A1(new_n872), .A2(new_n1754), .B(new_n3816), .C(\a[14] ), .Y(new_n3819));
  AOI21xp33_ASAP7_75t_L     g03563(.A1(new_n3818), .A2(\a[14] ), .B(new_n3819), .Y(new_n3820));
  OAI21xp33_ASAP7_75t_L     g03564(.A1(new_n3814), .A2(new_n3811), .B(new_n3820), .Y(new_n3821));
  NOR2xp33_ASAP7_75t_L      g03565(.A(new_n3587), .B(new_n3591), .Y(new_n3822));
  A2O1A1Ixp33_ASAP7_75t_L   g03566(.A1(\a[14] ), .A2(new_n3605), .B(new_n3606), .C(new_n3822), .Y(new_n3823));
  NOR3xp33_ASAP7_75t_L      g03567(.A(new_n3811), .B(new_n3814), .C(new_n3820), .Y(new_n3824));
  INVx1_ASAP7_75t_L         g03568(.A(new_n3824), .Y(new_n3825));
  AOI22xp33_ASAP7_75t_L     g03569(.A1(new_n3825), .A2(new_n3821), .B1(new_n3823), .B2(new_n3615), .Y(new_n3826));
  NAND2xp33_ASAP7_75t_L     g03570(.A(new_n3604), .B(new_n3601), .Y(new_n3827));
  O2A1O1Ixp33_ASAP7_75t_L   g03571(.A1(new_n3594), .A2(new_n867), .B(new_n3596), .C(new_n3827), .Y(new_n3828));
  A2O1A1O1Ixp25_ASAP7_75t_L g03572(.A1(new_n3613), .A2(new_n3614), .B(new_n3828), .C(new_n3821), .D(new_n3824), .Y(new_n3829));
  NOR2xp33_ASAP7_75t_L      g03573(.A(new_n2188), .B(new_n710), .Y(new_n3830));
  AOI221xp5_ASAP7_75t_L     g03574(.A1(\b[22] ), .A2(new_n635), .B1(\b[21] ), .B2(new_n713), .C(new_n3830), .Y(new_n3831));
  O2A1O1Ixp33_ASAP7_75t_L   g03575(.A1(new_n641), .A2(new_n2194), .B(new_n3831), .C(new_n637), .Y(new_n3832));
  OAI21xp33_ASAP7_75t_L     g03576(.A1(new_n641), .A2(new_n2194), .B(new_n3831), .Y(new_n3833));
  NAND2xp33_ASAP7_75t_L     g03577(.A(new_n637), .B(new_n3833), .Y(new_n3834));
  OAI21xp33_ASAP7_75t_L     g03578(.A1(new_n637), .A2(new_n3832), .B(new_n3834), .Y(new_n3835));
  AOI211xp5_ASAP7_75t_L     g03579(.A1(new_n3829), .A2(new_n3821), .B(new_n3835), .C(new_n3826), .Y(new_n3836));
  A2O1A1Ixp33_ASAP7_75t_L   g03580(.A1(new_n3476), .A2(new_n3409), .B(new_n3609), .C(new_n3823), .Y(new_n3837));
  INVx1_ASAP7_75t_L         g03581(.A(new_n3837), .Y(new_n3838));
  INVx1_ASAP7_75t_L         g03582(.A(new_n3603), .Y(new_n3839));
  O2A1O1Ixp33_ASAP7_75t_L   g03583(.A1(new_n3588), .A2(new_n3582), .B(new_n3586), .C(new_n3839), .Y(new_n3840));
  NAND2xp33_ASAP7_75t_L     g03584(.A(new_n3813), .B(new_n3840), .Y(new_n3841));
  A2O1A1Ixp33_ASAP7_75t_L   g03585(.A1(new_n3584), .A2(new_n3586), .B(new_n3839), .C(new_n3809), .Y(new_n3842));
  INVx1_ASAP7_75t_L         g03586(.A(new_n3820), .Y(new_n3843));
  AOI21xp33_ASAP7_75t_L     g03587(.A1(new_n3841), .A2(new_n3842), .B(new_n3843), .Y(new_n3844));
  A2O1A1O1Ixp25_ASAP7_75t_L g03588(.A1(new_n3476), .A2(new_n3409), .B(new_n3609), .C(new_n3823), .D(new_n3844), .Y(new_n3845));
  NAND4xp25_ASAP7_75t_L     g03589(.A(new_n3615), .B(new_n3825), .C(new_n3821), .D(new_n3823), .Y(new_n3846));
  OA21x2_ASAP7_75t_L        g03590(.A1(new_n637), .A2(new_n3832), .B(new_n3834), .Y(new_n3847));
  A2O1A1O1Ixp25_ASAP7_75t_L g03591(.A1(new_n3825), .A2(new_n3845), .B(new_n3838), .C(new_n3846), .D(new_n3847), .Y(new_n3848));
  NOR3xp33_ASAP7_75t_L      g03592(.A(new_n3697), .B(new_n3848), .C(new_n3836), .Y(new_n3849));
  INVx1_ASAP7_75t_L         g03593(.A(new_n3849), .Y(new_n3850));
  OAI21xp33_ASAP7_75t_L     g03594(.A1(new_n3848), .A2(new_n3836), .B(new_n3697), .Y(new_n3851));
  OAI22xp33_ASAP7_75t_L     g03595(.A1(new_n513), .A2(new_n2377), .B1(new_n2205), .B2(new_n506), .Y(new_n3852));
  AOI221xp5_ASAP7_75t_L     g03596(.A1(new_n475), .A2(\b[26] ), .B1(new_n483), .B2(new_n2709), .C(new_n3852), .Y(new_n3853));
  XNOR2x2_ASAP7_75t_L       g03597(.A(new_n466), .B(new_n3853), .Y(new_n3854));
  NAND3xp33_ASAP7_75t_L     g03598(.A(new_n3850), .B(new_n3851), .C(new_n3854), .Y(new_n3855));
  NAND2xp33_ASAP7_75t_L     g03599(.A(new_n3615), .B(new_n3610), .Y(new_n3856));
  O2A1O1Ixp33_ASAP7_75t_L   g03600(.A1(new_n3618), .A2(new_n637), .B(new_n3620), .C(new_n3856), .Y(new_n3857));
  OAI21xp33_ASAP7_75t_L     g03601(.A1(new_n3824), .A2(new_n3844), .B(new_n3837), .Y(new_n3858));
  NAND3xp33_ASAP7_75t_L     g03602(.A(new_n3858), .B(new_n3846), .C(new_n3847), .Y(new_n3859));
  A2O1A1Ixp33_ASAP7_75t_L   g03603(.A1(new_n3829), .A2(new_n3821), .B(new_n3826), .C(new_n3835), .Y(new_n3860));
  AOI211xp5_ASAP7_75t_L     g03604(.A1(new_n3860), .A2(new_n3859), .B(new_n3857), .C(new_n3641), .Y(new_n3861));
  XNOR2x2_ASAP7_75t_L       g03605(.A(\a[8] ), .B(new_n3853), .Y(new_n3862));
  OAI21xp33_ASAP7_75t_L     g03606(.A1(new_n3849), .A2(new_n3861), .B(new_n3862), .Y(new_n3863));
  NAND2xp33_ASAP7_75t_L     g03607(.A(new_n3632), .B(new_n3628), .Y(new_n3864));
  O2A1O1Ixp33_ASAP7_75t_L   g03608(.A1(new_n3635), .A2(new_n466), .B(new_n3642), .C(new_n3864), .Y(new_n3865));
  INVx1_ASAP7_75t_L         g03609(.A(new_n3639), .Y(new_n3866));
  O2A1O1Ixp33_ASAP7_75t_L   g03610(.A1(new_n3643), .A2(new_n3866), .B(new_n3646), .C(new_n3865), .Y(new_n3867));
  NAND3xp33_ASAP7_75t_L     g03611(.A(new_n3867), .B(new_n3863), .C(new_n3855), .Y(new_n3868));
  NOR3xp33_ASAP7_75t_L      g03612(.A(new_n3862), .B(new_n3861), .C(new_n3849), .Y(new_n3869));
  INVx1_ASAP7_75t_L         g03613(.A(new_n3863), .Y(new_n3870));
  MAJIxp5_ASAP7_75t_L       g03614(.A(new_n3648), .B(new_n3864), .C(new_n3638), .Y(new_n3871));
  OAI21xp33_ASAP7_75t_L     g03615(.A1(new_n3869), .A2(new_n3870), .B(new_n3871), .Y(new_n3872));
  AND2x2_ASAP7_75t_L        g03616(.A(new_n3101), .B(new_n3103), .Y(new_n3873));
  OAI22xp33_ASAP7_75t_L     g03617(.A1(new_n350), .A2(new_n3079), .B1(new_n2879), .B2(new_n375), .Y(new_n3874));
  AOI221xp5_ASAP7_75t_L     g03618(.A1(new_n361), .A2(\b[29] ), .B1(new_n359), .B2(new_n3873), .C(new_n3874), .Y(new_n3875));
  XNOR2x2_ASAP7_75t_L       g03619(.A(\a[5] ), .B(new_n3875), .Y(new_n3876));
  AO21x2_ASAP7_75t_L        g03620(.A1(new_n3868), .A2(new_n3872), .B(new_n3876), .Y(new_n3877));
  NOR3xp33_ASAP7_75t_L      g03621(.A(new_n3647), .B(new_n3649), .C(new_n3656), .Y(new_n3878));
  INVx1_ASAP7_75t_L         g03622(.A(new_n3878), .Y(new_n3879));
  NAND3xp33_ASAP7_75t_L     g03623(.A(new_n3876), .B(new_n3872), .C(new_n3868), .Y(new_n3880));
  AOI22xp33_ASAP7_75t_L     g03624(.A1(new_n3880), .A2(new_n3877), .B1(new_n3879), .B2(new_n3668), .Y(new_n3881));
  NOR2xp33_ASAP7_75t_L      g03625(.A(new_n346), .B(new_n3446), .Y(new_n3882));
  NOR3xp33_ASAP7_75t_L      g03626(.A(new_n3445), .B(new_n3448), .C(new_n3444), .Y(new_n3883));
  O2A1O1Ixp33_ASAP7_75t_L   g03627(.A1(new_n3882), .A2(new_n3440), .B(new_n3660), .C(new_n3883), .Y(new_n3884));
  OAI21xp33_ASAP7_75t_L     g03628(.A1(new_n3884), .A2(new_n3451), .B(new_n3660), .Y(new_n3885));
  AND3x1_ASAP7_75t_L        g03629(.A(new_n3876), .B(new_n3872), .C(new_n3868), .Y(new_n3886));
  A2O1A1O1Ixp25_ASAP7_75t_L g03630(.A1(new_n3667), .A2(new_n3885), .B(new_n3878), .C(new_n3877), .D(new_n3886), .Y(new_n3887));
  NOR2xp33_ASAP7_75t_L      g03631(.A(new_n3456), .B(new_n287), .Y(new_n3888));
  AOI221xp5_ASAP7_75t_L     g03632(.A1(\b[31] ), .A2(new_n264), .B1(\b[32] ), .B2(new_n283), .C(new_n3888), .Y(new_n3889));
  NOR2xp33_ASAP7_75t_L      g03633(.A(\b[31] ), .B(\b[32] ), .Y(new_n3890));
  INVx1_ASAP7_75t_L         g03634(.A(\b[32] ), .Y(new_n3891));
  NOR2xp33_ASAP7_75t_L      g03635(.A(new_n3674), .B(new_n3891), .Y(new_n3892));
  NOR2xp33_ASAP7_75t_L      g03636(.A(new_n3890), .B(new_n3892), .Y(new_n3893));
  A2O1A1Ixp33_ASAP7_75t_L   g03637(.A1(\b[31] ), .A2(\b[30] ), .B(new_n3678), .C(new_n3893), .Y(new_n3894));
  O2A1O1Ixp33_ASAP7_75t_L   g03638(.A1(new_n3457), .A2(new_n3460), .B(new_n3676), .C(new_n3675), .Y(new_n3895));
  OAI21xp33_ASAP7_75t_L     g03639(.A1(new_n3890), .A2(new_n3892), .B(new_n3895), .Y(new_n3896));
  NAND2xp33_ASAP7_75t_L     g03640(.A(new_n3894), .B(new_n3896), .Y(new_n3897));
  O2A1O1Ixp33_ASAP7_75t_L   g03641(.A1(new_n279), .A2(new_n3897), .B(new_n3889), .C(new_n257), .Y(new_n3898));
  INVx1_ASAP7_75t_L         g03642(.A(new_n3889), .Y(new_n3899));
  INVx1_ASAP7_75t_L         g03643(.A(new_n3897), .Y(new_n3900));
  A2O1A1Ixp33_ASAP7_75t_L   g03644(.A1(new_n3900), .A2(new_n273), .B(new_n3899), .C(new_n257), .Y(new_n3901));
  OAI21xp33_ASAP7_75t_L     g03645(.A1(new_n257), .A2(new_n3898), .B(new_n3901), .Y(new_n3902));
  INVx1_ASAP7_75t_L         g03646(.A(new_n3902), .Y(new_n3903));
  A2O1A1Ixp33_ASAP7_75t_L   g03647(.A1(new_n3887), .A2(new_n3877), .B(new_n3881), .C(new_n3903), .Y(new_n3904));
  A2O1A1Ixp33_ASAP7_75t_L   g03648(.A1(new_n3273), .A2(new_n3659), .B(new_n3260), .C(new_n3450), .Y(new_n3905));
  A2O1A1Ixp33_ASAP7_75t_L   g03649(.A1(new_n3905), .A2(new_n3660), .B(new_n3658), .C(new_n3879), .Y(new_n3906));
  AOI21xp33_ASAP7_75t_L     g03650(.A1(new_n3872), .A2(new_n3868), .B(new_n3876), .Y(new_n3907));
  OAI21xp33_ASAP7_75t_L     g03651(.A1(new_n3886), .A2(new_n3907), .B(new_n3906), .Y(new_n3908));
  NAND4xp25_ASAP7_75t_L     g03652(.A(new_n3668), .B(new_n3880), .C(new_n3877), .D(new_n3879), .Y(new_n3909));
  NAND3xp33_ASAP7_75t_L     g03653(.A(new_n3908), .B(new_n3909), .C(new_n3902), .Y(new_n3910));
  NAND2xp33_ASAP7_75t_L     g03654(.A(new_n3910), .B(new_n3904), .Y(new_n3911));
  XOR2x2_ASAP7_75t_L        g03655(.A(new_n3911), .B(new_n3695), .Y(\f[32] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03656(.A1(new_n3872), .A2(new_n3868), .B(new_n3876), .C(new_n3887), .D(new_n3881), .Y(new_n3913));
  A2O1A1Ixp33_ASAP7_75t_L   g03657(.A1(new_n3690), .A2(new_n3691), .B(new_n3685), .C(new_n3911), .Y(new_n3914));
  A2O1A1Ixp33_ASAP7_75t_L   g03658(.A1(new_n3668), .A2(new_n3879), .B(new_n3907), .C(new_n3880), .Y(new_n3915));
  INVx1_ASAP7_75t_L         g03659(.A(new_n3618), .Y(new_n3916));
  A2O1A1Ixp33_ASAP7_75t_L   g03660(.A1(\a[11] ), .A2(new_n3916), .B(new_n3619), .C(new_n3696), .Y(new_n3917));
  A2O1A1Ixp33_ASAP7_75t_L   g03661(.A1(new_n3632), .A2(new_n3917), .B(new_n3836), .C(new_n3860), .Y(new_n3918));
  NAND2xp33_ASAP7_75t_L     g03662(.A(new_n3796), .B(new_n3790), .Y(new_n3919));
  O2A1O1Ixp33_ASAP7_75t_L   g03663(.A1(new_n3806), .A2(new_n1206), .B(new_n3802), .C(new_n3919), .Y(new_n3920));
  INVx1_ASAP7_75t_L         g03664(.A(new_n3920), .Y(new_n3921));
  A2O1A1O1Ixp25_ASAP7_75t_L g03665(.A1(new_n3563), .A2(new_n3568), .B(new_n3571), .C(new_n3783), .D(new_n3795), .Y(new_n3922));
  INVx1_ASAP7_75t_L         g03666(.A(\a[33] ), .Y(new_n3923));
  NAND2xp33_ASAP7_75t_L     g03667(.A(\a[32] ), .B(new_n3923), .Y(new_n3924));
  NAND2xp33_ASAP7_75t_L     g03668(.A(\a[33] ), .B(new_n3493), .Y(new_n3925));
  AND2x2_ASAP7_75t_L        g03669(.A(new_n3924), .B(new_n3925), .Y(new_n3926));
  NOR2xp33_ASAP7_75t_L      g03670(.A(new_n284), .B(new_n3926), .Y(new_n3927));
  A2O1A1Ixp33_ASAP7_75t_L   g03671(.A1(new_n3727), .A2(new_n3728), .B(new_n3520), .C(new_n3927), .Y(new_n3928));
  INVx1_ASAP7_75t_L         g03672(.A(new_n3927), .Y(new_n3929));
  NAND2xp33_ASAP7_75t_L     g03673(.A(new_n3929), .B(new_n3714), .Y(new_n3930));
  NAND2xp33_ASAP7_75t_L     g03674(.A(\b[3] ), .B(new_n3503), .Y(new_n3931));
  NAND2xp33_ASAP7_75t_L     g03675(.A(\b[1] ), .B(new_n3708), .Y(new_n3932));
  NAND2xp33_ASAP7_75t_L     g03676(.A(\b[2] ), .B(new_n3499), .Y(new_n3933));
  NAND2xp33_ASAP7_75t_L     g03677(.A(new_n3505), .B(new_n312), .Y(new_n3934));
  NAND4xp25_ASAP7_75t_L     g03678(.A(new_n3934), .B(new_n3931), .C(new_n3932), .D(new_n3933), .Y(new_n3935));
  OAI211xp5_ASAP7_75t_L     g03679(.A1(new_n3703), .A2(new_n262), .B(new_n3931), .C(new_n3933), .Y(new_n3936));
  A2O1A1Ixp33_ASAP7_75t_L   g03680(.A1(new_n312), .A2(new_n3505), .B(new_n3936), .C(\a[32] ), .Y(new_n3937));
  AOI211xp5_ASAP7_75t_L     g03681(.A1(new_n312), .A2(new_n3505), .B(new_n3493), .C(new_n3936), .Y(new_n3938));
  AOI21xp33_ASAP7_75t_L     g03682(.A1(new_n3937), .A2(new_n3935), .B(new_n3938), .Y(new_n3939));
  AOI21xp33_ASAP7_75t_L     g03683(.A1(new_n3930), .A2(new_n3928), .B(new_n3939), .Y(new_n3940));
  A2O1A1O1Ixp25_ASAP7_75t_L g03684(.A1(\a[32] ), .A2(new_n3706), .B(new_n3710), .C(new_n3508), .D(new_n3929), .Y(new_n3941));
  NOR2xp33_ASAP7_75t_L      g03685(.A(new_n3927), .B(new_n3730), .Y(new_n3942));
  NAND5xp2_ASAP7_75t_L      g03686(.A(new_n3934), .B(new_n3933), .C(new_n3932), .D(new_n3931), .E(\a[32] ), .Y(new_n3943));
  A2O1A1Ixp33_ASAP7_75t_L   g03687(.A1(new_n312), .A2(new_n3505), .B(new_n3936), .C(new_n3493), .Y(new_n3944));
  NAND2xp33_ASAP7_75t_L     g03688(.A(new_n3943), .B(new_n3944), .Y(new_n3945));
  NOR3xp33_ASAP7_75t_L      g03689(.A(new_n3941), .B(new_n3942), .C(new_n3945), .Y(new_n3946));
  NOR2xp33_ASAP7_75t_L      g03690(.A(new_n427), .B(new_n2930), .Y(new_n3947));
  AOI221xp5_ASAP7_75t_L     g03691(.A1(\b[4] ), .A2(new_n3129), .B1(\b[5] ), .B2(new_n2936), .C(new_n3947), .Y(new_n3948));
  O2A1O1Ixp33_ASAP7_75t_L   g03692(.A1(new_n2940), .A2(new_n434), .B(new_n3948), .C(new_n2928), .Y(new_n3949));
  OAI31xp33_ASAP7_75t_L     g03693(.A1(new_n433), .A2(new_n431), .A3(new_n2940), .B(new_n3948), .Y(new_n3950));
  NAND2xp33_ASAP7_75t_L     g03694(.A(new_n2928), .B(new_n3950), .Y(new_n3951));
  OAI21xp33_ASAP7_75t_L     g03695(.A1(new_n2928), .A2(new_n3949), .B(new_n3951), .Y(new_n3952));
  NOR3xp33_ASAP7_75t_L      g03696(.A(new_n3946), .B(new_n3940), .C(new_n3952), .Y(new_n3953));
  OAI21xp33_ASAP7_75t_L     g03697(.A1(new_n3942), .A2(new_n3941), .B(new_n3945), .Y(new_n3954));
  NAND3xp33_ASAP7_75t_L     g03698(.A(new_n3930), .B(new_n3928), .C(new_n3939), .Y(new_n3955));
  OA21x2_ASAP7_75t_L        g03699(.A1(new_n2928), .A2(new_n3949), .B(new_n3951), .Y(new_n3956));
  AOI21xp33_ASAP7_75t_L     g03700(.A1(new_n3954), .A2(new_n3955), .B(new_n3956), .Y(new_n3957));
  NOR3xp33_ASAP7_75t_L      g03701(.A(new_n3766), .B(new_n3953), .C(new_n3957), .Y(new_n3958));
  NAND3xp33_ASAP7_75t_L     g03702(.A(new_n3954), .B(new_n3956), .C(new_n3955), .Y(new_n3959));
  OAI21xp33_ASAP7_75t_L     g03703(.A1(new_n3940), .A2(new_n3946), .B(new_n3952), .Y(new_n3960));
  AOI211xp5_ASAP7_75t_L     g03704(.A1(new_n3960), .A2(new_n3959), .B(new_n3726), .C(new_n3750), .Y(new_n3961));
  NOR2xp33_ASAP7_75t_L      g03705(.A(new_n534), .B(new_n2410), .Y(new_n3962));
  AOI221xp5_ASAP7_75t_L     g03706(.A1(\b[7] ), .A2(new_n2577), .B1(\b[9] ), .B2(new_n2423), .C(new_n3962), .Y(new_n3963));
  O2A1O1Ixp33_ASAP7_75t_L   g03707(.A1(new_n2425), .A2(new_n1066), .B(new_n3963), .C(new_n2413), .Y(new_n3964));
  INVx1_ASAP7_75t_L         g03708(.A(new_n3963), .Y(new_n3965));
  A2O1A1Ixp33_ASAP7_75t_L   g03709(.A1(new_n602), .A2(new_n2417), .B(new_n3965), .C(new_n2413), .Y(new_n3966));
  OAI21xp33_ASAP7_75t_L     g03710(.A1(new_n2413), .A2(new_n3964), .B(new_n3966), .Y(new_n3967));
  OAI21xp33_ASAP7_75t_L     g03711(.A1(new_n3961), .A2(new_n3958), .B(new_n3967), .Y(new_n3968));
  OAI211xp5_ASAP7_75t_L     g03712(.A1(new_n3726), .A2(new_n3750), .B(new_n3959), .C(new_n3960), .Y(new_n3969));
  OAI21xp33_ASAP7_75t_L     g03713(.A1(new_n3953), .A2(new_n3957), .B(new_n3766), .Y(new_n3970));
  A2O1A1Ixp33_ASAP7_75t_L   g03714(.A1(new_n602), .A2(new_n2417), .B(new_n3965), .C(\a[26] ), .Y(new_n3971));
  NAND2xp33_ASAP7_75t_L     g03715(.A(\a[26] ), .B(new_n3971), .Y(new_n3972));
  NAND4xp25_ASAP7_75t_L     g03716(.A(new_n3969), .B(new_n3970), .C(new_n3966), .D(new_n3972), .Y(new_n3973));
  AOI221xp5_ASAP7_75t_L     g03717(.A1(new_n3968), .A2(new_n3973), .B1(new_n3747), .B2(new_n3746), .C(new_n3751), .Y(new_n3974));
  INVx1_ASAP7_75t_L         g03718(.A(new_n3974), .Y(new_n3975));
  A2O1A1Ixp33_ASAP7_75t_L   g03719(.A1(new_n3738), .A2(new_n3739), .B(new_n3752), .C(new_n3767), .Y(new_n3976));
  NAND3xp33_ASAP7_75t_L     g03720(.A(new_n3976), .B(new_n3968), .C(new_n3973), .Y(new_n3977));
  NOR2xp33_ASAP7_75t_L      g03721(.A(new_n748), .B(new_n1962), .Y(new_n3978));
  AOI221xp5_ASAP7_75t_L     g03722(.A1(new_n1955), .A2(\b[12] ), .B1(new_n2093), .B2(\b[10] ), .C(new_n3978), .Y(new_n3979));
  O2A1O1Ixp33_ASAP7_75t_L   g03723(.A1(new_n1956), .A2(new_n841), .B(new_n3979), .C(new_n1952), .Y(new_n3980));
  INVx1_ASAP7_75t_L         g03724(.A(new_n3980), .Y(new_n3981));
  O2A1O1Ixp33_ASAP7_75t_L   g03725(.A1(new_n1956), .A2(new_n841), .B(new_n3979), .C(\a[23] ), .Y(new_n3982));
  AO21x2_ASAP7_75t_L        g03726(.A1(\a[23] ), .A2(new_n3981), .B(new_n3982), .Y(new_n3983));
  AOI21xp33_ASAP7_75t_L     g03727(.A1(new_n3977), .A2(new_n3975), .B(new_n3983), .Y(new_n3984));
  O2A1O1Ixp33_ASAP7_75t_L   g03728(.A1(new_n3736), .A2(new_n3737), .B(new_n3767), .C(new_n3768), .Y(new_n3985));
  NAND2xp33_ASAP7_75t_L     g03729(.A(new_n3973), .B(new_n3968), .Y(new_n3986));
  O2A1O1Ixp33_ASAP7_75t_L   g03730(.A1(new_n3985), .A2(new_n3752), .B(new_n3767), .C(new_n3986), .Y(new_n3987));
  AOI21xp33_ASAP7_75t_L     g03731(.A1(new_n3981), .A2(\a[23] ), .B(new_n3982), .Y(new_n3988));
  NOR3xp33_ASAP7_75t_L      g03732(.A(new_n3987), .B(new_n3988), .C(new_n3974), .Y(new_n3989));
  NOR3xp33_ASAP7_75t_L      g03733(.A(new_n3787), .B(new_n3984), .C(new_n3989), .Y(new_n3990));
  OAI21xp33_ASAP7_75t_L     g03734(.A1(new_n3974), .A2(new_n3987), .B(new_n3988), .Y(new_n3991));
  NAND3xp33_ASAP7_75t_L     g03735(.A(new_n3977), .B(new_n3975), .C(new_n3983), .Y(new_n3992));
  AOI211xp5_ASAP7_75t_L     g03736(.A1(new_n3992), .A2(new_n3991), .B(new_n3761), .C(new_n3794), .Y(new_n3993));
  NOR2xp33_ASAP7_75t_L      g03737(.A(new_n960), .B(new_n1517), .Y(new_n3994));
  AOI221xp5_ASAP7_75t_L     g03738(.A1(\b[13] ), .A2(new_n1659), .B1(\b[15] ), .B2(new_n1511), .C(new_n3994), .Y(new_n3995));
  O2A1O1Ixp33_ASAP7_75t_L   g03739(.A1(new_n1521), .A2(new_n1774), .B(new_n3995), .C(new_n1501), .Y(new_n3996));
  INVx1_ASAP7_75t_L         g03740(.A(new_n3995), .Y(new_n3997));
  A2O1A1Ixp33_ASAP7_75t_L   g03741(.A1(new_n1052), .A2(new_n1513), .B(new_n3997), .C(new_n1501), .Y(new_n3998));
  OAI21xp33_ASAP7_75t_L     g03742(.A1(new_n1501), .A2(new_n3996), .B(new_n3998), .Y(new_n3999));
  NOR3xp33_ASAP7_75t_L      g03743(.A(new_n3990), .B(new_n3993), .C(new_n3999), .Y(new_n4000));
  OAI211xp5_ASAP7_75t_L     g03744(.A1(new_n3761), .A2(new_n3794), .B(new_n3991), .C(new_n3992), .Y(new_n4001));
  OAI21xp33_ASAP7_75t_L     g03745(.A1(new_n3984), .A2(new_n3989), .B(new_n3787), .Y(new_n4002));
  A2O1A1Ixp33_ASAP7_75t_L   g03746(.A1(new_n1052), .A2(new_n1513), .B(new_n3997), .C(\a[20] ), .Y(new_n4003));
  O2A1O1Ixp33_ASAP7_75t_L   g03747(.A1(new_n1521), .A2(new_n1774), .B(new_n3995), .C(\a[20] ), .Y(new_n4004));
  AOI21xp33_ASAP7_75t_L     g03748(.A1(new_n4003), .A2(\a[20] ), .B(new_n4004), .Y(new_n4005));
  AOI21xp33_ASAP7_75t_L     g03749(.A1(new_n4001), .A2(new_n4002), .B(new_n4005), .Y(new_n4006));
  NOR3xp33_ASAP7_75t_L      g03750(.A(new_n3922), .B(new_n4000), .C(new_n4006), .Y(new_n4007));
  NAND3xp33_ASAP7_75t_L     g03751(.A(new_n4001), .B(new_n4005), .C(new_n4002), .Y(new_n4008));
  OAI21xp33_ASAP7_75t_L     g03752(.A1(new_n3993), .A2(new_n3990), .B(new_n3999), .Y(new_n4009));
  AOI221xp5_ASAP7_75t_L     g03753(.A1(new_n3698), .A2(new_n3783), .B1(new_n4008), .B2(new_n4009), .C(new_n3795), .Y(new_n4010));
  NOR2xp33_ASAP7_75t_L      g03754(.A(new_n1349), .B(new_n2118), .Y(new_n4011));
  AOI221xp5_ASAP7_75t_L     g03755(.A1(\b[16] ), .A2(new_n1290), .B1(\b[18] ), .B2(new_n1209), .C(new_n4011), .Y(new_n4012));
  O2A1O1Ixp33_ASAP7_75t_L   g03756(.A1(new_n1210), .A2(new_n1464), .B(new_n4012), .C(new_n1206), .Y(new_n4013));
  INVx1_ASAP7_75t_L         g03757(.A(new_n4012), .Y(new_n4014));
  A2O1A1Ixp33_ASAP7_75t_L   g03758(.A1(new_n2329), .A2(new_n1216), .B(new_n4014), .C(new_n1206), .Y(new_n4015));
  OAI21xp33_ASAP7_75t_L     g03759(.A1(new_n1206), .A2(new_n4013), .B(new_n4015), .Y(new_n4016));
  OAI21xp33_ASAP7_75t_L     g03760(.A1(new_n4010), .A2(new_n4007), .B(new_n4016), .Y(new_n4017));
  OAI21xp33_ASAP7_75t_L     g03761(.A1(new_n3792), .A2(new_n3791), .B(new_n3789), .Y(new_n4018));
  NAND3xp33_ASAP7_75t_L     g03762(.A(new_n4018), .B(new_n4008), .C(new_n4009), .Y(new_n4019));
  OAI21xp33_ASAP7_75t_L     g03763(.A1(new_n4000), .A2(new_n4006), .B(new_n3922), .Y(new_n4020));
  A2O1A1Ixp33_ASAP7_75t_L   g03764(.A1(new_n2329), .A2(new_n1216), .B(new_n4014), .C(\a[17] ), .Y(new_n4021));
  O2A1O1Ixp33_ASAP7_75t_L   g03765(.A1(new_n1210), .A2(new_n1464), .B(new_n4012), .C(\a[17] ), .Y(new_n4022));
  AOI21xp33_ASAP7_75t_L     g03766(.A1(new_n4021), .A2(\a[17] ), .B(new_n4022), .Y(new_n4023));
  NAND3xp33_ASAP7_75t_L     g03767(.A(new_n4019), .B(new_n4020), .C(new_n4023), .Y(new_n4024));
  NAND2xp33_ASAP7_75t_L     g03768(.A(new_n4024), .B(new_n4017), .Y(new_n4025));
  NAND3xp33_ASAP7_75t_L     g03769(.A(new_n3842), .B(new_n4025), .C(new_n3921), .Y(new_n4026));
  AOI21xp33_ASAP7_75t_L     g03770(.A1(new_n4019), .A2(new_n4020), .B(new_n4023), .Y(new_n4027));
  NOR3xp33_ASAP7_75t_L      g03771(.A(new_n4007), .B(new_n4016), .C(new_n4010), .Y(new_n4028));
  NOR2xp33_ASAP7_75t_L      g03772(.A(new_n4027), .B(new_n4028), .Y(new_n4029));
  A2O1A1Ixp33_ASAP7_75t_L   g03773(.A1(new_n3809), .A2(new_n3810), .B(new_n3920), .C(new_n4029), .Y(new_n4030));
  NOR2xp33_ASAP7_75t_L      g03774(.A(new_n1745), .B(new_n864), .Y(new_n4031));
  AOI221xp5_ASAP7_75t_L     g03775(.A1(\b[19] ), .A2(new_n985), .B1(\b[21] ), .B2(new_n886), .C(new_n4031), .Y(new_n4032));
  INVx1_ASAP7_75t_L         g03776(.A(new_n4032), .Y(new_n4033));
  A2O1A1Ixp33_ASAP7_75t_L   g03777(.A1(new_n2836), .A2(new_n873), .B(new_n4033), .C(\a[14] ), .Y(new_n4034));
  O2A1O1Ixp33_ASAP7_75t_L   g03778(.A1(new_n872), .A2(new_n1901), .B(new_n4032), .C(\a[14] ), .Y(new_n4035));
  AOI21xp33_ASAP7_75t_L     g03779(.A1(new_n4034), .A2(\a[14] ), .B(new_n4035), .Y(new_n4036));
  NAND3xp33_ASAP7_75t_L     g03780(.A(new_n4030), .B(new_n4026), .C(new_n4036), .Y(new_n4037));
  AOI221xp5_ASAP7_75t_L     g03781(.A1(new_n4024), .A2(new_n4017), .B1(new_n3809), .B2(new_n3810), .C(new_n3920), .Y(new_n4038));
  O2A1O1Ixp33_ASAP7_75t_L   g03782(.A1(new_n3813), .A2(new_n3840), .B(new_n3921), .C(new_n4025), .Y(new_n4039));
  O2A1O1Ixp33_ASAP7_75t_L   g03783(.A1(new_n872), .A2(new_n1901), .B(new_n4032), .C(new_n867), .Y(new_n4040));
  INVx1_ASAP7_75t_L         g03784(.A(new_n4035), .Y(new_n4041));
  OAI21xp33_ASAP7_75t_L     g03785(.A1(new_n867), .A2(new_n4040), .B(new_n4041), .Y(new_n4042));
  OAI21xp33_ASAP7_75t_L     g03786(.A1(new_n4038), .A2(new_n4039), .B(new_n4042), .Y(new_n4043));
  OAI211xp5_ASAP7_75t_L     g03787(.A1(new_n3824), .A2(new_n3845), .B(new_n4037), .C(new_n4043), .Y(new_n4044));
  NAND2xp33_ASAP7_75t_L     g03788(.A(new_n4043), .B(new_n4037), .Y(new_n4045));
  NAND2xp33_ASAP7_75t_L     g03789(.A(new_n3829), .B(new_n4045), .Y(new_n4046));
  NOR2xp33_ASAP7_75t_L      g03790(.A(new_n2188), .B(new_n1550), .Y(new_n4047));
  AOI221xp5_ASAP7_75t_L     g03791(.A1(\b[22] ), .A2(new_n713), .B1(\b[24] ), .B2(new_n640), .C(new_n4047), .Y(new_n4048));
  O2A1O1Ixp33_ASAP7_75t_L   g03792(.A1(new_n641), .A2(new_n2853), .B(new_n4048), .C(new_n637), .Y(new_n4049));
  INVx1_ASAP7_75t_L         g03793(.A(new_n4049), .Y(new_n4050));
  O2A1O1Ixp33_ASAP7_75t_L   g03794(.A1(new_n641), .A2(new_n2853), .B(new_n4048), .C(\a[11] ), .Y(new_n4051));
  AOI21xp33_ASAP7_75t_L     g03795(.A1(new_n4050), .A2(\a[11] ), .B(new_n4051), .Y(new_n4052));
  NAND3xp33_ASAP7_75t_L     g03796(.A(new_n4044), .B(new_n4046), .C(new_n4052), .Y(new_n4053));
  NOR2xp33_ASAP7_75t_L      g03797(.A(new_n3829), .B(new_n4045), .Y(new_n4054));
  AOI211xp5_ASAP7_75t_L     g03798(.A1(new_n4043), .A2(new_n4037), .B(new_n3824), .C(new_n3845), .Y(new_n4055));
  NOR2xp33_ASAP7_75t_L      g03799(.A(new_n637), .B(new_n4049), .Y(new_n4056));
  OAI22xp33_ASAP7_75t_L     g03800(.A1(new_n4055), .A2(new_n4054), .B1(new_n4051), .B2(new_n4056), .Y(new_n4057));
  NAND3xp33_ASAP7_75t_L     g03801(.A(new_n3918), .B(new_n4053), .C(new_n4057), .Y(new_n4058));
  NAND2xp33_ASAP7_75t_L     g03802(.A(new_n3622), .B(new_n3626), .Y(new_n4059));
  A2O1A1O1Ixp25_ASAP7_75t_L g03803(.A1(new_n3631), .A2(new_n4059), .B(new_n3857), .C(new_n3859), .D(new_n3848), .Y(new_n4060));
  NAND2xp33_ASAP7_75t_L     g03804(.A(new_n4053), .B(new_n4057), .Y(new_n4061));
  NAND2xp33_ASAP7_75t_L     g03805(.A(new_n4060), .B(new_n4061), .Y(new_n4062));
  NOR2xp33_ASAP7_75t_L      g03806(.A(new_n2703), .B(new_n513), .Y(new_n4063));
  AOI221xp5_ASAP7_75t_L     g03807(.A1(\b[25] ), .A2(new_n560), .B1(\b[27] ), .B2(new_n475), .C(new_n4063), .Y(new_n4064));
  O2A1O1Ixp33_ASAP7_75t_L   g03808(.A1(new_n477), .A2(new_n2889), .B(new_n4064), .C(new_n466), .Y(new_n4065));
  INVx1_ASAP7_75t_L         g03809(.A(new_n4065), .Y(new_n4066));
  O2A1O1Ixp33_ASAP7_75t_L   g03810(.A1(new_n477), .A2(new_n2889), .B(new_n4064), .C(\a[8] ), .Y(new_n4067));
  AOI21xp33_ASAP7_75t_L     g03811(.A1(new_n4066), .A2(\a[8] ), .B(new_n4067), .Y(new_n4068));
  NAND3xp33_ASAP7_75t_L     g03812(.A(new_n4068), .B(new_n4062), .C(new_n4058), .Y(new_n4069));
  NOR2xp33_ASAP7_75t_L      g03813(.A(new_n4060), .B(new_n4061), .Y(new_n4070));
  AOI21xp33_ASAP7_75t_L     g03814(.A1(new_n4057), .A2(new_n4053), .B(new_n3918), .Y(new_n4071));
  NOR2xp33_ASAP7_75t_L      g03815(.A(new_n466), .B(new_n4065), .Y(new_n4072));
  OAI22xp33_ASAP7_75t_L     g03816(.A1(new_n4070), .A2(new_n4071), .B1(new_n4067), .B2(new_n4072), .Y(new_n4073));
  NOR3xp33_ASAP7_75t_L      g03817(.A(new_n3854), .B(new_n3861), .C(new_n3849), .Y(new_n4074));
  O2A1O1Ixp33_ASAP7_75t_L   g03818(.A1(new_n3869), .A2(new_n3862), .B(new_n3871), .C(new_n4074), .Y(new_n4075));
  NAND3xp33_ASAP7_75t_L     g03819(.A(new_n4075), .B(new_n4073), .C(new_n4069), .Y(new_n4076));
  NAND2xp33_ASAP7_75t_L     g03820(.A(new_n4069), .B(new_n4073), .Y(new_n4077));
  NOR2xp33_ASAP7_75t_L      g03821(.A(new_n3849), .B(new_n3861), .Y(new_n4078));
  NAND2xp33_ASAP7_75t_L     g03822(.A(new_n3862), .B(new_n4078), .Y(new_n4079));
  A2O1A1Ixp33_ASAP7_75t_L   g03823(.A1(new_n3854), .A2(new_n3855), .B(new_n3867), .C(new_n4079), .Y(new_n4080));
  NAND2xp33_ASAP7_75t_L     g03824(.A(new_n4080), .B(new_n4077), .Y(new_n4081));
  NOR2xp33_ASAP7_75t_L      g03825(.A(new_n3079), .B(new_n375), .Y(new_n4082));
  AOI221xp5_ASAP7_75t_L     g03826(.A1(\b[30] ), .A2(new_n361), .B1(new_n349), .B2(\b[29] ), .C(new_n4082), .Y(new_n4083));
  O2A1O1Ixp33_ASAP7_75t_L   g03827(.A1(new_n356), .A2(new_n3464), .B(new_n4083), .C(new_n346), .Y(new_n4084));
  O2A1O1Ixp33_ASAP7_75t_L   g03828(.A1(new_n356), .A2(new_n3464), .B(new_n4083), .C(\a[5] ), .Y(new_n4085));
  INVx1_ASAP7_75t_L         g03829(.A(new_n4085), .Y(new_n4086));
  OA21x2_ASAP7_75t_L        g03830(.A1(new_n346), .A2(new_n4084), .B(new_n4086), .Y(new_n4087));
  NAND3xp33_ASAP7_75t_L     g03831(.A(new_n4076), .B(new_n4081), .C(new_n4087), .Y(new_n4088));
  NOR2xp33_ASAP7_75t_L      g03832(.A(new_n4080), .B(new_n4077), .Y(new_n4089));
  AOI21xp33_ASAP7_75t_L     g03833(.A1(new_n4073), .A2(new_n4069), .B(new_n4075), .Y(new_n4090));
  OAI21xp33_ASAP7_75t_L     g03834(.A1(new_n346), .A2(new_n4084), .B(new_n4086), .Y(new_n4091));
  OAI21xp33_ASAP7_75t_L     g03835(.A1(new_n4090), .A2(new_n4089), .B(new_n4091), .Y(new_n4092));
  NAND3xp33_ASAP7_75t_L     g03836(.A(new_n3915), .B(new_n4088), .C(new_n4092), .Y(new_n4093));
  NAND3xp33_ASAP7_75t_L     g03837(.A(new_n4076), .B(new_n4081), .C(new_n4091), .Y(new_n4094));
  NOR3xp33_ASAP7_75t_L      g03838(.A(new_n4089), .B(new_n4090), .C(new_n4091), .Y(new_n4095));
  A2O1A1Ixp33_ASAP7_75t_L   g03839(.A1(new_n4091), .A2(new_n4094), .B(new_n4095), .C(new_n3887), .Y(new_n4096));
  NOR2xp33_ASAP7_75t_L      g03840(.A(new_n3674), .B(new_n287), .Y(new_n4097));
  AOI221xp5_ASAP7_75t_L     g03841(.A1(\b[32] ), .A2(new_n264), .B1(\b[33] ), .B2(new_n283), .C(new_n4097), .Y(new_n4098));
  INVx1_ASAP7_75t_L         g03842(.A(new_n3895), .Y(new_n4099));
  NOR2xp33_ASAP7_75t_L      g03843(.A(\b[32] ), .B(\b[33] ), .Y(new_n4100));
  INVx1_ASAP7_75t_L         g03844(.A(\b[33] ), .Y(new_n4101));
  NOR2xp33_ASAP7_75t_L      g03845(.A(new_n3891), .B(new_n4101), .Y(new_n4102));
  NOR2xp33_ASAP7_75t_L      g03846(.A(new_n4100), .B(new_n4102), .Y(new_n4103));
  A2O1A1Ixp33_ASAP7_75t_L   g03847(.A1(new_n4099), .A2(new_n3893), .B(new_n3892), .C(new_n4103), .Y(new_n4104));
  O2A1O1Ixp33_ASAP7_75t_L   g03848(.A1(new_n3675), .A2(new_n3678), .B(new_n3893), .C(new_n3892), .Y(new_n4105));
  INVx1_ASAP7_75t_L         g03849(.A(new_n4103), .Y(new_n4106));
  NAND2xp33_ASAP7_75t_L     g03850(.A(new_n4106), .B(new_n4105), .Y(new_n4107));
  NAND2xp33_ASAP7_75t_L     g03851(.A(new_n4107), .B(new_n4104), .Y(new_n4108));
  OAI21xp33_ASAP7_75t_L     g03852(.A1(new_n279), .A2(new_n4108), .B(new_n4098), .Y(new_n4109));
  NOR2xp33_ASAP7_75t_L      g03853(.A(new_n257), .B(new_n4109), .Y(new_n4110));
  O2A1O1Ixp33_ASAP7_75t_L   g03854(.A1(new_n279), .A2(new_n4108), .B(new_n4098), .C(\a[2] ), .Y(new_n4111));
  NOR2xp33_ASAP7_75t_L      g03855(.A(new_n4111), .B(new_n4110), .Y(new_n4112));
  AOI21xp33_ASAP7_75t_L     g03856(.A1(new_n4093), .A2(new_n4096), .B(new_n4112), .Y(new_n4113));
  INVx1_ASAP7_75t_L         g03857(.A(new_n4113), .Y(new_n4114));
  NAND3xp33_ASAP7_75t_L     g03858(.A(new_n4093), .B(new_n4096), .C(new_n4112), .Y(new_n4115));
  NAND2xp33_ASAP7_75t_L     g03859(.A(new_n4115), .B(new_n4114), .Y(new_n4116));
  O2A1O1Ixp33_ASAP7_75t_L   g03860(.A1(new_n3913), .A2(new_n3903), .B(new_n3914), .C(new_n4116), .Y(new_n4117));
  A2O1A1Ixp33_ASAP7_75t_L   g03861(.A1(new_n3909), .A2(new_n3908), .B(new_n3903), .C(new_n3914), .Y(new_n4118));
  AOI21xp33_ASAP7_75t_L     g03862(.A1(new_n4115), .A2(new_n4114), .B(new_n4118), .Y(new_n4119));
  NOR2xp33_ASAP7_75t_L      g03863(.A(new_n4117), .B(new_n4119), .Y(\f[33] ));
  O2A1O1Ixp33_ASAP7_75t_L   g03864(.A1(new_n3907), .A2(new_n3915), .B(new_n3908), .C(new_n3903), .Y(new_n4121));
  A2O1A1O1Ixp25_ASAP7_75t_L g03865(.A1(new_n3691), .A2(new_n3690), .B(new_n3685), .C(new_n3911), .D(new_n4121), .Y(new_n4122));
  NAND2xp33_ASAP7_75t_L     g03866(.A(new_n4026), .B(new_n4030), .Y(new_n4123));
  O2A1O1Ixp33_ASAP7_75t_L   g03867(.A1(new_n4040), .A2(new_n867), .B(new_n4041), .C(new_n4123), .Y(new_n4124));
  NAND3xp33_ASAP7_75t_L     g03868(.A(new_n3954), .B(new_n3955), .C(new_n3952), .Y(new_n4125));
  A2O1A1Ixp33_ASAP7_75t_L   g03869(.A1(new_n3959), .A2(new_n3960), .B(new_n3766), .C(new_n4125), .Y(new_n4126));
  NOR2xp33_ASAP7_75t_L      g03870(.A(new_n448), .B(new_n2930), .Y(new_n4127));
  AOI221xp5_ASAP7_75t_L     g03871(.A1(\b[5] ), .A2(new_n3129), .B1(\b[6] ), .B2(new_n2936), .C(new_n4127), .Y(new_n4128));
  NAND2xp33_ASAP7_75t_L     g03872(.A(new_n2932), .B(new_n1188), .Y(new_n4129));
  O2A1O1Ixp33_ASAP7_75t_L   g03873(.A1(new_n2940), .A2(new_n456), .B(new_n4128), .C(new_n2928), .Y(new_n4130));
  OAI211xp5_ASAP7_75t_L     g03874(.A1(new_n2940), .A2(new_n456), .B(\a[29] ), .C(new_n4128), .Y(new_n4131));
  A2O1A1Ixp33_ASAP7_75t_L   g03875(.A1(new_n4129), .A2(new_n4128), .B(new_n4130), .C(new_n4131), .Y(new_n4132));
  MAJIxp5_ASAP7_75t_L       g03876(.A(new_n3939), .B(new_n3730), .C(new_n3929), .Y(new_n4133));
  NAND2xp33_ASAP7_75t_L     g03877(.A(\b[3] ), .B(new_n3499), .Y(new_n4134));
  OAI221xp5_ASAP7_75t_L     g03878(.A1(new_n3510), .A2(new_n332), .B1(new_n289), .B2(new_n3703), .C(new_n4134), .Y(new_n4135));
  A2O1A1Ixp33_ASAP7_75t_L   g03879(.A1(new_n342), .A2(new_n3505), .B(new_n4135), .C(\a[32] ), .Y(new_n4136));
  AOI211xp5_ASAP7_75t_L     g03880(.A1(new_n342), .A2(new_n3505), .B(new_n3493), .C(new_n4135), .Y(new_n4137));
  A2O1A1O1Ixp25_ASAP7_75t_L g03881(.A1(new_n3505), .A2(new_n342), .B(new_n4135), .C(new_n4136), .D(new_n4137), .Y(new_n4138));
  INVx1_ASAP7_75t_L         g03882(.A(\a[34] ), .Y(new_n4139));
  NOR2xp33_ASAP7_75t_L      g03883(.A(\a[33] ), .B(new_n4139), .Y(new_n4140));
  NOR2xp33_ASAP7_75t_L      g03884(.A(\a[34] ), .B(new_n3923), .Y(new_n4141));
  OAI21xp33_ASAP7_75t_L     g03885(.A1(new_n4140), .A2(new_n4141), .B(new_n3926), .Y(new_n4142));
  NAND2xp33_ASAP7_75t_L     g03886(.A(new_n3925), .B(new_n3924), .Y(new_n4143));
  NAND2xp33_ASAP7_75t_L     g03887(.A(\a[35] ), .B(new_n4139), .Y(new_n4144));
  INVx1_ASAP7_75t_L         g03888(.A(\a[35] ), .Y(new_n4145));
  NAND2xp33_ASAP7_75t_L     g03889(.A(\a[34] ), .B(new_n4145), .Y(new_n4146));
  NAND3xp33_ASAP7_75t_L     g03890(.A(new_n4143), .B(new_n4144), .C(new_n4146), .Y(new_n4147));
  OAI22xp33_ASAP7_75t_L     g03891(.A1(new_n4142), .A2(new_n284), .B1(new_n262), .B2(new_n4147), .Y(new_n4148));
  NAND2xp33_ASAP7_75t_L     g03892(.A(new_n4146), .B(new_n4144), .Y(new_n4149));
  NAND2xp33_ASAP7_75t_L     g03893(.A(new_n4149), .B(new_n4143), .Y(new_n4150));
  INVx1_ASAP7_75t_L         g03894(.A(new_n4150), .Y(new_n4151));
  AOI21xp33_ASAP7_75t_L     g03895(.A1(new_n275), .A2(new_n4151), .B(new_n4148), .Y(new_n4152));
  NAND3xp33_ASAP7_75t_L     g03896(.A(new_n4152), .B(new_n3929), .C(\a[35] ), .Y(new_n4153));
  NOR2xp33_ASAP7_75t_L      g03897(.A(new_n4140), .B(new_n4141), .Y(new_n4154));
  NOR2xp33_ASAP7_75t_L      g03898(.A(new_n4143), .B(new_n4154), .Y(new_n4155));
  NOR2xp33_ASAP7_75t_L      g03899(.A(new_n4149), .B(new_n3926), .Y(new_n4156));
  AOI22xp33_ASAP7_75t_L     g03900(.A1(new_n4155), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n4156), .Y(new_n4157));
  O2A1O1Ixp33_ASAP7_75t_L   g03901(.A1(new_n4150), .A2(new_n274), .B(new_n4157), .C(new_n4145), .Y(new_n4158));
  A2O1A1Ixp33_ASAP7_75t_L   g03902(.A1(new_n4151), .A2(new_n275), .B(new_n4148), .C(new_n4145), .Y(new_n4159));
  A2O1A1Ixp33_ASAP7_75t_L   g03903(.A1(new_n4158), .A2(new_n3927), .B(new_n4145), .C(new_n4159), .Y(new_n4160));
  NAND2xp33_ASAP7_75t_L     g03904(.A(new_n4153), .B(new_n4160), .Y(new_n4161));
  NAND2xp33_ASAP7_75t_L     g03905(.A(new_n4138), .B(new_n4161), .Y(new_n4162));
  AOI21xp33_ASAP7_75t_L     g03906(.A1(new_n342), .A2(new_n3505), .B(new_n4135), .Y(new_n4163));
  NOR2xp33_ASAP7_75t_L      g03907(.A(\a[32] ), .B(new_n4163), .Y(new_n4164));
  OAI211xp5_ASAP7_75t_L     g03908(.A1(new_n4137), .A2(new_n4164), .B(new_n4153), .C(new_n4160), .Y(new_n4165));
  NAND3xp33_ASAP7_75t_L     g03909(.A(new_n4162), .B(new_n4133), .C(new_n4165), .Y(new_n4166));
  MAJIxp5_ASAP7_75t_L       g03910(.A(new_n3945), .B(new_n3927), .C(new_n3714), .Y(new_n4167));
  AOI211xp5_ASAP7_75t_L     g03911(.A1(new_n4160), .A2(new_n4153), .B(new_n4137), .C(new_n4164), .Y(new_n4168));
  NOR2xp33_ASAP7_75t_L      g03912(.A(new_n4138), .B(new_n4161), .Y(new_n4169));
  OAI21xp33_ASAP7_75t_L     g03913(.A1(new_n4168), .A2(new_n4169), .B(new_n4167), .Y(new_n4170));
  AO21x2_ASAP7_75t_L        g03914(.A1(new_n4166), .A2(new_n4170), .B(new_n4132), .Y(new_n4171));
  NAND3xp33_ASAP7_75t_L     g03915(.A(new_n4170), .B(new_n4166), .C(new_n4132), .Y(new_n4172));
  NAND3xp33_ASAP7_75t_L     g03916(.A(new_n4126), .B(new_n4171), .C(new_n4172), .Y(new_n4173));
  INVx1_ASAP7_75t_L         g03917(.A(new_n4125), .Y(new_n4174));
  NAND2xp33_ASAP7_75t_L     g03918(.A(new_n3959), .B(new_n3960), .Y(new_n4175));
  O2A1O1Ixp33_ASAP7_75t_L   g03919(.A1(new_n3750), .A2(new_n3726), .B(new_n4175), .C(new_n4174), .Y(new_n4176));
  AOI21xp33_ASAP7_75t_L     g03920(.A1(new_n4170), .A2(new_n4166), .B(new_n4132), .Y(new_n4177));
  AND3x1_ASAP7_75t_L        g03921(.A(new_n4170), .B(new_n4166), .C(new_n4132), .Y(new_n4178));
  OAI21xp33_ASAP7_75t_L     g03922(.A1(new_n4177), .A2(new_n4178), .B(new_n4176), .Y(new_n4179));
  NOR2xp33_ASAP7_75t_L      g03923(.A(new_n680), .B(new_n2415), .Y(new_n4180));
  AOI221xp5_ASAP7_75t_L     g03924(.A1(\b[8] ), .A2(new_n2577), .B1(\b[9] ), .B2(new_n2421), .C(new_n4180), .Y(new_n4181));
  OA21x2_ASAP7_75t_L        g03925(.A1(new_n2425), .A2(new_n1175), .B(new_n4181), .Y(new_n4182));
  O2A1O1Ixp33_ASAP7_75t_L   g03926(.A1(new_n2425), .A2(new_n1175), .B(new_n4181), .C(new_n2413), .Y(new_n4183));
  NAND2xp33_ASAP7_75t_L     g03927(.A(\a[26] ), .B(new_n4182), .Y(new_n4184));
  OA21x2_ASAP7_75t_L        g03928(.A1(new_n4182), .A2(new_n4183), .B(new_n4184), .Y(new_n4185));
  NAND3xp33_ASAP7_75t_L     g03929(.A(new_n4179), .B(new_n4173), .C(new_n4185), .Y(new_n4186));
  AO21x2_ASAP7_75t_L        g03930(.A1(new_n4173), .A2(new_n4179), .B(new_n4185), .Y(new_n4187));
  AOI22xp33_ASAP7_75t_L     g03931(.A1(new_n3972), .A2(new_n3966), .B1(new_n3970), .B2(new_n3969), .Y(new_n4188));
  A2O1A1O1Ixp25_ASAP7_75t_L g03932(.A1(new_n3747), .A2(new_n3746), .B(new_n3751), .C(new_n3973), .D(new_n4188), .Y(new_n4189));
  AND3x1_ASAP7_75t_L        g03933(.A(new_n4189), .B(new_n4187), .C(new_n4186), .Y(new_n4190));
  AOI21xp33_ASAP7_75t_L     g03934(.A1(new_n4187), .A2(new_n4186), .B(new_n4189), .Y(new_n4191));
  NOR2xp33_ASAP7_75t_L      g03935(.A(new_n833), .B(new_n1962), .Y(new_n4192));
  AOI221xp5_ASAP7_75t_L     g03936(.A1(new_n1955), .A2(\b[13] ), .B1(new_n2093), .B2(\b[11] ), .C(new_n4192), .Y(new_n4193));
  O2A1O1Ixp33_ASAP7_75t_L   g03937(.A1(new_n1956), .A2(new_n942), .B(new_n4193), .C(new_n1952), .Y(new_n4194));
  INVx1_ASAP7_75t_L         g03938(.A(new_n4194), .Y(new_n4195));
  O2A1O1Ixp33_ASAP7_75t_L   g03939(.A1(new_n1956), .A2(new_n942), .B(new_n4193), .C(\a[23] ), .Y(new_n4196));
  AOI21xp33_ASAP7_75t_L     g03940(.A1(new_n4195), .A2(\a[23] ), .B(new_n4196), .Y(new_n4197));
  OAI21xp33_ASAP7_75t_L     g03941(.A1(new_n4191), .A2(new_n4190), .B(new_n4197), .Y(new_n4198));
  A2O1A1O1Ixp25_ASAP7_75t_L g03942(.A1(new_n3700), .A2(new_n3775), .B(new_n3761), .C(new_n3991), .D(new_n3989), .Y(new_n4199));
  NAND3xp33_ASAP7_75t_L     g03943(.A(new_n4189), .B(new_n4187), .C(new_n4186), .Y(new_n4200));
  AO21x2_ASAP7_75t_L        g03944(.A1(new_n4186), .A2(new_n4187), .B(new_n4189), .Y(new_n4201));
  AO21x2_ASAP7_75t_L        g03945(.A1(\a[23] ), .A2(new_n4195), .B(new_n4196), .Y(new_n4202));
  NAND3xp33_ASAP7_75t_L     g03946(.A(new_n4202), .B(new_n4201), .C(new_n4200), .Y(new_n4203));
  AOI21xp33_ASAP7_75t_L     g03947(.A1(new_n4198), .A2(new_n4203), .B(new_n4199), .Y(new_n4204));
  A2O1A1Ixp33_ASAP7_75t_L   g03948(.A1(new_n3565), .A2(new_n3793), .B(new_n3770), .C(new_n3774), .Y(new_n4205));
  NOR3xp33_ASAP7_75t_L      g03949(.A(new_n4197), .B(new_n4190), .C(new_n4191), .Y(new_n4206));
  A2O1A1O1Ixp25_ASAP7_75t_L g03950(.A1(new_n3991), .A2(new_n4205), .B(new_n3989), .C(new_n4198), .D(new_n4206), .Y(new_n4207));
  NOR2xp33_ASAP7_75t_L      g03951(.A(new_n1043), .B(new_n1517), .Y(new_n4208));
  AOI221xp5_ASAP7_75t_L     g03952(.A1(\b[14] ), .A2(new_n1659), .B1(\b[16] ), .B2(new_n1511), .C(new_n4208), .Y(new_n4209));
  OAI311xp33_ASAP7_75t_L    g03953(.A1(new_n1155), .A2(new_n1521), .A3(new_n1154), .B1(\a[20] ), .C1(new_n4209), .Y(new_n4210));
  INVx1_ASAP7_75t_L         g03954(.A(new_n4209), .Y(new_n4211));
  A2O1A1Ixp33_ASAP7_75t_L   g03955(.A1(new_n1156), .A2(new_n1513), .B(new_n4211), .C(new_n1501), .Y(new_n4212));
  NAND2xp33_ASAP7_75t_L     g03956(.A(new_n4210), .B(new_n4212), .Y(new_n4213));
  INVx1_ASAP7_75t_L         g03957(.A(new_n4213), .Y(new_n4214));
  A2O1A1Ixp33_ASAP7_75t_L   g03958(.A1(new_n4207), .A2(new_n4198), .B(new_n4204), .C(new_n4214), .Y(new_n4215));
  AOI21xp33_ASAP7_75t_L     g03959(.A1(new_n4201), .A2(new_n4200), .B(new_n4202), .Y(new_n4216));
  A2O1A1Ixp33_ASAP7_75t_L   g03960(.A1(new_n3786), .A2(new_n3551), .B(new_n3785), .C(new_n3775), .Y(new_n4217));
  A2O1A1Ixp33_ASAP7_75t_L   g03961(.A1(new_n4217), .A2(new_n3774), .B(new_n3984), .C(new_n3992), .Y(new_n4218));
  OAI21xp33_ASAP7_75t_L     g03962(.A1(new_n4206), .A2(new_n4216), .B(new_n4218), .Y(new_n4219));
  OAI21xp33_ASAP7_75t_L     g03963(.A1(new_n4216), .A2(new_n4199), .B(new_n4203), .Y(new_n4220));
  OAI211xp5_ASAP7_75t_L     g03964(.A1(new_n4216), .A2(new_n4220), .B(new_n4213), .C(new_n4219), .Y(new_n4221));
  NOR2xp33_ASAP7_75t_L      g03965(.A(new_n3993), .B(new_n3990), .Y(new_n4222));
  MAJIxp5_ASAP7_75t_L       g03966(.A(new_n4018), .B(new_n4222), .C(new_n3999), .Y(new_n4223));
  NAND3xp33_ASAP7_75t_L     g03967(.A(new_n4223), .B(new_n4221), .C(new_n4215), .Y(new_n4224));
  A2O1A1Ixp33_ASAP7_75t_L   g03968(.A1(new_n4207), .A2(new_n4198), .B(new_n4204), .C(new_n4213), .Y(new_n4225));
  O2A1O1Ixp33_ASAP7_75t_L   g03969(.A1(new_n4216), .A2(new_n4220), .B(new_n4219), .C(new_n4213), .Y(new_n4226));
  NAND2xp33_ASAP7_75t_L     g03970(.A(new_n4002), .B(new_n4001), .Y(new_n4227));
  MAJIxp5_ASAP7_75t_L       g03971(.A(new_n3922), .B(new_n4227), .C(new_n4005), .Y(new_n4228));
  A2O1A1Ixp33_ASAP7_75t_L   g03972(.A1(new_n4225), .A2(new_n4213), .B(new_n4226), .C(new_n4228), .Y(new_n4229));
  NOR2xp33_ASAP7_75t_L      g03973(.A(new_n1458), .B(new_n2118), .Y(new_n4230));
  AOI221xp5_ASAP7_75t_L     g03974(.A1(\b[17] ), .A2(new_n1290), .B1(\b[19] ), .B2(new_n1209), .C(new_n4230), .Y(new_n4231));
  INVx1_ASAP7_75t_L         g03975(.A(new_n4231), .Y(new_n4232));
  A2O1A1Ixp33_ASAP7_75t_L   g03976(.A1(new_n1607), .A2(new_n1216), .B(new_n4232), .C(\a[17] ), .Y(new_n4233));
  O2A1O1Ixp33_ASAP7_75t_L   g03977(.A1(new_n1210), .A2(new_n1628), .B(new_n4231), .C(\a[17] ), .Y(new_n4234));
  AOI21xp33_ASAP7_75t_L     g03978(.A1(new_n4233), .A2(\a[17] ), .B(new_n4234), .Y(new_n4235));
  NAND3xp33_ASAP7_75t_L     g03979(.A(new_n4224), .B(new_n4229), .C(new_n4235), .Y(new_n4236));
  NAND2xp33_ASAP7_75t_L     g03980(.A(new_n4221), .B(new_n4215), .Y(new_n4237));
  NOR2xp33_ASAP7_75t_L      g03981(.A(new_n4228), .B(new_n4237), .Y(new_n4238));
  O2A1O1Ixp33_ASAP7_75t_L   g03982(.A1(new_n4216), .A2(new_n4220), .B(new_n4219), .C(new_n4214), .Y(new_n4239));
  O2A1O1Ixp33_ASAP7_75t_L   g03983(.A1(new_n4214), .A2(new_n4239), .B(new_n4215), .C(new_n4223), .Y(new_n4240));
  OAI211xp5_ASAP7_75t_L     g03984(.A1(new_n1210), .A2(new_n1628), .B(\a[17] ), .C(new_n4231), .Y(new_n4241));
  A2O1A1Ixp33_ASAP7_75t_L   g03985(.A1(new_n1607), .A2(new_n1216), .B(new_n4232), .C(new_n1206), .Y(new_n4242));
  NAND2xp33_ASAP7_75t_L     g03986(.A(new_n4241), .B(new_n4242), .Y(new_n4243));
  OAI21xp33_ASAP7_75t_L     g03987(.A1(new_n4240), .A2(new_n4238), .B(new_n4243), .Y(new_n4244));
  NAND2xp33_ASAP7_75t_L     g03988(.A(new_n4236), .B(new_n4244), .Y(new_n4245));
  A2O1A1Ixp33_ASAP7_75t_L   g03989(.A1(new_n3842), .A2(new_n3921), .B(new_n4028), .C(new_n4017), .Y(new_n4246));
  NOR2xp33_ASAP7_75t_L      g03990(.A(new_n4245), .B(new_n4246), .Y(new_n4247));
  NAND2xp33_ASAP7_75t_L     g03991(.A(new_n4229), .B(new_n4224), .Y(new_n4248));
  NAND3xp33_ASAP7_75t_L     g03992(.A(new_n4224), .B(new_n4229), .C(new_n4243), .Y(new_n4249));
  INVx1_ASAP7_75t_L         g03993(.A(new_n4249), .Y(new_n4250));
  A2O1A1O1Ixp25_ASAP7_75t_L g03994(.A1(new_n3809), .A2(new_n3810), .B(new_n3920), .C(new_n4024), .D(new_n4027), .Y(new_n4251));
  O2A1O1Ixp33_ASAP7_75t_L   g03995(.A1(new_n4248), .A2(new_n4250), .B(new_n4244), .C(new_n4251), .Y(new_n4252));
  NOR2xp33_ASAP7_75t_L      g03996(.A(new_n1895), .B(new_n864), .Y(new_n4253));
  AOI221xp5_ASAP7_75t_L     g03997(.A1(\b[20] ), .A2(new_n985), .B1(\b[22] ), .B2(new_n886), .C(new_n4253), .Y(new_n4254));
  O2A1O1Ixp33_ASAP7_75t_L   g03998(.A1(new_n872), .A2(new_n2522), .B(new_n4254), .C(new_n867), .Y(new_n4255));
  O2A1O1Ixp33_ASAP7_75t_L   g03999(.A1(new_n872), .A2(new_n2522), .B(new_n4254), .C(\a[14] ), .Y(new_n4256));
  INVx1_ASAP7_75t_L         g04000(.A(new_n4256), .Y(new_n4257));
  OAI21xp33_ASAP7_75t_L     g04001(.A1(new_n867), .A2(new_n4255), .B(new_n4257), .Y(new_n4258));
  NOR3xp33_ASAP7_75t_L      g04002(.A(new_n4247), .B(new_n4252), .C(new_n4258), .Y(new_n4259));
  NOR2xp33_ASAP7_75t_L      g04003(.A(new_n4240), .B(new_n4238), .Y(new_n4260));
  AOI21xp33_ASAP7_75t_L     g04004(.A1(new_n4224), .A2(new_n4229), .B(new_n4235), .Y(new_n4261));
  AOI21xp33_ASAP7_75t_L     g04005(.A1(new_n4249), .A2(new_n4260), .B(new_n4261), .Y(new_n4262));
  NAND2xp33_ASAP7_75t_L     g04006(.A(new_n4251), .B(new_n4262), .Y(new_n4263));
  OAI21xp33_ASAP7_75t_L     g04007(.A1(new_n4027), .A2(new_n4039), .B(new_n4245), .Y(new_n4264));
  INVx1_ASAP7_75t_L         g04008(.A(new_n4254), .Y(new_n4265));
  A2O1A1Ixp33_ASAP7_75t_L   g04009(.A1(new_n2056), .A2(new_n873), .B(new_n4265), .C(\a[14] ), .Y(new_n4266));
  AOI21xp33_ASAP7_75t_L     g04010(.A1(new_n4266), .A2(\a[14] ), .B(new_n4256), .Y(new_n4267));
  AOI21xp33_ASAP7_75t_L     g04011(.A1(new_n4263), .A2(new_n4264), .B(new_n4267), .Y(new_n4268));
  A2O1A1Ixp33_ASAP7_75t_L   g04012(.A1(new_n3614), .A2(new_n3613), .B(new_n3828), .C(new_n3821), .Y(new_n4269));
  AOI22xp33_ASAP7_75t_L     g04013(.A1(new_n4037), .A2(new_n4043), .B1(new_n3825), .B2(new_n4269), .Y(new_n4270));
  NOR4xp25_ASAP7_75t_L      g04014(.A(new_n4270), .B(new_n4124), .C(new_n4259), .D(new_n4268), .Y(new_n4271));
  INVx1_ASAP7_75t_L         g04015(.A(new_n4124), .Y(new_n4272));
  NAND3xp33_ASAP7_75t_L     g04016(.A(new_n4263), .B(new_n4264), .C(new_n4267), .Y(new_n4273));
  OAI21xp33_ASAP7_75t_L     g04017(.A1(new_n4252), .A2(new_n4247), .B(new_n4258), .Y(new_n4274));
  OAI21xp33_ASAP7_75t_L     g04018(.A1(new_n3824), .A2(new_n3845), .B(new_n4045), .Y(new_n4275));
  AOI22xp33_ASAP7_75t_L     g04019(.A1(new_n4274), .A2(new_n4273), .B1(new_n4272), .B2(new_n4275), .Y(new_n4276));
  NOR2xp33_ASAP7_75t_L      g04020(.A(new_n2205), .B(new_n1550), .Y(new_n4277));
  AOI221xp5_ASAP7_75t_L     g04021(.A1(\b[23] ), .A2(new_n713), .B1(\b[25] ), .B2(new_n640), .C(new_n4277), .Y(new_n4278));
  O2A1O1Ixp33_ASAP7_75t_L   g04022(.A1(new_n641), .A2(new_n2385), .B(new_n4278), .C(new_n637), .Y(new_n4279));
  INVx1_ASAP7_75t_L         g04023(.A(new_n4279), .Y(new_n4280));
  O2A1O1Ixp33_ASAP7_75t_L   g04024(.A1(new_n641), .A2(new_n2385), .B(new_n4278), .C(\a[11] ), .Y(new_n4281));
  AOI21xp33_ASAP7_75t_L     g04025(.A1(new_n4280), .A2(\a[11] ), .B(new_n4281), .Y(new_n4282));
  OAI21xp33_ASAP7_75t_L     g04026(.A1(new_n4271), .A2(new_n4276), .B(new_n4282), .Y(new_n4283));
  INVx1_ASAP7_75t_L         g04027(.A(new_n4057), .Y(new_n4284));
  AOI21xp33_ASAP7_75t_L     g04028(.A1(new_n3918), .A2(new_n4053), .B(new_n4284), .Y(new_n4285));
  NAND4xp25_ASAP7_75t_L     g04029(.A(new_n4275), .B(new_n4272), .C(new_n4273), .D(new_n4274), .Y(new_n4286));
  NAND2xp33_ASAP7_75t_L     g04030(.A(new_n4273), .B(new_n4274), .Y(new_n4287));
  MAJIxp5_ASAP7_75t_L       g04031(.A(new_n3829), .B(new_n4123), .C(new_n4036), .Y(new_n4288));
  NAND2xp33_ASAP7_75t_L     g04032(.A(new_n4288), .B(new_n4287), .Y(new_n4289));
  AO21x2_ASAP7_75t_L        g04033(.A1(\a[11] ), .A2(new_n4280), .B(new_n4281), .Y(new_n4290));
  NAND3xp33_ASAP7_75t_L     g04034(.A(new_n4289), .B(new_n4286), .C(new_n4290), .Y(new_n4291));
  AOI21xp33_ASAP7_75t_L     g04035(.A1(new_n4283), .A2(new_n4291), .B(new_n4285), .Y(new_n4292));
  NOR3xp33_ASAP7_75t_L      g04036(.A(new_n4276), .B(new_n4271), .C(new_n4282), .Y(new_n4293));
  A2O1A1O1Ixp25_ASAP7_75t_L g04037(.A1(new_n4053), .A2(new_n3918), .B(new_n4284), .C(new_n4283), .D(new_n4293), .Y(new_n4294));
  NOR2xp33_ASAP7_75t_L      g04038(.A(new_n2879), .B(new_n513), .Y(new_n4295));
  AOI221xp5_ASAP7_75t_L     g04039(.A1(\b[26] ), .A2(new_n560), .B1(\b[28] ), .B2(new_n475), .C(new_n4295), .Y(new_n4296));
  INVx1_ASAP7_75t_L         g04040(.A(new_n4296), .Y(new_n4297));
  A2O1A1Ixp33_ASAP7_75t_L   g04041(.A1(new_n3085), .A2(new_n483), .B(new_n4297), .C(\a[8] ), .Y(new_n4298));
  O2A1O1Ixp33_ASAP7_75t_L   g04042(.A1(new_n477), .A2(new_n3087), .B(new_n4296), .C(\a[8] ), .Y(new_n4299));
  AOI21xp33_ASAP7_75t_L     g04043(.A1(new_n4298), .A2(\a[8] ), .B(new_n4299), .Y(new_n4300));
  A2O1A1Ixp33_ASAP7_75t_L   g04044(.A1(new_n4294), .A2(new_n4283), .B(new_n4292), .C(new_n4300), .Y(new_n4301));
  INVx1_ASAP7_75t_L         g04045(.A(new_n4053), .Y(new_n4302));
  OAI21xp33_ASAP7_75t_L     g04046(.A1(new_n4302), .A2(new_n4060), .B(new_n4057), .Y(new_n4303));
  AOI21xp33_ASAP7_75t_L     g04047(.A1(new_n4289), .A2(new_n4286), .B(new_n4290), .Y(new_n4304));
  OAI21xp33_ASAP7_75t_L     g04048(.A1(new_n4293), .A2(new_n4304), .B(new_n4303), .Y(new_n4305));
  NAND3xp33_ASAP7_75t_L     g04049(.A(new_n4285), .B(new_n4291), .C(new_n4283), .Y(new_n4306));
  INVx1_ASAP7_75t_L         g04050(.A(new_n4300), .Y(new_n4307));
  NAND3xp33_ASAP7_75t_L     g04051(.A(new_n4307), .B(new_n4306), .C(new_n4305), .Y(new_n4308));
  NAND2xp33_ASAP7_75t_L     g04052(.A(new_n4308), .B(new_n4301), .Y(new_n4309));
  NAND2xp33_ASAP7_75t_L     g04053(.A(new_n4058), .B(new_n4062), .Y(new_n4310));
  MAJIxp5_ASAP7_75t_L       g04054(.A(new_n4075), .B(new_n4310), .C(new_n4068), .Y(new_n4311));
  NOR2xp33_ASAP7_75t_L      g04055(.A(new_n4309), .B(new_n4311), .Y(new_n4312));
  AOI21xp33_ASAP7_75t_L     g04056(.A1(new_n4306), .A2(new_n4305), .B(new_n4307), .Y(new_n4313));
  AOI211xp5_ASAP7_75t_L     g04057(.A1(new_n4294), .A2(new_n4283), .B(new_n4300), .C(new_n4292), .Y(new_n4314));
  NOR2xp33_ASAP7_75t_L      g04058(.A(new_n4313), .B(new_n4314), .Y(new_n4315));
  O2A1O1Ixp33_ASAP7_75t_L   g04059(.A1(new_n4310), .A2(new_n4068), .B(new_n4081), .C(new_n4315), .Y(new_n4316));
  INVx1_ASAP7_75t_L         g04060(.A(new_n3681), .Y(new_n4317));
  NAND2xp33_ASAP7_75t_L     g04061(.A(\b[31] ), .B(new_n361), .Y(new_n4318));
  OAI221xp5_ASAP7_75t_L     g04062(.A1(new_n350), .A2(new_n3456), .B1(new_n3098), .B2(new_n375), .C(new_n4318), .Y(new_n4319));
  A2O1A1Ixp33_ASAP7_75t_L   g04063(.A1(new_n4317), .A2(new_n359), .B(new_n4319), .C(\a[5] ), .Y(new_n4320));
  AOI211xp5_ASAP7_75t_L     g04064(.A1(new_n4317), .A2(new_n359), .B(new_n4319), .C(new_n346), .Y(new_n4321));
  A2O1A1O1Ixp25_ASAP7_75t_L g04065(.A1(new_n4317), .A2(new_n359), .B(new_n4319), .C(new_n4320), .D(new_n4321), .Y(new_n4322));
  OAI21xp33_ASAP7_75t_L     g04066(.A1(new_n4312), .A2(new_n4316), .B(new_n4322), .Y(new_n4323));
  O2A1O1Ixp33_ASAP7_75t_L   g04067(.A1(new_n3658), .A2(new_n3662), .B(new_n3879), .C(new_n3907), .Y(new_n4324));
  INVx1_ASAP7_75t_L         g04068(.A(new_n4094), .Y(new_n4325));
  NAND2xp33_ASAP7_75t_L     g04069(.A(new_n4088), .B(new_n4092), .Y(new_n4326));
  O2A1O1Ixp33_ASAP7_75t_L   g04070(.A1(new_n4324), .A2(new_n3886), .B(new_n4326), .C(new_n4325), .Y(new_n4327));
  INVx1_ASAP7_75t_L         g04071(.A(new_n4067), .Y(new_n4328));
  O2A1O1Ixp33_ASAP7_75t_L   g04072(.A1(new_n4065), .A2(new_n466), .B(new_n4328), .C(new_n4310), .Y(new_n4329));
  AOI21xp33_ASAP7_75t_L     g04073(.A1(new_n4077), .A2(new_n4080), .B(new_n4329), .Y(new_n4330));
  NAND2xp33_ASAP7_75t_L     g04074(.A(new_n4315), .B(new_n4330), .Y(new_n4331));
  A2O1A1Ixp33_ASAP7_75t_L   g04075(.A1(new_n4077), .A2(new_n4080), .B(new_n4329), .C(new_n4309), .Y(new_n4332));
  INVx1_ASAP7_75t_L         g04076(.A(new_n4321), .Y(new_n4333));
  A2O1A1Ixp33_ASAP7_75t_L   g04077(.A1(new_n4317), .A2(new_n359), .B(new_n4319), .C(new_n346), .Y(new_n4334));
  NAND2xp33_ASAP7_75t_L     g04078(.A(new_n4334), .B(new_n4333), .Y(new_n4335));
  NAND3xp33_ASAP7_75t_L     g04079(.A(new_n4335), .B(new_n4332), .C(new_n4331), .Y(new_n4336));
  AOI21xp33_ASAP7_75t_L     g04080(.A1(new_n4323), .A2(new_n4336), .B(new_n4327), .Y(new_n4337));
  NOR3xp33_ASAP7_75t_L      g04081(.A(new_n4316), .B(new_n4322), .C(new_n4312), .Y(new_n4338));
  A2O1A1O1Ixp25_ASAP7_75t_L g04082(.A1(new_n4326), .A2(new_n3915), .B(new_n4325), .C(new_n4323), .D(new_n4338), .Y(new_n4339));
  NOR2xp33_ASAP7_75t_L      g04083(.A(new_n3891), .B(new_n287), .Y(new_n4340));
  AOI221xp5_ASAP7_75t_L     g04084(.A1(\b[33] ), .A2(new_n264), .B1(\b[34] ), .B2(new_n283), .C(new_n4340), .Y(new_n4341));
  INVx1_ASAP7_75t_L         g04085(.A(new_n4102), .Y(new_n4342));
  NOR2xp33_ASAP7_75t_L      g04086(.A(\b[33] ), .B(\b[34] ), .Y(new_n4343));
  INVx1_ASAP7_75t_L         g04087(.A(\b[34] ), .Y(new_n4344));
  NOR2xp33_ASAP7_75t_L      g04088(.A(new_n4101), .B(new_n4344), .Y(new_n4345));
  NOR2xp33_ASAP7_75t_L      g04089(.A(new_n4343), .B(new_n4345), .Y(new_n4346));
  INVx1_ASAP7_75t_L         g04090(.A(new_n4346), .Y(new_n4347));
  O2A1O1Ixp33_ASAP7_75t_L   g04091(.A1(new_n4106), .A2(new_n4105), .B(new_n4342), .C(new_n4347), .Y(new_n4348));
  INVx1_ASAP7_75t_L         g04092(.A(new_n4348), .Y(new_n4349));
  A2O1A1O1Ixp25_ASAP7_75t_L g04093(.A1(new_n3893), .A2(new_n4099), .B(new_n3892), .C(new_n4103), .D(new_n4102), .Y(new_n4350));
  NAND2xp33_ASAP7_75t_L     g04094(.A(new_n4347), .B(new_n4350), .Y(new_n4351));
  NAND2xp33_ASAP7_75t_L     g04095(.A(new_n4349), .B(new_n4351), .Y(new_n4352));
  O2A1O1Ixp33_ASAP7_75t_L   g04096(.A1(new_n279), .A2(new_n4352), .B(new_n4341), .C(new_n257), .Y(new_n4353));
  OAI21xp33_ASAP7_75t_L     g04097(.A1(new_n279), .A2(new_n4352), .B(new_n4341), .Y(new_n4354));
  NAND2xp33_ASAP7_75t_L     g04098(.A(new_n257), .B(new_n4354), .Y(new_n4355));
  OA21x2_ASAP7_75t_L        g04099(.A1(new_n257), .A2(new_n4353), .B(new_n4355), .Y(new_n4356));
  A2O1A1Ixp33_ASAP7_75t_L   g04100(.A1(new_n4339), .A2(new_n4323), .B(new_n4337), .C(new_n4356), .Y(new_n4357));
  AOI21xp33_ASAP7_75t_L     g04101(.A1(new_n4323), .A2(new_n4339), .B(new_n4337), .Y(new_n4358));
  INVx1_ASAP7_75t_L         g04102(.A(new_n4356), .Y(new_n4359));
  NAND2xp33_ASAP7_75t_L     g04103(.A(new_n4359), .B(new_n4358), .Y(new_n4360));
  AND2x2_ASAP7_75t_L        g04104(.A(new_n4357), .B(new_n4360), .Y(new_n4361));
  O2A1O1Ixp33_ASAP7_75t_L   g04105(.A1(new_n4122), .A2(new_n4116), .B(new_n4114), .C(new_n4361), .Y(new_n4362));
  A2O1A1O1Ixp25_ASAP7_75t_L g04106(.A1(new_n3911), .A2(new_n3695), .B(new_n4121), .C(new_n4115), .D(new_n4113), .Y(new_n4363));
  AND2x2_ASAP7_75t_L        g04107(.A(new_n4363), .B(new_n4361), .Y(new_n4364));
  NOR2xp33_ASAP7_75t_L      g04108(.A(new_n4362), .B(new_n4364), .Y(\f[34] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04109(.A1(new_n4339), .A2(new_n4323), .B(new_n4337), .C(new_n4359), .Y(new_n4366));
  O2A1O1Ixp33_ASAP7_75t_L   g04110(.A1(new_n4302), .A2(new_n4060), .B(new_n4057), .C(new_n4304), .Y(new_n4367));
  A2O1A1O1Ixp25_ASAP7_75t_L g04111(.A1(new_n4291), .A2(new_n4367), .B(new_n4285), .C(new_n4306), .D(new_n4300), .Y(new_n4368));
  NOR2xp33_ASAP7_75t_L      g04112(.A(new_n2703), .B(new_n710), .Y(new_n4369));
  AOI221xp5_ASAP7_75t_L     g04113(.A1(\b[25] ), .A2(new_n635), .B1(\b[24] ), .B2(new_n713), .C(new_n4369), .Y(new_n4370));
  O2A1O1Ixp33_ASAP7_75t_L   g04114(.A1(new_n641), .A2(new_n2708), .B(new_n4370), .C(new_n637), .Y(new_n4371));
  OAI21xp33_ASAP7_75t_L     g04115(.A1(new_n641), .A2(new_n2708), .B(new_n4370), .Y(new_n4372));
  NAND2xp33_ASAP7_75t_L     g04116(.A(new_n637), .B(new_n4372), .Y(new_n4373));
  OAI21xp33_ASAP7_75t_L     g04117(.A1(new_n637), .A2(new_n4371), .B(new_n4373), .Y(new_n4374));
  INVx1_ASAP7_75t_L         g04118(.A(new_n4374), .Y(new_n4375));
  NOR2xp33_ASAP7_75t_L      g04119(.A(new_n4252), .B(new_n4247), .Y(new_n4376));
  MAJIxp5_ASAP7_75t_L       g04120(.A(new_n4288), .B(new_n4376), .C(new_n4258), .Y(new_n4377));
  A2O1A1Ixp33_ASAP7_75t_L   g04121(.A1(new_n4248), .A2(new_n4244), .B(new_n4251), .C(new_n4249), .Y(new_n4378));
  NAND2xp33_ASAP7_75t_L     g04122(.A(new_n2417), .B(new_n690), .Y(new_n4379));
  A2O1A1Ixp33_ASAP7_75t_L   g04123(.A1(new_n4379), .A2(new_n4181), .B(new_n4183), .C(new_n4184), .Y(new_n4380));
  NAND3xp33_ASAP7_75t_L     g04124(.A(new_n4179), .B(new_n4173), .C(new_n4380), .Y(new_n4381));
  A2O1A1Ixp33_ASAP7_75t_L   g04125(.A1(new_n4185), .A2(new_n4186), .B(new_n4189), .C(new_n4381), .Y(new_n4382));
  NOR2xp33_ASAP7_75t_L      g04126(.A(new_n680), .B(new_n2410), .Y(new_n4383));
  AOI221xp5_ASAP7_75t_L     g04127(.A1(\b[9] ), .A2(new_n2577), .B1(\b[11] ), .B2(new_n2423), .C(new_n4383), .Y(new_n4384));
  O2A1O1Ixp33_ASAP7_75t_L   g04128(.A1(new_n2425), .A2(new_n754), .B(new_n4384), .C(new_n2413), .Y(new_n4385));
  INVx1_ASAP7_75t_L         g04129(.A(new_n4385), .Y(new_n4386));
  O2A1O1Ixp33_ASAP7_75t_L   g04130(.A1(new_n2425), .A2(new_n754), .B(new_n4384), .C(\a[26] ), .Y(new_n4387));
  AOI21xp33_ASAP7_75t_L     g04131(.A1(new_n4386), .A2(\a[26] ), .B(new_n4387), .Y(new_n4388));
  OAI22xp33_ASAP7_75t_L     g04132(.A1(new_n3750), .A2(new_n3726), .B1(new_n3957), .B2(new_n3953), .Y(new_n4389));
  A2O1A1Ixp33_ASAP7_75t_L   g04133(.A1(new_n4389), .A2(new_n4125), .B(new_n4177), .C(new_n4172), .Y(new_n4390));
  NOR2xp33_ASAP7_75t_L      g04134(.A(new_n534), .B(new_n2930), .Y(new_n4391));
  AOI221xp5_ASAP7_75t_L     g04135(.A1(\b[6] ), .A2(new_n3129), .B1(\b[7] ), .B2(new_n2936), .C(new_n4391), .Y(new_n4392));
  O2A1O1Ixp33_ASAP7_75t_L   g04136(.A1(new_n2940), .A2(new_n540), .B(new_n4392), .C(new_n2928), .Y(new_n4393));
  OAI21xp33_ASAP7_75t_L     g04137(.A1(new_n2940), .A2(new_n540), .B(new_n4392), .Y(new_n4394));
  NAND2xp33_ASAP7_75t_L     g04138(.A(new_n2928), .B(new_n4394), .Y(new_n4395));
  OAI21xp33_ASAP7_75t_L     g04139(.A1(new_n2928), .A2(new_n4393), .B(new_n4395), .Y(new_n4396));
  NAND3xp33_ASAP7_75t_L     g04140(.A(new_n3926), .B(new_n4154), .C(new_n4149), .Y(new_n4397));
  NAND2xp33_ASAP7_75t_L     g04141(.A(\b[1] ), .B(new_n4155), .Y(new_n4398));
  OAI221xp5_ASAP7_75t_L     g04142(.A1(new_n4147), .A2(new_n289), .B1(new_n284), .B2(new_n4397), .C(new_n4398), .Y(new_n4399));
  A2O1A1Ixp33_ASAP7_75t_L   g04143(.A1(new_n294), .A2(new_n4151), .B(new_n4399), .C(\a[35] ), .Y(new_n4400));
  NOR2xp33_ASAP7_75t_L      g04144(.A(new_n289), .B(new_n4147), .Y(new_n4401));
  AND3x1_ASAP7_75t_L        g04145(.A(new_n3926), .B(new_n4149), .C(new_n4154), .Y(new_n4402));
  AOI221xp5_ASAP7_75t_L     g04146(.A1(new_n4155), .A2(\b[1] ), .B1(new_n4402), .B2(\b[0] ), .C(new_n4401), .Y(new_n4403));
  O2A1O1Ixp33_ASAP7_75t_L   g04147(.A1(new_n509), .A2(new_n4150), .B(new_n4403), .C(\a[35] ), .Y(new_n4404));
  A2O1A1O1Ixp25_ASAP7_75t_L g04148(.A1(new_n4152), .A2(new_n3929), .B(new_n4400), .C(\a[35] ), .D(new_n4404), .Y(new_n4405));
  OAI21xp33_ASAP7_75t_L     g04149(.A1(new_n4150), .A2(new_n274), .B(new_n4157), .Y(new_n4406));
  NOR2xp33_ASAP7_75t_L      g04150(.A(new_n4150), .B(new_n509), .Y(new_n4407));
  NOR5xp2_ASAP7_75t_L       g04151(.A(new_n4406), .B(new_n4399), .C(new_n4407), .D(new_n3927), .E(new_n4145), .Y(new_n4408));
  NAND2xp33_ASAP7_75t_L     g04152(.A(\b[4] ), .B(new_n3499), .Y(new_n4409));
  OAI221xp5_ASAP7_75t_L     g04153(.A1(new_n3510), .A2(new_n384), .B1(new_n301), .B2(new_n3703), .C(new_n4409), .Y(new_n4410));
  A2O1A1Ixp33_ASAP7_75t_L   g04154(.A1(new_n394), .A2(new_n3505), .B(new_n4410), .C(\a[32] ), .Y(new_n4411));
  NOR2xp33_ASAP7_75t_L      g04155(.A(new_n384), .B(new_n3510), .Y(new_n4412));
  AOI221xp5_ASAP7_75t_L     g04156(.A1(\b[3] ), .A2(new_n3708), .B1(\b[4] ), .B2(new_n3499), .C(new_n4412), .Y(new_n4413));
  O2A1O1Ixp33_ASAP7_75t_L   g04157(.A1(new_n3513), .A2(new_n728), .B(new_n4413), .C(\a[32] ), .Y(new_n4414));
  AOI21xp33_ASAP7_75t_L     g04158(.A1(new_n4411), .A2(\a[32] ), .B(new_n4414), .Y(new_n4415));
  OAI21xp33_ASAP7_75t_L     g04159(.A1(new_n4408), .A2(new_n4405), .B(new_n4415), .Y(new_n4416));
  AOI21xp33_ASAP7_75t_L     g04160(.A1(new_n4162), .A2(new_n4133), .B(new_n4169), .Y(new_n4417));
  NOR2xp33_ASAP7_75t_L      g04161(.A(new_n4408), .B(new_n4405), .Y(new_n4418));
  A2O1A1Ixp33_ASAP7_75t_L   g04162(.A1(\a[32] ), .A2(new_n4411), .B(new_n4414), .C(new_n4418), .Y(new_n4419));
  AOI21xp33_ASAP7_75t_L     g04163(.A1(new_n4416), .A2(new_n4419), .B(new_n4417), .Y(new_n4420));
  NOR3xp33_ASAP7_75t_L      g04164(.A(new_n4415), .B(new_n4405), .C(new_n4408), .Y(new_n4421));
  A2O1A1O1Ixp25_ASAP7_75t_L g04165(.A1(new_n4133), .A2(new_n4162), .B(new_n4169), .C(new_n4416), .D(new_n4421), .Y(new_n4422));
  A2O1A1Ixp33_ASAP7_75t_L   g04166(.A1(new_n4422), .A2(new_n4416), .B(new_n4420), .C(new_n4396), .Y(new_n4423));
  INVx1_ASAP7_75t_L         g04167(.A(new_n4407), .Y(new_n4424));
  NAND3xp33_ASAP7_75t_L     g04168(.A(new_n4403), .B(\a[35] ), .C(new_n4424), .Y(new_n4425));
  A2O1A1Ixp33_ASAP7_75t_L   g04169(.A1(new_n294), .A2(new_n4151), .B(new_n4399), .C(new_n4145), .Y(new_n4426));
  NAND3xp33_ASAP7_75t_L     g04170(.A(new_n4153), .B(new_n4425), .C(new_n4426), .Y(new_n4427));
  NAND5xp2_ASAP7_75t_L      g04171(.A(\a[35] ), .B(new_n4152), .C(new_n4403), .D(new_n4424), .E(new_n3929), .Y(new_n4428));
  AOI221xp5_ASAP7_75t_L     g04172(.A1(new_n4411), .A2(\a[32] ), .B1(new_n4428), .B2(new_n4427), .C(new_n4414), .Y(new_n4429));
  OAI21xp33_ASAP7_75t_L     g04173(.A1(new_n4168), .A2(new_n4167), .B(new_n4165), .Y(new_n4430));
  OAI21xp33_ASAP7_75t_L     g04174(.A1(new_n4421), .A2(new_n4429), .B(new_n4430), .Y(new_n4431));
  INVx1_ASAP7_75t_L         g04175(.A(new_n4422), .Y(new_n4432));
  O2A1O1Ixp33_ASAP7_75t_L   g04176(.A1(new_n4429), .A2(new_n4432), .B(new_n4431), .C(new_n4396), .Y(new_n4433));
  A2O1A1Ixp33_ASAP7_75t_L   g04177(.A1(new_n4396), .A2(new_n4423), .B(new_n4433), .C(new_n4390), .Y(new_n4434));
  A2O1A1Ixp33_ASAP7_75t_L   g04178(.A1(new_n3525), .A2(new_n3702), .B(new_n3731), .C(new_n3721), .Y(new_n4435));
  A2O1A1O1Ixp25_ASAP7_75t_L g04179(.A1(new_n4175), .A2(new_n4435), .B(new_n4174), .C(new_n4171), .D(new_n4178), .Y(new_n4436));
  NOR3xp33_ASAP7_75t_L      g04180(.A(new_n4430), .B(new_n4421), .C(new_n4429), .Y(new_n4437));
  OA21x2_ASAP7_75t_L        g04181(.A1(new_n2928), .A2(new_n4393), .B(new_n4395), .Y(new_n4438));
  OAI21xp33_ASAP7_75t_L     g04182(.A1(new_n4437), .A2(new_n4420), .B(new_n4438), .Y(new_n4439));
  O2A1O1Ixp33_ASAP7_75t_L   g04183(.A1(new_n4167), .A2(new_n4168), .B(new_n4165), .C(new_n4429), .Y(new_n4440));
  OAI311xp33_ASAP7_75t_L    g04184(.A1(new_n4440), .A2(new_n4429), .A3(new_n4421), .B1(new_n4396), .C1(new_n4431), .Y(new_n4441));
  NAND3xp33_ASAP7_75t_L     g04185(.A(new_n4436), .B(new_n4439), .C(new_n4441), .Y(new_n4442));
  AOI21xp33_ASAP7_75t_L     g04186(.A1(new_n4434), .A2(new_n4442), .B(new_n4388), .Y(new_n4443));
  INVx1_ASAP7_75t_L         g04187(.A(new_n4387), .Y(new_n4444));
  OAI21xp33_ASAP7_75t_L     g04188(.A1(new_n2413), .A2(new_n4385), .B(new_n4444), .Y(new_n4445));
  AOI21xp33_ASAP7_75t_L     g04189(.A1(new_n4441), .A2(new_n4439), .B(new_n4436), .Y(new_n4446));
  NAND2xp33_ASAP7_75t_L     g04190(.A(new_n4441), .B(new_n4439), .Y(new_n4447));
  NOR2xp33_ASAP7_75t_L      g04191(.A(new_n4390), .B(new_n4447), .Y(new_n4448));
  NOR3xp33_ASAP7_75t_L      g04192(.A(new_n4448), .B(new_n4445), .C(new_n4446), .Y(new_n4449));
  NOR2xp33_ASAP7_75t_L      g04193(.A(new_n4443), .B(new_n4449), .Y(new_n4450));
  NAND2xp33_ASAP7_75t_L     g04194(.A(new_n4382), .B(new_n4450), .Y(new_n4451));
  AOI21xp33_ASAP7_75t_L     g04195(.A1(new_n4179), .A2(new_n4173), .B(new_n4185), .Y(new_n4452));
  AOI31xp33_ASAP7_75t_L     g04196(.A1(new_n4381), .A2(new_n4173), .A3(new_n4179), .B(new_n4452), .Y(new_n4453));
  OAI221xp5_ASAP7_75t_L     g04197(.A1(new_n4443), .A2(new_n4449), .B1(new_n4189), .B2(new_n4453), .C(new_n4381), .Y(new_n4454));
  NOR2xp33_ASAP7_75t_L      g04198(.A(new_n936), .B(new_n1962), .Y(new_n4455));
  AOI221xp5_ASAP7_75t_L     g04199(.A1(new_n1955), .A2(\b[14] ), .B1(new_n2093), .B2(\b[12] ), .C(new_n4455), .Y(new_n4456));
  INVx1_ASAP7_75t_L         g04200(.A(new_n4456), .Y(new_n4457));
  A2O1A1Ixp33_ASAP7_75t_L   g04201(.A1(new_n971), .A2(new_n1964), .B(new_n4457), .C(\a[23] ), .Y(new_n4458));
  O2A1O1Ixp33_ASAP7_75t_L   g04202(.A1(new_n1956), .A2(new_n1268), .B(new_n4456), .C(\a[23] ), .Y(new_n4459));
  AOI21xp33_ASAP7_75t_L     g04203(.A1(new_n4458), .A2(\a[23] ), .B(new_n4459), .Y(new_n4460));
  NAND3xp33_ASAP7_75t_L     g04204(.A(new_n4451), .B(new_n4454), .C(new_n4460), .Y(new_n4461));
  OAI21xp33_ASAP7_75t_L     g04205(.A1(new_n4443), .A2(new_n4449), .B(new_n4382), .Y(new_n4462));
  NOR2xp33_ASAP7_75t_L      g04206(.A(new_n4382), .B(new_n4450), .Y(new_n4463));
  AO21x2_ASAP7_75t_L        g04207(.A1(\a[23] ), .A2(new_n4458), .B(new_n4459), .Y(new_n4464));
  A2O1A1Ixp33_ASAP7_75t_L   g04208(.A1(new_n4462), .A2(new_n4382), .B(new_n4463), .C(new_n4464), .Y(new_n4465));
  NAND3xp33_ASAP7_75t_L     g04209(.A(new_n4220), .B(new_n4461), .C(new_n4465), .Y(new_n4466));
  OAI21xp33_ASAP7_75t_L     g04210(.A1(new_n4446), .A2(new_n4448), .B(new_n4445), .Y(new_n4467));
  NAND3xp33_ASAP7_75t_L     g04211(.A(new_n4434), .B(new_n4388), .C(new_n4442), .Y(new_n4468));
  NAND2xp33_ASAP7_75t_L     g04212(.A(new_n4468), .B(new_n4467), .Y(new_n4469));
  O2A1O1Ixp33_ASAP7_75t_L   g04213(.A1(new_n4453), .A2(new_n4189), .B(new_n4381), .C(new_n4469), .Y(new_n4470));
  NOR3xp33_ASAP7_75t_L      g04214(.A(new_n4470), .B(new_n4463), .C(new_n4464), .Y(new_n4471));
  AOI21xp33_ASAP7_75t_L     g04215(.A1(new_n4451), .A2(new_n4454), .B(new_n4460), .Y(new_n4472));
  OAI21xp33_ASAP7_75t_L     g04216(.A1(new_n4472), .A2(new_n4471), .B(new_n4207), .Y(new_n4473));
  NOR2xp33_ASAP7_75t_L      g04217(.A(new_n1150), .B(new_n1517), .Y(new_n4474));
  AOI221xp5_ASAP7_75t_L     g04218(.A1(\b[15] ), .A2(new_n1659), .B1(\b[17] ), .B2(new_n1511), .C(new_n4474), .Y(new_n4475));
  INVx1_ASAP7_75t_L         g04219(.A(new_n4475), .Y(new_n4476));
  A2O1A1Ixp33_ASAP7_75t_L   g04220(.A1(new_n1633), .A2(new_n1513), .B(new_n4476), .C(\a[20] ), .Y(new_n4477));
  O2A1O1Ixp33_ASAP7_75t_L   g04221(.A1(new_n1521), .A2(new_n1356), .B(new_n4475), .C(\a[20] ), .Y(new_n4478));
  AOI21xp33_ASAP7_75t_L     g04222(.A1(new_n4477), .A2(\a[20] ), .B(new_n4478), .Y(new_n4479));
  NAND3xp33_ASAP7_75t_L     g04223(.A(new_n4466), .B(new_n4473), .C(new_n4479), .Y(new_n4480));
  NOR3xp33_ASAP7_75t_L      g04224(.A(new_n4207), .B(new_n4471), .C(new_n4472), .Y(new_n4481));
  AOI21xp33_ASAP7_75t_L     g04225(.A1(new_n4465), .A2(new_n4461), .B(new_n4220), .Y(new_n4482));
  O2A1O1Ixp33_ASAP7_75t_L   g04226(.A1(new_n1521), .A2(new_n1356), .B(new_n4475), .C(new_n1501), .Y(new_n4483));
  A2O1A1Ixp33_ASAP7_75t_L   g04227(.A1(new_n1633), .A2(new_n1513), .B(new_n4476), .C(new_n1501), .Y(new_n4484));
  OAI21xp33_ASAP7_75t_L     g04228(.A1(new_n1501), .A2(new_n4483), .B(new_n4484), .Y(new_n4485));
  OAI21xp33_ASAP7_75t_L     g04229(.A1(new_n4482), .A2(new_n4481), .B(new_n4485), .Y(new_n4486));
  NAND2xp33_ASAP7_75t_L     g04230(.A(new_n4480), .B(new_n4486), .Y(new_n4487));
  A2O1A1O1Ixp25_ASAP7_75t_L g04231(.A1(new_n4201), .A2(new_n4200), .B(new_n4202), .C(new_n4207), .D(new_n4204), .Y(new_n4488));
  MAJIxp5_ASAP7_75t_L       g04232(.A(new_n4223), .B(new_n4488), .C(new_n4214), .Y(new_n4489));
  NOR2xp33_ASAP7_75t_L      g04233(.A(new_n4487), .B(new_n4489), .Y(new_n4490));
  NOR2xp33_ASAP7_75t_L      g04234(.A(new_n4482), .B(new_n4481), .Y(new_n4491));
  NAND3xp33_ASAP7_75t_L     g04235(.A(new_n4466), .B(new_n4473), .C(new_n4485), .Y(new_n4492));
  AOI21xp33_ASAP7_75t_L     g04236(.A1(new_n4466), .A2(new_n4473), .B(new_n4479), .Y(new_n4493));
  AOI21xp33_ASAP7_75t_L     g04237(.A1(new_n4492), .A2(new_n4491), .B(new_n4493), .Y(new_n4494));
  O2A1O1Ixp33_ASAP7_75t_L   g04238(.A1(new_n4488), .A2(new_n4214), .B(new_n4229), .C(new_n4494), .Y(new_n4495));
  OAI22xp33_ASAP7_75t_L     g04239(.A1(new_n1285), .A2(new_n1458), .B1(new_n1599), .B2(new_n2118), .Y(new_n4496));
  AOI221xp5_ASAP7_75t_L     g04240(.A1(new_n1209), .A2(\b[20] ), .B1(new_n1216), .B2(new_n1752), .C(new_n4496), .Y(new_n4497));
  XNOR2x2_ASAP7_75t_L       g04241(.A(new_n1206), .B(new_n4497), .Y(new_n4498));
  NOR3xp33_ASAP7_75t_L      g04242(.A(new_n4495), .B(new_n4498), .C(new_n4490), .Y(new_n4499));
  O2A1O1Ixp33_ASAP7_75t_L   g04243(.A1(new_n4226), .A2(new_n4213), .B(new_n4228), .C(new_n4239), .Y(new_n4500));
  NAND2xp33_ASAP7_75t_L     g04244(.A(new_n4494), .B(new_n4500), .Y(new_n4501));
  A2O1A1Ixp33_ASAP7_75t_L   g04245(.A1(new_n4237), .A2(new_n4228), .B(new_n4239), .C(new_n4487), .Y(new_n4502));
  XNOR2x2_ASAP7_75t_L       g04246(.A(\a[17] ), .B(new_n4497), .Y(new_n4503));
  AOI21xp33_ASAP7_75t_L     g04247(.A1(new_n4502), .A2(new_n4501), .B(new_n4503), .Y(new_n4504));
  OAI21xp33_ASAP7_75t_L     g04248(.A1(new_n4499), .A2(new_n4504), .B(new_n4378), .Y(new_n4505));
  INVx1_ASAP7_75t_L         g04249(.A(new_n4499), .Y(new_n4506));
  OAI21xp33_ASAP7_75t_L     g04250(.A1(new_n4490), .A2(new_n4495), .B(new_n4498), .Y(new_n4507));
  NAND4xp25_ASAP7_75t_L     g04251(.A(new_n4264), .B(new_n4506), .C(new_n4507), .D(new_n4249), .Y(new_n4508));
  NOR2xp33_ASAP7_75t_L      g04252(.A(new_n2188), .B(new_n869), .Y(new_n4509));
  AOI221xp5_ASAP7_75t_L     g04253(.A1(\b[21] ), .A2(new_n985), .B1(\b[22] ), .B2(new_n885), .C(new_n4509), .Y(new_n4510));
  OAI21xp33_ASAP7_75t_L     g04254(.A1(new_n872), .A2(new_n2194), .B(new_n4510), .Y(new_n4511));
  NOR2xp33_ASAP7_75t_L      g04255(.A(new_n867), .B(new_n4511), .Y(new_n4512));
  O2A1O1Ixp33_ASAP7_75t_L   g04256(.A1(new_n872), .A2(new_n2194), .B(new_n4510), .C(\a[14] ), .Y(new_n4513));
  NOR2xp33_ASAP7_75t_L      g04257(.A(new_n4513), .B(new_n4512), .Y(new_n4514));
  NAND3xp33_ASAP7_75t_L     g04258(.A(new_n4508), .B(new_n4514), .C(new_n4505), .Y(new_n4515));
  AOI22xp33_ASAP7_75t_L     g04259(.A1(new_n4506), .A2(new_n4507), .B1(new_n4249), .B2(new_n4264), .Y(new_n4516));
  A2O1A1O1Ixp25_ASAP7_75t_L g04260(.A1(new_n4245), .A2(new_n4246), .B(new_n4250), .C(new_n4507), .D(new_n4499), .Y(new_n4517));
  O2A1O1Ixp33_ASAP7_75t_L   g04261(.A1(new_n872), .A2(new_n2194), .B(new_n4510), .C(new_n867), .Y(new_n4518));
  INVx1_ASAP7_75t_L         g04262(.A(new_n4513), .Y(new_n4519));
  OAI21xp33_ASAP7_75t_L     g04263(.A1(new_n867), .A2(new_n4518), .B(new_n4519), .Y(new_n4520));
  A2O1A1Ixp33_ASAP7_75t_L   g04264(.A1(new_n4517), .A2(new_n4507), .B(new_n4516), .C(new_n4520), .Y(new_n4521));
  NAND2xp33_ASAP7_75t_L     g04265(.A(new_n4515), .B(new_n4521), .Y(new_n4522));
  NOR2xp33_ASAP7_75t_L      g04266(.A(new_n4377), .B(new_n4522), .Y(new_n4523));
  NAND2xp33_ASAP7_75t_L     g04267(.A(new_n4264), .B(new_n4263), .Y(new_n4524));
  O2A1O1Ixp33_ASAP7_75t_L   g04268(.A1(new_n4255), .A2(new_n867), .B(new_n4257), .C(new_n4524), .Y(new_n4525));
  AOI221xp5_ASAP7_75t_L     g04269(.A1(new_n4287), .A2(new_n4288), .B1(new_n4515), .B2(new_n4521), .C(new_n4525), .Y(new_n4526));
  OAI21xp33_ASAP7_75t_L     g04270(.A1(new_n4526), .A2(new_n4523), .B(new_n4375), .Y(new_n4527));
  A2O1A1Ixp33_ASAP7_75t_L   g04271(.A1(\a[14] ), .A2(new_n4266), .B(new_n4256), .C(new_n4376), .Y(new_n4528));
  O2A1O1Ixp33_ASAP7_75t_L   g04272(.A1(new_n3824), .A2(new_n3845), .B(new_n4045), .C(new_n4124), .Y(new_n4529));
  A2O1A1Ixp33_ASAP7_75t_L   g04273(.A1(new_n4273), .A2(new_n4274), .B(new_n4529), .C(new_n4528), .Y(new_n4530));
  NOR3xp33_ASAP7_75t_L      g04274(.A(new_n4378), .B(new_n4499), .C(new_n4504), .Y(new_n4531));
  NOR3xp33_ASAP7_75t_L      g04275(.A(new_n4531), .B(new_n4516), .C(new_n4520), .Y(new_n4532));
  AOI21xp33_ASAP7_75t_L     g04276(.A1(new_n4508), .A2(new_n4505), .B(new_n4514), .Y(new_n4533));
  NOR2xp33_ASAP7_75t_L      g04277(.A(new_n4533), .B(new_n4532), .Y(new_n4534));
  NAND2xp33_ASAP7_75t_L     g04278(.A(new_n4530), .B(new_n4534), .Y(new_n4535));
  NAND2xp33_ASAP7_75t_L     g04279(.A(new_n4377), .B(new_n4522), .Y(new_n4536));
  NAND3xp33_ASAP7_75t_L     g04280(.A(new_n4535), .B(new_n4536), .C(new_n4374), .Y(new_n4537));
  OAI211xp5_ASAP7_75t_L     g04281(.A1(new_n4293), .A2(new_n4367), .B(new_n4527), .C(new_n4537), .Y(new_n4538));
  AOI21xp33_ASAP7_75t_L     g04282(.A1(new_n4535), .A2(new_n4536), .B(new_n4374), .Y(new_n4539));
  NOR3xp33_ASAP7_75t_L      g04283(.A(new_n4523), .B(new_n4526), .C(new_n4375), .Y(new_n4540));
  OAI21xp33_ASAP7_75t_L     g04284(.A1(new_n4540), .A2(new_n4539), .B(new_n4294), .Y(new_n4541));
  NOR2xp33_ASAP7_75t_L      g04285(.A(new_n3079), .B(new_n513), .Y(new_n4542));
  AOI221xp5_ASAP7_75t_L     g04286(.A1(\b[27] ), .A2(new_n560), .B1(\b[29] ), .B2(new_n475), .C(new_n4542), .Y(new_n4543));
  O2A1O1Ixp33_ASAP7_75t_L   g04287(.A1(new_n477), .A2(new_n3104), .B(new_n4543), .C(new_n466), .Y(new_n4544));
  INVx1_ASAP7_75t_L         g04288(.A(new_n4544), .Y(new_n4545));
  O2A1O1Ixp33_ASAP7_75t_L   g04289(.A1(new_n477), .A2(new_n3104), .B(new_n4543), .C(\a[8] ), .Y(new_n4546));
  AOI21xp33_ASAP7_75t_L     g04290(.A1(new_n4545), .A2(\a[8] ), .B(new_n4546), .Y(new_n4547));
  NAND3xp33_ASAP7_75t_L     g04291(.A(new_n4538), .B(new_n4547), .C(new_n4541), .Y(new_n4548));
  NOR3xp33_ASAP7_75t_L      g04292(.A(new_n4294), .B(new_n4539), .C(new_n4540), .Y(new_n4549));
  AOI211xp5_ASAP7_75t_L     g04293(.A1(new_n4537), .A2(new_n4527), .B(new_n4293), .C(new_n4367), .Y(new_n4550));
  INVx1_ASAP7_75t_L         g04294(.A(new_n4546), .Y(new_n4551));
  OAI21xp33_ASAP7_75t_L     g04295(.A1(new_n466), .A2(new_n4544), .B(new_n4551), .Y(new_n4552));
  OAI21xp33_ASAP7_75t_L     g04296(.A1(new_n4549), .A2(new_n4550), .B(new_n4552), .Y(new_n4553));
  NAND2xp33_ASAP7_75t_L     g04297(.A(new_n4548), .B(new_n4553), .Y(new_n4554));
  AOI211xp5_ASAP7_75t_L     g04298(.A1(new_n4309), .A2(new_n4311), .B(new_n4368), .C(new_n4554), .Y(new_n4555));
  INVx1_ASAP7_75t_L         g04299(.A(new_n4368), .Y(new_n4556));
  NOR2xp33_ASAP7_75t_L      g04300(.A(new_n4549), .B(new_n4550), .Y(new_n4557));
  NAND3xp33_ASAP7_75t_L     g04301(.A(new_n4538), .B(new_n4541), .C(new_n4552), .Y(new_n4558));
  AOI21xp33_ASAP7_75t_L     g04302(.A1(new_n4538), .A2(new_n4541), .B(new_n4547), .Y(new_n4559));
  AOI21xp33_ASAP7_75t_L     g04303(.A1(new_n4557), .A2(new_n4558), .B(new_n4559), .Y(new_n4560));
  O2A1O1Ixp33_ASAP7_75t_L   g04304(.A1(new_n4315), .A2(new_n4330), .B(new_n4556), .C(new_n4560), .Y(new_n4561));
  NOR2xp33_ASAP7_75t_L      g04305(.A(new_n3456), .B(new_n375), .Y(new_n4562));
  AOI221xp5_ASAP7_75t_L     g04306(.A1(\b[32] ), .A2(new_n361), .B1(new_n349), .B2(\b[31] ), .C(new_n4562), .Y(new_n4563));
  O2A1O1Ixp33_ASAP7_75t_L   g04307(.A1(new_n356), .A2(new_n3897), .B(new_n4563), .C(new_n346), .Y(new_n4564));
  INVx1_ASAP7_75t_L         g04308(.A(new_n4564), .Y(new_n4565));
  O2A1O1Ixp33_ASAP7_75t_L   g04309(.A1(new_n356), .A2(new_n3897), .B(new_n4563), .C(\a[5] ), .Y(new_n4566));
  AOI21xp33_ASAP7_75t_L     g04310(.A1(new_n4565), .A2(\a[5] ), .B(new_n4566), .Y(new_n4567));
  OAI21xp33_ASAP7_75t_L     g04311(.A1(new_n4561), .A2(new_n4555), .B(new_n4567), .Y(new_n4568));
  INVx1_ASAP7_75t_L         g04312(.A(new_n4555), .Y(new_n4569));
  A2O1A1Ixp33_ASAP7_75t_L   g04313(.A1(new_n4309), .A2(new_n4311), .B(new_n4368), .C(new_n4554), .Y(new_n4570));
  INVx1_ASAP7_75t_L         g04314(.A(new_n4567), .Y(new_n4571));
  NAND3xp33_ASAP7_75t_L     g04315(.A(new_n4569), .B(new_n4570), .C(new_n4571), .Y(new_n4572));
  AOI21xp33_ASAP7_75t_L     g04316(.A1(new_n4572), .A2(new_n4568), .B(new_n4339), .Y(new_n4573));
  NAND2xp33_ASAP7_75t_L     g04317(.A(new_n4081), .B(new_n4076), .Y(new_n4574));
  MAJIxp5_ASAP7_75t_L       g04318(.A(new_n3887), .B(new_n4574), .C(new_n4087), .Y(new_n4575));
  NOR3xp33_ASAP7_75t_L      g04319(.A(new_n4555), .B(new_n4561), .C(new_n4567), .Y(new_n4576));
  A2O1A1O1Ixp25_ASAP7_75t_L g04320(.A1(new_n4323), .A2(new_n4575), .B(new_n4338), .C(new_n4568), .D(new_n4576), .Y(new_n4577));
  NOR2xp33_ASAP7_75t_L      g04321(.A(new_n4101), .B(new_n287), .Y(new_n4578));
  AOI221xp5_ASAP7_75t_L     g04322(.A1(\b[34] ), .A2(new_n264), .B1(\b[35] ), .B2(new_n283), .C(new_n4578), .Y(new_n4579));
  NOR2xp33_ASAP7_75t_L      g04323(.A(\b[34] ), .B(\b[35] ), .Y(new_n4580));
  INVx1_ASAP7_75t_L         g04324(.A(\b[35] ), .Y(new_n4581));
  NOR2xp33_ASAP7_75t_L      g04325(.A(new_n4344), .B(new_n4581), .Y(new_n4582));
  NOR2xp33_ASAP7_75t_L      g04326(.A(new_n4580), .B(new_n4582), .Y(new_n4583));
  A2O1A1Ixp33_ASAP7_75t_L   g04327(.A1(\b[34] ), .A2(\b[33] ), .B(new_n4348), .C(new_n4583), .Y(new_n4584));
  O2A1O1Ixp33_ASAP7_75t_L   g04328(.A1(new_n3674), .A2(new_n3891), .B(new_n3894), .C(new_n4106), .Y(new_n4585));
  O2A1O1Ixp33_ASAP7_75t_L   g04329(.A1(new_n4102), .A2(new_n4585), .B(new_n4346), .C(new_n4345), .Y(new_n4586));
  INVx1_ASAP7_75t_L         g04330(.A(new_n4583), .Y(new_n4587));
  NAND2xp33_ASAP7_75t_L     g04331(.A(new_n4587), .B(new_n4586), .Y(new_n4588));
  NAND2xp33_ASAP7_75t_L     g04332(.A(new_n4584), .B(new_n4588), .Y(new_n4589));
  O2A1O1Ixp33_ASAP7_75t_L   g04333(.A1(new_n279), .A2(new_n4589), .B(new_n4579), .C(new_n257), .Y(new_n4590));
  INVx1_ASAP7_75t_L         g04334(.A(new_n4590), .Y(new_n4591));
  O2A1O1Ixp33_ASAP7_75t_L   g04335(.A1(new_n279), .A2(new_n4589), .B(new_n4579), .C(\a[2] ), .Y(new_n4592));
  AOI21xp33_ASAP7_75t_L     g04336(.A1(new_n4591), .A2(\a[2] ), .B(new_n4592), .Y(new_n4593));
  A2O1A1Ixp33_ASAP7_75t_L   g04337(.A1(new_n4577), .A2(new_n4568), .B(new_n4573), .C(new_n4593), .Y(new_n4594));
  AOI21xp33_ASAP7_75t_L     g04338(.A1(new_n4076), .A2(new_n4081), .B(new_n4087), .Y(new_n4595));
  OAI22xp33_ASAP7_75t_L     g04339(.A1(new_n4324), .A2(new_n3886), .B1(new_n4595), .B2(new_n4095), .Y(new_n4596));
  AOI21xp33_ASAP7_75t_L     g04340(.A1(new_n4331), .A2(new_n4332), .B(new_n4335), .Y(new_n4597));
  A2O1A1Ixp33_ASAP7_75t_L   g04341(.A1(new_n4596), .A2(new_n4094), .B(new_n4597), .C(new_n4336), .Y(new_n4598));
  INVx1_ASAP7_75t_L         g04342(.A(new_n4568), .Y(new_n4599));
  OAI21xp33_ASAP7_75t_L     g04343(.A1(new_n4576), .A2(new_n4599), .B(new_n4598), .Y(new_n4600));
  NAND3xp33_ASAP7_75t_L     g04344(.A(new_n4339), .B(new_n4572), .C(new_n4568), .Y(new_n4601));
  INVx1_ASAP7_75t_L         g04345(.A(new_n4593), .Y(new_n4602));
  NAND3xp33_ASAP7_75t_L     g04346(.A(new_n4600), .B(new_n4601), .C(new_n4602), .Y(new_n4603));
  NAND2xp33_ASAP7_75t_L     g04347(.A(new_n4603), .B(new_n4594), .Y(new_n4604));
  INVx1_ASAP7_75t_L         g04348(.A(new_n4604), .Y(new_n4605));
  A2O1A1O1Ixp25_ASAP7_75t_L g04349(.A1(new_n4357), .A2(new_n4360), .B(new_n4363), .C(new_n4366), .D(new_n4605), .Y(new_n4606));
  MAJIxp5_ASAP7_75t_L       g04350(.A(new_n4363), .B(new_n4356), .C(new_n4358), .Y(new_n4607));
  NOR2xp33_ASAP7_75t_L      g04351(.A(new_n4604), .B(new_n4607), .Y(new_n4608));
  NOR2xp33_ASAP7_75t_L      g04352(.A(new_n4608), .B(new_n4606), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g04353(.A(new_n4344), .B(new_n287), .Y(new_n4610));
  AOI221xp5_ASAP7_75t_L     g04354(.A1(\b[35] ), .A2(new_n264), .B1(\b[36] ), .B2(new_n283), .C(new_n4610), .Y(new_n4611));
  NOR2xp33_ASAP7_75t_L      g04355(.A(\b[35] ), .B(\b[36] ), .Y(new_n4612));
  INVx1_ASAP7_75t_L         g04356(.A(\b[36] ), .Y(new_n4613));
  NOR2xp33_ASAP7_75t_L      g04357(.A(new_n4581), .B(new_n4613), .Y(new_n4614));
  NOR2xp33_ASAP7_75t_L      g04358(.A(new_n4612), .B(new_n4614), .Y(new_n4615));
  INVx1_ASAP7_75t_L         g04359(.A(new_n4615), .Y(new_n4616));
  O2A1O1Ixp33_ASAP7_75t_L   g04360(.A1(new_n4344), .A2(new_n4581), .B(new_n4584), .C(new_n4616), .Y(new_n4617));
  O2A1O1Ixp33_ASAP7_75t_L   g04361(.A1(new_n4345), .A2(new_n4348), .B(new_n4583), .C(new_n4582), .Y(new_n4618));
  INVx1_ASAP7_75t_L         g04362(.A(new_n4618), .Y(new_n4619));
  NOR2xp33_ASAP7_75t_L      g04363(.A(new_n4615), .B(new_n4619), .Y(new_n4620));
  NOR2xp33_ASAP7_75t_L      g04364(.A(new_n4617), .B(new_n4620), .Y(new_n4621));
  INVx1_ASAP7_75t_L         g04365(.A(new_n4621), .Y(new_n4622));
  O2A1O1Ixp33_ASAP7_75t_L   g04366(.A1(new_n279), .A2(new_n4622), .B(new_n4611), .C(new_n257), .Y(new_n4623));
  OAI21xp33_ASAP7_75t_L     g04367(.A1(new_n279), .A2(new_n4622), .B(new_n4611), .Y(new_n4624));
  NAND2xp33_ASAP7_75t_L     g04368(.A(new_n257), .B(new_n4624), .Y(new_n4625));
  OA21x2_ASAP7_75t_L        g04369(.A1(new_n257), .A2(new_n4623), .B(new_n4625), .Y(new_n4626));
  NOR2xp33_ASAP7_75t_L      g04370(.A(new_n3674), .B(new_n375), .Y(new_n4627));
  AOI221xp5_ASAP7_75t_L     g04371(.A1(\b[33] ), .A2(new_n361), .B1(new_n349), .B2(\b[32] ), .C(new_n4627), .Y(new_n4628));
  OA21x2_ASAP7_75t_L        g04372(.A1(new_n356), .A2(new_n4108), .B(new_n4628), .Y(new_n4629));
  O2A1O1Ixp33_ASAP7_75t_L   g04373(.A1(new_n356), .A2(new_n4108), .B(new_n4628), .C(new_n346), .Y(new_n4630));
  NAND2xp33_ASAP7_75t_L     g04374(.A(\a[5] ), .B(new_n4629), .Y(new_n4631));
  OA21x2_ASAP7_75t_L        g04375(.A1(new_n4629), .A2(new_n4630), .B(new_n4631), .Y(new_n4632));
  AOI21xp33_ASAP7_75t_L     g04376(.A1(new_n4311), .A2(new_n4309), .B(new_n4368), .Y(new_n4633));
  A2O1A1Ixp33_ASAP7_75t_L   g04377(.A1(new_n4053), .A2(new_n3918), .B(new_n4284), .C(new_n4283), .Y(new_n4634));
  A2O1A1Ixp33_ASAP7_75t_L   g04378(.A1(new_n4634), .A2(new_n4291), .B(new_n4539), .C(new_n4537), .Y(new_n4635));
  INVx1_ASAP7_75t_L         g04379(.A(new_n4492), .Y(new_n4636));
  A2O1A1O1Ixp25_ASAP7_75t_L g04380(.A1(new_n4218), .A2(new_n4198), .B(new_n4206), .C(new_n4461), .D(new_n4472), .Y(new_n4637));
  NAND2xp33_ASAP7_75t_L     g04381(.A(new_n4442), .B(new_n4434), .Y(new_n4638));
  INVx1_ASAP7_75t_L         g04382(.A(new_n4423), .Y(new_n4639));
  NOR2xp33_ASAP7_75t_L      g04383(.A(new_n427), .B(new_n3510), .Y(new_n4640));
  AOI221xp5_ASAP7_75t_L     g04384(.A1(\b[4] ), .A2(new_n3708), .B1(\b[5] ), .B2(new_n3499), .C(new_n4640), .Y(new_n4641));
  O2A1O1Ixp33_ASAP7_75t_L   g04385(.A1(new_n3513), .A2(new_n434), .B(new_n4641), .C(new_n3493), .Y(new_n4642));
  OAI31xp33_ASAP7_75t_L     g04386(.A1(new_n433), .A2(new_n431), .A3(new_n3513), .B(new_n4641), .Y(new_n4643));
  NAND2xp33_ASAP7_75t_L     g04387(.A(new_n3493), .B(new_n4643), .Y(new_n4644));
  OAI21xp33_ASAP7_75t_L     g04388(.A1(new_n3493), .A2(new_n4642), .B(new_n4644), .Y(new_n4645));
  INVx1_ASAP7_75t_L         g04389(.A(\a[36] ), .Y(new_n4646));
  NAND2xp33_ASAP7_75t_L     g04390(.A(\a[35] ), .B(new_n4646), .Y(new_n4647));
  NAND2xp33_ASAP7_75t_L     g04391(.A(\a[36] ), .B(new_n4145), .Y(new_n4648));
  AND2x2_ASAP7_75t_L        g04392(.A(new_n4647), .B(new_n4648), .Y(new_n4649));
  NOR2xp33_ASAP7_75t_L      g04393(.A(new_n284), .B(new_n4649), .Y(new_n4650));
  INVx1_ASAP7_75t_L         g04394(.A(new_n4650), .Y(new_n4651));
  NOR2xp33_ASAP7_75t_L      g04395(.A(new_n4651), .B(new_n4408), .Y(new_n4652));
  NOR2xp33_ASAP7_75t_L      g04396(.A(new_n4650), .B(new_n4428), .Y(new_n4653));
  NAND2xp33_ASAP7_75t_L     g04397(.A(\b[3] ), .B(new_n4156), .Y(new_n4654));
  NAND2xp33_ASAP7_75t_L     g04398(.A(\b[1] ), .B(new_n4402), .Y(new_n4655));
  NAND2xp33_ASAP7_75t_L     g04399(.A(\b[2] ), .B(new_n4155), .Y(new_n4656));
  NAND2xp33_ASAP7_75t_L     g04400(.A(new_n4151), .B(new_n312), .Y(new_n4657));
  NAND5xp2_ASAP7_75t_L      g04401(.A(new_n4657), .B(new_n4656), .C(new_n4655), .D(new_n4654), .E(\a[35] ), .Y(new_n4658));
  OAI211xp5_ASAP7_75t_L     g04402(.A1(new_n4397), .A2(new_n262), .B(new_n4654), .C(new_n4656), .Y(new_n4659));
  A2O1A1Ixp33_ASAP7_75t_L   g04403(.A1(new_n312), .A2(new_n4151), .B(new_n4659), .C(new_n4145), .Y(new_n4660));
  NAND2xp33_ASAP7_75t_L     g04404(.A(new_n4658), .B(new_n4660), .Y(new_n4661));
  OAI21xp33_ASAP7_75t_L     g04405(.A1(new_n4653), .A2(new_n4652), .B(new_n4661), .Y(new_n4662));
  A2O1A1Ixp33_ASAP7_75t_L   g04406(.A1(new_n4425), .A2(new_n4426), .B(new_n4153), .C(new_n4650), .Y(new_n4663));
  NAND2xp33_ASAP7_75t_L     g04407(.A(new_n4651), .B(new_n4408), .Y(new_n4664));
  INVx1_ASAP7_75t_L         g04408(.A(new_n4657), .Y(new_n4665));
  A2O1A1Ixp33_ASAP7_75t_L   g04409(.A1(new_n312), .A2(new_n4151), .B(new_n4659), .C(\a[35] ), .Y(new_n4666));
  AOI211xp5_ASAP7_75t_L     g04410(.A1(new_n312), .A2(new_n4151), .B(new_n4145), .C(new_n4659), .Y(new_n4667));
  O2A1O1Ixp33_ASAP7_75t_L   g04411(.A1(new_n4659), .A2(new_n4665), .B(new_n4666), .C(new_n4667), .Y(new_n4668));
  NAND3xp33_ASAP7_75t_L     g04412(.A(new_n4664), .B(new_n4668), .C(new_n4663), .Y(new_n4669));
  NAND3xp33_ASAP7_75t_L     g04413(.A(new_n4662), .B(new_n4669), .C(new_n4645), .Y(new_n4670));
  AOI21xp33_ASAP7_75t_L     g04414(.A1(new_n4664), .A2(new_n4663), .B(new_n4668), .Y(new_n4671));
  NOR3xp33_ASAP7_75t_L      g04415(.A(new_n4652), .B(new_n4653), .C(new_n4661), .Y(new_n4672));
  NOR3xp33_ASAP7_75t_L      g04416(.A(new_n4672), .B(new_n4671), .C(new_n4645), .Y(new_n4673));
  AOI211xp5_ASAP7_75t_L     g04417(.A1(new_n4645), .A2(new_n4670), .B(new_n4673), .C(new_n4422), .Y(new_n4674));
  OAI211xp5_ASAP7_75t_L     g04418(.A1(new_n3513), .A2(new_n434), .B(\a[32] ), .C(new_n4641), .Y(new_n4675));
  NAND4xp25_ASAP7_75t_L     g04419(.A(new_n4662), .B(new_n4669), .C(new_n4644), .D(new_n4675), .Y(new_n4676));
  OAI21xp33_ASAP7_75t_L     g04420(.A1(new_n4671), .A2(new_n4672), .B(new_n4645), .Y(new_n4677));
  AOI211xp5_ASAP7_75t_L     g04421(.A1(new_n4677), .A2(new_n4676), .B(new_n4421), .C(new_n4440), .Y(new_n4678));
  NOR2xp33_ASAP7_75t_L      g04422(.A(new_n534), .B(new_n2925), .Y(new_n4679));
  AOI221xp5_ASAP7_75t_L     g04423(.A1(\b[7] ), .A2(new_n3129), .B1(\b[9] ), .B2(new_n2938), .C(new_n4679), .Y(new_n4680));
  O2A1O1Ixp33_ASAP7_75t_L   g04424(.A1(new_n2940), .A2(new_n1066), .B(new_n4680), .C(new_n2928), .Y(new_n4681));
  INVx1_ASAP7_75t_L         g04425(.A(new_n4680), .Y(new_n4682));
  A2O1A1Ixp33_ASAP7_75t_L   g04426(.A1(new_n602), .A2(new_n2932), .B(new_n4682), .C(new_n2928), .Y(new_n4683));
  OAI21xp33_ASAP7_75t_L     g04427(.A1(new_n2928), .A2(new_n4681), .B(new_n4683), .Y(new_n4684));
  OAI21xp33_ASAP7_75t_L     g04428(.A1(new_n4678), .A2(new_n4674), .B(new_n4684), .Y(new_n4685));
  OAI211xp5_ASAP7_75t_L     g04429(.A1(new_n4421), .A2(new_n4440), .B(new_n4676), .C(new_n4677), .Y(new_n4686));
  A2O1A1Ixp33_ASAP7_75t_L   g04430(.A1(new_n4645), .A2(new_n4670), .B(new_n4673), .C(new_n4422), .Y(new_n4687));
  A2O1A1Ixp33_ASAP7_75t_L   g04431(.A1(new_n602), .A2(new_n2932), .B(new_n4682), .C(\a[29] ), .Y(new_n4688));
  O2A1O1Ixp33_ASAP7_75t_L   g04432(.A1(new_n2940), .A2(new_n1066), .B(new_n4680), .C(\a[29] ), .Y(new_n4689));
  AOI21xp33_ASAP7_75t_L     g04433(.A1(new_n4688), .A2(\a[29] ), .B(new_n4689), .Y(new_n4690));
  NAND3xp33_ASAP7_75t_L     g04434(.A(new_n4687), .B(new_n4690), .C(new_n4686), .Y(new_n4691));
  AOI221xp5_ASAP7_75t_L     g04435(.A1(new_n4685), .A2(new_n4691), .B1(new_n4390), .B2(new_n4447), .C(new_n4639), .Y(new_n4692));
  NOR3xp33_ASAP7_75t_L      g04436(.A(new_n4438), .B(new_n4420), .C(new_n4437), .Y(new_n4693));
  O2A1O1Ixp33_ASAP7_75t_L   g04437(.A1(new_n4420), .A2(new_n4437), .B(new_n4423), .C(new_n4693), .Y(new_n4694));
  NAND2xp33_ASAP7_75t_L     g04438(.A(new_n4691), .B(new_n4685), .Y(new_n4695));
  O2A1O1Ixp33_ASAP7_75t_L   g04439(.A1(new_n4436), .A2(new_n4694), .B(new_n4423), .C(new_n4695), .Y(new_n4696));
  NOR2xp33_ASAP7_75t_L      g04440(.A(new_n748), .B(new_n2410), .Y(new_n4697));
  AOI221xp5_ASAP7_75t_L     g04441(.A1(\b[10] ), .A2(new_n2577), .B1(\b[12] ), .B2(new_n2423), .C(new_n4697), .Y(new_n4698));
  O2A1O1Ixp33_ASAP7_75t_L   g04442(.A1(new_n2425), .A2(new_n841), .B(new_n4698), .C(new_n2413), .Y(new_n4699));
  INVx1_ASAP7_75t_L         g04443(.A(new_n4699), .Y(new_n4700));
  O2A1O1Ixp33_ASAP7_75t_L   g04444(.A1(new_n2425), .A2(new_n841), .B(new_n4698), .C(\a[26] ), .Y(new_n4701));
  AOI21xp33_ASAP7_75t_L     g04445(.A1(new_n4700), .A2(\a[26] ), .B(new_n4701), .Y(new_n4702));
  OAI21xp33_ASAP7_75t_L     g04446(.A1(new_n4692), .A2(new_n4696), .B(new_n4702), .Y(new_n4703));
  O2A1O1Ixp33_ASAP7_75t_L   g04447(.A1(new_n4396), .A2(new_n4433), .B(new_n4390), .C(new_n4639), .Y(new_n4704));
  NAND2xp33_ASAP7_75t_L     g04448(.A(new_n4695), .B(new_n4704), .Y(new_n4705));
  AOI21xp33_ASAP7_75t_L     g04449(.A1(new_n4687), .A2(new_n4686), .B(new_n4690), .Y(new_n4706));
  NOR3xp33_ASAP7_75t_L      g04450(.A(new_n4674), .B(new_n4678), .C(new_n4684), .Y(new_n4707));
  NOR2xp33_ASAP7_75t_L      g04451(.A(new_n4706), .B(new_n4707), .Y(new_n4708));
  A2O1A1Ixp33_ASAP7_75t_L   g04452(.A1(new_n4447), .A2(new_n4390), .B(new_n4639), .C(new_n4708), .Y(new_n4709));
  INVx1_ASAP7_75t_L         g04453(.A(new_n4701), .Y(new_n4710));
  OAI21xp33_ASAP7_75t_L     g04454(.A1(new_n2413), .A2(new_n4699), .B(new_n4710), .Y(new_n4711));
  NAND3xp33_ASAP7_75t_L     g04455(.A(new_n4705), .B(new_n4709), .C(new_n4711), .Y(new_n4712));
  NAND2xp33_ASAP7_75t_L     g04456(.A(new_n4703), .B(new_n4712), .Y(new_n4713));
  O2A1O1Ixp33_ASAP7_75t_L   g04457(.A1(new_n4388), .A2(new_n4638), .B(new_n4462), .C(new_n4713), .Y(new_n4714));
  O2A1O1Ixp33_ASAP7_75t_L   g04458(.A1(new_n2413), .A2(new_n4385), .B(new_n4444), .C(new_n4638), .Y(new_n4715));
  AOI221xp5_ASAP7_75t_L     g04459(.A1(new_n4469), .A2(new_n4382), .B1(new_n4712), .B2(new_n4703), .C(new_n4715), .Y(new_n4716));
  NOR2xp33_ASAP7_75t_L      g04460(.A(new_n960), .B(new_n1962), .Y(new_n4717));
  AOI221xp5_ASAP7_75t_L     g04461(.A1(new_n1955), .A2(\b[15] ), .B1(new_n2093), .B2(\b[13] ), .C(new_n4717), .Y(new_n4718));
  O2A1O1Ixp33_ASAP7_75t_L   g04462(.A1(new_n1956), .A2(new_n1774), .B(new_n4718), .C(new_n1952), .Y(new_n4719));
  INVx1_ASAP7_75t_L         g04463(.A(new_n4718), .Y(new_n4720));
  A2O1A1Ixp33_ASAP7_75t_L   g04464(.A1(new_n1052), .A2(new_n1964), .B(new_n4720), .C(new_n1952), .Y(new_n4721));
  OAI21xp33_ASAP7_75t_L     g04465(.A1(new_n1952), .A2(new_n4719), .B(new_n4721), .Y(new_n4722));
  NOR3xp33_ASAP7_75t_L      g04466(.A(new_n4714), .B(new_n4716), .C(new_n4722), .Y(new_n4723));
  AOI21xp33_ASAP7_75t_L     g04467(.A1(new_n4705), .A2(new_n4709), .B(new_n4711), .Y(new_n4724));
  NOR3xp33_ASAP7_75t_L      g04468(.A(new_n4696), .B(new_n4702), .C(new_n4692), .Y(new_n4725));
  NOR2xp33_ASAP7_75t_L      g04469(.A(new_n4725), .B(new_n4724), .Y(new_n4726));
  A2O1A1Ixp33_ASAP7_75t_L   g04470(.A1(new_n4469), .A2(new_n4382), .B(new_n4715), .C(new_n4726), .Y(new_n4727));
  O2A1O1Ixp33_ASAP7_75t_L   g04471(.A1(new_n4449), .A2(new_n4445), .B(new_n4382), .C(new_n4715), .Y(new_n4728));
  NAND2xp33_ASAP7_75t_L     g04472(.A(new_n4713), .B(new_n4728), .Y(new_n4729));
  A2O1A1Ixp33_ASAP7_75t_L   g04473(.A1(new_n1052), .A2(new_n1964), .B(new_n4720), .C(\a[23] ), .Y(new_n4730));
  O2A1O1Ixp33_ASAP7_75t_L   g04474(.A1(new_n1956), .A2(new_n1774), .B(new_n4718), .C(\a[23] ), .Y(new_n4731));
  AOI21xp33_ASAP7_75t_L     g04475(.A1(new_n4730), .A2(\a[23] ), .B(new_n4731), .Y(new_n4732));
  AOI21xp33_ASAP7_75t_L     g04476(.A1(new_n4727), .A2(new_n4729), .B(new_n4732), .Y(new_n4733));
  NOR3xp33_ASAP7_75t_L      g04477(.A(new_n4637), .B(new_n4733), .C(new_n4723), .Y(new_n4734));
  A2O1A1Ixp33_ASAP7_75t_L   g04478(.A1(new_n4205), .A2(new_n3991), .B(new_n3989), .C(new_n4198), .Y(new_n4735));
  A2O1A1Ixp33_ASAP7_75t_L   g04479(.A1(new_n4735), .A2(new_n4203), .B(new_n4471), .C(new_n4465), .Y(new_n4736));
  NAND3xp33_ASAP7_75t_L     g04480(.A(new_n4727), .B(new_n4729), .C(new_n4732), .Y(new_n4737));
  OAI21xp33_ASAP7_75t_L     g04481(.A1(new_n4716), .A2(new_n4714), .B(new_n4722), .Y(new_n4738));
  AOI21xp33_ASAP7_75t_L     g04482(.A1(new_n4738), .A2(new_n4737), .B(new_n4736), .Y(new_n4739));
  NOR2xp33_ASAP7_75t_L      g04483(.A(new_n1349), .B(new_n1517), .Y(new_n4740));
  AOI221xp5_ASAP7_75t_L     g04484(.A1(\b[16] ), .A2(new_n1659), .B1(\b[18] ), .B2(new_n1511), .C(new_n4740), .Y(new_n4741));
  O2A1O1Ixp33_ASAP7_75t_L   g04485(.A1(new_n1521), .A2(new_n1464), .B(new_n4741), .C(new_n1501), .Y(new_n4742));
  INVx1_ASAP7_75t_L         g04486(.A(new_n4741), .Y(new_n4743));
  A2O1A1Ixp33_ASAP7_75t_L   g04487(.A1(new_n2329), .A2(new_n1513), .B(new_n4743), .C(new_n1501), .Y(new_n4744));
  OAI21xp33_ASAP7_75t_L     g04488(.A1(new_n1501), .A2(new_n4742), .B(new_n4744), .Y(new_n4745));
  OAI21xp33_ASAP7_75t_L     g04489(.A1(new_n4739), .A2(new_n4734), .B(new_n4745), .Y(new_n4746));
  NAND3xp33_ASAP7_75t_L     g04490(.A(new_n4736), .B(new_n4737), .C(new_n4738), .Y(new_n4747));
  OAI21xp33_ASAP7_75t_L     g04491(.A1(new_n4723), .A2(new_n4733), .B(new_n4637), .Y(new_n4748));
  A2O1A1Ixp33_ASAP7_75t_L   g04492(.A1(new_n2329), .A2(new_n1513), .B(new_n4743), .C(\a[20] ), .Y(new_n4749));
  O2A1O1Ixp33_ASAP7_75t_L   g04493(.A1(new_n1521), .A2(new_n1464), .B(new_n4741), .C(\a[20] ), .Y(new_n4750));
  AOI21xp33_ASAP7_75t_L     g04494(.A1(new_n4749), .A2(\a[20] ), .B(new_n4750), .Y(new_n4751));
  NAND3xp33_ASAP7_75t_L     g04495(.A(new_n4747), .B(new_n4751), .C(new_n4748), .Y(new_n4752));
  AOI221xp5_ASAP7_75t_L     g04496(.A1(new_n4746), .A2(new_n4752), .B1(new_n4487), .B2(new_n4489), .C(new_n4636), .Y(new_n4753));
  NAND2xp33_ASAP7_75t_L     g04497(.A(new_n4752), .B(new_n4746), .Y(new_n4754));
  O2A1O1Ixp33_ASAP7_75t_L   g04498(.A1(new_n4494), .A2(new_n4500), .B(new_n4492), .C(new_n4754), .Y(new_n4755));
  NOR2xp33_ASAP7_75t_L      g04499(.A(new_n1745), .B(new_n2118), .Y(new_n4756));
  AOI221xp5_ASAP7_75t_L     g04500(.A1(\b[19] ), .A2(new_n1290), .B1(\b[21] ), .B2(new_n1209), .C(new_n4756), .Y(new_n4757));
  O2A1O1Ixp33_ASAP7_75t_L   g04501(.A1(new_n1210), .A2(new_n1901), .B(new_n4757), .C(new_n1206), .Y(new_n4758));
  O2A1O1Ixp33_ASAP7_75t_L   g04502(.A1(new_n1210), .A2(new_n1901), .B(new_n4757), .C(\a[17] ), .Y(new_n4759));
  INVx1_ASAP7_75t_L         g04503(.A(new_n4759), .Y(new_n4760));
  OAI21xp33_ASAP7_75t_L     g04504(.A1(new_n1206), .A2(new_n4758), .B(new_n4760), .Y(new_n4761));
  NOR3xp33_ASAP7_75t_L      g04505(.A(new_n4755), .B(new_n4761), .C(new_n4753), .Y(new_n4762));
  OAI211xp5_ASAP7_75t_L     g04506(.A1(new_n4494), .A2(new_n4500), .B(new_n4754), .C(new_n4492), .Y(new_n4763));
  AOI21xp33_ASAP7_75t_L     g04507(.A1(new_n4747), .A2(new_n4748), .B(new_n4751), .Y(new_n4764));
  NOR3xp33_ASAP7_75t_L      g04508(.A(new_n4734), .B(new_n4739), .C(new_n4745), .Y(new_n4765));
  NOR2xp33_ASAP7_75t_L      g04509(.A(new_n4764), .B(new_n4765), .Y(new_n4766));
  A2O1A1Ixp33_ASAP7_75t_L   g04510(.A1(new_n4487), .A2(new_n4489), .B(new_n4636), .C(new_n4766), .Y(new_n4767));
  INVx1_ASAP7_75t_L         g04511(.A(new_n4757), .Y(new_n4768));
  A2O1A1Ixp33_ASAP7_75t_L   g04512(.A1(new_n2836), .A2(new_n1216), .B(new_n4768), .C(\a[17] ), .Y(new_n4769));
  AOI21xp33_ASAP7_75t_L     g04513(.A1(new_n4769), .A2(\a[17] ), .B(new_n4759), .Y(new_n4770));
  AOI21xp33_ASAP7_75t_L     g04514(.A1(new_n4767), .A2(new_n4763), .B(new_n4770), .Y(new_n4771));
  NOR3xp33_ASAP7_75t_L      g04515(.A(new_n4517), .B(new_n4762), .C(new_n4771), .Y(new_n4772));
  A2O1A1O1Ixp25_ASAP7_75t_L g04516(.A1(new_n4244), .A2(new_n4248), .B(new_n4251), .C(new_n4249), .D(new_n4504), .Y(new_n4773));
  NAND3xp33_ASAP7_75t_L     g04517(.A(new_n4767), .B(new_n4763), .C(new_n4770), .Y(new_n4774));
  OAI21xp33_ASAP7_75t_L     g04518(.A1(new_n4753), .A2(new_n4755), .B(new_n4761), .Y(new_n4775));
  AOI211xp5_ASAP7_75t_L     g04519(.A1(new_n4775), .A2(new_n4774), .B(new_n4499), .C(new_n4773), .Y(new_n4776));
  NOR2xp33_ASAP7_75t_L      g04520(.A(new_n2188), .B(new_n864), .Y(new_n4777));
  AOI221xp5_ASAP7_75t_L     g04521(.A1(\b[22] ), .A2(new_n985), .B1(\b[24] ), .B2(new_n886), .C(new_n4777), .Y(new_n4778));
  O2A1O1Ixp33_ASAP7_75t_L   g04522(.A1(new_n872), .A2(new_n2853), .B(new_n4778), .C(new_n867), .Y(new_n4779));
  O2A1O1Ixp33_ASAP7_75t_L   g04523(.A1(new_n872), .A2(new_n2853), .B(new_n4778), .C(\a[14] ), .Y(new_n4780));
  INVx1_ASAP7_75t_L         g04524(.A(new_n4780), .Y(new_n4781));
  OAI21xp33_ASAP7_75t_L     g04525(.A1(new_n867), .A2(new_n4779), .B(new_n4781), .Y(new_n4782));
  NOR3xp33_ASAP7_75t_L      g04526(.A(new_n4772), .B(new_n4776), .C(new_n4782), .Y(new_n4783));
  OAI211xp5_ASAP7_75t_L     g04527(.A1(new_n4499), .A2(new_n4773), .B(new_n4774), .C(new_n4775), .Y(new_n4784));
  OAI21xp33_ASAP7_75t_L     g04528(.A1(new_n4762), .A2(new_n4771), .B(new_n4517), .Y(new_n4785));
  OA21x2_ASAP7_75t_L        g04529(.A1(new_n867), .A2(new_n4779), .B(new_n4781), .Y(new_n4786));
  AOI21xp33_ASAP7_75t_L     g04530(.A1(new_n4784), .A2(new_n4785), .B(new_n4786), .Y(new_n4787));
  NOR2xp33_ASAP7_75t_L      g04531(.A(new_n4787), .B(new_n4783), .Y(new_n4788));
  A2O1A1Ixp33_ASAP7_75t_L   g04532(.A1(new_n4534), .A2(new_n4530), .B(new_n4533), .C(new_n4788), .Y(new_n4789));
  A2O1A1O1Ixp25_ASAP7_75t_L g04533(.A1(new_n4288), .A2(new_n4287), .B(new_n4525), .C(new_n4515), .D(new_n4533), .Y(new_n4790));
  NAND3xp33_ASAP7_75t_L     g04534(.A(new_n4786), .B(new_n4785), .C(new_n4784), .Y(new_n4791));
  OAI21xp33_ASAP7_75t_L     g04535(.A1(new_n4776), .A2(new_n4772), .B(new_n4782), .Y(new_n4792));
  NAND2xp33_ASAP7_75t_L     g04536(.A(new_n4791), .B(new_n4792), .Y(new_n4793));
  NAND2xp33_ASAP7_75t_L     g04537(.A(new_n4790), .B(new_n4793), .Y(new_n4794));
  NOR2xp33_ASAP7_75t_L      g04538(.A(new_n2703), .B(new_n1550), .Y(new_n4795));
  AOI221xp5_ASAP7_75t_L     g04539(.A1(\b[25] ), .A2(new_n713), .B1(\b[27] ), .B2(new_n640), .C(new_n4795), .Y(new_n4796));
  INVx1_ASAP7_75t_L         g04540(.A(new_n4796), .Y(new_n4797));
  A2O1A1Ixp33_ASAP7_75t_L   g04541(.A1(new_n2887), .A2(new_n718), .B(new_n4797), .C(\a[11] ), .Y(new_n4798));
  O2A1O1Ixp33_ASAP7_75t_L   g04542(.A1(new_n641), .A2(new_n2889), .B(new_n4796), .C(\a[11] ), .Y(new_n4799));
  AOI21xp33_ASAP7_75t_L     g04543(.A1(new_n4798), .A2(\a[11] ), .B(new_n4799), .Y(new_n4800));
  NAND3xp33_ASAP7_75t_L     g04544(.A(new_n4789), .B(new_n4794), .C(new_n4800), .Y(new_n4801));
  O2A1O1Ixp33_ASAP7_75t_L   g04545(.A1(new_n4377), .A2(new_n4522), .B(new_n4521), .C(new_n4793), .Y(new_n4802));
  AOI221xp5_ASAP7_75t_L     g04546(.A1(new_n4792), .A2(new_n4791), .B1(new_n4515), .B2(new_n4530), .C(new_n4533), .Y(new_n4803));
  O2A1O1Ixp33_ASAP7_75t_L   g04547(.A1(new_n641), .A2(new_n2889), .B(new_n4796), .C(new_n637), .Y(new_n4804));
  INVx1_ASAP7_75t_L         g04548(.A(new_n4799), .Y(new_n4805));
  OAI21xp33_ASAP7_75t_L     g04549(.A1(new_n637), .A2(new_n4804), .B(new_n4805), .Y(new_n4806));
  OAI21xp33_ASAP7_75t_L     g04550(.A1(new_n4803), .A2(new_n4802), .B(new_n4806), .Y(new_n4807));
  NAND3xp33_ASAP7_75t_L     g04551(.A(new_n4635), .B(new_n4801), .C(new_n4807), .Y(new_n4808));
  A2O1A1O1Ixp25_ASAP7_75t_L g04552(.A1(new_n4283), .A2(new_n4303), .B(new_n4293), .C(new_n4527), .D(new_n4540), .Y(new_n4809));
  NOR3xp33_ASAP7_75t_L      g04553(.A(new_n4802), .B(new_n4803), .C(new_n4806), .Y(new_n4810));
  AOI21xp33_ASAP7_75t_L     g04554(.A1(new_n4789), .A2(new_n4794), .B(new_n4800), .Y(new_n4811));
  OAI21xp33_ASAP7_75t_L     g04555(.A1(new_n4810), .A2(new_n4811), .B(new_n4809), .Y(new_n4812));
  AND2x2_ASAP7_75t_L        g04556(.A(new_n3463), .B(new_n3461), .Y(new_n4813));
  NOR2xp33_ASAP7_75t_L      g04557(.A(new_n3098), .B(new_n513), .Y(new_n4814));
  AOI221xp5_ASAP7_75t_L     g04558(.A1(\b[28] ), .A2(new_n560), .B1(\b[30] ), .B2(new_n475), .C(new_n4814), .Y(new_n4815));
  INVx1_ASAP7_75t_L         g04559(.A(new_n4815), .Y(new_n4816));
  A2O1A1Ixp33_ASAP7_75t_L   g04560(.A1(new_n4813), .A2(new_n483), .B(new_n4816), .C(\a[8] ), .Y(new_n4817));
  O2A1O1Ixp33_ASAP7_75t_L   g04561(.A1(new_n477), .A2(new_n3464), .B(new_n4815), .C(\a[8] ), .Y(new_n4818));
  AOI21xp33_ASAP7_75t_L     g04562(.A1(new_n4817), .A2(\a[8] ), .B(new_n4818), .Y(new_n4819));
  NAND3xp33_ASAP7_75t_L     g04563(.A(new_n4808), .B(new_n4812), .C(new_n4819), .Y(new_n4820));
  NOR3xp33_ASAP7_75t_L      g04564(.A(new_n4809), .B(new_n4810), .C(new_n4811), .Y(new_n4821));
  AOI21xp33_ASAP7_75t_L     g04565(.A1(new_n4807), .A2(new_n4801), .B(new_n4635), .Y(new_n4822));
  AO21x2_ASAP7_75t_L        g04566(.A1(\a[8] ), .A2(new_n4817), .B(new_n4818), .Y(new_n4823));
  OAI21xp33_ASAP7_75t_L     g04567(.A1(new_n4822), .A2(new_n4821), .B(new_n4823), .Y(new_n4824));
  NAND2xp33_ASAP7_75t_L     g04568(.A(new_n4820), .B(new_n4824), .Y(new_n4825));
  O2A1O1Ixp33_ASAP7_75t_L   g04569(.A1(new_n4560), .A2(new_n4633), .B(new_n4558), .C(new_n4825), .Y(new_n4826));
  INVx1_ASAP7_75t_L         g04570(.A(new_n4558), .Y(new_n4827));
  OAI21xp33_ASAP7_75t_L     g04571(.A1(new_n4315), .A2(new_n4330), .B(new_n4556), .Y(new_n4828));
  AOI221xp5_ASAP7_75t_L     g04572(.A1(new_n4824), .A2(new_n4820), .B1(new_n4554), .B2(new_n4828), .C(new_n4827), .Y(new_n4829));
  NOR3xp33_ASAP7_75t_L      g04573(.A(new_n4826), .B(new_n4632), .C(new_n4829), .Y(new_n4830));
  INVx1_ASAP7_75t_L         g04574(.A(new_n4108), .Y(new_n4831));
  NAND2xp33_ASAP7_75t_L     g04575(.A(new_n359), .B(new_n4831), .Y(new_n4832));
  A2O1A1Ixp33_ASAP7_75t_L   g04576(.A1(new_n4832), .A2(new_n4628), .B(new_n4630), .C(new_n4631), .Y(new_n4833));
  AND2x2_ASAP7_75t_L        g04577(.A(new_n4820), .B(new_n4824), .Y(new_n4834));
  A2O1A1Ixp33_ASAP7_75t_L   g04578(.A1(new_n4552), .A2(new_n4557), .B(new_n4561), .C(new_n4834), .Y(new_n4835));
  A2O1A1O1Ixp25_ASAP7_75t_L g04579(.A1(new_n4309), .A2(new_n4311), .B(new_n4368), .C(new_n4554), .D(new_n4827), .Y(new_n4836));
  NAND2xp33_ASAP7_75t_L     g04580(.A(new_n4825), .B(new_n4836), .Y(new_n4837));
  AOI21xp33_ASAP7_75t_L     g04581(.A1(new_n4835), .A2(new_n4837), .B(new_n4833), .Y(new_n4838));
  NOR3xp33_ASAP7_75t_L      g04582(.A(new_n4577), .B(new_n4830), .C(new_n4838), .Y(new_n4839));
  OAI21xp33_ASAP7_75t_L     g04583(.A1(new_n4830), .A2(new_n4838), .B(new_n4577), .Y(new_n4840));
  INVx1_ASAP7_75t_L         g04584(.A(new_n4840), .Y(new_n4841));
  NOR3xp33_ASAP7_75t_L      g04585(.A(new_n4841), .B(new_n4626), .C(new_n4839), .Y(new_n4842));
  INVx1_ASAP7_75t_L         g04586(.A(new_n4577), .Y(new_n4843));
  NOR2xp33_ASAP7_75t_L      g04587(.A(new_n4830), .B(new_n4838), .Y(new_n4844));
  NAND2xp33_ASAP7_75t_L     g04588(.A(new_n4843), .B(new_n4844), .Y(new_n4845));
  NAND3xp33_ASAP7_75t_L     g04589(.A(new_n4845), .B(new_n4626), .C(new_n4840), .Y(new_n4846));
  O2A1O1Ixp33_ASAP7_75t_L   g04590(.A1(new_n4599), .A2(new_n4843), .B(new_n4600), .C(new_n4593), .Y(new_n4847));
  AO21x2_ASAP7_75t_L        g04591(.A1(new_n4604), .A2(new_n4607), .B(new_n4847), .Y(new_n4848));
  INVx1_ASAP7_75t_L         g04592(.A(new_n4848), .Y(new_n4849));
  O2A1O1Ixp33_ASAP7_75t_L   g04593(.A1(new_n4626), .A2(new_n4842), .B(new_n4846), .C(new_n4849), .Y(new_n4850));
  NOR2xp33_ASAP7_75t_L      g04594(.A(new_n257), .B(new_n4624), .Y(new_n4851));
  O2A1O1Ixp33_ASAP7_75t_L   g04595(.A1(new_n279), .A2(new_n4622), .B(new_n4611), .C(\a[2] ), .Y(new_n4852));
  OAI22xp33_ASAP7_75t_L     g04596(.A1(new_n4841), .A2(new_n4839), .B1(new_n4852), .B2(new_n4851), .Y(new_n4853));
  NAND2xp33_ASAP7_75t_L     g04597(.A(new_n4846), .B(new_n4853), .Y(new_n4854));
  NOR2xp33_ASAP7_75t_L      g04598(.A(new_n4854), .B(new_n4848), .Y(new_n4855));
  NOR2xp33_ASAP7_75t_L      g04599(.A(new_n4855), .B(new_n4850), .Y(\f[36] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g04600(.A1(new_n4607), .A2(new_n4604), .B(new_n4847), .C(new_n4854), .D(new_n4842), .Y(new_n4857));
  INVx1_ASAP7_75t_L         g04601(.A(new_n4824), .Y(new_n4858));
  NOR2xp33_ASAP7_75t_L      g04602(.A(new_n3456), .B(new_n513), .Y(new_n4859));
  AOI221xp5_ASAP7_75t_L     g04603(.A1(\b[29] ), .A2(new_n560), .B1(\b[31] ), .B2(new_n475), .C(new_n4859), .Y(new_n4860));
  O2A1O1Ixp33_ASAP7_75t_L   g04604(.A1(new_n477), .A2(new_n3681), .B(new_n4860), .C(new_n466), .Y(new_n4861));
  O2A1O1Ixp33_ASAP7_75t_L   g04605(.A1(new_n477), .A2(new_n3681), .B(new_n4860), .C(\a[8] ), .Y(new_n4862));
  INVx1_ASAP7_75t_L         g04606(.A(new_n4862), .Y(new_n4863));
  OAI21xp33_ASAP7_75t_L     g04607(.A1(new_n466), .A2(new_n4861), .B(new_n4863), .Y(new_n4864));
  NAND2xp33_ASAP7_75t_L     g04608(.A(new_n4794), .B(new_n4789), .Y(new_n4865));
  MAJIxp5_ASAP7_75t_L       g04609(.A(new_n4809), .B(new_n4865), .C(new_n4800), .Y(new_n4866));
  OAI21xp33_ASAP7_75t_L     g04610(.A1(new_n4783), .A2(new_n4790), .B(new_n4792), .Y(new_n4867));
  NOR2xp33_ASAP7_75t_L      g04611(.A(new_n1895), .B(new_n2118), .Y(new_n4868));
  AOI221xp5_ASAP7_75t_L     g04612(.A1(\b[20] ), .A2(new_n1290), .B1(\b[22] ), .B2(new_n1209), .C(new_n4868), .Y(new_n4869));
  O2A1O1Ixp33_ASAP7_75t_L   g04613(.A1(new_n1210), .A2(new_n2522), .B(new_n4869), .C(new_n1206), .Y(new_n4870));
  INVx1_ASAP7_75t_L         g04614(.A(new_n4869), .Y(new_n4871));
  A2O1A1Ixp33_ASAP7_75t_L   g04615(.A1(new_n2056), .A2(new_n1216), .B(new_n4871), .C(new_n1206), .Y(new_n4872));
  OAI21xp33_ASAP7_75t_L     g04616(.A1(new_n1206), .A2(new_n4870), .B(new_n4872), .Y(new_n4873));
  A2O1A1O1Ixp25_ASAP7_75t_L g04617(.A1(new_n4382), .A2(new_n4469), .B(new_n4715), .C(new_n4703), .D(new_n4725), .Y(new_n4874));
  OAI22xp33_ASAP7_75t_L     g04618(.A1(new_n2572), .A2(new_n748), .B1(new_n833), .B2(new_n2410), .Y(new_n4875));
  AOI221xp5_ASAP7_75t_L     g04619(.A1(new_n2423), .A2(\b[13] ), .B1(new_n2417), .B2(new_n1166), .C(new_n4875), .Y(new_n4876));
  XNOR2x2_ASAP7_75t_L       g04620(.A(\a[26] ), .B(new_n4876), .Y(new_n4877));
  A2O1A1O1Ixp25_ASAP7_75t_L g04621(.A1(new_n4390), .A2(new_n4447), .B(new_n4639), .C(new_n4691), .D(new_n4706), .Y(new_n4878));
  NOR2xp33_ASAP7_75t_L      g04622(.A(new_n590), .B(new_n2925), .Y(new_n4879));
  AOI221xp5_ASAP7_75t_L     g04623(.A1(\b[8] ), .A2(new_n3129), .B1(\b[10] ), .B2(new_n2938), .C(new_n4879), .Y(new_n4880));
  O2A1O1Ixp33_ASAP7_75t_L   g04624(.A1(new_n2940), .A2(new_n1175), .B(new_n4880), .C(new_n2928), .Y(new_n4881));
  INVx1_ASAP7_75t_L         g04625(.A(new_n4880), .Y(new_n4882));
  A2O1A1Ixp33_ASAP7_75t_L   g04626(.A1(new_n690), .A2(new_n2932), .B(new_n4882), .C(new_n2928), .Y(new_n4883));
  OAI21xp33_ASAP7_75t_L     g04627(.A1(new_n2928), .A2(new_n4881), .B(new_n4883), .Y(new_n4884));
  A2O1A1Ixp33_ASAP7_75t_L   g04628(.A1(new_n4676), .A2(new_n4677), .B(new_n4422), .C(new_n4670), .Y(new_n4885));
  NOR2xp33_ASAP7_75t_L      g04629(.A(new_n448), .B(new_n3510), .Y(new_n4886));
  AOI221xp5_ASAP7_75t_L     g04630(.A1(\b[5] ), .A2(new_n3708), .B1(\b[6] ), .B2(new_n3499), .C(new_n4886), .Y(new_n4887));
  O2A1O1Ixp33_ASAP7_75t_L   g04631(.A1(new_n3513), .A2(new_n456), .B(new_n4887), .C(new_n3493), .Y(new_n4888));
  OAI21xp33_ASAP7_75t_L     g04632(.A1(new_n3513), .A2(new_n456), .B(new_n4887), .Y(new_n4889));
  NAND2xp33_ASAP7_75t_L     g04633(.A(new_n3493), .B(new_n4889), .Y(new_n4890));
  OAI21xp33_ASAP7_75t_L     g04634(.A1(new_n3493), .A2(new_n4888), .B(new_n4890), .Y(new_n4891));
  INVx1_ASAP7_75t_L         g04635(.A(new_n4891), .Y(new_n4892));
  MAJIxp5_ASAP7_75t_L       g04636(.A(new_n4661), .B(new_n4650), .C(new_n4408), .Y(new_n4893));
  NAND2xp33_ASAP7_75t_L     g04637(.A(\b[3] ), .B(new_n4155), .Y(new_n4894));
  OAI221xp5_ASAP7_75t_L     g04638(.A1(new_n4147), .A2(new_n332), .B1(new_n289), .B2(new_n4397), .C(new_n4894), .Y(new_n4895));
  A2O1A1Ixp33_ASAP7_75t_L   g04639(.A1(new_n342), .A2(new_n4151), .B(new_n4895), .C(\a[35] ), .Y(new_n4896));
  NOR2xp33_ASAP7_75t_L      g04640(.A(new_n332), .B(new_n4147), .Y(new_n4897));
  AOI221xp5_ASAP7_75t_L     g04641(.A1(\b[2] ), .A2(new_n4402), .B1(\b[3] ), .B2(new_n4155), .C(new_n4897), .Y(new_n4898));
  O2A1O1Ixp33_ASAP7_75t_L   g04642(.A1(new_n4150), .A2(new_n1497), .B(new_n4898), .C(\a[35] ), .Y(new_n4899));
  INVx1_ASAP7_75t_L         g04643(.A(\a[37] ), .Y(new_n4900));
  NOR2xp33_ASAP7_75t_L      g04644(.A(\a[36] ), .B(new_n4900), .Y(new_n4901));
  NOR2xp33_ASAP7_75t_L      g04645(.A(\a[37] ), .B(new_n4646), .Y(new_n4902));
  OAI21xp33_ASAP7_75t_L     g04646(.A1(new_n4901), .A2(new_n4902), .B(new_n4649), .Y(new_n4903));
  NAND2xp33_ASAP7_75t_L     g04647(.A(new_n4648), .B(new_n4647), .Y(new_n4904));
  NAND2xp33_ASAP7_75t_L     g04648(.A(\a[38] ), .B(new_n4900), .Y(new_n4905));
  INVx1_ASAP7_75t_L         g04649(.A(\a[38] ), .Y(new_n4906));
  NAND2xp33_ASAP7_75t_L     g04650(.A(\a[37] ), .B(new_n4906), .Y(new_n4907));
  NAND3xp33_ASAP7_75t_L     g04651(.A(new_n4904), .B(new_n4905), .C(new_n4907), .Y(new_n4908));
  OAI22xp33_ASAP7_75t_L     g04652(.A1(new_n4903), .A2(new_n284), .B1(new_n262), .B2(new_n4908), .Y(new_n4909));
  NAND2xp33_ASAP7_75t_L     g04653(.A(new_n4907), .B(new_n4905), .Y(new_n4910));
  NAND2xp33_ASAP7_75t_L     g04654(.A(new_n4910), .B(new_n4904), .Y(new_n4911));
  INVx1_ASAP7_75t_L         g04655(.A(new_n4911), .Y(new_n4912));
  AOI21xp33_ASAP7_75t_L     g04656(.A1(new_n275), .A2(new_n4912), .B(new_n4909), .Y(new_n4913));
  NAND3xp33_ASAP7_75t_L     g04657(.A(new_n4913), .B(new_n4651), .C(\a[38] ), .Y(new_n4914));
  NOR2xp33_ASAP7_75t_L      g04658(.A(new_n4901), .B(new_n4902), .Y(new_n4915));
  NOR2xp33_ASAP7_75t_L      g04659(.A(new_n4904), .B(new_n4915), .Y(new_n4916));
  NOR2xp33_ASAP7_75t_L      g04660(.A(new_n4910), .B(new_n4649), .Y(new_n4917));
  AOI22xp33_ASAP7_75t_L     g04661(.A1(new_n4916), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n4917), .Y(new_n4918));
  O2A1O1Ixp33_ASAP7_75t_L   g04662(.A1(new_n4911), .A2(new_n274), .B(new_n4918), .C(new_n4906), .Y(new_n4919));
  A2O1A1Ixp33_ASAP7_75t_L   g04663(.A1(new_n4912), .A2(new_n275), .B(new_n4909), .C(new_n4906), .Y(new_n4920));
  A2O1A1Ixp33_ASAP7_75t_L   g04664(.A1(new_n4919), .A2(new_n4650), .B(new_n4906), .C(new_n4920), .Y(new_n4921));
  AOI221xp5_ASAP7_75t_L     g04665(.A1(\a[35] ), .A2(new_n4896), .B1(new_n4914), .B2(new_n4921), .C(new_n4899), .Y(new_n4922));
  O2A1O1Ixp33_ASAP7_75t_L   g04666(.A1(new_n4150), .A2(new_n1497), .B(new_n4898), .C(new_n4145), .Y(new_n4923));
  INVx1_ASAP7_75t_L         g04667(.A(new_n4899), .Y(new_n4924));
  NAND2xp33_ASAP7_75t_L     g04668(.A(new_n4914), .B(new_n4921), .Y(new_n4925));
  O2A1O1Ixp33_ASAP7_75t_L   g04669(.A1(new_n4145), .A2(new_n4923), .B(new_n4924), .C(new_n4925), .Y(new_n4926));
  NOR3xp33_ASAP7_75t_L      g04670(.A(new_n4926), .B(new_n4922), .C(new_n4893), .Y(new_n4927));
  MAJIxp5_ASAP7_75t_L       g04671(.A(new_n4668), .B(new_n4428), .C(new_n4651), .Y(new_n4928));
  NAND2xp33_ASAP7_75t_L     g04672(.A(\a[35] ), .B(new_n4896), .Y(new_n4929));
  INVx1_ASAP7_75t_L         g04673(.A(new_n4914), .Y(new_n4930));
  A2O1A1Ixp33_ASAP7_75t_L   g04674(.A1(new_n4912), .A2(new_n275), .B(new_n4909), .C(\a[38] ), .Y(new_n4931));
  INVx1_ASAP7_75t_L         g04675(.A(new_n4920), .Y(new_n4932));
  O2A1O1Ixp33_ASAP7_75t_L   g04676(.A1(new_n4651), .A2(new_n4931), .B(\a[38] ), .C(new_n4932), .Y(new_n4933));
  OAI211xp5_ASAP7_75t_L     g04677(.A1(new_n4930), .A2(new_n4933), .B(new_n4929), .C(new_n4924), .Y(new_n4934));
  NOR2xp33_ASAP7_75t_L      g04678(.A(new_n4145), .B(new_n4923), .Y(new_n4935));
  OAI211xp5_ASAP7_75t_L     g04679(.A1(new_n4899), .A2(new_n4935), .B(new_n4914), .C(new_n4921), .Y(new_n4936));
  AOI21xp33_ASAP7_75t_L     g04680(.A1(new_n4936), .A2(new_n4934), .B(new_n4928), .Y(new_n4937));
  OAI21xp33_ASAP7_75t_L     g04681(.A1(new_n4937), .A2(new_n4927), .B(new_n4892), .Y(new_n4938));
  NAND3xp33_ASAP7_75t_L     g04682(.A(new_n4928), .B(new_n4936), .C(new_n4934), .Y(new_n4939));
  OAI21xp33_ASAP7_75t_L     g04683(.A1(new_n4922), .A2(new_n4926), .B(new_n4893), .Y(new_n4940));
  NAND3xp33_ASAP7_75t_L     g04684(.A(new_n4940), .B(new_n4939), .C(new_n4891), .Y(new_n4941));
  NAND3xp33_ASAP7_75t_L     g04685(.A(new_n4885), .B(new_n4938), .C(new_n4941), .Y(new_n4942));
  AO21x2_ASAP7_75t_L        g04686(.A1(new_n4941), .A2(new_n4938), .B(new_n4885), .Y(new_n4943));
  AOI21xp33_ASAP7_75t_L     g04687(.A1(new_n4943), .A2(new_n4942), .B(new_n4884), .Y(new_n4944));
  AND3x1_ASAP7_75t_L        g04688(.A(new_n4943), .B(new_n4942), .C(new_n4884), .Y(new_n4945));
  OR3x1_ASAP7_75t_L         g04689(.A(new_n4878), .B(new_n4944), .C(new_n4945), .Y(new_n4946));
  OAI21xp33_ASAP7_75t_L     g04690(.A1(new_n4944), .A2(new_n4945), .B(new_n4878), .Y(new_n4947));
  AOI21xp33_ASAP7_75t_L     g04691(.A1(new_n4946), .A2(new_n4947), .B(new_n4877), .Y(new_n4948));
  XNOR2x2_ASAP7_75t_L       g04692(.A(new_n2413), .B(new_n4876), .Y(new_n4949));
  NOR3xp33_ASAP7_75t_L      g04693(.A(new_n4878), .B(new_n4944), .C(new_n4945), .Y(new_n4950));
  AO21x2_ASAP7_75t_L        g04694(.A1(new_n4942), .A2(new_n4943), .B(new_n4884), .Y(new_n4951));
  NAND3xp33_ASAP7_75t_L     g04695(.A(new_n4943), .B(new_n4942), .C(new_n4884), .Y(new_n4952));
  AOI211xp5_ASAP7_75t_L     g04696(.A1(new_n4952), .A2(new_n4951), .B(new_n4706), .C(new_n4696), .Y(new_n4953));
  NOR3xp33_ASAP7_75t_L      g04697(.A(new_n4949), .B(new_n4953), .C(new_n4950), .Y(new_n4954));
  NOR3xp33_ASAP7_75t_L      g04698(.A(new_n4874), .B(new_n4948), .C(new_n4954), .Y(new_n4955));
  INVx1_ASAP7_75t_L         g04699(.A(new_n4955), .Y(new_n4956));
  OAI21xp33_ASAP7_75t_L     g04700(.A1(new_n4948), .A2(new_n4954), .B(new_n4874), .Y(new_n4957));
  OAI22xp33_ASAP7_75t_L     g04701(.A1(new_n2089), .A2(new_n960), .B1(new_n1043), .B2(new_n1962), .Y(new_n4958));
  AOI221xp5_ASAP7_75t_L     g04702(.A1(new_n1955), .A2(\b[16] ), .B1(new_n1964), .B2(new_n1156), .C(new_n4958), .Y(new_n4959));
  XNOR2x2_ASAP7_75t_L       g04703(.A(new_n1952), .B(new_n4959), .Y(new_n4960));
  NAND3xp33_ASAP7_75t_L     g04704(.A(new_n4956), .B(new_n4957), .C(new_n4960), .Y(new_n4961));
  NOR2xp33_ASAP7_75t_L      g04705(.A(new_n4446), .B(new_n4448), .Y(new_n4962));
  A2O1A1Ixp33_ASAP7_75t_L   g04706(.A1(new_n4386), .A2(\a[26] ), .B(new_n4387), .C(new_n4962), .Y(new_n4963));
  A2O1A1Ixp33_ASAP7_75t_L   g04707(.A1(new_n4201), .A2(new_n4381), .B(new_n4450), .C(new_n4963), .Y(new_n4964));
  OAI21xp33_ASAP7_75t_L     g04708(.A1(new_n4950), .A2(new_n4953), .B(new_n4949), .Y(new_n4965));
  NAND3xp33_ASAP7_75t_L     g04709(.A(new_n4877), .B(new_n4946), .C(new_n4947), .Y(new_n4966));
  AOI221xp5_ASAP7_75t_L     g04710(.A1(new_n4964), .A2(new_n4726), .B1(new_n4965), .B2(new_n4966), .C(new_n4725), .Y(new_n4967));
  XNOR2x2_ASAP7_75t_L       g04711(.A(\a[23] ), .B(new_n4959), .Y(new_n4968));
  OAI21xp33_ASAP7_75t_L     g04712(.A1(new_n4967), .A2(new_n4955), .B(new_n4968), .Y(new_n4969));
  NOR2xp33_ASAP7_75t_L      g04713(.A(new_n4716), .B(new_n4714), .Y(new_n4970));
  MAJIxp5_ASAP7_75t_L       g04714(.A(new_n4736), .B(new_n4722), .C(new_n4970), .Y(new_n4971));
  NAND3xp33_ASAP7_75t_L     g04715(.A(new_n4971), .B(new_n4969), .C(new_n4961), .Y(new_n4972));
  NOR3xp33_ASAP7_75t_L      g04716(.A(new_n4968), .B(new_n4967), .C(new_n4955), .Y(new_n4973));
  AOI21xp33_ASAP7_75t_L     g04717(.A1(new_n4956), .A2(new_n4957), .B(new_n4960), .Y(new_n4974));
  XNOR2x2_ASAP7_75t_L       g04718(.A(new_n4713), .B(new_n4728), .Y(new_n4975));
  MAJIxp5_ASAP7_75t_L       g04719(.A(new_n4637), .B(new_n4732), .C(new_n4975), .Y(new_n4976));
  OAI21xp33_ASAP7_75t_L     g04720(.A1(new_n4973), .A2(new_n4974), .B(new_n4976), .Y(new_n4977));
  NOR2xp33_ASAP7_75t_L      g04721(.A(new_n1458), .B(new_n1517), .Y(new_n4978));
  AOI221xp5_ASAP7_75t_L     g04722(.A1(\b[17] ), .A2(new_n1659), .B1(\b[19] ), .B2(new_n1511), .C(new_n4978), .Y(new_n4979));
  INVx1_ASAP7_75t_L         g04723(.A(new_n4979), .Y(new_n4980));
  A2O1A1Ixp33_ASAP7_75t_L   g04724(.A1(new_n1607), .A2(new_n1513), .B(new_n4980), .C(\a[20] ), .Y(new_n4981));
  O2A1O1Ixp33_ASAP7_75t_L   g04725(.A1(new_n1521), .A2(new_n1628), .B(new_n4979), .C(\a[20] ), .Y(new_n4982));
  AOI21xp33_ASAP7_75t_L     g04726(.A1(new_n4981), .A2(\a[20] ), .B(new_n4982), .Y(new_n4983));
  NAND3xp33_ASAP7_75t_L     g04727(.A(new_n4972), .B(new_n4977), .C(new_n4983), .Y(new_n4984));
  AO21x2_ASAP7_75t_L        g04728(.A1(new_n4977), .A2(new_n4972), .B(new_n4983), .Y(new_n4985));
  A2O1A1O1Ixp25_ASAP7_75t_L g04729(.A1(new_n4487), .A2(new_n4489), .B(new_n4636), .C(new_n4752), .D(new_n4764), .Y(new_n4986));
  NAND3xp33_ASAP7_75t_L     g04730(.A(new_n4986), .B(new_n4985), .C(new_n4984), .Y(new_n4987));
  AO21x2_ASAP7_75t_L        g04731(.A1(new_n4984), .A2(new_n4985), .B(new_n4986), .Y(new_n4988));
  NAND3xp33_ASAP7_75t_L     g04732(.A(new_n4988), .B(new_n4987), .C(new_n4873), .Y(new_n4989));
  AND3x1_ASAP7_75t_L        g04733(.A(new_n4986), .B(new_n4985), .C(new_n4984), .Y(new_n4990));
  AOI21xp33_ASAP7_75t_L     g04734(.A1(new_n4985), .A2(new_n4984), .B(new_n4986), .Y(new_n4991));
  NOR3xp33_ASAP7_75t_L      g04735(.A(new_n4990), .B(new_n4991), .C(new_n4873), .Y(new_n4992));
  AOI21xp33_ASAP7_75t_L     g04736(.A1(new_n4989), .A2(new_n4873), .B(new_n4992), .Y(new_n4993));
  NAND2xp33_ASAP7_75t_L     g04737(.A(new_n4763), .B(new_n4767), .Y(new_n4994));
  O2A1O1Ixp33_ASAP7_75t_L   g04738(.A1(new_n4758), .A2(new_n1206), .B(new_n4760), .C(new_n4994), .Y(new_n4995));
  NAND2xp33_ASAP7_75t_L     g04739(.A(new_n4775), .B(new_n4774), .Y(new_n4996));
  O2A1O1Ixp33_ASAP7_75t_L   g04740(.A1(new_n4773), .A2(new_n4499), .B(new_n4996), .C(new_n4995), .Y(new_n4997));
  NAND2xp33_ASAP7_75t_L     g04741(.A(new_n4993), .B(new_n4997), .Y(new_n4998));
  MAJIxp5_ASAP7_75t_L       g04742(.A(new_n4517), .B(new_n4994), .C(new_n4770), .Y(new_n4999));
  A2O1A1Ixp33_ASAP7_75t_L   g04743(.A1(new_n4989), .A2(new_n4873), .B(new_n4992), .C(new_n4999), .Y(new_n5000));
  AND2x2_ASAP7_75t_L        g04744(.A(new_n2384), .B(new_n2382), .Y(new_n5001));
  NAND2xp33_ASAP7_75t_L     g04745(.A(\b[24] ), .B(new_n885), .Y(new_n5002));
  OAI221xp5_ASAP7_75t_L     g04746(.A1(new_n869), .A2(new_n2377), .B1(new_n2188), .B2(new_n980), .C(new_n5002), .Y(new_n5003));
  AOI211xp5_ASAP7_75t_L     g04747(.A1(new_n5001), .A2(new_n873), .B(new_n5003), .C(new_n867), .Y(new_n5004));
  INVx1_ASAP7_75t_L         g04748(.A(new_n5004), .Y(new_n5005));
  A2O1A1Ixp33_ASAP7_75t_L   g04749(.A1(new_n5001), .A2(new_n873), .B(new_n5003), .C(new_n867), .Y(new_n5006));
  NAND2xp33_ASAP7_75t_L     g04750(.A(new_n5006), .B(new_n5005), .Y(new_n5007));
  NAND3xp33_ASAP7_75t_L     g04751(.A(new_n4998), .B(new_n5007), .C(new_n5000), .Y(new_n5008));
  INVx1_ASAP7_75t_L         g04752(.A(new_n5008), .Y(new_n5009));
  AOI21xp33_ASAP7_75t_L     g04753(.A1(new_n4998), .A2(new_n5000), .B(new_n5007), .Y(new_n5010));
  OAI21xp33_ASAP7_75t_L     g04754(.A1(new_n5010), .A2(new_n5009), .B(new_n4867), .Y(new_n5011));
  A2O1A1O1Ixp25_ASAP7_75t_L g04755(.A1(new_n4515), .A2(new_n4530), .B(new_n4533), .C(new_n4791), .D(new_n4787), .Y(new_n5012));
  AO21x2_ASAP7_75t_L        g04756(.A1(new_n5000), .A2(new_n4998), .B(new_n5007), .Y(new_n5013));
  NAND3xp33_ASAP7_75t_L     g04757(.A(new_n5012), .B(new_n5008), .C(new_n5013), .Y(new_n5014));
  NOR2xp33_ASAP7_75t_L      g04758(.A(new_n3079), .B(new_n710), .Y(new_n5015));
  AOI221xp5_ASAP7_75t_L     g04759(.A1(\b[27] ), .A2(new_n635), .B1(\b[26] ), .B2(new_n713), .C(new_n5015), .Y(new_n5016));
  OAI21xp33_ASAP7_75t_L     g04760(.A1(new_n641), .A2(new_n3087), .B(new_n5016), .Y(new_n5017));
  NOR2xp33_ASAP7_75t_L      g04761(.A(new_n637), .B(new_n5017), .Y(new_n5018));
  O2A1O1Ixp33_ASAP7_75t_L   g04762(.A1(new_n641), .A2(new_n3087), .B(new_n5016), .C(\a[11] ), .Y(new_n5019));
  NOR2xp33_ASAP7_75t_L      g04763(.A(new_n5019), .B(new_n5018), .Y(new_n5020));
  NAND3xp33_ASAP7_75t_L     g04764(.A(new_n5020), .B(new_n5011), .C(new_n5014), .Y(new_n5021));
  AOI21xp33_ASAP7_75t_L     g04765(.A1(new_n5008), .A2(new_n5013), .B(new_n5012), .Y(new_n5022));
  OAI21xp33_ASAP7_75t_L     g04766(.A1(new_n4532), .A2(new_n4377), .B(new_n4521), .Y(new_n5023));
  A2O1A1O1Ixp25_ASAP7_75t_L g04767(.A1(new_n5023), .A2(new_n4788), .B(new_n4787), .C(new_n5013), .D(new_n5009), .Y(new_n5024));
  O2A1O1Ixp33_ASAP7_75t_L   g04768(.A1(new_n641), .A2(new_n3087), .B(new_n5016), .C(new_n637), .Y(new_n5025));
  INVx1_ASAP7_75t_L         g04769(.A(new_n5019), .Y(new_n5026));
  OAI21xp33_ASAP7_75t_L     g04770(.A1(new_n637), .A2(new_n5025), .B(new_n5026), .Y(new_n5027));
  A2O1A1Ixp33_ASAP7_75t_L   g04771(.A1(new_n5024), .A2(new_n5013), .B(new_n5022), .C(new_n5027), .Y(new_n5028));
  NAND3xp33_ASAP7_75t_L     g04772(.A(new_n4866), .B(new_n5021), .C(new_n5028), .Y(new_n5029));
  NOR2xp33_ASAP7_75t_L      g04773(.A(new_n4803), .B(new_n4802), .Y(new_n5030));
  MAJIxp5_ASAP7_75t_L       g04774(.A(new_n4635), .B(new_n4806), .C(new_n5030), .Y(new_n5031));
  AND3x1_ASAP7_75t_L        g04775(.A(new_n5020), .B(new_n5011), .C(new_n5014), .Y(new_n5032));
  O2A1O1Ixp33_ASAP7_75t_L   g04776(.A1(new_n4790), .A2(new_n4793), .B(new_n4792), .C(new_n5010), .Y(new_n5033));
  A2O1A1O1Ixp25_ASAP7_75t_L g04777(.A1(new_n5008), .A2(new_n5033), .B(new_n5012), .C(new_n5014), .D(new_n5020), .Y(new_n5034));
  OAI21xp33_ASAP7_75t_L     g04778(.A1(new_n5032), .A2(new_n5034), .B(new_n5031), .Y(new_n5035));
  AOI21xp33_ASAP7_75t_L     g04779(.A1(new_n5029), .A2(new_n5035), .B(new_n4864), .Y(new_n5036));
  INVx1_ASAP7_75t_L         g04780(.A(new_n4861), .Y(new_n5037));
  AOI21xp33_ASAP7_75t_L     g04781(.A1(new_n5037), .A2(\a[8] ), .B(new_n4862), .Y(new_n5038));
  NOR3xp33_ASAP7_75t_L      g04782(.A(new_n5031), .B(new_n5032), .C(new_n5034), .Y(new_n5039));
  AOI21xp33_ASAP7_75t_L     g04783(.A1(new_n5028), .A2(new_n5021), .B(new_n4866), .Y(new_n5040));
  NOR3xp33_ASAP7_75t_L      g04784(.A(new_n5039), .B(new_n5038), .C(new_n5040), .Y(new_n5041));
  NOR2xp33_ASAP7_75t_L      g04785(.A(new_n5036), .B(new_n5041), .Y(new_n5042));
  OAI21xp33_ASAP7_75t_L     g04786(.A1(new_n4858), .A2(new_n4826), .B(new_n5042), .Y(new_n5043));
  A2O1A1O1Ixp25_ASAP7_75t_L g04787(.A1(new_n4554), .A2(new_n4828), .B(new_n4827), .C(new_n4820), .D(new_n4858), .Y(new_n5044));
  OAI21xp33_ASAP7_75t_L     g04788(.A1(new_n5040), .A2(new_n5039), .B(new_n5038), .Y(new_n5045));
  NAND3xp33_ASAP7_75t_L     g04789(.A(new_n5029), .B(new_n4864), .C(new_n5035), .Y(new_n5046));
  NAND2xp33_ASAP7_75t_L     g04790(.A(new_n5046), .B(new_n5045), .Y(new_n5047));
  NAND2xp33_ASAP7_75t_L     g04791(.A(new_n5047), .B(new_n5044), .Y(new_n5048));
  NOR2xp33_ASAP7_75t_L      g04792(.A(new_n3891), .B(new_n375), .Y(new_n5049));
  AOI221xp5_ASAP7_75t_L     g04793(.A1(\b[34] ), .A2(new_n361), .B1(new_n349), .B2(\b[33] ), .C(new_n5049), .Y(new_n5050));
  O2A1O1Ixp33_ASAP7_75t_L   g04794(.A1(new_n356), .A2(new_n4352), .B(new_n5050), .C(new_n346), .Y(new_n5051));
  O2A1O1Ixp33_ASAP7_75t_L   g04795(.A1(new_n356), .A2(new_n4352), .B(new_n5050), .C(\a[5] ), .Y(new_n5052));
  INVx1_ASAP7_75t_L         g04796(.A(new_n5052), .Y(new_n5053));
  OA21x2_ASAP7_75t_L        g04797(.A1(new_n346), .A2(new_n5051), .B(new_n5053), .Y(new_n5054));
  NAND3xp33_ASAP7_75t_L     g04798(.A(new_n5043), .B(new_n5048), .C(new_n5054), .Y(new_n5055));
  NOR2xp33_ASAP7_75t_L      g04799(.A(new_n5047), .B(new_n5044), .Y(new_n5056));
  OAI21xp33_ASAP7_75t_L     g04800(.A1(new_n4560), .A2(new_n4633), .B(new_n4558), .Y(new_n5057));
  AOI221xp5_ASAP7_75t_L     g04801(.A1(new_n5046), .A2(new_n5045), .B1(new_n4834), .B2(new_n5057), .C(new_n4858), .Y(new_n5058));
  OAI21xp33_ASAP7_75t_L     g04802(.A1(new_n346), .A2(new_n5051), .B(new_n5053), .Y(new_n5059));
  OAI21xp33_ASAP7_75t_L     g04803(.A1(new_n5058), .A2(new_n5056), .B(new_n5059), .Y(new_n5060));
  NAND2xp33_ASAP7_75t_L     g04804(.A(new_n5060), .B(new_n5055), .Y(new_n5061));
  A2O1A1Ixp33_ASAP7_75t_L   g04805(.A1(new_n4575), .A2(new_n4323), .B(new_n4338), .C(new_n4568), .Y(new_n5062));
  NAND3xp33_ASAP7_75t_L     g04806(.A(new_n4835), .B(new_n4833), .C(new_n4837), .Y(new_n5063));
  A2O1A1Ixp33_ASAP7_75t_L   g04807(.A1(new_n5062), .A2(new_n4572), .B(new_n4838), .C(new_n5063), .Y(new_n5064));
  NOR2xp33_ASAP7_75t_L      g04808(.A(new_n5064), .B(new_n5061), .Y(new_n5065));
  NAND2xp33_ASAP7_75t_L     g04809(.A(new_n5048), .B(new_n5043), .Y(new_n5066));
  O2A1O1Ixp33_ASAP7_75t_L   g04810(.A1(new_n5051), .A2(new_n346), .B(new_n5053), .C(new_n5066), .Y(new_n5067));
  OAI21xp33_ASAP7_75t_L     g04811(.A1(new_n4829), .A2(new_n4826), .B(new_n4632), .Y(new_n5068));
  A2O1A1O1Ixp25_ASAP7_75t_L g04812(.A1(new_n4568), .A2(new_n4598), .B(new_n4576), .C(new_n5068), .D(new_n4830), .Y(new_n5069));
  O2A1O1Ixp33_ASAP7_75t_L   g04813(.A1(new_n5054), .A2(new_n5067), .B(new_n5055), .C(new_n5069), .Y(new_n5070));
  NOR2xp33_ASAP7_75t_L      g04814(.A(new_n4581), .B(new_n287), .Y(new_n5071));
  AOI221xp5_ASAP7_75t_L     g04815(.A1(\b[36] ), .A2(new_n264), .B1(\b[37] ), .B2(new_n283), .C(new_n5071), .Y(new_n5072));
  NOR2xp33_ASAP7_75t_L      g04816(.A(\b[36] ), .B(\b[37] ), .Y(new_n5073));
  INVx1_ASAP7_75t_L         g04817(.A(\b[37] ), .Y(new_n5074));
  NOR2xp33_ASAP7_75t_L      g04818(.A(new_n4613), .B(new_n5074), .Y(new_n5075));
  NOR2xp33_ASAP7_75t_L      g04819(.A(new_n5073), .B(new_n5075), .Y(new_n5076));
  A2O1A1Ixp33_ASAP7_75t_L   g04820(.A1(new_n4619), .A2(new_n4615), .B(new_n4614), .C(new_n5076), .Y(new_n5077));
  INVx1_ASAP7_75t_L         g04821(.A(new_n4345), .Y(new_n5078));
  A2O1A1Ixp33_ASAP7_75t_L   g04822(.A1(new_n4104), .A2(new_n4342), .B(new_n4347), .C(new_n5078), .Y(new_n5079));
  A2O1A1O1Ixp25_ASAP7_75t_L g04823(.A1(new_n4583), .A2(new_n5079), .B(new_n4582), .C(new_n4615), .D(new_n4614), .Y(new_n5080));
  INVx1_ASAP7_75t_L         g04824(.A(new_n5076), .Y(new_n5081));
  NAND2xp33_ASAP7_75t_L     g04825(.A(new_n5081), .B(new_n5080), .Y(new_n5082));
  NAND2xp33_ASAP7_75t_L     g04826(.A(new_n5077), .B(new_n5082), .Y(new_n5083));
  OAI21xp33_ASAP7_75t_L     g04827(.A1(new_n279), .A2(new_n5083), .B(new_n5072), .Y(new_n5084));
  NOR2xp33_ASAP7_75t_L      g04828(.A(new_n257), .B(new_n5084), .Y(new_n5085));
  O2A1O1Ixp33_ASAP7_75t_L   g04829(.A1(new_n279), .A2(new_n5083), .B(new_n5072), .C(\a[2] ), .Y(new_n5086));
  NOR2xp33_ASAP7_75t_L      g04830(.A(new_n5086), .B(new_n5085), .Y(new_n5087));
  OAI21xp33_ASAP7_75t_L     g04831(.A1(new_n5065), .A2(new_n5070), .B(new_n5087), .Y(new_n5088));
  NOR3xp33_ASAP7_75t_L      g04832(.A(new_n5070), .B(new_n5087), .C(new_n5065), .Y(new_n5089));
  INVx1_ASAP7_75t_L         g04833(.A(new_n5089), .Y(new_n5090));
  NAND2xp33_ASAP7_75t_L     g04834(.A(new_n5088), .B(new_n5090), .Y(new_n5091));
  XOR2x2_ASAP7_75t_L        g04835(.A(new_n4857), .B(new_n5091), .Y(\f[37] ));
  NOR2xp33_ASAP7_75t_L      g04836(.A(new_n5058), .B(new_n5056), .Y(new_n5093));
  MAJIxp5_ASAP7_75t_L       g04837(.A(new_n5064), .B(new_n5093), .C(new_n5059), .Y(new_n5094));
  NOR2xp33_ASAP7_75t_L      g04838(.A(new_n4101), .B(new_n375), .Y(new_n5095));
  AOI221xp5_ASAP7_75t_L     g04839(.A1(\b[35] ), .A2(new_n361), .B1(new_n349), .B2(\b[34] ), .C(new_n5095), .Y(new_n5096));
  O2A1O1Ixp33_ASAP7_75t_L   g04840(.A1(new_n356), .A2(new_n4589), .B(new_n5096), .C(new_n346), .Y(new_n5097));
  INVx1_ASAP7_75t_L         g04841(.A(new_n5097), .Y(new_n5098));
  O2A1O1Ixp33_ASAP7_75t_L   g04842(.A1(new_n356), .A2(new_n4589), .B(new_n5096), .C(\a[5] ), .Y(new_n5099));
  AOI21xp33_ASAP7_75t_L     g04843(.A1(new_n5098), .A2(\a[5] ), .B(new_n5099), .Y(new_n5100));
  INVx1_ASAP7_75t_L         g04844(.A(new_n5100), .Y(new_n5101));
  A2O1A1Ixp33_ASAP7_75t_L   g04845(.A1(new_n4570), .A2(new_n4558), .B(new_n4825), .C(new_n4824), .Y(new_n5102));
  NOR2xp33_ASAP7_75t_L      g04846(.A(new_n3674), .B(new_n513), .Y(new_n5103));
  AOI221xp5_ASAP7_75t_L     g04847(.A1(\b[30] ), .A2(new_n560), .B1(\b[32] ), .B2(new_n475), .C(new_n5103), .Y(new_n5104));
  O2A1O1Ixp33_ASAP7_75t_L   g04848(.A1(new_n477), .A2(new_n3897), .B(new_n5104), .C(new_n466), .Y(new_n5105));
  INVx1_ASAP7_75t_L         g04849(.A(new_n5104), .Y(new_n5106));
  A2O1A1Ixp33_ASAP7_75t_L   g04850(.A1(new_n3900), .A2(new_n483), .B(new_n5106), .C(new_n466), .Y(new_n5107));
  OAI21xp33_ASAP7_75t_L     g04851(.A1(new_n466), .A2(new_n5105), .B(new_n5107), .Y(new_n5108));
  A2O1A1Ixp33_ASAP7_75t_L   g04852(.A1(\a[11] ), .A2(new_n4798), .B(new_n4799), .C(new_n5030), .Y(new_n5109));
  OAI21xp33_ASAP7_75t_L     g04853(.A1(new_n4810), .A2(new_n4811), .B(new_n4635), .Y(new_n5110));
  A2O1A1Ixp33_ASAP7_75t_L   g04854(.A1(new_n5110), .A2(new_n5109), .B(new_n5032), .C(new_n5028), .Y(new_n5111));
  NOR2xp33_ASAP7_75t_L      g04855(.A(new_n3079), .B(new_n1550), .Y(new_n5112));
  AOI221xp5_ASAP7_75t_L     g04856(.A1(\b[27] ), .A2(new_n713), .B1(\b[29] ), .B2(new_n640), .C(new_n5112), .Y(new_n5113));
  O2A1O1Ixp33_ASAP7_75t_L   g04857(.A1(new_n641), .A2(new_n3104), .B(new_n5113), .C(new_n637), .Y(new_n5114));
  INVx1_ASAP7_75t_L         g04858(.A(new_n5113), .Y(new_n5115));
  A2O1A1Ixp33_ASAP7_75t_L   g04859(.A1(new_n3873), .A2(new_n718), .B(new_n5115), .C(new_n637), .Y(new_n5116));
  OAI21xp33_ASAP7_75t_L     g04860(.A1(new_n637), .A2(new_n5114), .B(new_n5116), .Y(new_n5117));
  INVx1_ASAP7_75t_L         g04861(.A(new_n4989), .Y(new_n5118));
  NOR2xp33_ASAP7_75t_L      g04862(.A(new_n4753), .B(new_n4755), .Y(new_n5119));
  A2O1A1Ixp33_ASAP7_75t_L   g04863(.A1(\a[17] ), .A2(new_n4769), .B(new_n4759), .C(new_n5119), .Y(new_n5120));
  A2O1A1Ixp33_ASAP7_75t_L   g04864(.A1(new_n2056), .A2(new_n1216), .B(new_n4871), .C(\a[17] ), .Y(new_n5121));
  NAND2xp33_ASAP7_75t_L     g04865(.A(\a[17] ), .B(new_n5121), .Y(new_n5122));
  NAND4xp25_ASAP7_75t_L     g04866(.A(new_n4988), .B(new_n5122), .C(new_n4872), .D(new_n4987), .Y(new_n5123));
  OAI21xp33_ASAP7_75t_L     g04867(.A1(new_n4991), .A2(new_n4990), .B(new_n4873), .Y(new_n5124));
  OAI22xp33_ASAP7_75t_L     g04868(.A1(new_n4773), .A2(new_n4499), .B1(new_n4771), .B2(new_n4762), .Y(new_n5125));
  AOI22xp33_ASAP7_75t_L     g04869(.A1(new_n5124), .A2(new_n5123), .B1(new_n5120), .B2(new_n5125), .Y(new_n5126));
  OAI21xp33_ASAP7_75t_L     g04870(.A1(new_n4948), .A2(new_n4874), .B(new_n4966), .Y(new_n5127));
  OAI21xp33_ASAP7_75t_L     g04871(.A1(new_n4944), .A2(new_n4878), .B(new_n4952), .Y(new_n5128));
  NOR2xp33_ASAP7_75t_L      g04872(.A(new_n680), .B(new_n2925), .Y(new_n5129));
  AOI221xp5_ASAP7_75t_L     g04873(.A1(\b[9] ), .A2(new_n3129), .B1(\b[11] ), .B2(new_n2938), .C(new_n5129), .Y(new_n5130));
  O2A1O1Ixp33_ASAP7_75t_L   g04874(.A1(new_n2940), .A2(new_n754), .B(new_n5130), .C(new_n2928), .Y(new_n5131));
  O2A1O1Ixp33_ASAP7_75t_L   g04875(.A1(new_n2940), .A2(new_n754), .B(new_n5130), .C(\a[29] ), .Y(new_n5132));
  INVx1_ASAP7_75t_L         g04876(.A(new_n5132), .Y(new_n5133));
  OAI21xp33_ASAP7_75t_L     g04877(.A1(new_n2928), .A2(new_n5131), .B(new_n5133), .Y(new_n5134));
  NOR3xp33_ASAP7_75t_L      g04878(.A(new_n4892), .B(new_n4927), .C(new_n4937), .Y(new_n5135));
  AOI21xp33_ASAP7_75t_L     g04879(.A1(new_n4885), .A2(new_n4938), .B(new_n5135), .Y(new_n5136));
  OAI21xp33_ASAP7_75t_L     g04880(.A1(new_n4922), .A2(new_n4893), .B(new_n4936), .Y(new_n5137));
  NOR2xp33_ASAP7_75t_L      g04881(.A(new_n289), .B(new_n4908), .Y(new_n5138));
  AND3x1_ASAP7_75t_L        g04882(.A(new_n4649), .B(new_n4910), .C(new_n4915), .Y(new_n5139));
  AOI221xp5_ASAP7_75t_L     g04883(.A1(new_n4916), .A2(\b[1] ), .B1(new_n5139), .B2(\b[0] ), .C(new_n5138), .Y(new_n5140));
  NOR2xp33_ASAP7_75t_L      g04884(.A(new_n4911), .B(new_n509), .Y(new_n5141));
  INVx1_ASAP7_75t_L         g04885(.A(new_n5141), .Y(new_n5142));
  NAND3xp33_ASAP7_75t_L     g04886(.A(new_n5140), .B(\a[38] ), .C(new_n5142), .Y(new_n5143));
  NAND3xp33_ASAP7_75t_L     g04887(.A(new_n4649), .B(new_n4915), .C(new_n4910), .Y(new_n5144));
  NAND2xp33_ASAP7_75t_L     g04888(.A(\b[1] ), .B(new_n4916), .Y(new_n5145));
  OAI221xp5_ASAP7_75t_L     g04889(.A1(new_n4908), .A2(new_n289), .B1(new_n284), .B2(new_n5144), .C(new_n5145), .Y(new_n5146));
  A2O1A1Ixp33_ASAP7_75t_L   g04890(.A1(new_n294), .A2(new_n4912), .B(new_n5146), .C(new_n4906), .Y(new_n5147));
  NAND3xp33_ASAP7_75t_L     g04891(.A(new_n4914), .B(new_n5143), .C(new_n5147), .Y(new_n5148));
  NAND5xp2_ASAP7_75t_L      g04892(.A(\a[38] ), .B(new_n4913), .C(new_n5140), .D(new_n5142), .E(new_n4651), .Y(new_n5149));
  NOR2xp33_ASAP7_75t_L      g04893(.A(new_n332), .B(new_n4142), .Y(new_n5150));
  AOI221xp5_ASAP7_75t_L     g04894(.A1(\b[3] ), .A2(new_n4402), .B1(\b[5] ), .B2(new_n4156), .C(new_n5150), .Y(new_n5151));
  OAI211xp5_ASAP7_75t_L     g04895(.A1(new_n728), .A2(new_n4150), .B(new_n5151), .C(\a[35] ), .Y(new_n5152));
  O2A1O1Ixp33_ASAP7_75t_L   g04896(.A1(new_n728), .A2(new_n4150), .B(new_n5151), .C(\a[35] ), .Y(new_n5153));
  INVx1_ASAP7_75t_L         g04897(.A(new_n5153), .Y(new_n5154));
  NAND4xp25_ASAP7_75t_L     g04898(.A(new_n5148), .B(new_n5154), .C(new_n5152), .D(new_n5149), .Y(new_n5155));
  AOI22xp33_ASAP7_75t_L     g04899(.A1(new_n5152), .A2(new_n5154), .B1(new_n5149), .B2(new_n5148), .Y(new_n5156));
  INVx1_ASAP7_75t_L         g04900(.A(new_n5156), .Y(new_n5157));
  NAND3xp33_ASAP7_75t_L     g04901(.A(new_n5137), .B(new_n5155), .C(new_n5157), .Y(new_n5158));
  A2O1A1Ixp33_ASAP7_75t_L   g04902(.A1(new_n294), .A2(new_n4912), .B(new_n5146), .C(\a[38] ), .Y(new_n5159));
  O2A1O1Ixp33_ASAP7_75t_L   g04903(.A1(new_n509), .A2(new_n4911), .B(new_n5140), .C(\a[38] ), .Y(new_n5160));
  A2O1A1O1Ixp25_ASAP7_75t_L g04904(.A1(new_n4913), .A2(new_n4651), .B(new_n5159), .C(\a[38] ), .D(new_n5160), .Y(new_n5161));
  OAI21xp33_ASAP7_75t_L     g04905(.A1(new_n4911), .A2(new_n274), .B(new_n4918), .Y(new_n5162));
  NOR5xp2_ASAP7_75t_L       g04906(.A(new_n5162), .B(new_n5146), .C(new_n5141), .D(new_n4650), .E(new_n4906), .Y(new_n5163));
  NAND2xp33_ASAP7_75t_L     g04907(.A(new_n4151), .B(new_n394), .Y(new_n5164));
  O2A1O1Ixp33_ASAP7_75t_L   g04908(.A1(new_n728), .A2(new_n4150), .B(new_n5151), .C(new_n4145), .Y(new_n5165));
  A2O1A1Ixp33_ASAP7_75t_L   g04909(.A1(new_n5164), .A2(new_n5151), .B(new_n5165), .C(new_n5152), .Y(new_n5166));
  NOR3xp33_ASAP7_75t_L      g04910(.A(new_n5166), .B(new_n5161), .C(new_n5163), .Y(new_n5167));
  OAI221xp5_ASAP7_75t_L     g04911(.A1(new_n4922), .A2(new_n4893), .B1(new_n5156), .B2(new_n5167), .C(new_n4936), .Y(new_n5168));
  NOR2xp33_ASAP7_75t_L      g04912(.A(new_n448), .B(new_n3509), .Y(new_n5169));
  AOI221xp5_ASAP7_75t_L     g04913(.A1(\b[6] ), .A2(new_n3708), .B1(\b[8] ), .B2(new_n3503), .C(new_n5169), .Y(new_n5170));
  INVx1_ASAP7_75t_L         g04914(.A(new_n5170), .Y(new_n5171));
  A2O1A1Ixp33_ASAP7_75t_L   g04915(.A1(new_n1684), .A2(new_n3505), .B(new_n5171), .C(\a[32] ), .Y(new_n5172));
  O2A1O1Ixp33_ASAP7_75t_L   g04916(.A1(new_n3513), .A2(new_n540), .B(new_n5170), .C(\a[32] ), .Y(new_n5173));
  AOI21xp33_ASAP7_75t_L     g04917(.A1(new_n5172), .A2(\a[32] ), .B(new_n5173), .Y(new_n5174));
  AOI21xp33_ASAP7_75t_L     g04918(.A1(new_n5158), .A2(new_n5168), .B(new_n5174), .Y(new_n5175));
  AND3x1_ASAP7_75t_L        g04919(.A(new_n5158), .B(new_n5174), .C(new_n5168), .Y(new_n5176));
  NOR3xp33_ASAP7_75t_L      g04920(.A(new_n5136), .B(new_n5175), .C(new_n5176), .Y(new_n5177));
  AO21x2_ASAP7_75t_L        g04921(.A1(new_n4938), .A2(new_n4885), .B(new_n5135), .Y(new_n5178));
  NOR2xp33_ASAP7_75t_L      g04922(.A(new_n5175), .B(new_n5176), .Y(new_n5179));
  NOR2xp33_ASAP7_75t_L      g04923(.A(new_n5178), .B(new_n5179), .Y(new_n5180));
  OAI21xp33_ASAP7_75t_L     g04924(.A1(new_n5177), .A2(new_n5180), .B(new_n5134), .Y(new_n5181));
  INVx1_ASAP7_75t_L         g04925(.A(new_n5131), .Y(new_n5182));
  AOI21xp33_ASAP7_75t_L     g04926(.A1(new_n5182), .A2(\a[29] ), .B(new_n5132), .Y(new_n5183));
  NAND2xp33_ASAP7_75t_L     g04927(.A(new_n5178), .B(new_n5179), .Y(new_n5184));
  OAI21xp33_ASAP7_75t_L     g04928(.A1(new_n5175), .A2(new_n5176), .B(new_n5136), .Y(new_n5185));
  NAND3xp33_ASAP7_75t_L     g04929(.A(new_n5184), .B(new_n5183), .C(new_n5185), .Y(new_n5186));
  NAND3xp33_ASAP7_75t_L     g04930(.A(new_n5128), .B(new_n5181), .C(new_n5186), .Y(new_n5187));
  A2O1A1Ixp33_ASAP7_75t_L   g04931(.A1(new_n4439), .A2(new_n4438), .B(new_n4436), .C(new_n4423), .Y(new_n5188));
  A2O1A1O1Ixp25_ASAP7_75t_L g04932(.A1(new_n4708), .A2(new_n5188), .B(new_n4706), .C(new_n4951), .D(new_n4945), .Y(new_n5189));
  AOI21xp33_ASAP7_75t_L     g04933(.A1(new_n5184), .A2(new_n5185), .B(new_n5183), .Y(new_n5190));
  NOR3xp33_ASAP7_75t_L      g04934(.A(new_n5180), .B(new_n5177), .C(new_n5134), .Y(new_n5191));
  OAI21xp33_ASAP7_75t_L     g04935(.A1(new_n5190), .A2(new_n5191), .B(new_n5189), .Y(new_n5192));
  NOR2xp33_ASAP7_75t_L      g04936(.A(new_n936), .B(new_n2410), .Y(new_n5193));
  AOI221xp5_ASAP7_75t_L     g04937(.A1(\b[12] ), .A2(new_n2577), .B1(\b[14] ), .B2(new_n2423), .C(new_n5193), .Y(new_n5194));
  INVx1_ASAP7_75t_L         g04938(.A(new_n5194), .Y(new_n5195));
  A2O1A1Ixp33_ASAP7_75t_L   g04939(.A1(new_n971), .A2(new_n2417), .B(new_n5195), .C(\a[26] ), .Y(new_n5196));
  O2A1O1Ixp33_ASAP7_75t_L   g04940(.A1(new_n2425), .A2(new_n1268), .B(new_n5194), .C(\a[26] ), .Y(new_n5197));
  AOI21xp33_ASAP7_75t_L     g04941(.A1(new_n5196), .A2(\a[26] ), .B(new_n5197), .Y(new_n5198));
  NAND3xp33_ASAP7_75t_L     g04942(.A(new_n5187), .B(new_n5198), .C(new_n5192), .Y(new_n5199));
  OAI21xp33_ASAP7_75t_L     g04943(.A1(new_n5190), .A2(new_n5191), .B(new_n5128), .Y(new_n5200));
  AOI21xp33_ASAP7_75t_L     g04944(.A1(new_n5186), .A2(new_n5181), .B(new_n5128), .Y(new_n5201));
  O2A1O1Ixp33_ASAP7_75t_L   g04945(.A1(new_n2425), .A2(new_n1268), .B(new_n5194), .C(new_n2413), .Y(new_n5202));
  A2O1A1Ixp33_ASAP7_75t_L   g04946(.A1(new_n971), .A2(new_n2417), .B(new_n5195), .C(new_n2413), .Y(new_n5203));
  OAI21xp33_ASAP7_75t_L     g04947(.A1(new_n2413), .A2(new_n5202), .B(new_n5203), .Y(new_n5204));
  A2O1A1Ixp33_ASAP7_75t_L   g04948(.A1(new_n5200), .A2(new_n5128), .B(new_n5201), .C(new_n5204), .Y(new_n5205));
  NAND3xp33_ASAP7_75t_L     g04949(.A(new_n5127), .B(new_n5199), .C(new_n5205), .Y(new_n5206));
  A2O1A1O1Ixp25_ASAP7_75t_L g04950(.A1(new_n4726), .A2(new_n4964), .B(new_n4725), .C(new_n4965), .D(new_n4954), .Y(new_n5207));
  NAND2xp33_ASAP7_75t_L     g04951(.A(new_n5199), .B(new_n5205), .Y(new_n5208));
  NAND2xp33_ASAP7_75t_L     g04952(.A(new_n5208), .B(new_n5207), .Y(new_n5209));
  NOR2xp33_ASAP7_75t_L      g04953(.A(new_n1150), .B(new_n1962), .Y(new_n5210));
  AOI221xp5_ASAP7_75t_L     g04954(.A1(new_n1955), .A2(\b[17] ), .B1(new_n2093), .B2(\b[15] ), .C(new_n5210), .Y(new_n5211));
  INVx1_ASAP7_75t_L         g04955(.A(new_n5211), .Y(new_n5212));
  A2O1A1Ixp33_ASAP7_75t_L   g04956(.A1(new_n1633), .A2(new_n1964), .B(new_n5212), .C(\a[23] ), .Y(new_n5213));
  O2A1O1Ixp33_ASAP7_75t_L   g04957(.A1(new_n1956), .A2(new_n1356), .B(new_n5211), .C(\a[23] ), .Y(new_n5214));
  AOI21xp33_ASAP7_75t_L     g04958(.A1(new_n5213), .A2(\a[23] ), .B(new_n5214), .Y(new_n5215));
  NAND3xp33_ASAP7_75t_L     g04959(.A(new_n5209), .B(new_n5206), .C(new_n5215), .Y(new_n5216));
  NOR2xp33_ASAP7_75t_L      g04960(.A(new_n5208), .B(new_n5207), .Y(new_n5217));
  AOI21xp33_ASAP7_75t_L     g04961(.A1(new_n5205), .A2(new_n5199), .B(new_n5127), .Y(new_n5218));
  INVx1_ASAP7_75t_L         g04962(.A(new_n5215), .Y(new_n5219));
  OAI21xp33_ASAP7_75t_L     g04963(.A1(new_n5218), .A2(new_n5217), .B(new_n5219), .Y(new_n5220));
  NAND2xp33_ASAP7_75t_L     g04964(.A(new_n5216), .B(new_n5220), .Y(new_n5221));
  NOR2xp33_ASAP7_75t_L      g04965(.A(new_n4955), .B(new_n4967), .Y(new_n5222));
  NAND2xp33_ASAP7_75t_L     g04966(.A(new_n4968), .B(new_n5222), .Y(new_n5223));
  A2O1A1Ixp33_ASAP7_75t_L   g04967(.A1(new_n4960), .A2(new_n4961), .B(new_n4971), .C(new_n5223), .Y(new_n5224));
  NOR2xp33_ASAP7_75t_L      g04968(.A(new_n5224), .B(new_n5221), .Y(new_n5225));
  NOR3xp33_ASAP7_75t_L      g04969(.A(new_n4960), .B(new_n4967), .C(new_n4955), .Y(new_n5226));
  O2A1O1Ixp33_ASAP7_75t_L   g04970(.A1(new_n4973), .A2(new_n4968), .B(new_n4976), .C(new_n5226), .Y(new_n5227));
  AOI21xp33_ASAP7_75t_L     g04971(.A1(new_n5220), .A2(new_n5216), .B(new_n5227), .Y(new_n5228));
  NOR2xp33_ASAP7_75t_L      g04972(.A(new_n1745), .B(new_n1518), .Y(new_n5229));
  AOI221xp5_ASAP7_75t_L     g04973(.A1(\b[18] ), .A2(new_n1659), .B1(\b[19] ), .B2(new_n1507), .C(new_n5229), .Y(new_n5230));
  O2A1O1Ixp33_ASAP7_75t_L   g04974(.A1(new_n1521), .A2(new_n1754), .B(new_n5230), .C(new_n1501), .Y(new_n5231));
  OAI21xp33_ASAP7_75t_L     g04975(.A1(new_n1521), .A2(new_n1754), .B(new_n5230), .Y(new_n5232));
  NAND2xp33_ASAP7_75t_L     g04976(.A(new_n1501), .B(new_n5232), .Y(new_n5233));
  OAI21xp33_ASAP7_75t_L     g04977(.A1(new_n1501), .A2(new_n5231), .B(new_n5233), .Y(new_n5234));
  NOR3xp33_ASAP7_75t_L      g04978(.A(new_n5225), .B(new_n5228), .C(new_n5234), .Y(new_n5235));
  OA21x2_ASAP7_75t_L        g04979(.A1(new_n5228), .A2(new_n5225), .B(new_n5234), .Y(new_n5236));
  NAND2xp33_ASAP7_75t_L     g04980(.A(new_n4977), .B(new_n4972), .Y(new_n5237));
  MAJIxp5_ASAP7_75t_L       g04981(.A(new_n4986), .B(new_n5237), .C(new_n4983), .Y(new_n5238));
  NOR3xp33_ASAP7_75t_L      g04982(.A(new_n5238), .B(new_n5236), .C(new_n5235), .Y(new_n5239));
  OA21x2_ASAP7_75t_L        g04983(.A1(new_n5235), .A2(new_n5236), .B(new_n5238), .Y(new_n5240));
  NOR2xp33_ASAP7_75t_L      g04984(.A(new_n2188), .B(new_n1284), .Y(new_n5241));
  AOI221xp5_ASAP7_75t_L     g04985(.A1(\b[21] ), .A2(new_n1290), .B1(\b[22] ), .B2(new_n1204), .C(new_n5241), .Y(new_n5242));
  OAI21xp33_ASAP7_75t_L     g04986(.A1(new_n1210), .A2(new_n2194), .B(new_n5242), .Y(new_n5243));
  NOR2xp33_ASAP7_75t_L      g04987(.A(new_n1206), .B(new_n5243), .Y(new_n5244));
  O2A1O1Ixp33_ASAP7_75t_L   g04988(.A1(new_n1210), .A2(new_n2194), .B(new_n5242), .C(\a[17] ), .Y(new_n5245));
  NOR2xp33_ASAP7_75t_L      g04989(.A(new_n5245), .B(new_n5244), .Y(new_n5246));
  NOR3xp33_ASAP7_75t_L      g04990(.A(new_n5240), .B(new_n5246), .C(new_n5239), .Y(new_n5247));
  INVx1_ASAP7_75t_L         g04991(.A(new_n5237), .Y(new_n5248));
  A2O1A1Ixp33_ASAP7_75t_L   g04992(.A1(\a[20] ), .A2(new_n4981), .B(new_n4982), .C(new_n5248), .Y(new_n5249));
  INVx1_ASAP7_75t_L         g04993(.A(new_n5235), .Y(new_n5250));
  OAI21xp33_ASAP7_75t_L     g04994(.A1(new_n5228), .A2(new_n5225), .B(new_n5234), .Y(new_n5251));
  NAND4xp25_ASAP7_75t_L     g04995(.A(new_n5250), .B(new_n4988), .C(new_n5249), .D(new_n5251), .Y(new_n5252));
  OAI21xp33_ASAP7_75t_L     g04996(.A1(new_n5235), .A2(new_n5236), .B(new_n5238), .Y(new_n5253));
  O2A1O1Ixp33_ASAP7_75t_L   g04997(.A1(new_n1210), .A2(new_n2194), .B(new_n5242), .C(new_n1206), .Y(new_n5254));
  INVx1_ASAP7_75t_L         g04998(.A(new_n5245), .Y(new_n5255));
  OAI21xp33_ASAP7_75t_L     g04999(.A1(new_n1206), .A2(new_n5254), .B(new_n5255), .Y(new_n5256));
  AOI21xp33_ASAP7_75t_L     g05000(.A1(new_n5252), .A2(new_n5253), .B(new_n5256), .Y(new_n5257));
  OAI22xp33_ASAP7_75t_L     g05001(.A1(new_n5126), .A2(new_n5118), .B1(new_n5257), .B2(new_n5247), .Y(new_n5258));
  NAND3xp33_ASAP7_75t_L     g05002(.A(new_n5252), .B(new_n5256), .C(new_n5253), .Y(new_n5259));
  OAI21xp33_ASAP7_75t_L     g05003(.A1(new_n5239), .A2(new_n5240), .B(new_n5246), .Y(new_n5260));
  NAND4xp25_ASAP7_75t_L     g05004(.A(new_n5000), .B(new_n5259), .C(new_n5260), .D(new_n4989), .Y(new_n5261));
  NOR2xp33_ASAP7_75t_L      g05005(.A(new_n2703), .B(new_n869), .Y(new_n5262));
  AOI221xp5_ASAP7_75t_L     g05006(.A1(\b[24] ), .A2(new_n985), .B1(\b[25] ), .B2(new_n885), .C(new_n5262), .Y(new_n5263));
  O2A1O1Ixp33_ASAP7_75t_L   g05007(.A1(new_n872), .A2(new_n2708), .B(new_n5263), .C(new_n867), .Y(new_n5264));
  NOR2xp33_ASAP7_75t_L      g05008(.A(new_n867), .B(new_n5264), .Y(new_n5265));
  O2A1O1Ixp33_ASAP7_75t_L   g05009(.A1(new_n872), .A2(new_n2708), .B(new_n5263), .C(\a[14] ), .Y(new_n5266));
  NOR2xp33_ASAP7_75t_L      g05010(.A(new_n5266), .B(new_n5265), .Y(new_n5267));
  NAND3xp33_ASAP7_75t_L     g05011(.A(new_n5261), .B(new_n5258), .C(new_n5267), .Y(new_n5268));
  AO21x2_ASAP7_75t_L        g05012(.A1(new_n5258), .A2(new_n5261), .B(new_n5267), .Y(new_n5269));
  OAI211xp5_ASAP7_75t_L     g05013(.A1(new_n5009), .A2(new_n5033), .B(new_n5268), .C(new_n5269), .Y(new_n5270));
  A2O1A1Ixp33_ASAP7_75t_L   g05014(.A1(new_n5023), .A2(new_n4788), .B(new_n4787), .C(new_n5013), .Y(new_n5271));
  AND3x1_ASAP7_75t_L        g05015(.A(new_n5261), .B(new_n5258), .C(new_n5267), .Y(new_n5272));
  AOI21xp33_ASAP7_75t_L     g05016(.A1(new_n5261), .A2(new_n5258), .B(new_n5267), .Y(new_n5273));
  OAI211xp5_ASAP7_75t_L     g05017(.A1(new_n5273), .A2(new_n5272), .B(new_n5271), .C(new_n5008), .Y(new_n5274));
  AO21x2_ASAP7_75t_L        g05018(.A1(new_n5270), .A2(new_n5274), .B(new_n5117), .Y(new_n5275));
  AND3x1_ASAP7_75t_L        g05019(.A(new_n5274), .B(new_n5270), .C(new_n5117), .Y(new_n5276));
  INVx1_ASAP7_75t_L         g05020(.A(new_n5276), .Y(new_n5277));
  NAND3xp33_ASAP7_75t_L     g05021(.A(new_n5111), .B(new_n5277), .C(new_n5275), .Y(new_n5278));
  O2A1O1Ixp33_ASAP7_75t_L   g05022(.A1(new_n4804), .A2(new_n637), .B(new_n4805), .C(new_n4865), .Y(new_n5279));
  NAND2xp33_ASAP7_75t_L     g05023(.A(new_n4807), .B(new_n4801), .Y(new_n5280));
  A2O1A1O1Ixp25_ASAP7_75t_L g05024(.A1(new_n4635), .A2(new_n5280), .B(new_n5279), .C(new_n5021), .D(new_n5034), .Y(new_n5281));
  AOI21xp33_ASAP7_75t_L     g05025(.A1(new_n5274), .A2(new_n5270), .B(new_n5117), .Y(new_n5282));
  OAI21xp33_ASAP7_75t_L     g05026(.A1(new_n5282), .A2(new_n5276), .B(new_n5281), .Y(new_n5283));
  AOI21xp33_ASAP7_75t_L     g05027(.A1(new_n5278), .A2(new_n5283), .B(new_n5108), .Y(new_n5284));
  INVx1_ASAP7_75t_L         g05028(.A(new_n5108), .Y(new_n5285));
  NOR3xp33_ASAP7_75t_L      g05029(.A(new_n5281), .B(new_n5282), .C(new_n5276), .Y(new_n5286));
  AOI21xp33_ASAP7_75t_L     g05030(.A1(new_n5277), .A2(new_n5275), .B(new_n5111), .Y(new_n5287));
  NOR3xp33_ASAP7_75t_L      g05031(.A(new_n5287), .B(new_n5285), .C(new_n5286), .Y(new_n5288));
  NOR2xp33_ASAP7_75t_L      g05032(.A(new_n5284), .B(new_n5288), .Y(new_n5289));
  A2O1A1Ixp33_ASAP7_75t_L   g05033(.A1(new_n5042), .A2(new_n5102), .B(new_n5041), .C(new_n5289), .Y(new_n5290));
  A2O1A1O1Ixp25_ASAP7_75t_L g05034(.A1(new_n4834), .A2(new_n5057), .B(new_n4858), .C(new_n5045), .D(new_n5041), .Y(new_n5291));
  OAI21xp33_ASAP7_75t_L     g05035(.A1(new_n5286), .A2(new_n5287), .B(new_n5285), .Y(new_n5292));
  NAND3xp33_ASAP7_75t_L     g05036(.A(new_n5278), .B(new_n5108), .C(new_n5283), .Y(new_n5293));
  NAND2xp33_ASAP7_75t_L     g05037(.A(new_n5293), .B(new_n5292), .Y(new_n5294));
  NAND2xp33_ASAP7_75t_L     g05038(.A(new_n5294), .B(new_n5291), .Y(new_n5295));
  AOI21xp33_ASAP7_75t_L     g05039(.A1(new_n5290), .A2(new_n5295), .B(new_n5101), .Y(new_n5296));
  O2A1O1Ixp33_ASAP7_75t_L   g05040(.A1(new_n5044), .A2(new_n5047), .B(new_n5046), .C(new_n5294), .Y(new_n5297));
  OAI21xp33_ASAP7_75t_L     g05041(.A1(new_n5047), .A2(new_n5044), .B(new_n5046), .Y(new_n5298));
  NOR2xp33_ASAP7_75t_L      g05042(.A(new_n5289), .B(new_n5298), .Y(new_n5299));
  NOR3xp33_ASAP7_75t_L      g05043(.A(new_n5299), .B(new_n5297), .C(new_n5100), .Y(new_n5300));
  NOR3xp33_ASAP7_75t_L      g05044(.A(new_n5094), .B(new_n5296), .C(new_n5300), .Y(new_n5301));
  MAJIxp5_ASAP7_75t_L       g05045(.A(new_n5069), .B(new_n5054), .C(new_n5066), .Y(new_n5302));
  OAI21xp33_ASAP7_75t_L     g05046(.A1(new_n5297), .A2(new_n5299), .B(new_n5100), .Y(new_n5303));
  NAND3xp33_ASAP7_75t_L     g05047(.A(new_n5290), .B(new_n5295), .C(new_n5101), .Y(new_n5304));
  AOI21xp33_ASAP7_75t_L     g05048(.A1(new_n5304), .A2(new_n5303), .B(new_n5302), .Y(new_n5305));
  NOR2xp33_ASAP7_75t_L      g05049(.A(new_n4613), .B(new_n287), .Y(new_n5306));
  AOI221xp5_ASAP7_75t_L     g05050(.A1(\b[37] ), .A2(new_n264), .B1(\b[38] ), .B2(new_n283), .C(new_n5306), .Y(new_n5307));
  A2O1A1Ixp33_ASAP7_75t_L   g05051(.A1(new_n5079), .A2(new_n4583), .B(new_n4582), .C(new_n4615), .Y(new_n5308));
  O2A1O1Ixp33_ASAP7_75t_L   g05052(.A1(new_n4581), .A2(new_n4613), .B(new_n5308), .C(new_n5081), .Y(new_n5309));
  NOR2xp33_ASAP7_75t_L      g05053(.A(\b[37] ), .B(\b[38] ), .Y(new_n5310));
  INVx1_ASAP7_75t_L         g05054(.A(\b[38] ), .Y(new_n5311));
  NOR2xp33_ASAP7_75t_L      g05055(.A(new_n5074), .B(new_n5311), .Y(new_n5312));
  NOR2xp33_ASAP7_75t_L      g05056(.A(new_n5310), .B(new_n5312), .Y(new_n5313));
  A2O1A1Ixp33_ASAP7_75t_L   g05057(.A1(\b[37] ), .A2(\b[36] ), .B(new_n5309), .C(new_n5313), .Y(new_n5314));
  A2O1A1O1Ixp25_ASAP7_75t_L g05058(.A1(new_n4615), .A2(new_n4619), .B(new_n4614), .C(new_n5076), .D(new_n5075), .Y(new_n5315));
  INVx1_ASAP7_75t_L         g05059(.A(new_n5313), .Y(new_n5316));
  NAND2xp33_ASAP7_75t_L     g05060(.A(new_n5316), .B(new_n5315), .Y(new_n5317));
  NAND2xp33_ASAP7_75t_L     g05061(.A(new_n5317), .B(new_n5314), .Y(new_n5318));
  O2A1O1Ixp33_ASAP7_75t_L   g05062(.A1(new_n279), .A2(new_n5318), .B(new_n5307), .C(new_n257), .Y(new_n5319));
  INVx1_ASAP7_75t_L         g05063(.A(new_n5319), .Y(new_n5320));
  O2A1O1Ixp33_ASAP7_75t_L   g05064(.A1(new_n279), .A2(new_n5318), .B(new_n5307), .C(\a[2] ), .Y(new_n5321));
  AO21x2_ASAP7_75t_L        g05065(.A1(\a[2] ), .A2(new_n5320), .B(new_n5321), .Y(new_n5322));
  NOR3xp33_ASAP7_75t_L      g05066(.A(new_n5301), .B(new_n5305), .C(new_n5322), .Y(new_n5323));
  NAND3xp33_ASAP7_75t_L     g05067(.A(new_n5302), .B(new_n5303), .C(new_n5304), .Y(new_n5324));
  OAI21xp33_ASAP7_75t_L     g05068(.A1(new_n5296), .A2(new_n5300), .B(new_n5094), .Y(new_n5325));
  AOI21xp33_ASAP7_75t_L     g05069(.A1(new_n5320), .A2(\a[2] ), .B(new_n5321), .Y(new_n5326));
  AOI21xp33_ASAP7_75t_L     g05070(.A1(new_n5324), .A2(new_n5325), .B(new_n5326), .Y(new_n5327));
  NOR2xp33_ASAP7_75t_L      g05071(.A(new_n5327), .B(new_n5323), .Y(new_n5328));
  O2A1O1Ixp33_ASAP7_75t_L   g05072(.A1(new_n4857), .A2(new_n5091), .B(new_n5090), .C(new_n5328), .Y(new_n5329));
  A2O1A1O1Ixp25_ASAP7_75t_L g05073(.A1(new_n4854), .A2(new_n4848), .B(new_n4842), .C(new_n5088), .D(new_n5089), .Y(new_n5330));
  AND2x2_ASAP7_75t_L        g05074(.A(new_n5328), .B(new_n5330), .Y(new_n5331));
  NOR2xp33_ASAP7_75t_L      g05075(.A(new_n5331), .B(new_n5329), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g05076(.A(new_n5305), .B(new_n5301), .Y(new_n5333));
  A2O1A1Ixp33_ASAP7_75t_L   g05077(.A1(\a[2] ), .A2(new_n5320), .B(new_n5321), .C(new_n5333), .Y(new_n5334));
  OAI21xp33_ASAP7_75t_L     g05078(.A1(new_n5296), .A2(new_n5094), .B(new_n5304), .Y(new_n5335));
  OAI21xp33_ASAP7_75t_L     g05079(.A1(new_n5282), .A2(new_n5281), .B(new_n5277), .Y(new_n5336));
  A2O1A1O1Ixp25_ASAP7_75t_L g05080(.A1(new_n5125), .A2(new_n5120), .B(new_n4993), .C(new_n4989), .D(new_n5257), .Y(new_n5337));
  NOR2xp33_ASAP7_75t_L      g05081(.A(new_n5228), .B(new_n5225), .Y(new_n5338));
  NAND2xp33_ASAP7_75t_L     g05082(.A(new_n5234), .B(new_n5338), .Y(new_n5339));
  NAND2xp33_ASAP7_75t_L     g05083(.A(new_n5206), .B(new_n5209), .Y(new_n5340));
  INVx1_ASAP7_75t_L         g05084(.A(new_n5213), .Y(new_n5341));
  INVx1_ASAP7_75t_L         g05085(.A(new_n5214), .Y(new_n5342));
  O2A1O1Ixp33_ASAP7_75t_L   g05086(.A1(new_n5341), .A2(new_n1952), .B(new_n5342), .C(new_n5340), .Y(new_n5343));
  O2A1O1Ixp33_ASAP7_75t_L   g05087(.A1(new_n4945), .A2(new_n4950), .B(new_n5200), .C(new_n5201), .Y(new_n5344));
  INVx1_ASAP7_75t_L         g05088(.A(\a[39] ), .Y(new_n5345));
  NAND2xp33_ASAP7_75t_L     g05089(.A(\a[38] ), .B(new_n5345), .Y(new_n5346));
  NAND2xp33_ASAP7_75t_L     g05090(.A(\a[39] ), .B(new_n4906), .Y(new_n5347));
  AND2x2_ASAP7_75t_L        g05091(.A(new_n5346), .B(new_n5347), .Y(new_n5348));
  NOR2xp33_ASAP7_75t_L      g05092(.A(new_n284), .B(new_n5348), .Y(new_n5349));
  A2O1A1Ixp33_ASAP7_75t_L   g05093(.A1(new_n5143), .A2(new_n5147), .B(new_n4914), .C(new_n5349), .Y(new_n5350));
  A2O1A1Ixp33_ASAP7_75t_L   g05094(.A1(new_n5346), .A2(new_n5347), .B(new_n284), .C(new_n5163), .Y(new_n5351));
  NAND2xp33_ASAP7_75t_L     g05095(.A(\b[3] ), .B(new_n4917), .Y(new_n5352));
  NAND2xp33_ASAP7_75t_L     g05096(.A(\b[1] ), .B(new_n5139), .Y(new_n5353));
  NAND2xp33_ASAP7_75t_L     g05097(.A(\b[2] ), .B(new_n4916), .Y(new_n5354));
  NAND2xp33_ASAP7_75t_L     g05098(.A(new_n4912), .B(new_n312), .Y(new_n5355));
  NAND4xp25_ASAP7_75t_L     g05099(.A(new_n5355), .B(new_n5352), .C(new_n5353), .D(new_n5354), .Y(new_n5356));
  OAI211xp5_ASAP7_75t_L     g05100(.A1(new_n5144), .A2(new_n262), .B(new_n5352), .C(new_n5354), .Y(new_n5357));
  A2O1A1Ixp33_ASAP7_75t_L   g05101(.A1(new_n312), .A2(new_n4912), .B(new_n5357), .C(\a[38] ), .Y(new_n5358));
  AOI211xp5_ASAP7_75t_L     g05102(.A1(new_n312), .A2(new_n4912), .B(new_n4906), .C(new_n5357), .Y(new_n5359));
  AOI21xp33_ASAP7_75t_L     g05103(.A1(new_n5358), .A2(new_n5356), .B(new_n5359), .Y(new_n5360));
  AO21x2_ASAP7_75t_L        g05104(.A1(new_n5350), .A2(new_n5351), .B(new_n5360), .Y(new_n5361));
  NAND3xp33_ASAP7_75t_L     g05105(.A(new_n5351), .B(new_n5350), .C(new_n5360), .Y(new_n5362));
  NOR2xp33_ASAP7_75t_L      g05106(.A(new_n431), .B(new_n433), .Y(new_n5363));
  NAND2xp33_ASAP7_75t_L     g05107(.A(\b[5] ), .B(new_n4155), .Y(new_n5364));
  OAI221xp5_ASAP7_75t_L     g05108(.A1(new_n4147), .A2(new_n427), .B1(new_n332), .B2(new_n4397), .C(new_n5364), .Y(new_n5365));
  A2O1A1Ixp33_ASAP7_75t_L   g05109(.A1(new_n5363), .A2(new_n4151), .B(new_n5365), .C(\a[35] ), .Y(new_n5366));
  AOI211xp5_ASAP7_75t_L     g05110(.A1(new_n5363), .A2(new_n4151), .B(new_n5365), .C(new_n4145), .Y(new_n5367));
  A2O1A1O1Ixp25_ASAP7_75t_L g05111(.A1(new_n4151), .A2(new_n5363), .B(new_n5365), .C(new_n5366), .D(new_n5367), .Y(new_n5368));
  NAND3xp33_ASAP7_75t_L     g05112(.A(new_n5361), .B(new_n5362), .C(new_n5368), .Y(new_n5369));
  AOI21xp33_ASAP7_75t_L     g05113(.A1(new_n5351), .A2(new_n5350), .B(new_n5360), .Y(new_n5370));
  AND3x1_ASAP7_75t_L        g05114(.A(new_n5351), .B(new_n5360), .C(new_n5350), .Y(new_n5371));
  INVx1_ASAP7_75t_L         g05115(.A(new_n5368), .Y(new_n5372));
  OAI21xp33_ASAP7_75t_L     g05116(.A1(new_n5370), .A2(new_n5371), .B(new_n5372), .Y(new_n5373));
  NOR2xp33_ASAP7_75t_L      g05117(.A(new_n5163), .B(new_n5161), .Y(new_n5374));
  MAJIxp5_ASAP7_75t_L       g05118(.A(new_n5137), .B(new_n5374), .C(new_n5166), .Y(new_n5375));
  NAND3xp33_ASAP7_75t_L     g05119(.A(new_n5375), .B(new_n5373), .C(new_n5369), .Y(new_n5376));
  NOR3xp33_ASAP7_75t_L      g05120(.A(new_n5371), .B(new_n5372), .C(new_n5370), .Y(new_n5377));
  AOI21xp33_ASAP7_75t_L     g05121(.A1(new_n5361), .A2(new_n5362), .B(new_n5368), .Y(new_n5378));
  AOI21xp33_ASAP7_75t_L     g05122(.A1(new_n4928), .A2(new_n4934), .B(new_n4926), .Y(new_n5379));
  INVx1_ASAP7_75t_L         g05123(.A(new_n5165), .Y(new_n5380));
  A2O1A1Ixp33_ASAP7_75t_L   g05124(.A1(\a[35] ), .A2(new_n5380), .B(new_n5153), .C(new_n5374), .Y(new_n5381));
  NOR2xp33_ASAP7_75t_L      g05125(.A(new_n5156), .B(new_n5167), .Y(new_n5382));
  OAI21xp33_ASAP7_75t_L     g05126(.A1(new_n5382), .A2(new_n5379), .B(new_n5381), .Y(new_n5383));
  OAI21xp33_ASAP7_75t_L     g05127(.A1(new_n5377), .A2(new_n5378), .B(new_n5383), .Y(new_n5384));
  NOR2xp33_ASAP7_75t_L      g05128(.A(new_n534), .B(new_n3509), .Y(new_n5385));
  AOI221xp5_ASAP7_75t_L     g05129(.A1(\b[7] ), .A2(new_n3708), .B1(\b[9] ), .B2(new_n3503), .C(new_n5385), .Y(new_n5386));
  INVx1_ASAP7_75t_L         g05130(.A(new_n5386), .Y(new_n5387));
  A2O1A1Ixp33_ASAP7_75t_L   g05131(.A1(new_n602), .A2(new_n3505), .B(new_n5387), .C(\a[32] ), .Y(new_n5388));
  O2A1O1Ixp33_ASAP7_75t_L   g05132(.A1(new_n3513), .A2(new_n1066), .B(new_n5386), .C(\a[32] ), .Y(new_n5389));
  AOI21xp33_ASAP7_75t_L     g05133(.A1(new_n5388), .A2(\a[32] ), .B(new_n5389), .Y(new_n5390));
  NAND3xp33_ASAP7_75t_L     g05134(.A(new_n5384), .B(new_n5376), .C(new_n5390), .Y(new_n5391));
  OAI21xp33_ASAP7_75t_L     g05135(.A1(new_n5167), .A2(new_n5156), .B(new_n5137), .Y(new_n5392));
  AND4x1_ASAP7_75t_L        g05136(.A(new_n5392), .B(new_n5373), .C(new_n5369), .D(new_n5381), .Y(new_n5393));
  AOI21xp33_ASAP7_75t_L     g05137(.A1(new_n5373), .A2(new_n5369), .B(new_n5375), .Y(new_n5394));
  AO21x2_ASAP7_75t_L        g05138(.A1(\a[32] ), .A2(new_n5388), .B(new_n5389), .Y(new_n5395));
  OAI21xp33_ASAP7_75t_L     g05139(.A1(new_n5394), .A2(new_n5393), .B(new_n5395), .Y(new_n5396));
  NAND3xp33_ASAP7_75t_L     g05140(.A(new_n5158), .B(new_n5168), .C(new_n5174), .Y(new_n5397));
  A2O1A1O1Ixp25_ASAP7_75t_L g05141(.A1(new_n4938), .A2(new_n4885), .B(new_n5135), .C(new_n5397), .D(new_n5175), .Y(new_n5398));
  NAND3xp33_ASAP7_75t_L     g05142(.A(new_n5398), .B(new_n5396), .C(new_n5391), .Y(new_n5399));
  AO21x2_ASAP7_75t_L        g05143(.A1(new_n5391), .A2(new_n5396), .B(new_n5398), .Y(new_n5400));
  NOR2xp33_ASAP7_75t_L      g05144(.A(new_n748), .B(new_n2925), .Y(new_n5401));
  AOI221xp5_ASAP7_75t_L     g05145(.A1(\b[10] ), .A2(new_n3129), .B1(\b[12] ), .B2(new_n2938), .C(new_n5401), .Y(new_n5402));
  O2A1O1Ixp33_ASAP7_75t_L   g05146(.A1(new_n2940), .A2(new_n841), .B(new_n5402), .C(new_n2928), .Y(new_n5403));
  INVx1_ASAP7_75t_L         g05147(.A(new_n5402), .Y(new_n5404));
  A2O1A1Ixp33_ASAP7_75t_L   g05148(.A1(new_n1057), .A2(new_n2932), .B(new_n5404), .C(new_n2928), .Y(new_n5405));
  OAI21xp33_ASAP7_75t_L     g05149(.A1(new_n2928), .A2(new_n5403), .B(new_n5405), .Y(new_n5406));
  AOI21xp33_ASAP7_75t_L     g05150(.A1(new_n5400), .A2(new_n5399), .B(new_n5406), .Y(new_n5407));
  AND3x1_ASAP7_75t_L        g05151(.A(new_n5398), .B(new_n5396), .C(new_n5391), .Y(new_n5408));
  AOI21xp33_ASAP7_75t_L     g05152(.A1(new_n5396), .A2(new_n5391), .B(new_n5398), .Y(new_n5409));
  A2O1A1Ixp33_ASAP7_75t_L   g05153(.A1(new_n1057), .A2(new_n2932), .B(new_n5404), .C(\a[29] ), .Y(new_n5410));
  O2A1O1Ixp33_ASAP7_75t_L   g05154(.A1(new_n2940), .A2(new_n841), .B(new_n5402), .C(\a[29] ), .Y(new_n5411));
  AOI21xp33_ASAP7_75t_L     g05155(.A1(new_n5410), .A2(\a[29] ), .B(new_n5411), .Y(new_n5412));
  NOR3xp33_ASAP7_75t_L      g05156(.A(new_n5408), .B(new_n5409), .C(new_n5412), .Y(new_n5413));
  NOR2xp33_ASAP7_75t_L      g05157(.A(new_n5407), .B(new_n5413), .Y(new_n5414));
  NAND2xp33_ASAP7_75t_L     g05158(.A(new_n5185), .B(new_n5184), .Y(new_n5415));
  MAJIxp5_ASAP7_75t_L       g05159(.A(new_n5189), .B(new_n5183), .C(new_n5415), .Y(new_n5416));
  NAND2xp33_ASAP7_75t_L     g05160(.A(new_n5414), .B(new_n5416), .Y(new_n5417));
  NOR2xp33_ASAP7_75t_L      g05161(.A(new_n5177), .B(new_n5180), .Y(new_n5418));
  A2O1A1Ixp33_ASAP7_75t_L   g05162(.A1(new_n5182), .A2(\a[29] ), .B(new_n5132), .C(new_n5418), .Y(new_n5419));
  NOR2xp33_ASAP7_75t_L      g05163(.A(new_n5190), .B(new_n5191), .Y(new_n5420));
  OAI221xp5_ASAP7_75t_L     g05164(.A1(new_n5407), .A2(new_n5413), .B1(new_n5189), .B2(new_n5420), .C(new_n5419), .Y(new_n5421));
  NOR2xp33_ASAP7_75t_L      g05165(.A(new_n960), .B(new_n2410), .Y(new_n5422));
  AOI221xp5_ASAP7_75t_L     g05166(.A1(\b[13] ), .A2(new_n2577), .B1(\b[15] ), .B2(new_n2423), .C(new_n5422), .Y(new_n5423));
  INVx1_ASAP7_75t_L         g05167(.A(new_n5423), .Y(new_n5424));
  A2O1A1Ixp33_ASAP7_75t_L   g05168(.A1(new_n1052), .A2(new_n2417), .B(new_n5424), .C(\a[26] ), .Y(new_n5425));
  O2A1O1Ixp33_ASAP7_75t_L   g05169(.A1(new_n2425), .A2(new_n1774), .B(new_n5423), .C(\a[26] ), .Y(new_n5426));
  AOI21xp33_ASAP7_75t_L     g05170(.A1(new_n5425), .A2(\a[26] ), .B(new_n5426), .Y(new_n5427));
  NAND3xp33_ASAP7_75t_L     g05171(.A(new_n5417), .B(new_n5427), .C(new_n5421), .Y(new_n5428));
  OAI21xp33_ASAP7_75t_L     g05172(.A1(new_n5409), .A2(new_n5408), .B(new_n5412), .Y(new_n5429));
  NAND3xp33_ASAP7_75t_L     g05173(.A(new_n5400), .B(new_n5399), .C(new_n5406), .Y(new_n5430));
  NAND2xp33_ASAP7_75t_L     g05174(.A(new_n5430), .B(new_n5429), .Y(new_n5431));
  O2A1O1Ixp33_ASAP7_75t_L   g05175(.A1(new_n5189), .A2(new_n5420), .B(new_n5419), .C(new_n5431), .Y(new_n5432));
  NOR2xp33_ASAP7_75t_L      g05176(.A(new_n5414), .B(new_n5416), .Y(new_n5433));
  O2A1O1Ixp33_ASAP7_75t_L   g05177(.A1(new_n2425), .A2(new_n1774), .B(new_n5423), .C(new_n2413), .Y(new_n5434));
  A2O1A1Ixp33_ASAP7_75t_L   g05178(.A1(new_n1052), .A2(new_n2417), .B(new_n5424), .C(new_n2413), .Y(new_n5435));
  OAI21xp33_ASAP7_75t_L     g05179(.A1(new_n2413), .A2(new_n5434), .B(new_n5435), .Y(new_n5436));
  OAI21xp33_ASAP7_75t_L     g05180(.A1(new_n5432), .A2(new_n5433), .B(new_n5436), .Y(new_n5437));
  NAND2xp33_ASAP7_75t_L     g05181(.A(new_n5428), .B(new_n5437), .Y(new_n5438));
  O2A1O1Ixp33_ASAP7_75t_L   g05182(.A1(new_n5344), .A2(new_n5198), .B(new_n5206), .C(new_n5438), .Y(new_n5439));
  OAI21xp33_ASAP7_75t_L     g05183(.A1(new_n5207), .A2(new_n5208), .B(new_n5205), .Y(new_n5440));
  NAND2xp33_ASAP7_75t_L     g05184(.A(new_n5421), .B(new_n5417), .Y(new_n5441));
  O2A1O1Ixp33_ASAP7_75t_L   g05185(.A1(new_n5434), .A2(new_n2413), .B(new_n5435), .C(new_n5441), .Y(new_n5442));
  O2A1O1Ixp33_ASAP7_75t_L   g05186(.A1(new_n5427), .A2(new_n5442), .B(new_n5428), .C(new_n5440), .Y(new_n5443));
  NOR2xp33_ASAP7_75t_L      g05187(.A(new_n1349), .B(new_n1962), .Y(new_n5444));
  AOI221xp5_ASAP7_75t_L     g05188(.A1(new_n1955), .A2(\b[18] ), .B1(new_n2093), .B2(\b[16] ), .C(new_n5444), .Y(new_n5445));
  INVx1_ASAP7_75t_L         g05189(.A(new_n5445), .Y(new_n5446));
  A2O1A1Ixp33_ASAP7_75t_L   g05190(.A1(new_n2329), .A2(new_n1964), .B(new_n5446), .C(\a[23] ), .Y(new_n5447));
  O2A1O1Ixp33_ASAP7_75t_L   g05191(.A1(new_n1956), .A2(new_n1464), .B(new_n5445), .C(\a[23] ), .Y(new_n5448));
  AOI21xp33_ASAP7_75t_L     g05192(.A1(new_n5447), .A2(\a[23] ), .B(new_n5448), .Y(new_n5449));
  INVx1_ASAP7_75t_L         g05193(.A(new_n5449), .Y(new_n5450));
  OAI21xp33_ASAP7_75t_L     g05194(.A1(new_n5439), .A2(new_n5443), .B(new_n5450), .Y(new_n5451));
  NAND3xp33_ASAP7_75t_L     g05195(.A(new_n5440), .B(new_n5428), .C(new_n5437), .Y(new_n5452));
  A2O1A1Ixp33_ASAP7_75t_L   g05196(.A1(new_n4462), .A2(new_n4963), .B(new_n4724), .C(new_n4712), .Y(new_n5453));
  AOI21xp33_ASAP7_75t_L     g05197(.A1(new_n5187), .A2(new_n5192), .B(new_n5198), .Y(new_n5454));
  A2O1A1O1Ixp25_ASAP7_75t_L g05198(.A1(new_n4965), .A2(new_n5453), .B(new_n4954), .C(new_n5199), .D(new_n5454), .Y(new_n5455));
  NAND2xp33_ASAP7_75t_L     g05199(.A(new_n5455), .B(new_n5438), .Y(new_n5456));
  NAND3xp33_ASAP7_75t_L     g05200(.A(new_n5452), .B(new_n5456), .C(new_n5449), .Y(new_n5457));
  AO221x2_ASAP7_75t_L       g05201(.A1(new_n5221), .A2(new_n5224), .B1(new_n5451), .B2(new_n5457), .C(new_n5343), .Y(new_n5458));
  NOR2xp33_ASAP7_75t_L      g05202(.A(new_n5218), .B(new_n5217), .Y(new_n5459));
  A2O1A1Ixp33_ASAP7_75t_L   g05203(.A1(\a[23] ), .A2(new_n5213), .B(new_n5214), .C(new_n5459), .Y(new_n5460));
  A2O1A1Ixp33_ASAP7_75t_L   g05204(.A1(new_n5215), .A2(new_n5216), .B(new_n5227), .C(new_n5460), .Y(new_n5461));
  NAND3xp33_ASAP7_75t_L     g05205(.A(new_n5461), .B(new_n5451), .C(new_n5457), .Y(new_n5462));
  NOR2xp33_ASAP7_75t_L      g05206(.A(new_n1745), .B(new_n1517), .Y(new_n5463));
  AOI221xp5_ASAP7_75t_L     g05207(.A1(\b[19] ), .A2(new_n1659), .B1(\b[21] ), .B2(new_n1511), .C(new_n5463), .Y(new_n5464));
  O2A1O1Ixp33_ASAP7_75t_L   g05208(.A1(new_n1521), .A2(new_n1901), .B(new_n5464), .C(new_n1501), .Y(new_n5465));
  INVx1_ASAP7_75t_L         g05209(.A(new_n5465), .Y(new_n5466));
  O2A1O1Ixp33_ASAP7_75t_L   g05210(.A1(new_n1521), .A2(new_n1901), .B(new_n5464), .C(\a[20] ), .Y(new_n5467));
  AOI21xp33_ASAP7_75t_L     g05211(.A1(new_n5466), .A2(\a[20] ), .B(new_n5467), .Y(new_n5468));
  NAND3xp33_ASAP7_75t_L     g05212(.A(new_n5462), .B(new_n5458), .C(new_n5468), .Y(new_n5469));
  AOI21xp33_ASAP7_75t_L     g05213(.A1(new_n5457), .A2(new_n5451), .B(new_n5461), .Y(new_n5470));
  NAND2xp33_ASAP7_75t_L     g05214(.A(new_n5224), .B(new_n5221), .Y(new_n5471));
  NAND2xp33_ASAP7_75t_L     g05215(.A(new_n5457), .B(new_n5451), .Y(new_n5472));
  O2A1O1Ixp33_ASAP7_75t_L   g05216(.A1(new_n5340), .A2(new_n5215), .B(new_n5471), .C(new_n5472), .Y(new_n5473));
  AO21x2_ASAP7_75t_L        g05217(.A1(\a[20] ), .A2(new_n5466), .B(new_n5467), .Y(new_n5474));
  OAI21xp33_ASAP7_75t_L     g05218(.A1(new_n5470), .A2(new_n5473), .B(new_n5474), .Y(new_n5475));
  AND4x1_ASAP7_75t_L        g05219(.A(new_n5253), .B(new_n5339), .C(new_n5475), .D(new_n5469), .Y(new_n5476));
  MAJIxp5_ASAP7_75t_L       g05220(.A(new_n5238), .B(new_n5234), .C(new_n5338), .Y(new_n5477));
  AOI21xp33_ASAP7_75t_L     g05221(.A1(new_n5475), .A2(new_n5469), .B(new_n5477), .Y(new_n5478));
  NOR2xp33_ASAP7_75t_L      g05222(.A(new_n2205), .B(new_n1284), .Y(new_n5479));
  AOI221xp5_ASAP7_75t_L     g05223(.A1(\b[22] ), .A2(new_n1290), .B1(\b[23] ), .B2(new_n1204), .C(new_n5479), .Y(new_n5480));
  OA21x2_ASAP7_75t_L        g05224(.A1(new_n1210), .A2(new_n2853), .B(new_n5480), .Y(new_n5481));
  O2A1O1Ixp33_ASAP7_75t_L   g05225(.A1(new_n1210), .A2(new_n2853), .B(new_n5480), .C(new_n1206), .Y(new_n5482));
  NAND2xp33_ASAP7_75t_L     g05226(.A(\a[17] ), .B(new_n5481), .Y(new_n5483));
  OA21x2_ASAP7_75t_L        g05227(.A1(new_n5481), .A2(new_n5482), .B(new_n5483), .Y(new_n5484));
  OAI21xp33_ASAP7_75t_L     g05228(.A1(new_n5478), .A2(new_n5476), .B(new_n5484), .Y(new_n5485));
  NAND3xp33_ASAP7_75t_L     g05229(.A(new_n5477), .B(new_n5475), .C(new_n5469), .Y(new_n5486));
  AO22x1_ASAP7_75t_L        g05230(.A1(new_n5469), .A2(new_n5475), .B1(new_n5339), .B2(new_n5253), .Y(new_n5487));
  NAND2xp33_ASAP7_75t_L     g05231(.A(new_n1216), .B(new_n2216), .Y(new_n5488));
  A2O1A1Ixp33_ASAP7_75t_L   g05232(.A1(new_n5488), .A2(new_n5480), .B(new_n5482), .C(new_n5483), .Y(new_n5489));
  NAND3xp33_ASAP7_75t_L     g05233(.A(new_n5487), .B(new_n5486), .C(new_n5489), .Y(new_n5490));
  OAI211xp5_ASAP7_75t_L     g05234(.A1(new_n5247), .A2(new_n5337), .B(new_n5485), .C(new_n5490), .Y(new_n5491));
  NAND2xp33_ASAP7_75t_L     g05235(.A(new_n5123), .B(new_n5124), .Y(new_n5492));
  A2O1A1O1Ixp25_ASAP7_75t_L g05236(.A1(new_n4999), .A2(new_n5492), .B(new_n5118), .C(new_n5260), .D(new_n5247), .Y(new_n5493));
  AOI21xp33_ASAP7_75t_L     g05237(.A1(new_n5487), .A2(new_n5486), .B(new_n5489), .Y(new_n5494));
  NOR3xp33_ASAP7_75t_L      g05238(.A(new_n5476), .B(new_n5484), .C(new_n5478), .Y(new_n5495));
  OAI21xp33_ASAP7_75t_L     g05239(.A1(new_n5494), .A2(new_n5495), .B(new_n5493), .Y(new_n5496));
  NOR2xp33_ASAP7_75t_L      g05240(.A(new_n2703), .B(new_n864), .Y(new_n5497));
  AOI221xp5_ASAP7_75t_L     g05241(.A1(\b[25] ), .A2(new_n985), .B1(\b[27] ), .B2(new_n886), .C(new_n5497), .Y(new_n5498));
  INVx1_ASAP7_75t_L         g05242(.A(new_n5498), .Y(new_n5499));
  A2O1A1Ixp33_ASAP7_75t_L   g05243(.A1(new_n2887), .A2(new_n873), .B(new_n5499), .C(\a[14] ), .Y(new_n5500));
  O2A1O1Ixp33_ASAP7_75t_L   g05244(.A1(new_n872), .A2(new_n2889), .B(new_n5498), .C(\a[14] ), .Y(new_n5501));
  AOI21xp33_ASAP7_75t_L     g05245(.A1(new_n5500), .A2(\a[14] ), .B(new_n5501), .Y(new_n5502));
  NAND3xp33_ASAP7_75t_L     g05246(.A(new_n5491), .B(new_n5496), .C(new_n5502), .Y(new_n5503));
  NOR3xp33_ASAP7_75t_L      g05247(.A(new_n5493), .B(new_n5494), .C(new_n5495), .Y(new_n5504));
  AOI211xp5_ASAP7_75t_L     g05248(.A1(new_n5490), .A2(new_n5485), .B(new_n5247), .C(new_n5337), .Y(new_n5505));
  O2A1O1Ixp33_ASAP7_75t_L   g05249(.A1(new_n872), .A2(new_n2889), .B(new_n5498), .C(new_n867), .Y(new_n5506));
  INVx1_ASAP7_75t_L         g05250(.A(new_n5501), .Y(new_n5507));
  OAI21xp33_ASAP7_75t_L     g05251(.A1(new_n867), .A2(new_n5506), .B(new_n5507), .Y(new_n5508));
  OAI21xp33_ASAP7_75t_L     g05252(.A1(new_n5504), .A2(new_n5505), .B(new_n5508), .Y(new_n5509));
  NAND2xp33_ASAP7_75t_L     g05253(.A(new_n5509), .B(new_n5503), .Y(new_n5510));
  O2A1O1Ixp33_ASAP7_75t_L   g05254(.A1(new_n5024), .A2(new_n5272), .B(new_n5269), .C(new_n5510), .Y(new_n5511));
  A2O1A1Ixp33_ASAP7_75t_L   g05255(.A1(new_n5271), .A2(new_n5008), .B(new_n5272), .C(new_n5269), .Y(new_n5512));
  NAND3xp33_ASAP7_75t_L     g05256(.A(new_n5491), .B(new_n5508), .C(new_n5496), .Y(new_n5513));
  INVx1_ASAP7_75t_L         g05257(.A(new_n5513), .Y(new_n5514));
  O2A1O1Ixp33_ASAP7_75t_L   g05258(.A1(new_n5502), .A2(new_n5514), .B(new_n5503), .C(new_n5512), .Y(new_n5515));
  NOR2xp33_ASAP7_75t_L      g05259(.A(new_n3098), .B(new_n1550), .Y(new_n5516));
  AOI221xp5_ASAP7_75t_L     g05260(.A1(\b[28] ), .A2(new_n713), .B1(\b[30] ), .B2(new_n640), .C(new_n5516), .Y(new_n5517));
  O2A1O1Ixp33_ASAP7_75t_L   g05261(.A1(new_n641), .A2(new_n3464), .B(new_n5517), .C(new_n637), .Y(new_n5518));
  NOR2xp33_ASAP7_75t_L      g05262(.A(new_n637), .B(new_n5518), .Y(new_n5519));
  O2A1O1Ixp33_ASAP7_75t_L   g05263(.A1(new_n641), .A2(new_n3464), .B(new_n5517), .C(\a[11] ), .Y(new_n5520));
  OAI22xp33_ASAP7_75t_L     g05264(.A1(new_n5515), .A2(new_n5511), .B1(new_n5520), .B2(new_n5519), .Y(new_n5521));
  NAND3xp33_ASAP7_75t_L     g05265(.A(new_n5512), .B(new_n5503), .C(new_n5509), .Y(new_n5522));
  A2O1A1O1Ixp25_ASAP7_75t_L g05266(.A1(new_n5013), .A2(new_n4867), .B(new_n5009), .C(new_n5268), .D(new_n5273), .Y(new_n5523));
  NOR3xp33_ASAP7_75t_L      g05267(.A(new_n5508), .B(new_n5505), .C(new_n5504), .Y(new_n5524));
  A2O1A1Ixp33_ASAP7_75t_L   g05268(.A1(new_n5508), .A2(new_n5513), .B(new_n5524), .C(new_n5523), .Y(new_n5525));
  NOR2xp33_ASAP7_75t_L      g05269(.A(new_n5520), .B(new_n5519), .Y(new_n5526));
  NAND3xp33_ASAP7_75t_L     g05270(.A(new_n5522), .B(new_n5526), .C(new_n5525), .Y(new_n5527));
  NAND3xp33_ASAP7_75t_L     g05271(.A(new_n5336), .B(new_n5521), .C(new_n5527), .Y(new_n5528));
  A2O1A1O1Ixp25_ASAP7_75t_L g05272(.A1(new_n5021), .A2(new_n4866), .B(new_n5034), .C(new_n5275), .D(new_n5276), .Y(new_n5529));
  AOI21xp33_ASAP7_75t_L     g05273(.A1(new_n5522), .A2(new_n5525), .B(new_n5526), .Y(new_n5530));
  AND3x1_ASAP7_75t_L        g05274(.A(new_n5522), .B(new_n5526), .C(new_n5525), .Y(new_n5531));
  OAI21xp33_ASAP7_75t_L     g05275(.A1(new_n5530), .A2(new_n5531), .B(new_n5529), .Y(new_n5532));
  NOR2xp33_ASAP7_75t_L      g05276(.A(new_n3891), .B(new_n513), .Y(new_n5533));
  AOI221xp5_ASAP7_75t_L     g05277(.A1(\b[31] ), .A2(new_n560), .B1(\b[33] ), .B2(new_n475), .C(new_n5533), .Y(new_n5534));
  O2A1O1Ixp33_ASAP7_75t_L   g05278(.A1(new_n477), .A2(new_n4108), .B(new_n5534), .C(new_n466), .Y(new_n5535));
  INVx1_ASAP7_75t_L         g05279(.A(new_n5535), .Y(new_n5536));
  O2A1O1Ixp33_ASAP7_75t_L   g05280(.A1(new_n477), .A2(new_n4108), .B(new_n5534), .C(\a[8] ), .Y(new_n5537));
  AOI21xp33_ASAP7_75t_L     g05281(.A1(new_n5536), .A2(\a[8] ), .B(new_n5537), .Y(new_n5538));
  NAND3xp33_ASAP7_75t_L     g05282(.A(new_n5528), .B(new_n5538), .C(new_n5532), .Y(new_n5539));
  NOR3xp33_ASAP7_75t_L      g05283(.A(new_n5529), .B(new_n5531), .C(new_n5530), .Y(new_n5540));
  AOI21xp33_ASAP7_75t_L     g05284(.A1(new_n5527), .A2(new_n5521), .B(new_n5336), .Y(new_n5541));
  AO21x2_ASAP7_75t_L        g05285(.A1(\a[8] ), .A2(new_n5536), .B(new_n5537), .Y(new_n5542));
  OAI21xp33_ASAP7_75t_L     g05286(.A1(new_n5540), .A2(new_n5541), .B(new_n5542), .Y(new_n5543));
  AND2x2_ASAP7_75t_L        g05287(.A(new_n5539), .B(new_n5543), .Y(new_n5544));
  A2O1A1Ixp33_ASAP7_75t_L   g05288(.A1(new_n5292), .A2(new_n5298), .B(new_n5288), .C(new_n5544), .Y(new_n5545));
  A2O1A1O1Ixp25_ASAP7_75t_L g05289(.A1(new_n5045), .A2(new_n5102), .B(new_n5041), .C(new_n5292), .D(new_n5288), .Y(new_n5546));
  NAND2xp33_ASAP7_75t_L     g05290(.A(new_n5539), .B(new_n5543), .Y(new_n5547));
  NAND2xp33_ASAP7_75t_L     g05291(.A(new_n5546), .B(new_n5547), .Y(new_n5548));
  OAI22xp33_ASAP7_75t_L     g05292(.A1(new_n350), .A2(new_n4581), .B1(new_n4344), .B2(new_n375), .Y(new_n5549));
  AOI221xp5_ASAP7_75t_L     g05293(.A1(new_n361), .A2(\b[36] ), .B1(new_n359), .B2(new_n4621), .C(new_n5549), .Y(new_n5550));
  XNOR2x2_ASAP7_75t_L       g05294(.A(new_n346), .B(new_n5550), .Y(new_n5551));
  NAND3xp33_ASAP7_75t_L     g05295(.A(new_n5545), .B(new_n5548), .C(new_n5551), .Y(new_n5552));
  O2A1O1Ixp33_ASAP7_75t_L   g05296(.A1(new_n5291), .A2(new_n5284), .B(new_n5293), .C(new_n5547), .Y(new_n5553));
  OAI21xp33_ASAP7_75t_L     g05297(.A1(new_n5294), .A2(new_n5291), .B(new_n5293), .Y(new_n5554));
  NAND2xp33_ASAP7_75t_L     g05298(.A(new_n5532), .B(new_n5528), .Y(new_n5555));
  INVx1_ASAP7_75t_L         g05299(.A(new_n5537), .Y(new_n5556));
  O2A1O1Ixp33_ASAP7_75t_L   g05300(.A1(new_n5535), .A2(new_n466), .B(new_n5556), .C(new_n5555), .Y(new_n5557));
  O2A1O1Ixp33_ASAP7_75t_L   g05301(.A1(new_n5555), .A2(new_n5557), .B(new_n5543), .C(new_n5554), .Y(new_n5558));
  INVx1_ASAP7_75t_L         g05302(.A(new_n5551), .Y(new_n5559));
  OAI21xp33_ASAP7_75t_L     g05303(.A1(new_n5553), .A2(new_n5558), .B(new_n5559), .Y(new_n5560));
  NAND3xp33_ASAP7_75t_L     g05304(.A(new_n5335), .B(new_n5552), .C(new_n5560), .Y(new_n5561));
  A2O1A1O1Ixp25_ASAP7_75t_L g05305(.A1(new_n5064), .A2(new_n5061), .B(new_n5067), .C(new_n5303), .D(new_n5300), .Y(new_n5562));
  NOR3xp33_ASAP7_75t_L      g05306(.A(new_n5558), .B(new_n5559), .C(new_n5553), .Y(new_n5563));
  AOI21xp33_ASAP7_75t_L     g05307(.A1(new_n5545), .A2(new_n5548), .B(new_n5551), .Y(new_n5564));
  OAI21xp33_ASAP7_75t_L     g05308(.A1(new_n5564), .A2(new_n5563), .B(new_n5562), .Y(new_n5565));
  NOR2xp33_ASAP7_75t_L      g05309(.A(new_n5074), .B(new_n287), .Y(new_n5566));
  AOI221xp5_ASAP7_75t_L     g05310(.A1(\b[38] ), .A2(new_n264), .B1(\b[39] ), .B2(new_n283), .C(new_n5566), .Y(new_n5567));
  INVx1_ASAP7_75t_L         g05311(.A(new_n5312), .Y(new_n5568));
  NOR2xp33_ASAP7_75t_L      g05312(.A(\b[38] ), .B(\b[39] ), .Y(new_n5569));
  INVx1_ASAP7_75t_L         g05313(.A(\b[39] ), .Y(new_n5570));
  NOR2xp33_ASAP7_75t_L      g05314(.A(new_n5311), .B(new_n5570), .Y(new_n5571));
  NOR2xp33_ASAP7_75t_L      g05315(.A(new_n5569), .B(new_n5571), .Y(new_n5572));
  INVx1_ASAP7_75t_L         g05316(.A(new_n5572), .Y(new_n5573));
  O2A1O1Ixp33_ASAP7_75t_L   g05317(.A1(new_n5316), .A2(new_n5315), .B(new_n5568), .C(new_n5573), .Y(new_n5574));
  INVx1_ASAP7_75t_L         g05318(.A(new_n5574), .Y(new_n5575));
  O2A1O1Ixp33_ASAP7_75t_L   g05319(.A1(new_n5075), .A2(new_n5309), .B(new_n5313), .C(new_n5312), .Y(new_n5576));
  NAND2xp33_ASAP7_75t_L     g05320(.A(new_n5573), .B(new_n5576), .Y(new_n5577));
  NAND2xp33_ASAP7_75t_L     g05321(.A(new_n5575), .B(new_n5577), .Y(new_n5578));
  O2A1O1Ixp33_ASAP7_75t_L   g05322(.A1(new_n279), .A2(new_n5578), .B(new_n5567), .C(new_n257), .Y(new_n5579));
  NOR2xp33_ASAP7_75t_L      g05323(.A(new_n257), .B(new_n5579), .Y(new_n5580));
  O2A1O1Ixp33_ASAP7_75t_L   g05324(.A1(new_n279), .A2(new_n5578), .B(new_n5567), .C(\a[2] ), .Y(new_n5581));
  NOR2xp33_ASAP7_75t_L      g05325(.A(new_n5581), .B(new_n5580), .Y(new_n5582));
  NAND3xp33_ASAP7_75t_L     g05326(.A(new_n5561), .B(new_n5565), .C(new_n5582), .Y(new_n5583));
  NOR3xp33_ASAP7_75t_L      g05327(.A(new_n5562), .B(new_n5563), .C(new_n5564), .Y(new_n5584));
  AOI21xp33_ASAP7_75t_L     g05328(.A1(new_n5560), .A2(new_n5552), .B(new_n5335), .Y(new_n5585));
  OAI22xp33_ASAP7_75t_L     g05329(.A1(new_n5585), .A2(new_n5584), .B1(new_n5581), .B2(new_n5580), .Y(new_n5586));
  NAND2xp33_ASAP7_75t_L     g05330(.A(new_n5583), .B(new_n5586), .Y(new_n5587));
  INVx1_ASAP7_75t_L         g05331(.A(new_n5587), .Y(new_n5588));
  O2A1O1Ixp33_ASAP7_75t_L   g05332(.A1(new_n5328), .A2(new_n5330), .B(new_n5334), .C(new_n5588), .Y(new_n5589));
  OAI21xp33_ASAP7_75t_L     g05333(.A1(new_n5328), .A2(new_n5330), .B(new_n5334), .Y(new_n5590));
  NOR2xp33_ASAP7_75t_L      g05334(.A(new_n5587), .B(new_n5590), .Y(new_n5591));
  NOR2xp33_ASAP7_75t_L      g05335(.A(new_n5591), .B(new_n5589), .Y(\f[39] ));
  NOR3xp33_ASAP7_75t_L      g05336(.A(new_n5585), .B(new_n5584), .C(new_n5582), .Y(new_n5593));
  A2O1A1O1Ixp25_ASAP7_75t_L g05337(.A1(new_n5322), .A2(new_n5333), .B(new_n5329), .C(new_n5587), .D(new_n5593), .Y(new_n5594));
  OAI21xp33_ASAP7_75t_L     g05338(.A1(new_n5563), .A2(new_n5562), .B(new_n5560), .Y(new_n5595));
  NOR2xp33_ASAP7_75t_L      g05339(.A(new_n4101), .B(new_n513), .Y(new_n5596));
  AOI221xp5_ASAP7_75t_L     g05340(.A1(\b[32] ), .A2(new_n560), .B1(\b[34] ), .B2(new_n475), .C(new_n5596), .Y(new_n5597));
  O2A1O1Ixp33_ASAP7_75t_L   g05341(.A1(new_n477), .A2(new_n4352), .B(new_n5597), .C(new_n466), .Y(new_n5598));
  AND2x2_ASAP7_75t_L        g05342(.A(new_n4349), .B(new_n4351), .Y(new_n5599));
  INVx1_ASAP7_75t_L         g05343(.A(new_n5597), .Y(new_n5600));
  A2O1A1Ixp33_ASAP7_75t_L   g05344(.A1(new_n5599), .A2(new_n483), .B(new_n5600), .C(new_n466), .Y(new_n5601));
  OAI21xp33_ASAP7_75t_L     g05345(.A1(new_n466), .A2(new_n5598), .B(new_n5601), .Y(new_n5602));
  OAI21xp33_ASAP7_75t_L     g05346(.A1(new_n5531), .A2(new_n5529), .B(new_n5521), .Y(new_n5603));
  A2O1A1Ixp33_ASAP7_75t_L   g05347(.A1(new_n5503), .A2(new_n5502), .B(new_n5523), .C(new_n5513), .Y(new_n5604));
  OAI22xp33_ASAP7_75t_L     g05348(.A1(new_n980), .A2(new_n2703), .B1(new_n2879), .B2(new_n864), .Y(new_n5605));
  AOI221xp5_ASAP7_75t_L     g05349(.A1(new_n886), .A2(\b[28] ), .B1(new_n873), .B2(new_n3085), .C(new_n5605), .Y(new_n5606));
  XNOR2x2_ASAP7_75t_L       g05350(.A(new_n867), .B(new_n5606), .Y(new_n5607));
  O2A1O1Ixp33_ASAP7_75t_L   g05351(.A1(new_n2928), .A2(new_n5131), .B(new_n5133), .C(new_n5415), .Y(new_n5608));
  NAND2xp33_ASAP7_75t_L     g05352(.A(new_n5186), .B(new_n5181), .Y(new_n5609));
  A2O1A1O1Ixp25_ASAP7_75t_L g05353(.A1(new_n5128), .A2(new_n5609), .B(new_n5608), .C(new_n5429), .D(new_n5413), .Y(new_n5610));
  NAND3xp33_ASAP7_75t_L     g05354(.A(new_n5384), .B(new_n5376), .C(new_n5395), .Y(new_n5611));
  A2O1A1Ixp33_ASAP7_75t_L   g05355(.A1(new_n5391), .A2(new_n5390), .B(new_n5398), .C(new_n5611), .Y(new_n5612));
  INVx1_ASAP7_75t_L         g05356(.A(new_n5349), .Y(new_n5613));
  MAJIxp5_ASAP7_75t_L       g05357(.A(new_n5360), .B(new_n5149), .C(new_n5613), .Y(new_n5614));
  NOR2xp33_ASAP7_75t_L      g05358(.A(new_n332), .B(new_n4908), .Y(new_n5615));
  AOI221xp5_ASAP7_75t_L     g05359(.A1(\b[2] ), .A2(new_n5139), .B1(\b[3] ), .B2(new_n4916), .C(new_n5615), .Y(new_n5616));
  OAI211xp5_ASAP7_75t_L     g05360(.A1(new_n1497), .A2(new_n4911), .B(new_n5616), .C(\a[38] ), .Y(new_n5617));
  NAND2xp33_ASAP7_75t_L     g05361(.A(\b[3] ), .B(new_n4916), .Y(new_n5618));
  OAI221xp5_ASAP7_75t_L     g05362(.A1(new_n4908), .A2(new_n332), .B1(new_n289), .B2(new_n5144), .C(new_n5618), .Y(new_n5619));
  A2O1A1Ixp33_ASAP7_75t_L   g05363(.A1(new_n342), .A2(new_n4912), .B(new_n5619), .C(new_n4906), .Y(new_n5620));
  NAND2xp33_ASAP7_75t_L     g05364(.A(new_n5347), .B(new_n5346), .Y(new_n5621));
  XNOR2x2_ASAP7_75t_L       g05365(.A(\a[40] ), .B(\a[39] ), .Y(new_n5622));
  NOR2xp33_ASAP7_75t_L      g05366(.A(new_n5622), .B(new_n5621), .Y(new_n5623));
  INVx1_ASAP7_75t_L         g05367(.A(\a[40] ), .Y(new_n5624));
  NAND2xp33_ASAP7_75t_L     g05368(.A(\a[41] ), .B(new_n5624), .Y(new_n5625));
  INVx1_ASAP7_75t_L         g05369(.A(\a[41] ), .Y(new_n5626));
  NAND2xp33_ASAP7_75t_L     g05370(.A(\a[40] ), .B(new_n5626), .Y(new_n5627));
  NAND2xp33_ASAP7_75t_L     g05371(.A(new_n5627), .B(new_n5625), .Y(new_n5628));
  NOR2xp33_ASAP7_75t_L      g05372(.A(new_n5628), .B(new_n5348), .Y(new_n5629));
  NAND2xp33_ASAP7_75t_L     g05373(.A(new_n5628), .B(new_n5621), .Y(new_n5630));
  NOR2xp33_ASAP7_75t_L      g05374(.A(new_n274), .B(new_n5630), .Y(new_n5631));
  AOI221xp5_ASAP7_75t_L     g05375(.A1(\b[1] ), .A2(new_n5629), .B1(new_n5623), .B2(\b[0] ), .C(new_n5631), .Y(new_n5632));
  NAND3xp33_ASAP7_75t_L     g05376(.A(new_n5632), .B(new_n5613), .C(\a[41] ), .Y(new_n5633));
  INVx1_ASAP7_75t_L         g05377(.A(new_n5633), .Y(new_n5634));
  A2O1A1Ixp33_ASAP7_75t_L   g05378(.A1(new_n5346), .A2(new_n5347), .B(new_n284), .C(\a[41] ), .Y(new_n5635));
  AOI22xp33_ASAP7_75t_L     g05379(.A1(new_n5623), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n5629), .Y(new_n5636));
  AOI21xp33_ASAP7_75t_L     g05380(.A1(new_n5627), .A2(new_n5625), .B(new_n5348), .Y(new_n5637));
  NAND2xp33_ASAP7_75t_L     g05381(.A(new_n275), .B(new_n5637), .Y(new_n5638));
  NAND3xp33_ASAP7_75t_L     g05382(.A(new_n5636), .B(\a[41] ), .C(new_n5638), .Y(new_n5639));
  OR2x4_ASAP7_75t_L         g05383(.A(new_n5622), .B(new_n5621), .Y(new_n5640));
  NAND3xp33_ASAP7_75t_L     g05384(.A(new_n5621), .B(new_n5625), .C(new_n5627), .Y(new_n5641));
  OAI22xp33_ASAP7_75t_L     g05385(.A1(new_n5640), .A2(new_n284), .B1(new_n262), .B2(new_n5641), .Y(new_n5642));
  A2O1A1Ixp33_ASAP7_75t_L   g05386(.A1(new_n5637), .A2(new_n275), .B(new_n5642), .C(new_n5626), .Y(new_n5643));
  AND3x1_ASAP7_75t_L        g05387(.A(new_n5643), .B(new_n5639), .C(new_n5635), .Y(new_n5644));
  OAI211xp5_ASAP7_75t_L     g05388(.A1(new_n5634), .A2(new_n5644), .B(new_n5620), .C(new_n5617), .Y(new_n5645));
  NAND2xp33_ASAP7_75t_L     g05389(.A(new_n5620), .B(new_n5617), .Y(new_n5646));
  O2A1O1Ixp33_ASAP7_75t_L   g05390(.A1(new_n5630), .A2(new_n274), .B(new_n5636), .C(new_n5626), .Y(new_n5647));
  A2O1A1Ixp33_ASAP7_75t_L   g05391(.A1(new_n5647), .A2(new_n5349), .B(new_n5626), .C(new_n5643), .Y(new_n5648));
  NAND3xp33_ASAP7_75t_L     g05392(.A(new_n5646), .B(new_n5633), .C(new_n5648), .Y(new_n5649));
  NAND3xp33_ASAP7_75t_L     g05393(.A(new_n5614), .B(new_n5645), .C(new_n5649), .Y(new_n5650));
  NAND5xp2_ASAP7_75t_L      g05394(.A(new_n5355), .B(new_n5354), .C(new_n5353), .D(new_n5352), .E(\a[38] ), .Y(new_n5651));
  A2O1A1Ixp33_ASAP7_75t_L   g05395(.A1(new_n312), .A2(new_n4912), .B(new_n5357), .C(new_n4906), .Y(new_n5652));
  NAND2xp33_ASAP7_75t_L     g05396(.A(new_n5651), .B(new_n5652), .Y(new_n5653));
  MAJIxp5_ASAP7_75t_L       g05397(.A(new_n5653), .B(new_n5349), .C(new_n5163), .Y(new_n5654));
  AOI21xp33_ASAP7_75t_L     g05398(.A1(new_n5648), .A2(new_n5633), .B(new_n5646), .Y(new_n5655));
  AOI211xp5_ASAP7_75t_L     g05399(.A1(new_n5617), .A2(new_n5620), .B(new_n5634), .C(new_n5644), .Y(new_n5656));
  OAI21xp33_ASAP7_75t_L     g05400(.A1(new_n5656), .A2(new_n5655), .B(new_n5654), .Y(new_n5657));
  NOR2xp33_ASAP7_75t_L      g05401(.A(new_n427), .B(new_n4142), .Y(new_n5658));
  AOI221xp5_ASAP7_75t_L     g05402(.A1(\b[5] ), .A2(new_n4402), .B1(\b[7] ), .B2(new_n4156), .C(new_n5658), .Y(new_n5659));
  O2A1O1Ixp33_ASAP7_75t_L   g05403(.A1(new_n4150), .A2(new_n456), .B(new_n5659), .C(new_n4145), .Y(new_n5660));
  NOR2xp33_ASAP7_75t_L      g05404(.A(new_n4145), .B(new_n5660), .Y(new_n5661));
  INVx1_ASAP7_75t_L         g05405(.A(new_n5661), .Y(new_n5662));
  O2A1O1Ixp33_ASAP7_75t_L   g05406(.A1(new_n4150), .A2(new_n456), .B(new_n5659), .C(\a[35] ), .Y(new_n5663));
  INVx1_ASAP7_75t_L         g05407(.A(new_n5663), .Y(new_n5664));
  NAND4xp25_ASAP7_75t_L     g05408(.A(new_n5650), .B(new_n5664), .C(new_n5662), .D(new_n5657), .Y(new_n5665));
  NOR3xp33_ASAP7_75t_L      g05409(.A(new_n5654), .B(new_n5656), .C(new_n5655), .Y(new_n5666));
  AOI21xp33_ASAP7_75t_L     g05410(.A1(new_n5649), .A2(new_n5645), .B(new_n5614), .Y(new_n5667));
  OAI21xp33_ASAP7_75t_L     g05411(.A1(new_n4145), .A2(new_n5660), .B(new_n5664), .Y(new_n5668));
  OAI21xp33_ASAP7_75t_L     g05412(.A1(new_n5666), .A2(new_n5667), .B(new_n5668), .Y(new_n5669));
  NAND2xp33_ASAP7_75t_L     g05413(.A(new_n5669), .B(new_n5665), .Y(new_n5670));
  NAND2xp33_ASAP7_75t_L     g05414(.A(new_n5362), .B(new_n5361), .Y(new_n5671));
  MAJIxp5_ASAP7_75t_L       g05415(.A(new_n5375), .B(new_n5368), .C(new_n5671), .Y(new_n5672));
  NOR2xp33_ASAP7_75t_L      g05416(.A(new_n5670), .B(new_n5672), .Y(new_n5673));
  NAND3xp33_ASAP7_75t_L     g05417(.A(new_n5650), .B(new_n5657), .C(new_n5668), .Y(new_n5674));
  NOR3xp33_ASAP7_75t_L      g05418(.A(new_n5667), .B(new_n5666), .C(new_n5668), .Y(new_n5675));
  O2A1O1Ixp33_ASAP7_75t_L   g05419(.A1(new_n5661), .A2(new_n5663), .B(new_n5674), .C(new_n5675), .Y(new_n5676));
  O2A1O1Ixp33_ASAP7_75t_L   g05420(.A1(new_n5671), .A2(new_n5368), .B(new_n5384), .C(new_n5676), .Y(new_n5677));
  NOR2xp33_ASAP7_75t_L      g05421(.A(new_n590), .B(new_n3509), .Y(new_n5678));
  AOI221xp5_ASAP7_75t_L     g05422(.A1(\b[8] ), .A2(new_n3708), .B1(\b[10] ), .B2(new_n3503), .C(new_n5678), .Y(new_n5679));
  O2A1O1Ixp33_ASAP7_75t_L   g05423(.A1(new_n3513), .A2(new_n1175), .B(new_n5679), .C(new_n3493), .Y(new_n5680));
  INVx1_ASAP7_75t_L         g05424(.A(new_n5680), .Y(new_n5681));
  O2A1O1Ixp33_ASAP7_75t_L   g05425(.A1(new_n3513), .A2(new_n1175), .B(new_n5679), .C(\a[32] ), .Y(new_n5682));
  AOI21xp33_ASAP7_75t_L     g05426(.A1(new_n5681), .A2(\a[32] ), .B(new_n5682), .Y(new_n5683));
  NOR3xp33_ASAP7_75t_L      g05427(.A(new_n5677), .B(new_n5683), .C(new_n5673), .Y(new_n5684));
  NOR2xp33_ASAP7_75t_L      g05428(.A(new_n5370), .B(new_n5371), .Y(new_n5685));
  NOR2xp33_ASAP7_75t_L      g05429(.A(new_n5368), .B(new_n5671), .Y(new_n5686));
  O2A1O1Ixp33_ASAP7_75t_L   g05430(.A1(new_n5378), .A2(new_n5685), .B(new_n5383), .C(new_n5686), .Y(new_n5687));
  NAND2xp33_ASAP7_75t_L     g05431(.A(new_n5676), .B(new_n5687), .Y(new_n5688));
  A2O1A1Ixp33_ASAP7_75t_L   g05432(.A1(new_n5372), .A2(new_n5685), .B(new_n5394), .C(new_n5670), .Y(new_n5689));
  INVx1_ASAP7_75t_L         g05433(.A(new_n5683), .Y(new_n5690));
  AOI21xp33_ASAP7_75t_L     g05434(.A1(new_n5688), .A2(new_n5689), .B(new_n5690), .Y(new_n5691));
  OAI21xp33_ASAP7_75t_L     g05435(.A1(new_n5684), .A2(new_n5691), .B(new_n5612), .Y(new_n5692));
  NAND3xp33_ASAP7_75t_L     g05436(.A(new_n5688), .B(new_n5690), .C(new_n5689), .Y(new_n5693));
  OAI21xp33_ASAP7_75t_L     g05437(.A1(new_n5673), .A2(new_n5677), .B(new_n5683), .Y(new_n5694));
  NAND4xp25_ASAP7_75t_L     g05438(.A(new_n5400), .B(new_n5693), .C(new_n5694), .D(new_n5611), .Y(new_n5695));
  NOR2xp33_ASAP7_75t_L      g05439(.A(new_n833), .B(new_n2925), .Y(new_n5696));
  AOI221xp5_ASAP7_75t_L     g05440(.A1(\b[11] ), .A2(new_n3129), .B1(\b[13] ), .B2(new_n2938), .C(new_n5696), .Y(new_n5697));
  INVx1_ASAP7_75t_L         g05441(.A(new_n5697), .Y(new_n5698));
  A2O1A1Ixp33_ASAP7_75t_L   g05442(.A1(new_n1166), .A2(new_n2932), .B(new_n5698), .C(\a[29] ), .Y(new_n5699));
  O2A1O1Ixp33_ASAP7_75t_L   g05443(.A1(new_n2940), .A2(new_n942), .B(new_n5697), .C(\a[29] ), .Y(new_n5700));
  AOI21xp33_ASAP7_75t_L     g05444(.A1(new_n5699), .A2(\a[29] ), .B(new_n5700), .Y(new_n5701));
  NAND3xp33_ASAP7_75t_L     g05445(.A(new_n5695), .B(new_n5692), .C(new_n5701), .Y(new_n5702));
  AOI22xp33_ASAP7_75t_L     g05446(.A1(new_n5693), .A2(new_n5694), .B1(new_n5611), .B2(new_n5400), .Y(new_n5703));
  AOI21xp33_ASAP7_75t_L     g05447(.A1(new_n5612), .A2(new_n5694), .B(new_n5684), .Y(new_n5704));
  O2A1O1Ixp33_ASAP7_75t_L   g05448(.A1(new_n2940), .A2(new_n942), .B(new_n5697), .C(new_n2928), .Y(new_n5705));
  A2O1A1Ixp33_ASAP7_75t_L   g05449(.A1(new_n1166), .A2(new_n2932), .B(new_n5698), .C(new_n2928), .Y(new_n5706));
  OAI21xp33_ASAP7_75t_L     g05450(.A1(new_n2928), .A2(new_n5705), .B(new_n5706), .Y(new_n5707));
  A2O1A1Ixp33_ASAP7_75t_L   g05451(.A1(new_n5704), .A2(new_n5694), .B(new_n5703), .C(new_n5707), .Y(new_n5708));
  NAND2xp33_ASAP7_75t_L     g05452(.A(new_n5702), .B(new_n5708), .Y(new_n5709));
  NOR2xp33_ASAP7_75t_L      g05453(.A(new_n5610), .B(new_n5709), .Y(new_n5710));
  AOI221xp5_ASAP7_75t_L     g05454(.A1(new_n5414), .A2(new_n5416), .B1(new_n5702), .B2(new_n5708), .C(new_n5413), .Y(new_n5711));
  NOR2xp33_ASAP7_75t_L      g05455(.A(new_n1043), .B(new_n2410), .Y(new_n5712));
  AOI221xp5_ASAP7_75t_L     g05456(.A1(\b[14] ), .A2(new_n2577), .B1(\b[16] ), .B2(new_n2423), .C(new_n5712), .Y(new_n5713));
  OAI211xp5_ASAP7_75t_L     g05457(.A1(new_n2425), .A2(new_n1161), .B(\a[26] ), .C(new_n5713), .Y(new_n5714));
  INVx1_ASAP7_75t_L         g05458(.A(new_n5713), .Y(new_n5715));
  A2O1A1Ixp33_ASAP7_75t_L   g05459(.A1(new_n1156), .A2(new_n2417), .B(new_n5715), .C(new_n2413), .Y(new_n5716));
  NAND2xp33_ASAP7_75t_L     g05460(.A(new_n5716), .B(new_n5714), .Y(new_n5717));
  NOR3xp33_ASAP7_75t_L      g05461(.A(new_n5710), .B(new_n5711), .C(new_n5717), .Y(new_n5718));
  A2O1A1Ixp33_ASAP7_75t_L   g05462(.A1(new_n5200), .A2(new_n5419), .B(new_n5407), .C(new_n5430), .Y(new_n5719));
  NOR3xp33_ASAP7_75t_L      g05463(.A(new_n5612), .B(new_n5691), .C(new_n5684), .Y(new_n5720));
  NOR3xp33_ASAP7_75t_L      g05464(.A(new_n5703), .B(new_n5720), .C(new_n5707), .Y(new_n5721));
  AOI21xp33_ASAP7_75t_L     g05465(.A1(new_n5695), .A2(new_n5692), .B(new_n5701), .Y(new_n5722));
  NOR2xp33_ASAP7_75t_L      g05466(.A(new_n5722), .B(new_n5721), .Y(new_n5723));
  NAND2xp33_ASAP7_75t_L     g05467(.A(new_n5723), .B(new_n5719), .Y(new_n5724));
  NAND2xp33_ASAP7_75t_L     g05468(.A(new_n5610), .B(new_n5709), .Y(new_n5725));
  A2O1A1Ixp33_ASAP7_75t_L   g05469(.A1(new_n1156), .A2(new_n2417), .B(new_n5715), .C(\a[26] ), .Y(new_n5726));
  O2A1O1Ixp33_ASAP7_75t_L   g05470(.A1(new_n2425), .A2(new_n1161), .B(new_n5713), .C(\a[26] ), .Y(new_n5727));
  AOI21xp33_ASAP7_75t_L     g05471(.A1(new_n5726), .A2(\a[26] ), .B(new_n5727), .Y(new_n5728));
  AOI21xp33_ASAP7_75t_L     g05472(.A1(new_n5724), .A2(new_n5725), .B(new_n5728), .Y(new_n5729));
  NOR2xp33_ASAP7_75t_L      g05473(.A(new_n5718), .B(new_n5729), .Y(new_n5730));
  A2O1A1O1Ixp25_ASAP7_75t_L g05474(.A1(new_n5199), .A2(new_n5127), .B(new_n5454), .C(new_n5438), .D(new_n5442), .Y(new_n5731));
  NAND2xp33_ASAP7_75t_L     g05475(.A(new_n5730), .B(new_n5731), .Y(new_n5732));
  NAND3xp33_ASAP7_75t_L     g05476(.A(new_n5724), .B(new_n5725), .C(new_n5728), .Y(new_n5733));
  OAI21xp33_ASAP7_75t_L     g05477(.A1(new_n5711), .A2(new_n5710), .B(new_n5717), .Y(new_n5734));
  NAND2xp33_ASAP7_75t_L     g05478(.A(new_n5733), .B(new_n5734), .Y(new_n5735));
  A2O1A1Ixp33_ASAP7_75t_L   g05479(.A1(new_n5438), .A2(new_n5440), .B(new_n5442), .C(new_n5735), .Y(new_n5736));
  NOR2xp33_ASAP7_75t_L      g05480(.A(new_n1458), .B(new_n1962), .Y(new_n5737));
  AOI221xp5_ASAP7_75t_L     g05481(.A1(new_n1955), .A2(\b[19] ), .B1(new_n2093), .B2(\b[17] ), .C(new_n5737), .Y(new_n5738));
  INVx1_ASAP7_75t_L         g05482(.A(new_n5738), .Y(new_n5739));
  A2O1A1Ixp33_ASAP7_75t_L   g05483(.A1(new_n1607), .A2(new_n1964), .B(new_n5739), .C(\a[23] ), .Y(new_n5740));
  O2A1O1Ixp33_ASAP7_75t_L   g05484(.A1(new_n1956), .A2(new_n1628), .B(new_n5738), .C(\a[23] ), .Y(new_n5741));
  AOI21xp33_ASAP7_75t_L     g05485(.A1(new_n5740), .A2(\a[23] ), .B(new_n5741), .Y(new_n5742));
  NAND3xp33_ASAP7_75t_L     g05486(.A(new_n5732), .B(new_n5736), .C(new_n5742), .Y(new_n5743));
  AO21x2_ASAP7_75t_L        g05487(.A1(new_n5736), .A2(new_n5732), .B(new_n5742), .Y(new_n5744));
  AOI21xp33_ASAP7_75t_L     g05488(.A1(new_n5452), .A2(new_n5456), .B(new_n5449), .Y(new_n5745));
  A2O1A1O1Ixp25_ASAP7_75t_L g05489(.A1(new_n5224), .A2(new_n5221), .B(new_n5343), .C(new_n5457), .D(new_n5745), .Y(new_n5746));
  NAND3xp33_ASAP7_75t_L     g05490(.A(new_n5746), .B(new_n5743), .C(new_n5744), .Y(new_n5747));
  AO21x2_ASAP7_75t_L        g05491(.A1(new_n5743), .A2(new_n5744), .B(new_n5746), .Y(new_n5748));
  NOR2xp33_ASAP7_75t_L      g05492(.A(new_n1895), .B(new_n1517), .Y(new_n5749));
  AOI221xp5_ASAP7_75t_L     g05493(.A1(\b[20] ), .A2(new_n1659), .B1(\b[22] ), .B2(new_n1511), .C(new_n5749), .Y(new_n5750));
  INVx1_ASAP7_75t_L         g05494(.A(new_n5750), .Y(new_n5751));
  A2O1A1Ixp33_ASAP7_75t_L   g05495(.A1(new_n2056), .A2(new_n1513), .B(new_n5751), .C(\a[20] ), .Y(new_n5752));
  O2A1O1Ixp33_ASAP7_75t_L   g05496(.A1(new_n1521), .A2(new_n2522), .B(new_n5750), .C(\a[20] ), .Y(new_n5753));
  AOI21xp33_ASAP7_75t_L     g05497(.A1(new_n5752), .A2(\a[20] ), .B(new_n5753), .Y(new_n5754));
  NAND3xp33_ASAP7_75t_L     g05498(.A(new_n5748), .B(new_n5747), .C(new_n5754), .Y(new_n5755));
  AND3x1_ASAP7_75t_L        g05499(.A(new_n5746), .B(new_n5744), .C(new_n5743), .Y(new_n5756));
  AOI21xp33_ASAP7_75t_L     g05500(.A1(new_n5743), .A2(new_n5744), .B(new_n5746), .Y(new_n5757));
  O2A1O1Ixp33_ASAP7_75t_L   g05501(.A1(new_n1521), .A2(new_n2522), .B(new_n5750), .C(new_n1501), .Y(new_n5758));
  INVx1_ASAP7_75t_L         g05502(.A(new_n5753), .Y(new_n5759));
  OAI21xp33_ASAP7_75t_L     g05503(.A1(new_n1501), .A2(new_n5758), .B(new_n5759), .Y(new_n5760));
  OAI21xp33_ASAP7_75t_L     g05504(.A1(new_n5757), .A2(new_n5756), .B(new_n5760), .Y(new_n5761));
  NAND2xp33_ASAP7_75t_L     g05505(.A(new_n5755), .B(new_n5761), .Y(new_n5762));
  NAND2xp33_ASAP7_75t_L     g05506(.A(new_n5458), .B(new_n5462), .Y(new_n5763));
  MAJIxp5_ASAP7_75t_L       g05507(.A(new_n5477), .B(new_n5763), .C(new_n5468), .Y(new_n5764));
  NOR2xp33_ASAP7_75t_L      g05508(.A(new_n5764), .B(new_n5762), .Y(new_n5765));
  INVx1_ASAP7_75t_L         g05509(.A(new_n5763), .Y(new_n5766));
  A2O1A1Ixp33_ASAP7_75t_L   g05510(.A1(\a[20] ), .A2(new_n5466), .B(new_n5467), .C(new_n5766), .Y(new_n5767));
  NAND3xp33_ASAP7_75t_L     g05511(.A(new_n5748), .B(new_n5747), .C(new_n5760), .Y(new_n5768));
  NOR3xp33_ASAP7_75t_L      g05512(.A(new_n5756), .B(new_n5757), .C(new_n5760), .Y(new_n5769));
  AOI21xp33_ASAP7_75t_L     g05513(.A1(new_n5768), .A2(new_n5760), .B(new_n5769), .Y(new_n5770));
  AOI21xp33_ASAP7_75t_L     g05514(.A1(new_n5487), .A2(new_n5767), .B(new_n5770), .Y(new_n5771));
  NAND2xp33_ASAP7_75t_L     g05515(.A(\b[24] ), .B(new_n1204), .Y(new_n5772));
  OAI221xp5_ASAP7_75t_L     g05516(.A1(new_n1284), .A2(new_n2377), .B1(new_n2188), .B2(new_n1285), .C(new_n5772), .Y(new_n5773));
  A2O1A1Ixp33_ASAP7_75t_L   g05517(.A1(new_n5001), .A2(new_n1216), .B(new_n5773), .C(\a[17] ), .Y(new_n5774));
  AOI211xp5_ASAP7_75t_L     g05518(.A1(new_n5001), .A2(new_n1216), .B(new_n5773), .C(new_n1206), .Y(new_n5775));
  A2O1A1O1Ixp25_ASAP7_75t_L g05519(.A1(new_n5001), .A2(new_n1216), .B(new_n5773), .C(new_n5774), .D(new_n5775), .Y(new_n5776));
  INVx1_ASAP7_75t_L         g05520(.A(new_n5776), .Y(new_n5777));
  NOR3xp33_ASAP7_75t_L      g05521(.A(new_n5771), .B(new_n5777), .C(new_n5765), .Y(new_n5778));
  NAND3xp33_ASAP7_75t_L     g05522(.A(new_n5770), .B(new_n5487), .C(new_n5767), .Y(new_n5779));
  A2O1A1Ixp33_ASAP7_75t_L   g05523(.A1(new_n5768), .A2(new_n5760), .B(new_n5769), .C(new_n5764), .Y(new_n5780));
  AOI21xp33_ASAP7_75t_L     g05524(.A1(new_n5779), .A2(new_n5780), .B(new_n5776), .Y(new_n5781));
  A2O1A1Ixp33_ASAP7_75t_L   g05525(.A1(new_n5492), .A2(new_n4999), .B(new_n5118), .C(new_n5260), .Y(new_n5782));
  A2O1A1Ixp33_ASAP7_75t_L   g05526(.A1(new_n5782), .A2(new_n5259), .B(new_n5494), .C(new_n5490), .Y(new_n5783));
  OAI21xp33_ASAP7_75t_L     g05527(.A1(new_n5781), .A2(new_n5778), .B(new_n5783), .Y(new_n5784));
  NAND3xp33_ASAP7_75t_L     g05528(.A(new_n5779), .B(new_n5780), .C(new_n5776), .Y(new_n5785));
  OAI21xp33_ASAP7_75t_L     g05529(.A1(new_n5765), .A2(new_n5771), .B(new_n5777), .Y(new_n5786));
  A2O1A1Ixp33_ASAP7_75t_L   g05530(.A1(new_n5120), .A2(new_n5125), .B(new_n4993), .C(new_n4989), .Y(new_n5787));
  A2O1A1O1Ixp25_ASAP7_75t_L g05531(.A1(new_n5260), .A2(new_n5787), .B(new_n5247), .C(new_n5485), .D(new_n5495), .Y(new_n5788));
  NAND3xp33_ASAP7_75t_L     g05532(.A(new_n5788), .B(new_n5786), .C(new_n5785), .Y(new_n5789));
  AOI21xp33_ASAP7_75t_L     g05533(.A1(new_n5789), .A2(new_n5784), .B(new_n5607), .Y(new_n5790));
  XNOR2x2_ASAP7_75t_L       g05534(.A(\a[14] ), .B(new_n5606), .Y(new_n5791));
  AOI21xp33_ASAP7_75t_L     g05535(.A1(new_n5786), .A2(new_n5785), .B(new_n5788), .Y(new_n5792));
  NOR3xp33_ASAP7_75t_L      g05536(.A(new_n5783), .B(new_n5781), .C(new_n5778), .Y(new_n5793));
  NOR3xp33_ASAP7_75t_L      g05537(.A(new_n5792), .B(new_n5793), .C(new_n5791), .Y(new_n5794));
  NOR2xp33_ASAP7_75t_L      g05538(.A(new_n5794), .B(new_n5790), .Y(new_n5795));
  NAND2xp33_ASAP7_75t_L     g05539(.A(new_n5604), .B(new_n5795), .Y(new_n5796));
  AOI21xp33_ASAP7_75t_L     g05540(.A1(new_n5512), .A2(new_n5510), .B(new_n5514), .Y(new_n5797));
  OAI21xp33_ASAP7_75t_L     g05541(.A1(new_n5793), .A2(new_n5792), .B(new_n5791), .Y(new_n5798));
  NAND3xp33_ASAP7_75t_L     g05542(.A(new_n5789), .B(new_n5784), .C(new_n5607), .Y(new_n5799));
  NAND2xp33_ASAP7_75t_L     g05543(.A(new_n5799), .B(new_n5798), .Y(new_n5800));
  NAND2xp33_ASAP7_75t_L     g05544(.A(new_n5800), .B(new_n5797), .Y(new_n5801));
  NOR2xp33_ASAP7_75t_L      g05545(.A(new_n3456), .B(new_n1550), .Y(new_n5802));
  AOI221xp5_ASAP7_75t_L     g05546(.A1(\b[29] ), .A2(new_n713), .B1(\b[31] ), .B2(new_n640), .C(new_n5802), .Y(new_n5803));
  O2A1O1Ixp33_ASAP7_75t_L   g05547(.A1(new_n641), .A2(new_n3681), .B(new_n5803), .C(new_n637), .Y(new_n5804));
  INVx1_ASAP7_75t_L         g05548(.A(new_n5804), .Y(new_n5805));
  O2A1O1Ixp33_ASAP7_75t_L   g05549(.A1(new_n641), .A2(new_n3681), .B(new_n5803), .C(\a[11] ), .Y(new_n5806));
  AOI21xp33_ASAP7_75t_L     g05550(.A1(new_n5805), .A2(\a[11] ), .B(new_n5806), .Y(new_n5807));
  NAND3xp33_ASAP7_75t_L     g05551(.A(new_n5796), .B(new_n5801), .C(new_n5807), .Y(new_n5808));
  OAI21xp33_ASAP7_75t_L     g05552(.A1(new_n5790), .A2(new_n5794), .B(new_n5604), .Y(new_n5809));
  NOR3xp33_ASAP7_75t_L      g05553(.A(new_n5792), .B(new_n5793), .C(new_n5607), .Y(new_n5810));
  O2A1O1Ixp33_ASAP7_75t_L   g05554(.A1(new_n5607), .A2(new_n5810), .B(new_n5799), .C(new_n5604), .Y(new_n5811));
  INVx1_ASAP7_75t_L         g05555(.A(new_n5806), .Y(new_n5812));
  OAI21xp33_ASAP7_75t_L     g05556(.A1(new_n637), .A2(new_n5804), .B(new_n5812), .Y(new_n5813));
  A2O1A1Ixp33_ASAP7_75t_L   g05557(.A1(new_n5809), .A2(new_n5604), .B(new_n5811), .C(new_n5813), .Y(new_n5814));
  NAND3xp33_ASAP7_75t_L     g05558(.A(new_n5603), .B(new_n5808), .C(new_n5814), .Y(new_n5815));
  A2O1A1O1Ixp25_ASAP7_75t_L g05559(.A1(new_n5275), .A2(new_n5111), .B(new_n5276), .C(new_n5527), .D(new_n5530), .Y(new_n5816));
  A2O1A1O1Ixp25_ASAP7_75t_L g05560(.A1(new_n5500), .A2(\a[14] ), .B(new_n5501), .C(new_n5513), .D(new_n5524), .Y(new_n5817));
  O2A1O1Ixp33_ASAP7_75t_L   g05561(.A1(new_n5523), .A2(new_n5817), .B(new_n5513), .C(new_n5800), .Y(new_n5818));
  NOR3xp33_ASAP7_75t_L      g05562(.A(new_n5818), .B(new_n5811), .C(new_n5813), .Y(new_n5819));
  AOI21xp33_ASAP7_75t_L     g05563(.A1(new_n5796), .A2(new_n5801), .B(new_n5807), .Y(new_n5820));
  OAI21xp33_ASAP7_75t_L     g05564(.A1(new_n5819), .A2(new_n5820), .B(new_n5816), .Y(new_n5821));
  AOI21xp33_ASAP7_75t_L     g05565(.A1(new_n5815), .A2(new_n5821), .B(new_n5602), .Y(new_n5822));
  A2O1A1Ixp33_ASAP7_75t_L   g05566(.A1(new_n5599), .A2(new_n483), .B(new_n5600), .C(\a[8] ), .Y(new_n5823));
  O2A1O1Ixp33_ASAP7_75t_L   g05567(.A1(new_n477), .A2(new_n4352), .B(new_n5597), .C(\a[8] ), .Y(new_n5824));
  AOI21xp33_ASAP7_75t_L     g05568(.A1(new_n5823), .A2(\a[8] ), .B(new_n5824), .Y(new_n5825));
  NOR3xp33_ASAP7_75t_L      g05569(.A(new_n5816), .B(new_n5819), .C(new_n5820), .Y(new_n5826));
  AOI21xp33_ASAP7_75t_L     g05570(.A1(new_n5814), .A2(new_n5808), .B(new_n5603), .Y(new_n5827));
  NOR3xp33_ASAP7_75t_L      g05571(.A(new_n5826), .B(new_n5827), .C(new_n5825), .Y(new_n5828));
  NOR2xp33_ASAP7_75t_L      g05572(.A(new_n5822), .B(new_n5828), .Y(new_n5829));
  A2O1A1Ixp33_ASAP7_75t_L   g05573(.A1(new_n5547), .A2(new_n5554), .B(new_n5557), .C(new_n5829), .Y(new_n5830));
  NOR2xp33_ASAP7_75t_L      g05574(.A(new_n5540), .B(new_n5541), .Y(new_n5831));
  A2O1A1Ixp33_ASAP7_75t_L   g05575(.A1(\a[8] ), .A2(new_n5536), .B(new_n5537), .C(new_n5831), .Y(new_n5832));
  OAI221xp5_ASAP7_75t_L     g05576(.A1(new_n5822), .A2(new_n5828), .B1(new_n5546), .B2(new_n5544), .C(new_n5832), .Y(new_n5833));
  NOR2xp33_ASAP7_75t_L      g05577(.A(new_n4581), .B(new_n375), .Y(new_n5834));
  AOI221xp5_ASAP7_75t_L     g05578(.A1(\b[37] ), .A2(new_n361), .B1(new_n349), .B2(\b[36] ), .C(new_n5834), .Y(new_n5835));
  O2A1O1Ixp33_ASAP7_75t_L   g05579(.A1(new_n356), .A2(new_n5083), .B(new_n5835), .C(new_n346), .Y(new_n5836));
  O2A1O1Ixp33_ASAP7_75t_L   g05580(.A1(new_n356), .A2(new_n5083), .B(new_n5835), .C(\a[5] ), .Y(new_n5837));
  INVx1_ASAP7_75t_L         g05581(.A(new_n5837), .Y(new_n5838));
  OA21x2_ASAP7_75t_L        g05582(.A1(new_n346), .A2(new_n5836), .B(new_n5838), .Y(new_n5839));
  NAND3xp33_ASAP7_75t_L     g05583(.A(new_n5830), .B(new_n5833), .C(new_n5839), .Y(new_n5840));
  OAI21xp33_ASAP7_75t_L     g05584(.A1(new_n5827), .A2(new_n5826), .B(new_n5825), .Y(new_n5841));
  NAND3xp33_ASAP7_75t_L     g05585(.A(new_n5815), .B(new_n5602), .C(new_n5821), .Y(new_n5842));
  NAND2xp33_ASAP7_75t_L     g05586(.A(new_n5842), .B(new_n5841), .Y(new_n5843));
  O2A1O1Ixp33_ASAP7_75t_L   g05587(.A1(new_n5546), .A2(new_n5544), .B(new_n5832), .C(new_n5843), .Y(new_n5844));
  AOI221xp5_ASAP7_75t_L     g05588(.A1(new_n5842), .A2(new_n5841), .B1(new_n5547), .B2(new_n5554), .C(new_n5557), .Y(new_n5845));
  OAI21xp33_ASAP7_75t_L     g05589(.A1(new_n346), .A2(new_n5836), .B(new_n5838), .Y(new_n5846));
  OAI21xp33_ASAP7_75t_L     g05590(.A1(new_n5845), .A2(new_n5844), .B(new_n5846), .Y(new_n5847));
  NAND3xp33_ASAP7_75t_L     g05591(.A(new_n5595), .B(new_n5840), .C(new_n5847), .Y(new_n5848));
  A2O1A1O1Ixp25_ASAP7_75t_L g05592(.A1(new_n5303), .A2(new_n5302), .B(new_n5300), .C(new_n5552), .D(new_n5564), .Y(new_n5849));
  NAND2xp33_ASAP7_75t_L     g05593(.A(new_n5847), .B(new_n5840), .Y(new_n5850));
  NAND2xp33_ASAP7_75t_L     g05594(.A(new_n5849), .B(new_n5850), .Y(new_n5851));
  NOR2xp33_ASAP7_75t_L      g05595(.A(new_n5311), .B(new_n287), .Y(new_n5852));
  AOI221xp5_ASAP7_75t_L     g05596(.A1(\b[39] ), .A2(new_n264), .B1(\b[40] ), .B2(new_n283), .C(new_n5852), .Y(new_n5853));
  NOR2xp33_ASAP7_75t_L      g05597(.A(\b[39] ), .B(\b[40] ), .Y(new_n5854));
  INVx1_ASAP7_75t_L         g05598(.A(\b[40] ), .Y(new_n5855));
  NOR2xp33_ASAP7_75t_L      g05599(.A(new_n5570), .B(new_n5855), .Y(new_n5856));
  NOR2xp33_ASAP7_75t_L      g05600(.A(new_n5854), .B(new_n5856), .Y(new_n5857));
  A2O1A1Ixp33_ASAP7_75t_L   g05601(.A1(\b[39] ), .A2(\b[38] ), .B(new_n5574), .C(new_n5857), .Y(new_n5858));
  O2A1O1Ixp33_ASAP7_75t_L   g05602(.A1(new_n4613), .A2(new_n5074), .B(new_n5077), .C(new_n5316), .Y(new_n5859));
  O2A1O1Ixp33_ASAP7_75t_L   g05603(.A1(new_n5312), .A2(new_n5859), .B(new_n5572), .C(new_n5571), .Y(new_n5860));
  OAI21xp33_ASAP7_75t_L     g05604(.A1(new_n5854), .A2(new_n5856), .B(new_n5860), .Y(new_n5861));
  NAND2xp33_ASAP7_75t_L     g05605(.A(new_n5858), .B(new_n5861), .Y(new_n5862));
  O2A1O1Ixp33_ASAP7_75t_L   g05606(.A1(new_n279), .A2(new_n5862), .B(new_n5853), .C(new_n257), .Y(new_n5863));
  NOR2xp33_ASAP7_75t_L      g05607(.A(new_n257), .B(new_n5863), .Y(new_n5864));
  O2A1O1Ixp33_ASAP7_75t_L   g05608(.A1(new_n279), .A2(new_n5862), .B(new_n5853), .C(\a[2] ), .Y(new_n5865));
  NOR2xp33_ASAP7_75t_L      g05609(.A(new_n5865), .B(new_n5864), .Y(new_n5866));
  AOI21xp33_ASAP7_75t_L     g05610(.A1(new_n5848), .A2(new_n5851), .B(new_n5866), .Y(new_n5867));
  INVx1_ASAP7_75t_L         g05611(.A(new_n5867), .Y(new_n5868));
  NAND3xp33_ASAP7_75t_L     g05612(.A(new_n5848), .B(new_n5851), .C(new_n5866), .Y(new_n5869));
  NAND2xp33_ASAP7_75t_L     g05613(.A(new_n5869), .B(new_n5868), .Y(new_n5870));
  XOR2x2_ASAP7_75t_L        g05614(.A(new_n5870), .B(new_n5594), .Y(\f[40] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g05615(.A1(new_n5587), .A2(new_n5590), .B(new_n5593), .C(new_n5869), .D(new_n5867), .Y(new_n5872));
  NAND3xp33_ASAP7_75t_L     g05616(.A(new_n5830), .B(new_n5833), .C(new_n5846), .Y(new_n5873));
  A2O1A1Ixp33_ASAP7_75t_L   g05617(.A1(new_n5552), .A2(new_n5335), .B(new_n5564), .C(new_n5850), .Y(new_n5874));
  A2O1A1Ixp33_ASAP7_75t_L   g05618(.A1(new_n5543), .A2(new_n5555), .B(new_n5546), .C(new_n5832), .Y(new_n5875));
  A2O1A1O1Ixp25_ASAP7_75t_L g05619(.A1(new_n5527), .A2(new_n5336), .B(new_n5530), .C(new_n5808), .D(new_n5820), .Y(new_n5876));
  NOR2xp33_ASAP7_75t_L      g05620(.A(new_n3674), .B(new_n1550), .Y(new_n5877));
  AOI221xp5_ASAP7_75t_L     g05621(.A1(\b[30] ), .A2(new_n713), .B1(\b[32] ), .B2(new_n640), .C(new_n5877), .Y(new_n5878));
  O2A1O1Ixp33_ASAP7_75t_L   g05622(.A1(new_n641), .A2(new_n3897), .B(new_n5878), .C(new_n637), .Y(new_n5879));
  INVx1_ASAP7_75t_L         g05623(.A(new_n5878), .Y(new_n5880));
  A2O1A1Ixp33_ASAP7_75t_L   g05624(.A1(new_n3900), .A2(new_n718), .B(new_n5880), .C(new_n637), .Y(new_n5881));
  OAI21xp33_ASAP7_75t_L     g05625(.A1(new_n637), .A2(new_n5879), .B(new_n5881), .Y(new_n5882));
  INVx1_ASAP7_75t_L         g05626(.A(new_n5810), .Y(new_n5883));
  OAI21xp33_ASAP7_75t_L     g05627(.A1(new_n5797), .A2(new_n5795), .B(new_n5883), .Y(new_n5884));
  NOR2xp33_ASAP7_75t_L      g05628(.A(new_n3079), .B(new_n864), .Y(new_n5885));
  AOI221xp5_ASAP7_75t_L     g05629(.A1(\b[27] ), .A2(new_n985), .B1(\b[29] ), .B2(new_n886), .C(new_n5885), .Y(new_n5886));
  O2A1O1Ixp33_ASAP7_75t_L   g05630(.A1(new_n872), .A2(new_n3104), .B(new_n5886), .C(new_n867), .Y(new_n5887));
  INVx1_ASAP7_75t_L         g05631(.A(new_n5887), .Y(new_n5888));
  O2A1O1Ixp33_ASAP7_75t_L   g05632(.A1(new_n872), .A2(new_n3104), .B(new_n5886), .C(\a[14] ), .Y(new_n5889));
  AO21x2_ASAP7_75t_L        g05633(.A1(\a[14] ), .A2(new_n5888), .B(new_n5889), .Y(new_n5890));
  XOR2x2_ASAP7_75t_L        g05634(.A(new_n5764), .B(new_n5762), .Y(new_n5891));
  NAND2xp33_ASAP7_75t_L     g05635(.A(new_n5777), .B(new_n5891), .Y(new_n5892));
  A2O1A1Ixp33_ASAP7_75t_L   g05636(.A1(new_n5776), .A2(new_n5785), .B(new_n5788), .C(new_n5892), .Y(new_n5893));
  A2O1A1Ixp33_ASAP7_75t_L   g05637(.A1(new_n5487), .A2(new_n5767), .B(new_n5770), .C(new_n5768), .Y(new_n5894));
  NOR3xp33_ASAP7_75t_L      g05638(.A(new_n5710), .B(new_n5711), .C(new_n5728), .Y(new_n5895));
  INVx1_ASAP7_75t_L         g05639(.A(new_n5895), .Y(new_n5896));
  NOR2xp33_ASAP7_75t_L      g05640(.A(new_n1150), .B(new_n2410), .Y(new_n5897));
  AOI221xp5_ASAP7_75t_L     g05641(.A1(\b[15] ), .A2(new_n2577), .B1(\b[17] ), .B2(new_n2423), .C(new_n5897), .Y(new_n5898));
  INVx1_ASAP7_75t_L         g05642(.A(new_n5898), .Y(new_n5899));
  A2O1A1Ixp33_ASAP7_75t_L   g05643(.A1(new_n1633), .A2(new_n2417), .B(new_n5899), .C(\a[26] ), .Y(new_n5900));
  O2A1O1Ixp33_ASAP7_75t_L   g05644(.A1(new_n2425), .A2(new_n1356), .B(new_n5898), .C(\a[26] ), .Y(new_n5901));
  AOI21xp33_ASAP7_75t_L     g05645(.A1(new_n5900), .A2(\a[26] ), .B(new_n5901), .Y(new_n5902));
  A2O1A1O1Ixp25_ASAP7_75t_L g05646(.A1(new_n5429), .A2(new_n5416), .B(new_n5413), .C(new_n5702), .D(new_n5722), .Y(new_n5903));
  NOR2xp33_ASAP7_75t_L      g05647(.A(new_n960), .B(new_n2930), .Y(new_n5904));
  AOI221xp5_ASAP7_75t_L     g05648(.A1(\b[12] ), .A2(new_n3129), .B1(\b[13] ), .B2(new_n2936), .C(new_n5904), .Y(new_n5905));
  O2A1O1Ixp33_ASAP7_75t_L   g05649(.A1(new_n2940), .A2(new_n1268), .B(new_n5905), .C(new_n2928), .Y(new_n5906));
  O2A1O1Ixp33_ASAP7_75t_L   g05650(.A1(new_n2940), .A2(new_n1268), .B(new_n5905), .C(\a[29] ), .Y(new_n5907));
  INVx1_ASAP7_75t_L         g05651(.A(new_n5907), .Y(new_n5908));
  OAI21xp33_ASAP7_75t_L     g05652(.A1(new_n2928), .A2(new_n5906), .B(new_n5908), .Y(new_n5909));
  A2O1A1Ixp33_ASAP7_75t_L   g05653(.A1(new_n5400), .A2(new_n5611), .B(new_n5691), .C(new_n5693), .Y(new_n5910));
  INVx1_ASAP7_75t_L         g05654(.A(new_n5674), .Y(new_n5911));
  NOR2xp33_ASAP7_75t_L      g05655(.A(new_n448), .B(new_n4142), .Y(new_n5912));
  AOI221xp5_ASAP7_75t_L     g05656(.A1(\b[6] ), .A2(new_n4402), .B1(\b[8] ), .B2(new_n4156), .C(new_n5912), .Y(new_n5913));
  OAI211xp5_ASAP7_75t_L     g05657(.A1(new_n4150), .A2(new_n540), .B(\a[35] ), .C(new_n5913), .Y(new_n5914));
  INVx1_ASAP7_75t_L         g05658(.A(new_n5913), .Y(new_n5915));
  A2O1A1Ixp33_ASAP7_75t_L   g05659(.A1(new_n1684), .A2(new_n4151), .B(new_n5915), .C(new_n4145), .Y(new_n5916));
  NAND2xp33_ASAP7_75t_L     g05660(.A(new_n5914), .B(new_n5916), .Y(new_n5917));
  OAI21xp33_ASAP7_75t_L     g05661(.A1(new_n5655), .A2(new_n5654), .B(new_n5649), .Y(new_n5918));
  NOR2xp33_ASAP7_75t_L      g05662(.A(new_n289), .B(new_n5641), .Y(new_n5919));
  AND3x1_ASAP7_75t_L        g05663(.A(new_n5348), .B(new_n5628), .C(new_n5622), .Y(new_n5920));
  AOI221xp5_ASAP7_75t_L     g05664(.A1(new_n5623), .A2(\b[1] ), .B1(new_n5920), .B2(\b[0] ), .C(new_n5919), .Y(new_n5921));
  NOR2xp33_ASAP7_75t_L      g05665(.A(new_n5630), .B(new_n509), .Y(new_n5922));
  INVx1_ASAP7_75t_L         g05666(.A(new_n5922), .Y(new_n5923));
  NAND3xp33_ASAP7_75t_L     g05667(.A(new_n5921), .B(\a[41] ), .C(new_n5923), .Y(new_n5924));
  NAND3xp33_ASAP7_75t_L     g05668(.A(new_n5348), .B(new_n5622), .C(new_n5628), .Y(new_n5925));
  NAND2xp33_ASAP7_75t_L     g05669(.A(\b[1] ), .B(new_n5623), .Y(new_n5926));
  OAI221xp5_ASAP7_75t_L     g05670(.A1(new_n5641), .A2(new_n289), .B1(new_n284), .B2(new_n5925), .C(new_n5926), .Y(new_n5927));
  A2O1A1Ixp33_ASAP7_75t_L   g05671(.A1(new_n294), .A2(new_n5637), .B(new_n5927), .C(new_n5626), .Y(new_n5928));
  NAND3xp33_ASAP7_75t_L     g05672(.A(new_n5924), .B(new_n5633), .C(new_n5928), .Y(new_n5929));
  NAND5xp2_ASAP7_75t_L      g05673(.A(\a[41] ), .B(new_n5921), .C(new_n5632), .D(new_n5923), .E(new_n5613), .Y(new_n5930));
  NOR2xp33_ASAP7_75t_L      g05674(.A(new_n384), .B(new_n4908), .Y(new_n5931));
  AOI221xp5_ASAP7_75t_L     g05675(.A1(\b[3] ), .A2(new_n5139), .B1(\b[4] ), .B2(new_n4916), .C(new_n5931), .Y(new_n5932));
  OAI211xp5_ASAP7_75t_L     g05676(.A1(new_n4911), .A2(new_n728), .B(\a[38] ), .C(new_n5932), .Y(new_n5933));
  OAI21xp33_ASAP7_75t_L     g05677(.A1(new_n4911), .A2(new_n728), .B(new_n5932), .Y(new_n5934));
  NAND2xp33_ASAP7_75t_L     g05678(.A(new_n4906), .B(new_n5934), .Y(new_n5935));
  AND4x1_ASAP7_75t_L        g05679(.A(new_n5929), .B(new_n5935), .C(new_n5930), .D(new_n5933), .Y(new_n5936));
  AOI22xp33_ASAP7_75t_L     g05680(.A1(new_n5933), .A2(new_n5935), .B1(new_n5930), .B2(new_n5929), .Y(new_n5937));
  OAI21xp33_ASAP7_75t_L     g05681(.A1(new_n5936), .A2(new_n5937), .B(new_n5918), .Y(new_n5938));
  AOI21xp33_ASAP7_75t_L     g05682(.A1(new_n5614), .A2(new_n5645), .B(new_n5656), .Y(new_n5939));
  NOR2xp33_ASAP7_75t_L      g05683(.A(new_n5937), .B(new_n5936), .Y(new_n5940));
  NAND2xp33_ASAP7_75t_L     g05684(.A(new_n5940), .B(new_n5939), .Y(new_n5941));
  NAND3xp33_ASAP7_75t_L     g05685(.A(new_n5941), .B(new_n5917), .C(new_n5938), .Y(new_n5942));
  O2A1O1Ixp33_ASAP7_75t_L   g05686(.A1(new_n5654), .A2(new_n5655), .B(new_n5649), .C(new_n5940), .Y(new_n5943));
  NOR3xp33_ASAP7_75t_L      g05687(.A(new_n5918), .B(new_n5936), .C(new_n5937), .Y(new_n5944));
  NOR3xp33_ASAP7_75t_L      g05688(.A(new_n5943), .B(new_n5944), .C(new_n5917), .Y(new_n5945));
  AOI21xp33_ASAP7_75t_L     g05689(.A1(new_n5942), .A2(new_n5917), .B(new_n5945), .Y(new_n5946));
  A2O1A1Ixp33_ASAP7_75t_L   g05690(.A1(new_n5670), .A2(new_n5672), .B(new_n5911), .C(new_n5946), .Y(new_n5947));
  AOI21xp33_ASAP7_75t_L     g05691(.A1(new_n5672), .A2(new_n5670), .B(new_n5911), .Y(new_n5948));
  A2O1A1Ixp33_ASAP7_75t_L   g05692(.A1(new_n5917), .A2(new_n5942), .B(new_n5945), .C(new_n5948), .Y(new_n5949));
  NOR2xp33_ASAP7_75t_L      g05693(.A(new_n680), .B(new_n3509), .Y(new_n5950));
  AOI221xp5_ASAP7_75t_L     g05694(.A1(\b[9] ), .A2(new_n3708), .B1(\b[11] ), .B2(new_n3503), .C(new_n5950), .Y(new_n5951));
  O2A1O1Ixp33_ASAP7_75t_L   g05695(.A1(new_n3513), .A2(new_n754), .B(new_n5951), .C(new_n3493), .Y(new_n5952));
  INVx1_ASAP7_75t_L         g05696(.A(new_n5951), .Y(new_n5953));
  A2O1A1Ixp33_ASAP7_75t_L   g05697(.A1(new_n976), .A2(new_n3505), .B(new_n5953), .C(new_n3493), .Y(new_n5954));
  OAI21xp33_ASAP7_75t_L     g05698(.A1(new_n3493), .A2(new_n5952), .B(new_n5954), .Y(new_n5955));
  INVx1_ASAP7_75t_L         g05699(.A(new_n5955), .Y(new_n5956));
  NAND3xp33_ASAP7_75t_L     g05700(.A(new_n5949), .B(new_n5947), .C(new_n5956), .Y(new_n5957));
  OAI21xp33_ASAP7_75t_L     g05701(.A1(new_n5944), .A2(new_n5943), .B(new_n5917), .Y(new_n5958));
  NAND4xp25_ASAP7_75t_L     g05702(.A(new_n5941), .B(new_n5914), .C(new_n5916), .D(new_n5938), .Y(new_n5959));
  NAND2xp33_ASAP7_75t_L     g05703(.A(new_n5959), .B(new_n5958), .Y(new_n5960));
  A2O1A1Ixp33_ASAP7_75t_L   g05704(.A1(new_n5670), .A2(new_n5672), .B(new_n5911), .C(new_n5960), .Y(new_n5961));
  O2A1O1Ixp33_ASAP7_75t_L   g05705(.A1(new_n5676), .A2(new_n5687), .B(new_n5674), .C(new_n5960), .Y(new_n5962));
  A2O1A1Ixp33_ASAP7_75t_L   g05706(.A1(new_n5961), .A2(new_n5960), .B(new_n5962), .C(new_n5955), .Y(new_n5963));
  NAND3xp33_ASAP7_75t_L     g05707(.A(new_n5910), .B(new_n5957), .C(new_n5963), .Y(new_n5964));
  AOI211xp5_ASAP7_75t_L     g05708(.A1(new_n5961), .A2(new_n5960), .B(new_n5962), .C(new_n5955), .Y(new_n5965));
  AOI21xp33_ASAP7_75t_L     g05709(.A1(new_n5949), .A2(new_n5947), .B(new_n5956), .Y(new_n5966));
  OAI21xp33_ASAP7_75t_L     g05710(.A1(new_n5966), .A2(new_n5965), .B(new_n5704), .Y(new_n5967));
  AOI21xp33_ASAP7_75t_L     g05711(.A1(new_n5964), .A2(new_n5967), .B(new_n5909), .Y(new_n5968));
  OAI21xp33_ASAP7_75t_L     g05712(.A1(new_n2940), .A2(new_n1268), .B(new_n5905), .Y(new_n5969));
  NOR2xp33_ASAP7_75t_L      g05713(.A(new_n2928), .B(new_n5969), .Y(new_n5970));
  NOR2xp33_ASAP7_75t_L      g05714(.A(new_n5907), .B(new_n5970), .Y(new_n5971));
  NOR3xp33_ASAP7_75t_L      g05715(.A(new_n5704), .B(new_n5965), .C(new_n5966), .Y(new_n5972));
  AOI21xp33_ASAP7_75t_L     g05716(.A1(new_n5963), .A2(new_n5957), .B(new_n5910), .Y(new_n5973));
  NOR3xp33_ASAP7_75t_L      g05717(.A(new_n5971), .B(new_n5973), .C(new_n5972), .Y(new_n5974));
  NOR3xp33_ASAP7_75t_L      g05718(.A(new_n5903), .B(new_n5968), .C(new_n5974), .Y(new_n5975));
  OAI21xp33_ASAP7_75t_L     g05719(.A1(new_n5721), .A2(new_n5610), .B(new_n5708), .Y(new_n5976));
  OAI21xp33_ASAP7_75t_L     g05720(.A1(new_n5972), .A2(new_n5973), .B(new_n5971), .Y(new_n5977));
  NAND3xp33_ASAP7_75t_L     g05721(.A(new_n5909), .B(new_n5964), .C(new_n5967), .Y(new_n5978));
  AOI21xp33_ASAP7_75t_L     g05722(.A1(new_n5978), .A2(new_n5977), .B(new_n5976), .Y(new_n5979));
  OAI21xp33_ASAP7_75t_L     g05723(.A1(new_n5975), .A2(new_n5979), .B(new_n5902), .Y(new_n5980));
  INVx1_ASAP7_75t_L         g05724(.A(new_n5902), .Y(new_n5981));
  NAND3xp33_ASAP7_75t_L     g05725(.A(new_n5976), .B(new_n5977), .C(new_n5978), .Y(new_n5982));
  OAI21xp33_ASAP7_75t_L     g05726(.A1(new_n5968), .A2(new_n5974), .B(new_n5903), .Y(new_n5983));
  NAND3xp33_ASAP7_75t_L     g05727(.A(new_n5981), .B(new_n5982), .C(new_n5983), .Y(new_n5984));
  NAND2xp33_ASAP7_75t_L     g05728(.A(new_n5980), .B(new_n5984), .Y(new_n5985));
  O2A1O1Ixp33_ASAP7_75t_L   g05729(.A1(new_n5730), .A2(new_n5731), .B(new_n5896), .C(new_n5985), .Y(new_n5986));
  OAI21xp33_ASAP7_75t_L     g05730(.A1(new_n5730), .A2(new_n5731), .B(new_n5896), .Y(new_n5987));
  AOI21xp33_ASAP7_75t_L     g05731(.A1(new_n5982), .A2(new_n5983), .B(new_n5981), .Y(new_n5988));
  NOR3xp33_ASAP7_75t_L      g05732(.A(new_n5979), .B(new_n5975), .C(new_n5902), .Y(new_n5989));
  NOR2xp33_ASAP7_75t_L      g05733(.A(new_n5989), .B(new_n5988), .Y(new_n5990));
  NOR2xp33_ASAP7_75t_L      g05734(.A(new_n5990), .B(new_n5987), .Y(new_n5991));
  NOR2xp33_ASAP7_75t_L      g05735(.A(new_n1599), .B(new_n1962), .Y(new_n5992));
  AOI221xp5_ASAP7_75t_L     g05736(.A1(new_n1955), .A2(\b[20] ), .B1(new_n2093), .B2(\b[18] ), .C(new_n5992), .Y(new_n5993));
  O2A1O1Ixp33_ASAP7_75t_L   g05737(.A1(new_n1956), .A2(new_n1754), .B(new_n5993), .C(new_n1952), .Y(new_n5994));
  OAI21xp33_ASAP7_75t_L     g05738(.A1(new_n1956), .A2(new_n1754), .B(new_n5993), .Y(new_n5995));
  NAND2xp33_ASAP7_75t_L     g05739(.A(new_n1952), .B(new_n5995), .Y(new_n5996));
  OAI21xp33_ASAP7_75t_L     g05740(.A1(new_n1952), .A2(new_n5994), .B(new_n5996), .Y(new_n5997));
  NOR3xp33_ASAP7_75t_L      g05741(.A(new_n5991), .B(new_n5997), .C(new_n5986), .Y(new_n5998));
  MAJIxp5_ASAP7_75t_L       g05742(.A(new_n5455), .B(new_n5441), .C(new_n5427), .Y(new_n5999));
  A2O1A1Ixp33_ASAP7_75t_L   g05743(.A1(new_n5735), .A2(new_n5999), .B(new_n5895), .C(new_n5990), .Y(new_n6000));
  O2A1O1Ixp33_ASAP7_75t_L   g05744(.A1(new_n5718), .A2(new_n5729), .B(new_n5999), .C(new_n5895), .Y(new_n6001));
  NAND2xp33_ASAP7_75t_L     g05745(.A(new_n5985), .B(new_n6001), .Y(new_n6002));
  OA21x2_ASAP7_75t_L        g05746(.A1(new_n1952), .A2(new_n5994), .B(new_n5996), .Y(new_n6003));
  AOI21xp33_ASAP7_75t_L     g05747(.A1(new_n6000), .A2(new_n6002), .B(new_n6003), .Y(new_n6004));
  XNOR2x2_ASAP7_75t_L       g05748(.A(new_n5999), .B(new_n5735), .Y(new_n6005));
  MAJIxp5_ASAP7_75t_L       g05749(.A(new_n5746), .B(new_n6005), .C(new_n5742), .Y(new_n6006));
  NOR3xp33_ASAP7_75t_L      g05750(.A(new_n6006), .B(new_n6004), .C(new_n5998), .Y(new_n6007));
  OA21x2_ASAP7_75t_L        g05751(.A1(new_n5998), .A2(new_n6004), .B(new_n6006), .Y(new_n6008));
  NOR2xp33_ASAP7_75t_L      g05752(.A(new_n2045), .B(new_n1517), .Y(new_n6009));
  AOI221xp5_ASAP7_75t_L     g05753(.A1(\b[21] ), .A2(new_n1659), .B1(\b[23] ), .B2(new_n1511), .C(new_n6009), .Y(new_n6010));
  O2A1O1Ixp33_ASAP7_75t_L   g05754(.A1(new_n1521), .A2(new_n2194), .B(new_n6010), .C(new_n1501), .Y(new_n6011));
  INVx1_ASAP7_75t_L         g05755(.A(new_n6011), .Y(new_n6012));
  O2A1O1Ixp33_ASAP7_75t_L   g05756(.A1(new_n1521), .A2(new_n2194), .B(new_n6010), .C(\a[20] ), .Y(new_n6013));
  AOI21xp33_ASAP7_75t_L     g05757(.A1(new_n6012), .A2(\a[20] ), .B(new_n6013), .Y(new_n6014));
  NOR3xp33_ASAP7_75t_L      g05758(.A(new_n6014), .B(new_n6008), .C(new_n6007), .Y(new_n6015));
  OA21x2_ASAP7_75t_L        g05759(.A1(new_n6007), .A2(new_n6008), .B(new_n6014), .Y(new_n6016));
  OAI21xp33_ASAP7_75t_L     g05760(.A1(new_n6015), .A2(new_n6016), .B(new_n5894), .Y(new_n6017));
  INVx1_ASAP7_75t_L         g05761(.A(new_n5768), .Y(new_n6018));
  O2A1O1Ixp33_ASAP7_75t_L   g05762(.A1(new_n5769), .A2(new_n5760), .B(new_n5764), .C(new_n6018), .Y(new_n6019));
  INVx1_ASAP7_75t_L         g05763(.A(new_n6015), .Y(new_n6020));
  OAI21xp33_ASAP7_75t_L     g05764(.A1(new_n6007), .A2(new_n6008), .B(new_n6014), .Y(new_n6021));
  NAND3xp33_ASAP7_75t_L     g05765(.A(new_n6019), .B(new_n6020), .C(new_n6021), .Y(new_n6022));
  NOR2xp33_ASAP7_75t_L      g05766(.A(new_n2377), .B(new_n2118), .Y(new_n6023));
  AOI221xp5_ASAP7_75t_L     g05767(.A1(\b[24] ), .A2(new_n1290), .B1(\b[26] ), .B2(new_n1209), .C(new_n6023), .Y(new_n6024));
  O2A1O1Ixp33_ASAP7_75t_L   g05768(.A1(new_n1210), .A2(new_n2708), .B(new_n6024), .C(new_n1206), .Y(new_n6025));
  INVx1_ASAP7_75t_L         g05769(.A(new_n6025), .Y(new_n6026));
  O2A1O1Ixp33_ASAP7_75t_L   g05770(.A1(new_n1210), .A2(new_n2708), .B(new_n6024), .C(\a[17] ), .Y(new_n6027));
  AOI21xp33_ASAP7_75t_L     g05771(.A1(new_n6026), .A2(\a[17] ), .B(new_n6027), .Y(new_n6028));
  NAND3xp33_ASAP7_75t_L     g05772(.A(new_n6017), .B(new_n6022), .C(new_n6028), .Y(new_n6029));
  AOI21xp33_ASAP7_75t_L     g05773(.A1(new_n6021), .A2(new_n6020), .B(new_n6019), .Y(new_n6030));
  A2O1A1O1Ixp25_ASAP7_75t_L g05774(.A1(new_n5764), .A2(new_n5762), .B(new_n6018), .C(new_n6021), .D(new_n6015), .Y(new_n6031));
  INVx1_ASAP7_75t_L         g05775(.A(new_n6028), .Y(new_n6032));
  A2O1A1Ixp33_ASAP7_75t_L   g05776(.A1(new_n6031), .A2(new_n6021), .B(new_n6030), .C(new_n6032), .Y(new_n6033));
  NAND3xp33_ASAP7_75t_L     g05777(.A(new_n5893), .B(new_n6029), .C(new_n6033), .Y(new_n6034));
  NOR3xp33_ASAP7_75t_L      g05778(.A(new_n5771), .B(new_n5776), .C(new_n5765), .Y(new_n6035));
  O2A1O1Ixp33_ASAP7_75t_L   g05779(.A1(new_n5891), .A2(new_n5781), .B(new_n5783), .C(new_n6035), .Y(new_n6036));
  AOI211xp5_ASAP7_75t_L     g05780(.A1(new_n6031), .A2(new_n6021), .B(new_n6032), .C(new_n6030), .Y(new_n6037));
  A2O1A1O1Ixp25_ASAP7_75t_L g05781(.A1(new_n5487), .A2(new_n5767), .B(new_n5770), .C(new_n5768), .D(new_n6016), .Y(new_n6038));
  A2O1A1O1Ixp25_ASAP7_75t_L g05782(.A1(new_n6020), .A2(new_n6038), .B(new_n6019), .C(new_n6022), .D(new_n6028), .Y(new_n6039));
  OAI21xp33_ASAP7_75t_L     g05783(.A1(new_n6037), .A2(new_n6039), .B(new_n6036), .Y(new_n6040));
  AOI21xp33_ASAP7_75t_L     g05784(.A1(new_n6034), .A2(new_n6040), .B(new_n5890), .Y(new_n6041));
  AOI21xp33_ASAP7_75t_L     g05785(.A1(new_n5888), .A2(\a[14] ), .B(new_n5889), .Y(new_n6042));
  NOR3xp33_ASAP7_75t_L      g05786(.A(new_n6036), .B(new_n6037), .C(new_n6039), .Y(new_n6043));
  AOI21xp33_ASAP7_75t_L     g05787(.A1(new_n6033), .A2(new_n6029), .B(new_n5893), .Y(new_n6044));
  NOR3xp33_ASAP7_75t_L      g05788(.A(new_n6044), .B(new_n6043), .C(new_n6042), .Y(new_n6045));
  NOR2xp33_ASAP7_75t_L      g05789(.A(new_n6045), .B(new_n6041), .Y(new_n6046));
  NAND2xp33_ASAP7_75t_L     g05790(.A(new_n5884), .B(new_n6046), .Y(new_n6047));
  O2A1O1Ixp33_ASAP7_75t_L   g05791(.A1(new_n5790), .A2(new_n5794), .B(new_n5604), .C(new_n5810), .Y(new_n6048));
  OAI21xp33_ASAP7_75t_L     g05792(.A1(new_n6041), .A2(new_n6045), .B(new_n6048), .Y(new_n6049));
  AOI21xp33_ASAP7_75t_L     g05793(.A1(new_n6047), .A2(new_n6049), .B(new_n5882), .Y(new_n6050));
  INVx1_ASAP7_75t_L         g05794(.A(new_n5882), .Y(new_n6051));
  NOR3xp33_ASAP7_75t_L      g05795(.A(new_n6048), .B(new_n6041), .C(new_n6045), .Y(new_n6052));
  OAI21xp33_ASAP7_75t_L     g05796(.A1(new_n6043), .A2(new_n6044), .B(new_n6042), .Y(new_n6053));
  NAND3xp33_ASAP7_75t_L     g05797(.A(new_n6034), .B(new_n5890), .C(new_n6040), .Y(new_n6054));
  AOI221xp5_ASAP7_75t_L     g05798(.A1(new_n5800), .A2(new_n5604), .B1(new_n6054), .B2(new_n6053), .C(new_n5810), .Y(new_n6055));
  NOR3xp33_ASAP7_75t_L      g05799(.A(new_n6052), .B(new_n6051), .C(new_n6055), .Y(new_n6056));
  NOR3xp33_ASAP7_75t_L      g05800(.A(new_n5876), .B(new_n6050), .C(new_n6056), .Y(new_n6057));
  OAI21xp33_ASAP7_75t_L     g05801(.A1(new_n5819), .A2(new_n5816), .B(new_n5814), .Y(new_n6058));
  OAI21xp33_ASAP7_75t_L     g05802(.A1(new_n6055), .A2(new_n6052), .B(new_n6051), .Y(new_n6059));
  NAND3xp33_ASAP7_75t_L     g05803(.A(new_n6047), .B(new_n5882), .C(new_n6049), .Y(new_n6060));
  AOI21xp33_ASAP7_75t_L     g05804(.A1(new_n6060), .A2(new_n6059), .B(new_n6058), .Y(new_n6061));
  NOR2xp33_ASAP7_75t_L      g05805(.A(new_n4344), .B(new_n513), .Y(new_n6062));
  AOI221xp5_ASAP7_75t_L     g05806(.A1(\b[33] ), .A2(new_n560), .B1(\b[35] ), .B2(new_n475), .C(new_n6062), .Y(new_n6063));
  O2A1O1Ixp33_ASAP7_75t_L   g05807(.A1(new_n477), .A2(new_n4589), .B(new_n6063), .C(new_n466), .Y(new_n6064));
  O2A1O1Ixp33_ASAP7_75t_L   g05808(.A1(new_n477), .A2(new_n4589), .B(new_n6063), .C(\a[8] ), .Y(new_n6065));
  INVx1_ASAP7_75t_L         g05809(.A(new_n6065), .Y(new_n6066));
  OAI21xp33_ASAP7_75t_L     g05810(.A1(new_n466), .A2(new_n6064), .B(new_n6066), .Y(new_n6067));
  NOR3xp33_ASAP7_75t_L      g05811(.A(new_n6061), .B(new_n6057), .C(new_n6067), .Y(new_n6068));
  NAND3xp33_ASAP7_75t_L     g05812(.A(new_n6058), .B(new_n6059), .C(new_n6060), .Y(new_n6069));
  OAI21xp33_ASAP7_75t_L     g05813(.A1(new_n6056), .A2(new_n6050), .B(new_n5876), .Y(new_n6070));
  INVx1_ASAP7_75t_L         g05814(.A(new_n6064), .Y(new_n6071));
  AOI21xp33_ASAP7_75t_L     g05815(.A1(new_n6071), .A2(\a[8] ), .B(new_n6065), .Y(new_n6072));
  AOI21xp33_ASAP7_75t_L     g05816(.A1(new_n6069), .A2(new_n6070), .B(new_n6072), .Y(new_n6073));
  NOR2xp33_ASAP7_75t_L      g05817(.A(new_n6073), .B(new_n6068), .Y(new_n6074));
  A2O1A1Ixp33_ASAP7_75t_L   g05818(.A1(new_n5829), .A2(new_n5875), .B(new_n5828), .C(new_n6074), .Y(new_n6075));
  A2O1A1O1Ixp25_ASAP7_75t_L g05819(.A1(new_n5547), .A2(new_n5554), .B(new_n5557), .C(new_n5841), .D(new_n5828), .Y(new_n6076));
  NOR2xp33_ASAP7_75t_L      g05820(.A(new_n6057), .B(new_n6061), .Y(new_n6077));
  A2O1A1Ixp33_ASAP7_75t_L   g05821(.A1(\a[8] ), .A2(new_n6071), .B(new_n6065), .C(new_n6077), .Y(new_n6078));
  A2O1A1Ixp33_ASAP7_75t_L   g05822(.A1(new_n6078), .A2(new_n6077), .B(new_n6073), .C(new_n6076), .Y(new_n6079));
  NOR2xp33_ASAP7_75t_L      g05823(.A(new_n4613), .B(new_n375), .Y(new_n6080));
  AOI221xp5_ASAP7_75t_L     g05824(.A1(\b[38] ), .A2(new_n361), .B1(new_n349), .B2(\b[37] ), .C(new_n6080), .Y(new_n6081));
  O2A1O1Ixp33_ASAP7_75t_L   g05825(.A1(new_n356), .A2(new_n5318), .B(new_n6081), .C(new_n346), .Y(new_n6082));
  AND2x2_ASAP7_75t_L        g05826(.A(new_n5317), .B(new_n5314), .Y(new_n6083));
  INVx1_ASAP7_75t_L         g05827(.A(new_n6081), .Y(new_n6084));
  A2O1A1Ixp33_ASAP7_75t_L   g05828(.A1(new_n6083), .A2(new_n359), .B(new_n6084), .C(new_n346), .Y(new_n6085));
  OAI21xp33_ASAP7_75t_L     g05829(.A1(new_n346), .A2(new_n6082), .B(new_n6085), .Y(new_n6086));
  INVx1_ASAP7_75t_L         g05830(.A(new_n6086), .Y(new_n6087));
  AOI21xp33_ASAP7_75t_L     g05831(.A1(new_n6079), .A2(new_n6075), .B(new_n6087), .Y(new_n6088));
  A2O1A1O1Ixp25_ASAP7_75t_L g05832(.A1(new_n5298), .A2(new_n5289), .B(new_n5288), .C(new_n5547), .D(new_n5557), .Y(new_n6089));
  NAND3xp33_ASAP7_75t_L     g05833(.A(new_n6069), .B(new_n6072), .C(new_n6070), .Y(new_n6090));
  OAI21xp33_ASAP7_75t_L     g05834(.A1(new_n6057), .A2(new_n6061), .B(new_n6067), .Y(new_n6091));
  NAND2xp33_ASAP7_75t_L     g05835(.A(new_n6090), .B(new_n6091), .Y(new_n6092));
  O2A1O1Ixp33_ASAP7_75t_L   g05836(.A1(new_n6089), .A2(new_n5843), .B(new_n5842), .C(new_n6092), .Y(new_n6093));
  A2O1A1Ixp33_ASAP7_75t_L   g05837(.A1(new_n5292), .A2(new_n5298), .B(new_n5288), .C(new_n5547), .Y(new_n6094));
  A2O1A1Ixp33_ASAP7_75t_L   g05838(.A1(new_n6094), .A2(new_n5832), .B(new_n5843), .C(new_n5842), .Y(new_n6095));
  NAND2xp33_ASAP7_75t_L     g05839(.A(new_n6070), .B(new_n6069), .Y(new_n6096));
  O2A1O1Ixp33_ASAP7_75t_L   g05840(.A1(new_n6064), .A2(new_n466), .B(new_n6066), .C(new_n6096), .Y(new_n6097));
  O2A1O1Ixp33_ASAP7_75t_L   g05841(.A1(new_n6096), .A2(new_n6097), .B(new_n6091), .C(new_n6095), .Y(new_n6098));
  NOR3xp33_ASAP7_75t_L      g05842(.A(new_n6098), .B(new_n6086), .C(new_n6093), .Y(new_n6099));
  OAI211xp5_ASAP7_75t_L     g05843(.A1(new_n6088), .A2(new_n6099), .B(new_n5874), .C(new_n5873), .Y(new_n6100));
  NAND2xp33_ASAP7_75t_L     g05844(.A(new_n5833), .B(new_n5830), .Y(new_n6101));
  O2A1O1Ixp33_ASAP7_75t_L   g05845(.A1(new_n5836), .A2(new_n346), .B(new_n5838), .C(new_n6101), .Y(new_n6102));
  NOR2xp33_ASAP7_75t_L      g05846(.A(new_n6088), .B(new_n6099), .Y(new_n6103));
  A2O1A1Ixp33_ASAP7_75t_L   g05847(.A1(new_n5850), .A2(new_n5595), .B(new_n6102), .C(new_n6103), .Y(new_n6104));
  NOR2xp33_ASAP7_75t_L      g05848(.A(new_n5570), .B(new_n287), .Y(new_n6105));
  AOI221xp5_ASAP7_75t_L     g05849(.A1(\b[40] ), .A2(new_n264), .B1(\b[41] ), .B2(new_n283), .C(new_n6105), .Y(new_n6106));
  INVx1_ASAP7_75t_L         g05850(.A(new_n5571), .Y(new_n6107));
  A2O1A1Ixp33_ASAP7_75t_L   g05851(.A1(new_n5314), .A2(new_n5568), .B(new_n5569), .C(new_n6107), .Y(new_n6108));
  NOR2xp33_ASAP7_75t_L      g05852(.A(\b[40] ), .B(\b[41] ), .Y(new_n6109));
  INVx1_ASAP7_75t_L         g05853(.A(\b[41] ), .Y(new_n6110));
  NOR2xp33_ASAP7_75t_L      g05854(.A(new_n5855), .B(new_n6110), .Y(new_n6111));
  NOR2xp33_ASAP7_75t_L      g05855(.A(new_n6109), .B(new_n6111), .Y(new_n6112));
  A2O1A1Ixp33_ASAP7_75t_L   g05856(.A1(new_n6108), .A2(new_n5857), .B(new_n5856), .C(new_n6112), .Y(new_n6113));
  O2A1O1Ixp33_ASAP7_75t_L   g05857(.A1(new_n5571), .A2(new_n5574), .B(new_n5857), .C(new_n5856), .Y(new_n6114));
  INVx1_ASAP7_75t_L         g05858(.A(new_n6112), .Y(new_n6115));
  NAND2xp33_ASAP7_75t_L     g05859(.A(new_n6115), .B(new_n6114), .Y(new_n6116));
  NAND2xp33_ASAP7_75t_L     g05860(.A(new_n6116), .B(new_n6113), .Y(new_n6117));
  INVx1_ASAP7_75t_L         g05861(.A(new_n6117), .Y(new_n6118));
  NAND2xp33_ASAP7_75t_L     g05862(.A(new_n273), .B(new_n6118), .Y(new_n6119));
  O2A1O1Ixp33_ASAP7_75t_L   g05863(.A1(new_n279), .A2(new_n6117), .B(new_n6106), .C(new_n257), .Y(new_n6120));
  OAI211xp5_ASAP7_75t_L     g05864(.A1(new_n279), .A2(new_n6117), .B(new_n6106), .C(\a[2] ), .Y(new_n6121));
  A2O1A1Ixp33_ASAP7_75t_L   g05865(.A1(new_n6119), .A2(new_n6106), .B(new_n6120), .C(new_n6121), .Y(new_n6122));
  AOI21xp33_ASAP7_75t_L     g05866(.A1(new_n6104), .A2(new_n6100), .B(new_n6122), .Y(new_n6123));
  NAND3xp33_ASAP7_75t_L     g05867(.A(new_n6104), .B(new_n6100), .C(new_n6122), .Y(new_n6124));
  INVx1_ASAP7_75t_L         g05868(.A(new_n6124), .Y(new_n6125));
  NOR2xp33_ASAP7_75t_L      g05869(.A(new_n6123), .B(new_n6125), .Y(new_n6126));
  XNOR2x2_ASAP7_75t_L       g05870(.A(new_n5872), .B(new_n6126), .Y(\f[41] ));
  NAND3xp33_ASAP7_75t_L     g05871(.A(new_n6079), .B(new_n6075), .C(new_n6087), .Y(new_n6128));
  A2O1A1O1Ixp25_ASAP7_75t_L g05872(.A1(new_n5595), .A2(new_n5850), .B(new_n6102), .C(new_n6128), .D(new_n6088), .Y(new_n6129));
  NOR2xp33_ASAP7_75t_L      g05873(.A(new_n5074), .B(new_n375), .Y(new_n6130));
  AOI221xp5_ASAP7_75t_L     g05874(.A1(\b[39] ), .A2(new_n361), .B1(new_n349), .B2(\b[38] ), .C(new_n6130), .Y(new_n6131));
  O2A1O1Ixp33_ASAP7_75t_L   g05875(.A1(new_n356), .A2(new_n5578), .B(new_n6131), .C(new_n346), .Y(new_n6132));
  INVx1_ASAP7_75t_L         g05876(.A(new_n6132), .Y(new_n6133));
  O2A1O1Ixp33_ASAP7_75t_L   g05877(.A1(new_n356), .A2(new_n5578), .B(new_n6131), .C(\a[5] ), .Y(new_n6134));
  AOI21xp33_ASAP7_75t_L     g05878(.A1(new_n6133), .A2(\a[5] ), .B(new_n6134), .Y(new_n6135));
  A2O1A1O1Ixp25_ASAP7_75t_L g05879(.A1(new_n5808), .A2(new_n5603), .B(new_n5820), .C(new_n6059), .D(new_n6056), .Y(new_n6136));
  A2O1A1O1Ixp25_ASAP7_75t_L g05880(.A1(new_n5604), .A2(new_n5800), .B(new_n5810), .C(new_n6053), .D(new_n6045), .Y(new_n6137));
  A2O1A1Ixp33_ASAP7_75t_L   g05881(.A1(new_n5784), .A2(new_n5892), .B(new_n6037), .C(new_n6033), .Y(new_n6138));
  OAI21xp33_ASAP7_75t_L     g05882(.A1(new_n5968), .A2(new_n5903), .B(new_n5978), .Y(new_n6139));
  OAI21xp33_ASAP7_75t_L     g05883(.A1(new_n5965), .A2(new_n5704), .B(new_n5963), .Y(new_n6140));
  NOR2xp33_ASAP7_75t_L      g05884(.A(new_n833), .B(new_n3510), .Y(new_n6141));
  AOI221xp5_ASAP7_75t_L     g05885(.A1(\b[10] ), .A2(new_n3708), .B1(\b[11] ), .B2(new_n3499), .C(new_n6141), .Y(new_n6142));
  O2A1O1Ixp33_ASAP7_75t_L   g05886(.A1(new_n3513), .A2(new_n841), .B(new_n6142), .C(new_n3493), .Y(new_n6143));
  OAI21xp33_ASAP7_75t_L     g05887(.A1(new_n3513), .A2(new_n841), .B(new_n6142), .Y(new_n6144));
  NAND2xp33_ASAP7_75t_L     g05888(.A(new_n3493), .B(new_n6144), .Y(new_n6145));
  OA21x2_ASAP7_75t_L        g05889(.A1(new_n3493), .A2(new_n6143), .B(new_n6145), .Y(new_n6146));
  A2O1A1Ixp33_ASAP7_75t_L   g05890(.A1(new_n5665), .A2(new_n5669), .B(new_n5687), .C(new_n5674), .Y(new_n6147));
  INVx1_ASAP7_75t_L         g05891(.A(new_n5942), .Y(new_n6148));
  INVx1_ASAP7_75t_L         g05892(.A(\a[42] ), .Y(new_n6149));
  NAND2xp33_ASAP7_75t_L     g05893(.A(\a[41] ), .B(new_n6149), .Y(new_n6150));
  NAND2xp33_ASAP7_75t_L     g05894(.A(\a[42] ), .B(new_n5626), .Y(new_n6151));
  AND2x2_ASAP7_75t_L        g05895(.A(new_n6150), .B(new_n6151), .Y(new_n6152));
  NOR2xp33_ASAP7_75t_L      g05896(.A(new_n284), .B(new_n6152), .Y(new_n6153));
  A2O1A1Ixp33_ASAP7_75t_L   g05897(.A1(new_n5924), .A2(new_n5928), .B(new_n5633), .C(new_n6153), .Y(new_n6154));
  NAND2xp33_ASAP7_75t_L     g05898(.A(new_n5638), .B(new_n5636), .Y(new_n6155));
  NOR5xp2_ASAP7_75t_L       g05899(.A(new_n6155), .B(new_n5927), .C(new_n5922), .D(new_n5349), .E(new_n5626), .Y(new_n6156));
  A2O1A1Ixp33_ASAP7_75t_L   g05900(.A1(new_n6150), .A2(new_n6151), .B(new_n284), .C(new_n6156), .Y(new_n6157));
  NAND2xp33_ASAP7_75t_L     g05901(.A(\b[3] ), .B(new_n5629), .Y(new_n6158));
  NAND2xp33_ASAP7_75t_L     g05902(.A(\b[2] ), .B(new_n5623), .Y(new_n6159));
  OAI211xp5_ASAP7_75t_L     g05903(.A1(new_n5925), .A2(new_n262), .B(new_n6158), .C(new_n6159), .Y(new_n6160));
  NAND2xp33_ASAP7_75t_L     g05904(.A(new_n5637), .B(new_n312), .Y(new_n6161));
  INVx1_ASAP7_75t_L         g05905(.A(new_n6161), .Y(new_n6162));
  A2O1A1Ixp33_ASAP7_75t_L   g05906(.A1(new_n312), .A2(new_n5637), .B(new_n6160), .C(\a[41] ), .Y(new_n6163));
  AOI211xp5_ASAP7_75t_L     g05907(.A1(new_n312), .A2(new_n5637), .B(new_n5626), .C(new_n6160), .Y(new_n6164));
  O2A1O1Ixp33_ASAP7_75t_L   g05908(.A1(new_n6160), .A2(new_n6162), .B(new_n6163), .C(new_n6164), .Y(new_n6165));
  AO21x2_ASAP7_75t_L        g05909(.A1(new_n6154), .A2(new_n6157), .B(new_n6165), .Y(new_n6166));
  NAND3xp33_ASAP7_75t_L     g05910(.A(new_n6157), .B(new_n6154), .C(new_n6165), .Y(new_n6167));
  NAND2xp33_ASAP7_75t_L     g05911(.A(\b[5] ), .B(new_n4916), .Y(new_n6168));
  OAI221xp5_ASAP7_75t_L     g05912(.A1(new_n4908), .A2(new_n427), .B1(new_n332), .B2(new_n5144), .C(new_n6168), .Y(new_n6169));
  A2O1A1Ixp33_ASAP7_75t_L   g05913(.A1(new_n5363), .A2(new_n4912), .B(new_n6169), .C(\a[38] ), .Y(new_n6170));
  NAND2xp33_ASAP7_75t_L     g05914(.A(\a[38] ), .B(new_n6170), .Y(new_n6171));
  A2O1A1Ixp33_ASAP7_75t_L   g05915(.A1(new_n5363), .A2(new_n4912), .B(new_n6169), .C(new_n4906), .Y(new_n6172));
  NAND2xp33_ASAP7_75t_L     g05916(.A(new_n6172), .B(new_n6171), .Y(new_n6173));
  INVx1_ASAP7_75t_L         g05917(.A(new_n6173), .Y(new_n6174));
  NAND3xp33_ASAP7_75t_L     g05918(.A(new_n6174), .B(new_n6167), .C(new_n6166), .Y(new_n6175));
  AOI21xp33_ASAP7_75t_L     g05919(.A1(new_n6157), .A2(new_n6154), .B(new_n6165), .Y(new_n6176));
  AND3x1_ASAP7_75t_L        g05920(.A(new_n6157), .B(new_n6165), .C(new_n6154), .Y(new_n6177));
  OAI21xp33_ASAP7_75t_L     g05921(.A1(new_n6176), .A2(new_n6177), .B(new_n6173), .Y(new_n6178));
  NAND2xp33_ASAP7_75t_L     g05922(.A(new_n5930), .B(new_n5929), .Y(new_n6179));
  O2A1O1Ixp33_ASAP7_75t_L   g05923(.A1(new_n4911), .A2(new_n728), .B(new_n5932), .C(new_n4906), .Y(new_n6180));
  O2A1O1Ixp33_ASAP7_75t_L   g05924(.A1(new_n6180), .A2(new_n4906), .B(new_n5935), .C(new_n6179), .Y(new_n6181));
  O2A1O1Ixp33_ASAP7_75t_L   g05925(.A1(new_n5936), .A2(new_n5937), .B(new_n5918), .C(new_n6181), .Y(new_n6182));
  NAND3xp33_ASAP7_75t_L     g05926(.A(new_n6182), .B(new_n6178), .C(new_n6175), .Y(new_n6183));
  NOR3xp33_ASAP7_75t_L      g05927(.A(new_n6177), .B(new_n6173), .C(new_n6176), .Y(new_n6184));
  AOI21xp33_ASAP7_75t_L     g05928(.A1(new_n6167), .A2(new_n6166), .B(new_n6174), .Y(new_n6185));
  AO21x2_ASAP7_75t_L        g05929(.A1(new_n5935), .A2(new_n5933), .B(new_n6179), .Y(new_n6186));
  OAI21xp33_ASAP7_75t_L     g05930(.A1(new_n5940), .A2(new_n5939), .B(new_n6186), .Y(new_n6187));
  OAI21xp33_ASAP7_75t_L     g05931(.A1(new_n6184), .A2(new_n6185), .B(new_n6187), .Y(new_n6188));
  NOR2xp33_ASAP7_75t_L      g05932(.A(new_n590), .B(new_n4147), .Y(new_n6189));
  AOI221xp5_ASAP7_75t_L     g05933(.A1(\b[7] ), .A2(new_n4402), .B1(\b[8] ), .B2(new_n4155), .C(new_n6189), .Y(new_n6190));
  O2A1O1Ixp33_ASAP7_75t_L   g05934(.A1(new_n4150), .A2(new_n1066), .B(new_n6190), .C(new_n4145), .Y(new_n6191));
  O2A1O1Ixp33_ASAP7_75t_L   g05935(.A1(new_n4150), .A2(new_n1066), .B(new_n6190), .C(\a[35] ), .Y(new_n6192));
  INVx1_ASAP7_75t_L         g05936(.A(new_n6192), .Y(new_n6193));
  OAI21xp33_ASAP7_75t_L     g05937(.A1(new_n4145), .A2(new_n6191), .B(new_n6193), .Y(new_n6194));
  AOI21xp33_ASAP7_75t_L     g05938(.A1(new_n6188), .A2(new_n6183), .B(new_n6194), .Y(new_n6195));
  AND4x1_ASAP7_75t_L        g05939(.A(new_n5938), .B(new_n6175), .C(new_n6186), .D(new_n6178), .Y(new_n6196));
  AOI21xp33_ASAP7_75t_L     g05940(.A1(new_n6178), .A2(new_n6175), .B(new_n6182), .Y(new_n6197));
  OAI21xp33_ASAP7_75t_L     g05941(.A1(new_n4150), .A2(new_n1066), .B(new_n6190), .Y(new_n6198));
  NOR2xp33_ASAP7_75t_L      g05942(.A(new_n4145), .B(new_n6198), .Y(new_n6199));
  NOR2xp33_ASAP7_75t_L      g05943(.A(new_n6192), .B(new_n6199), .Y(new_n6200));
  NOR3xp33_ASAP7_75t_L      g05944(.A(new_n6196), .B(new_n6200), .C(new_n6197), .Y(new_n6201));
  NOR2xp33_ASAP7_75t_L      g05945(.A(new_n6195), .B(new_n6201), .Y(new_n6202));
  A2O1A1Ixp33_ASAP7_75t_L   g05946(.A1(new_n5960), .A2(new_n6147), .B(new_n6148), .C(new_n6202), .Y(new_n6203));
  A2O1A1O1Ixp25_ASAP7_75t_L g05947(.A1(new_n5670), .A2(new_n5672), .B(new_n5911), .C(new_n5960), .D(new_n6148), .Y(new_n6204));
  OAI21xp33_ASAP7_75t_L     g05948(.A1(new_n6197), .A2(new_n6196), .B(new_n6200), .Y(new_n6205));
  NAND3xp33_ASAP7_75t_L     g05949(.A(new_n6194), .B(new_n6188), .C(new_n6183), .Y(new_n6206));
  NAND2xp33_ASAP7_75t_L     g05950(.A(new_n6206), .B(new_n6205), .Y(new_n6207));
  NAND2xp33_ASAP7_75t_L     g05951(.A(new_n6207), .B(new_n6204), .Y(new_n6208));
  AOI21xp33_ASAP7_75t_L     g05952(.A1(new_n6203), .A2(new_n6208), .B(new_n6146), .Y(new_n6209));
  OAI21xp33_ASAP7_75t_L     g05953(.A1(new_n3493), .A2(new_n6143), .B(new_n6145), .Y(new_n6210));
  O2A1O1Ixp33_ASAP7_75t_L   g05954(.A1(new_n5948), .A2(new_n5946), .B(new_n5942), .C(new_n6207), .Y(new_n6211));
  AOI221xp5_ASAP7_75t_L     g05955(.A1(new_n6206), .A2(new_n6205), .B1(new_n5960), .B2(new_n6147), .C(new_n6148), .Y(new_n6212));
  NOR3xp33_ASAP7_75t_L      g05956(.A(new_n6211), .B(new_n6212), .C(new_n6210), .Y(new_n6213));
  OAI21xp33_ASAP7_75t_L     g05957(.A1(new_n6209), .A2(new_n6213), .B(new_n6140), .Y(new_n6214));
  OAI21xp33_ASAP7_75t_L     g05958(.A1(new_n6212), .A2(new_n6211), .B(new_n6210), .Y(new_n6215));
  NAND3xp33_ASAP7_75t_L     g05959(.A(new_n6203), .B(new_n6208), .C(new_n6146), .Y(new_n6216));
  AOI21xp33_ASAP7_75t_L     g05960(.A1(new_n6216), .A2(new_n6215), .B(new_n6140), .Y(new_n6217));
  NOR2xp33_ASAP7_75t_L      g05961(.A(new_n960), .B(new_n2925), .Y(new_n6218));
  AOI221xp5_ASAP7_75t_L     g05962(.A1(\b[13] ), .A2(new_n3129), .B1(\b[15] ), .B2(new_n2938), .C(new_n6218), .Y(new_n6219));
  INVx1_ASAP7_75t_L         g05963(.A(new_n6219), .Y(new_n6220));
  A2O1A1Ixp33_ASAP7_75t_L   g05964(.A1(new_n1052), .A2(new_n2932), .B(new_n6220), .C(\a[29] ), .Y(new_n6221));
  O2A1O1Ixp33_ASAP7_75t_L   g05965(.A1(new_n2940), .A2(new_n1774), .B(new_n6219), .C(\a[29] ), .Y(new_n6222));
  AOI21xp33_ASAP7_75t_L     g05966(.A1(new_n6221), .A2(\a[29] ), .B(new_n6222), .Y(new_n6223));
  A2O1A1Ixp33_ASAP7_75t_L   g05967(.A1(new_n6214), .A2(new_n6140), .B(new_n6217), .C(new_n6223), .Y(new_n6224));
  NAND3xp33_ASAP7_75t_L     g05968(.A(new_n6140), .B(new_n6215), .C(new_n6216), .Y(new_n6225));
  A2O1A1O1Ixp25_ASAP7_75t_L g05969(.A1(new_n5612), .A2(new_n5694), .B(new_n5684), .C(new_n5957), .D(new_n5966), .Y(new_n6226));
  OAI21xp33_ASAP7_75t_L     g05970(.A1(new_n6209), .A2(new_n6213), .B(new_n6226), .Y(new_n6227));
  AO21x2_ASAP7_75t_L        g05971(.A1(\a[29] ), .A2(new_n6221), .B(new_n6222), .Y(new_n6228));
  NAND3xp33_ASAP7_75t_L     g05972(.A(new_n6228), .B(new_n6227), .C(new_n6225), .Y(new_n6229));
  NAND3xp33_ASAP7_75t_L     g05973(.A(new_n6139), .B(new_n6224), .C(new_n6229), .Y(new_n6230));
  A2O1A1O1Ixp25_ASAP7_75t_L g05974(.A1(new_n5723), .A2(new_n5719), .B(new_n5722), .C(new_n5977), .D(new_n5974), .Y(new_n6231));
  NAND2xp33_ASAP7_75t_L     g05975(.A(new_n6227), .B(new_n6225), .Y(new_n6232));
  A2O1A1Ixp33_ASAP7_75t_L   g05976(.A1(new_n6214), .A2(new_n6140), .B(new_n6217), .C(new_n6228), .Y(new_n6233));
  AOI211xp5_ASAP7_75t_L     g05977(.A1(new_n6214), .A2(new_n6140), .B(new_n6217), .C(new_n6223), .Y(new_n6234));
  A2O1A1Ixp33_ASAP7_75t_L   g05978(.A1(new_n6232), .A2(new_n6233), .B(new_n6234), .C(new_n6231), .Y(new_n6235));
  NOR2xp33_ASAP7_75t_L      g05979(.A(new_n1349), .B(new_n2410), .Y(new_n6236));
  AOI221xp5_ASAP7_75t_L     g05980(.A1(\b[16] ), .A2(new_n2577), .B1(\b[18] ), .B2(new_n2423), .C(new_n6236), .Y(new_n6237));
  INVx1_ASAP7_75t_L         g05981(.A(new_n6237), .Y(new_n6238));
  A2O1A1Ixp33_ASAP7_75t_L   g05982(.A1(new_n2329), .A2(new_n2417), .B(new_n6238), .C(\a[26] ), .Y(new_n6239));
  O2A1O1Ixp33_ASAP7_75t_L   g05983(.A1(new_n2425), .A2(new_n1464), .B(new_n6237), .C(\a[26] ), .Y(new_n6240));
  AOI21xp33_ASAP7_75t_L     g05984(.A1(new_n6239), .A2(\a[26] ), .B(new_n6240), .Y(new_n6241));
  AOI21xp33_ASAP7_75t_L     g05985(.A1(new_n6235), .A2(new_n6230), .B(new_n6241), .Y(new_n6242));
  AOI21xp33_ASAP7_75t_L     g05986(.A1(new_n6225), .A2(new_n6227), .B(new_n6228), .Y(new_n6243));
  NOR3xp33_ASAP7_75t_L      g05987(.A(new_n6231), .B(new_n6243), .C(new_n6234), .Y(new_n6244));
  AOI21xp33_ASAP7_75t_L     g05988(.A1(new_n6229), .A2(new_n6224), .B(new_n6139), .Y(new_n6245));
  O2A1O1Ixp33_ASAP7_75t_L   g05989(.A1(new_n2425), .A2(new_n1464), .B(new_n6237), .C(new_n2413), .Y(new_n6246));
  A2O1A1Ixp33_ASAP7_75t_L   g05990(.A1(new_n2329), .A2(new_n2417), .B(new_n6238), .C(new_n2413), .Y(new_n6247));
  OAI21xp33_ASAP7_75t_L     g05991(.A1(new_n2413), .A2(new_n6246), .B(new_n6247), .Y(new_n6248));
  NOR3xp33_ASAP7_75t_L      g05992(.A(new_n6244), .B(new_n6245), .C(new_n6248), .Y(new_n6249));
  NOR2xp33_ASAP7_75t_L      g05993(.A(new_n6242), .B(new_n6249), .Y(new_n6250));
  A2O1A1Ixp33_ASAP7_75t_L   g05994(.A1(new_n5990), .A2(new_n5987), .B(new_n5989), .C(new_n6250), .Y(new_n6251));
  A2O1A1O1Ixp25_ASAP7_75t_L g05995(.A1(new_n5999), .A2(new_n5735), .B(new_n5895), .C(new_n5980), .D(new_n5989), .Y(new_n6252));
  OAI21xp33_ASAP7_75t_L     g05996(.A1(new_n6245), .A2(new_n6244), .B(new_n6248), .Y(new_n6253));
  NAND3xp33_ASAP7_75t_L     g05997(.A(new_n6235), .B(new_n6230), .C(new_n6241), .Y(new_n6254));
  NAND2xp33_ASAP7_75t_L     g05998(.A(new_n6254), .B(new_n6253), .Y(new_n6255));
  NAND2xp33_ASAP7_75t_L     g05999(.A(new_n6252), .B(new_n6255), .Y(new_n6256));
  NOR2xp33_ASAP7_75t_L      g06000(.A(new_n1745), .B(new_n1962), .Y(new_n6257));
  AOI221xp5_ASAP7_75t_L     g06001(.A1(new_n1955), .A2(\b[21] ), .B1(new_n2093), .B2(\b[19] ), .C(new_n6257), .Y(new_n6258));
  INVx1_ASAP7_75t_L         g06002(.A(new_n6258), .Y(new_n6259));
  A2O1A1Ixp33_ASAP7_75t_L   g06003(.A1(new_n2836), .A2(new_n1964), .B(new_n6259), .C(\a[23] ), .Y(new_n6260));
  O2A1O1Ixp33_ASAP7_75t_L   g06004(.A1(new_n1956), .A2(new_n1901), .B(new_n6258), .C(\a[23] ), .Y(new_n6261));
  AOI21xp33_ASAP7_75t_L     g06005(.A1(new_n6260), .A2(\a[23] ), .B(new_n6261), .Y(new_n6262));
  NAND3xp33_ASAP7_75t_L     g06006(.A(new_n6251), .B(new_n6256), .C(new_n6262), .Y(new_n6263));
  NOR2xp33_ASAP7_75t_L      g06007(.A(new_n6252), .B(new_n6255), .Y(new_n6264));
  AOI221xp5_ASAP7_75t_L     g06008(.A1(new_n6254), .A2(new_n6253), .B1(new_n5990), .B2(new_n5987), .C(new_n5989), .Y(new_n6265));
  O2A1O1Ixp33_ASAP7_75t_L   g06009(.A1(new_n1956), .A2(new_n1901), .B(new_n6258), .C(new_n1952), .Y(new_n6266));
  NOR2xp33_ASAP7_75t_L      g06010(.A(new_n1952), .B(new_n6266), .Y(new_n6267));
  OAI22xp33_ASAP7_75t_L     g06011(.A1(new_n6264), .A2(new_n6265), .B1(new_n6261), .B2(new_n6267), .Y(new_n6268));
  AND2x2_ASAP7_75t_L        g06012(.A(new_n6268), .B(new_n6263), .Y(new_n6269));
  NOR2xp33_ASAP7_75t_L      g06013(.A(new_n5986), .B(new_n5991), .Y(new_n6270));
  MAJIxp5_ASAP7_75t_L       g06014(.A(new_n6006), .B(new_n5997), .C(new_n6270), .Y(new_n6271));
  NAND2xp33_ASAP7_75t_L     g06015(.A(new_n6271), .B(new_n6269), .Y(new_n6272));
  NAND2xp33_ASAP7_75t_L     g06016(.A(new_n6002), .B(new_n6000), .Y(new_n6273));
  O2A1O1Ixp33_ASAP7_75t_L   g06017(.A1(new_n5994), .A2(new_n1952), .B(new_n5996), .C(new_n6273), .Y(new_n6274));
  NAND3xp33_ASAP7_75t_L     g06018(.A(new_n6003), .B(new_n6002), .C(new_n6000), .Y(new_n6275));
  OAI21xp33_ASAP7_75t_L     g06019(.A1(new_n5986), .A2(new_n5991), .B(new_n5997), .Y(new_n6276));
  NAND2xp33_ASAP7_75t_L     g06020(.A(new_n6276), .B(new_n6275), .Y(new_n6277));
  NAND2xp33_ASAP7_75t_L     g06021(.A(new_n6268), .B(new_n6263), .Y(new_n6278));
  A2O1A1Ixp33_ASAP7_75t_L   g06022(.A1(new_n6277), .A2(new_n6006), .B(new_n6274), .C(new_n6278), .Y(new_n6279));
  OAI22xp33_ASAP7_75t_L     g06023(.A1(new_n1654), .A2(new_n2045), .B1(new_n2188), .B2(new_n1517), .Y(new_n6280));
  AOI221xp5_ASAP7_75t_L     g06024(.A1(new_n1511), .A2(\b[24] ), .B1(new_n1513), .B2(new_n2216), .C(new_n6280), .Y(new_n6281));
  XNOR2x2_ASAP7_75t_L       g06025(.A(\a[20] ), .B(new_n6281), .Y(new_n6282));
  AOI21xp33_ASAP7_75t_L     g06026(.A1(new_n6272), .A2(new_n6279), .B(new_n6282), .Y(new_n6283));
  AND3x1_ASAP7_75t_L        g06027(.A(new_n6272), .B(new_n6279), .C(new_n6282), .Y(new_n6284));
  NOR3xp33_ASAP7_75t_L      g06028(.A(new_n6031), .B(new_n6284), .C(new_n6283), .Y(new_n6285));
  AO21x2_ASAP7_75t_L        g06029(.A1(new_n6279), .A2(new_n6272), .B(new_n6282), .Y(new_n6286));
  NAND3xp33_ASAP7_75t_L     g06030(.A(new_n6272), .B(new_n6279), .C(new_n6282), .Y(new_n6287));
  AOI211xp5_ASAP7_75t_L     g06031(.A1(new_n6286), .A2(new_n6287), .B(new_n6015), .C(new_n6038), .Y(new_n6288));
  NOR2xp33_ASAP7_75t_L      g06032(.A(new_n6285), .B(new_n6288), .Y(new_n6289));
  NOR2xp33_ASAP7_75t_L      g06033(.A(new_n2703), .B(new_n2118), .Y(new_n6290));
  AOI221xp5_ASAP7_75t_L     g06034(.A1(\b[25] ), .A2(new_n1290), .B1(\b[27] ), .B2(new_n1209), .C(new_n6290), .Y(new_n6291));
  INVx1_ASAP7_75t_L         g06035(.A(new_n6291), .Y(new_n6292));
  A2O1A1Ixp33_ASAP7_75t_L   g06036(.A1(new_n2887), .A2(new_n1216), .B(new_n6292), .C(\a[17] ), .Y(new_n6293));
  O2A1O1Ixp33_ASAP7_75t_L   g06037(.A1(new_n1210), .A2(new_n2889), .B(new_n6291), .C(new_n1206), .Y(new_n6294));
  NOR2xp33_ASAP7_75t_L      g06038(.A(new_n1206), .B(new_n6294), .Y(new_n6295));
  A2O1A1O1Ixp25_ASAP7_75t_L g06039(.A1(new_n2887), .A2(new_n1216), .B(new_n6292), .C(new_n6293), .D(new_n6295), .Y(new_n6296));
  NAND2xp33_ASAP7_75t_L     g06040(.A(new_n6296), .B(new_n6289), .Y(new_n6297));
  OAI211xp5_ASAP7_75t_L     g06041(.A1(new_n6015), .A2(new_n6038), .B(new_n6286), .C(new_n6287), .Y(new_n6298));
  OAI21xp33_ASAP7_75t_L     g06042(.A1(new_n6283), .A2(new_n6284), .B(new_n6031), .Y(new_n6299));
  NAND2xp33_ASAP7_75t_L     g06043(.A(new_n6299), .B(new_n6298), .Y(new_n6300));
  NAND2xp33_ASAP7_75t_L     g06044(.A(new_n1216), .B(new_n2887), .Y(new_n6301));
  NAND2xp33_ASAP7_75t_L     g06045(.A(\a[17] ), .B(new_n6293), .Y(new_n6302));
  A2O1A1Ixp33_ASAP7_75t_L   g06046(.A1(new_n6301), .A2(new_n6291), .B(new_n6294), .C(new_n6302), .Y(new_n6303));
  NAND2xp33_ASAP7_75t_L     g06047(.A(new_n6303), .B(new_n6300), .Y(new_n6304));
  NAND3xp33_ASAP7_75t_L     g06048(.A(new_n6304), .B(new_n6297), .C(new_n6138), .Y(new_n6305));
  NAND2xp33_ASAP7_75t_L     g06049(.A(new_n5785), .B(new_n5786), .Y(new_n6306));
  A2O1A1O1Ixp25_ASAP7_75t_L g06050(.A1(new_n5783), .A2(new_n6306), .B(new_n6035), .C(new_n6029), .D(new_n6039), .Y(new_n6307));
  NOR3xp33_ASAP7_75t_L      g06051(.A(new_n6303), .B(new_n6288), .C(new_n6285), .Y(new_n6308));
  AOI21xp33_ASAP7_75t_L     g06052(.A1(new_n6298), .A2(new_n6299), .B(new_n6296), .Y(new_n6309));
  OAI21xp33_ASAP7_75t_L     g06053(.A1(new_n6308), .A2(new_n6309), .B(new_n6307), .Y(new_n6310));
  NOR2xp33_ASAP7_75t_L      g06054(.A(new_n3098), .B(new_n864), .Y(new_n6311));
  AOI221xp5_ASAP7_75t_L     g06055(.A1(\b[28] ), .A2(new_n985), .B1(\b[30] ), .B2(new_n886), .C(new_n6311), .Y(new_n6312));
  O2A1O1Ixp33_ASAP7_75t_L   g06056(.A1(new_n872), .A2(new_n3464), .B(new_n6312), .C(new_n867), .Y(new_n6313));
  INVx1_ASAP7_75t_L         g06057(.A(new_n6313), .Y(new_n6314));
  O2A1O1Ixp33_ASAP7_75t_L   g06058(.A1(new_n872), .A2(new_n3464), .B(new_n6312), .C(\a[14] ), .Y(new_n6315));
  AOI21xp33_ASAP7_75t_L     g06059(.A1(new_n6314), .A2(\a[14] ), .B(new_n6315), .Y(new_n6316));
  AOI21xp33_ASAP7_75t_L     g06060(.A1(new_n6305), .A2(new_n6310), .B(new_n6316), .Y(new_n6317));
  NOR3xp33_ASAP7_75t_L      g06061(.A(new_n6307), .B(new_n6308), .C(new_n6309), .Y(new_n6318));
  AOI21xp33_ASAP7_75t_L     g06062(.A1(new_n6304), .A2(new_n6297), .B(new_n6138), .Y(new_n6319));
  AO21x2_ASAP7_75t_L        g06063(.A1(\a[14] ), .A2(new_n6314), .B(new_n6315), .Y(new_n6320));
  NOR3xp33_ASAP7_75t_L      g06064(.A(new_n6319), .B(new_n6320), .C(new_n6318), .Y(new_n6321));
  NOR3xp33_ASAP7_75t_L      g06065(.A(new_n6137), .B(new_n6317), .C(new_n6321), .Y(new_n6322));
  OAI21xp33_ASAP7_75t_L     g06066(.A1(new_n6318), .A2(new_n6319), .B(new_n6320), .Y(new_n6323));
  NAND3xp33_ASAP7_75t_L     g06067(.A(new_n6305), .B(new_n6310), .C(new_n6316), .Y(new_n6324));
  AOI221xp5_ASAP7_75t_L     g06068(.A1(new_n6046), .A2(new_n5884), .B1(new_n6324), .B2(new_n6323), .C(new_n6045), .Y(new_n6325));
  NOR2xp33_ASAP7_75t_L      g06069(.A(new_n3891), .B(new_n1550), .Y(new_n6326));
  AOI221xp5_ASAP7_75t_L     g06070(.A1(\b[31] ), .A2(new_n713), .B1(\b[33] ), .B2(new_n640), .C(new_n6326), .Y(new_n6327));
  O2A1O1Ixp33_ASAP7_75t_L   g06071(.A1(new_n641), .A2(new_n4108), .B(new_n6327), .C(new_n637), .Y(new_n6328));
  INVx1_ASAP7_75t_L         g06072(.A(new_n6327), .Y(new_n6329));
  A2O1A1Ixp33_ASAP7_75t_L   g06073(.A1(new_n4831), .A2(new_n718), .B(new_n6329), .C(new_n637), .Y(new_n6330));
  OAI21xp33_ASAP7_75t_L     g06074(.A1(new_n637), .A2(new_n6328), .B(new_n6330), .Y(new_n6331));
  NOR3xp33_ASAP7_75t_L      g06075(.A(new_n6325), .B(new_n6322), .C(new_n6331), .Y(new_n6332));
  A2O1A1Ixp33_ASAP7_75t_L   g06076(.A1(new_n5809), .A2(new_n5883), .B(new_n6041), .C(new_n6054), .Y(new_n6333));
  NAND3xp33_ASAP7_75t_L     g06077(.A(new_n6333), .B(new_n6323), .C(new_n6324), .Y(new_n6334));
  OAI21xp33_ASAP7_75t_L     g06078(.A1(new_n6317), .A2(new_n6321), .B(new_n6137), .Y(new_n6335));
  INVx1_ASAP7_75t_L         g06079(.A(new_n6331), .Y(new_n6336));
  AOI21xp33_ASAP7_75t_L     g06080(.A1(new_n6334), .A2(new_n6335), .B(new_n6336), .Y(new_n6337));
  NOR3xp33_ASAP7_75t_L      g06081(.A(new_n6136), .B(new_n6332), .C(new_n6337), .Y(new_n6338));
  OAI21xp33_ASAP7_75t_L     g06082(.A1(new_n6050), .A2(new_n5876), .B(new_n6060), .Y(new_n6339));
  NAND3xp33_ASAP7_75t_L     g06083(.A(new_n6336), .B(new_n6334), .C(new_n6335), .Y(new_n6340));
  OAI21xp33_ASAP7_75t_L     g06084(.A1(new_n6322), .A2(new_n6325), .B(new_n6331), .Y(new_n6341));
  AOI21xp33_ASAP7_75t_L     g06085(.A1(new_n6341), .A2(new_n6340), .B(new_n6339), .Y(new_n6342));
  NOR2xp33_ASAP7_75t_L      g06086(.A(new_n4581), .B(new_n513), .Y(new_n6343));
  AOI221xp5_ASAP7_75t_L     g06087(.A1(\b[34] ), .A2(new_n560), .B1(\b[36] ), .B2(new_n475), .C(new_n6343), .Y(new_n6344));
  INVx1_ASAP7_75t_L         g06088(.A(new_n6344), .Y(new_n6345));
  A2O1A1Ixp33_ASAP7_75t_L   g06089(.A1(new_n4621), .A2(new_n483), .B(new_n6345), .C(\a[8] ), .Y(new_n6346));
  NAND2xp33_ASAP7_75t_L     g06090(.A(\a[8] ), .B(new_n6346), .Y(new_n6347));
  A2O1A1Ixp33_ASAP7_75t_L   g06091(.A1(new_n4621), .A2(new_n483), .B(new_n6345), .C(new_n466), .Y(new_n6348));
  NAND2xp33_ASAP7_75t_L     g06092(.A(new_n6348), .B(new_n6347), .Y(new_n6349));
  NOR3xp33_ASAP7_75t_L      g06093(.A(new_n6338), .B(new_n6342), .C(new_n6349), .Y(new_n6350));
  NAND3xp33_ASAP7_75t_L     g06094(.A(new_n6339), .B(new_n6340), .C(new_n6341), .Y(new_n6351));
  OAI21xp33_ASAP7_75t_L     g06095(.A1(new_n6332), .A2(new_n6337), .B(new_n6136), .Y(new_n6352));
  INVx1_ASAP7_75t_L         g06096(.A(new_n6348), .Y(new_n6353));
  AOI21xp33_ASAP7_75t_L     g06097(.A1(new_n6346), .A2(\a[8] ), .B(new_n6353), .Y(new_n6354));
  AOI21xp33_ASAP7_75t_L     g06098(.A1(new_n6351), .A2(new_n6352), .B(new_n6354), .Y(new_n6355));
  NOR2xp33_ASAP7_75t_L      g06099(.A(new_n6355), .B(new_n6350), .Y(new_n6356));
  A2O1A1Ixp33_ASAP7_75t_L   g06100(.A1(new_n6092), .A2(new_n6095), .B(new_n6097), .C(new_n6356), .Y(new_n6357));
  A2O1A1Ixp33_ASAP7_75t_L   g06101(.A1(new_n5829), .A2(new_n5875), .B(new_n5828), .C(new_n6092), .Y(new_n6358));
  NAND3xp33_ASAP7_75t_L     g06102(.A(new_n6351), .B(new_n6354), .C(new_n6352), .Y(new_n6359));
  OAI21xp33_ASAP7_75t_L     g06103(.A1(new_n6342), .A2(new_n6338), .B(new_n6349), .Y(new_n6360));
  NAND2xp33_ASAP7_75t_L     g06104(.A(new_n6359), .B(new_n6360), .Y(new_n6361));
  NAND3xp33_ASAP7_75t_L     g06105(.A(new_n6358), .B(new_n6078), .C(new_n6361), .Y(new_n6362));
  AOI21xp33_ASAP7_75t_L     g06106(.A1(new_n6357), .A2(new_n6362), .B(new_n6135), .Y(new_n6363));
  INVx1_ASAP7_75t_L         g06107(.A(new_n6134), .Y(new_n6364));
  OAI21xp33_ASAP7_75t_L     g06108(.A1(new_n346), .A2(new_n6132), .B(new_n6364), .Y(new_n6365));
  O2A1O1Ixp33_ASAP7_75t_L   g06109(.A1(new_n6076), .A2(new_n6074), .B(new_n6078), .C(new_n6361), .Y(new_n6366));
  AOI221xp5_ASAP7_75t_L     g06110(.A1(new_n6360), .A2(new_n6359), .B1(new_n6092), .B2(new_n6095), .C(new_n6097), .Y(new_n6367));
  NOR3xp33_ASAP7_75t_L      g06111(.A(new_n6366), .B(new_n6367), .C(new_n6365), .Y(new_n6368));
  NOR3xp33_ASAP7_75t_L      g06112(.A(new_n6129), .B(new_n6363), .C(new_n6368), .Y(new_n6369));
  A2O1A1Ixp33_ASAP7_75t_L   g06113(.A1(new_n5847), .A2(new_n6101), .B(new_n5849), .C(new_n5873), .Y(new_n6370));
  OAI21xp33_ASAP7_75t_L     g06114(.A1(new_n6367), .A2(new_n6366), .B(new_n6365), .Y(new_n6371));
  NAND3xp33_ASAP7_75t_L     g06115(.A(new_n6357), .B(new_n6362), .C(new_n6135), .Y(new_n6372));
  AOI221xp5_ASAP7_75t_L     g06116(.A1(new_n6370), .A2(new_n6128), .B1(new_n6371), .B2(new_n6372), .C(new_n6088), .Y(new_n6373));
  NOR2xp33_ASAP7_75t_L      g06117(.A(new_n5855), .B(new_n287), .Y(new_n6374));
  AOI221xp5_ASAP7_75t_L     g06118(.A1(\b[41] ), .A2(new_n264), .B1(\b[42] ), .B2(new_n283), .C(new_n6374), .Y(new_n6375));
  INVx1_ASAP7_75t_L         g06119(.A(new_n6111), .Y(new_n6376));
  NOR2xp33_ASAP7_75t_L      g06120(.A(\b[41] ), .B(\b[42] ), .Y(new_n6377));
  INVx1_ASAP7_75t_L         g06121(.A(\b[42] ), .Y(new_n6378));
  NOR2xp33_ASAP7_75t_L      g06122(.A(new_n6110), .B(new_n6378), .Y(new_n6379));
  NOR2xp33_ASAP7_75t_L      g06123(.A(new_n6377), .B(new_n6379), .Y(new_n6380));
  INVx1_ASAP7_75t_L         g06124(.A(new_n6380), .Y(new_n6381));
  O2A1O1Ixp33_ASAP7_75t_L   g06125(.A1(new_n6115), .A2(new_n6114), .B(new_n6376), .C(new_n6381), .Y(new_n6382));
  INVx1_ASAP7_75t_L         g06126(.A(new_n6382), .Y(new_n6383));
  A2O1A1O1Ixp25_ASAP7_75t_L g06127(.A1(new_n5857), .A2(new_n6108), .B(new_n5856), .C(new_n6112), .D(new_n6111), .Y(new_n6384));
  NAND2xp33_ASAP7_75t_L     g06128(.A(new_n6381), .B(new_n6384), .Y(new_n6385));
  NAND2xp33_ASAP7_75t_L     g06129(.A(new_n6383), .B(new_n6385), .Y(new_n6386));
  O2A1O1Ixp33_ASAP7_75t_L   g06130(.A1(new_n279), .A2(new_n6386), .B(new_n6375), .C(new_n257), .Y(new_n6387));
  INVx1_ASAP7_75t_L         g06131(.A(new_n6375), .Y(new_n6388));
  AND2x2_ASAP7_75t_L        g06132(.A(new_n6383), .B(new_n6385), .Y(new_n6389));
  A2O1A1Ixp33_ASAP7_75t_L   g06133(.A1(new_n6389), .A2(new_n273), .B(new_n6388), .C(new_n257), .Y(new_n6390));
  OAI21xp33_ASAP7_75t_L     g06134(.A1(new_n257), .A2(new_n6387), .B(new_n6390), .Y(new_n6391));
  INVx1_ASAP7_75t_L         g06135(.A(new_n6391), .Y(new_n6392));
  OAI21xp33_ASAP7_75t_L     g06136(.A1(new_n6373), .A2(new_n6369), .B(new_n6392), .Y(new_n6393));
  AOI21xp33_ASAP7_75t_L     g06137(.A1(new_n6372), .A2(new_n6371), .B(new_n6129), .Y(new_n6394));
  NAND2xp33_ASAP7_75t_L     g06138(.A(new_n6371), .B(new_n6372), .Y(new_n6395));
  NAND2xp33_ASAP7_75t_L     g06139(.A(new_n6129), .B(new_n6395), .Y(new_n6396));
  OAI211xp5_ASAP7_75t_L     g06140(.A1(new_n6394), .A2(new_n6129), .B(new_n6396), .C(new_n6391), .Y(new_n6397));
  NAND2xp33_ASAP7_75t_L     g06141(.A(new_n6393), .B(new_n6397), .Y(new_n6398));
  INVx1_ASAP7_75t_L         g06142(.A(new_n6398), .Y(new_n6399));
  O2A1O1Ixp33_ASAP7_75t_L   g06143(.A1(new_n5872), .A2(new_n6123), .B(new_n6124), .C(new_n6399), .Y(new_n6400));
  OAI21xp33_ASAP7_75t_L     g06144(.A1(new_n6123), .A2(new_n5872), .B(new_n6124), .Y(new_n6401));
  NOR2xp33_ASAP7_75t_L      g06145(.A(new_n6398), .B(new_n6401), .Y(new_n6402));
  NOR2xp33_ASAP7_75t_L      g06146(.A(new_n6402), .B(new_n6400), .Y(\f[42] ));
  NAND2xp33_ASAP7_75t_L     g06147(.A(new_n6362), .B(new_n6357), .Y(new_n6404));
  MAJIxp5_ASAP7_75t_L       g06148(.A(new_n6129), .B(new_n6135), .C(new_n6404), .Y(new_n6405));
  OAI21xp33_ASAP7_75t_L     g06149(.A1(new_n6321), .A2(new_n6137), .B(new_n6323), .Y(new_n6406));
  MAJIxp5_ASAP7_75t_L       g06150(.A(new_n6307), .B(new_n6300), .C(new_n6296), .Y(new_n6407));
  NOR2xp33_ASAP7_75t_L      g06151(.A(new_n3079), .B(new_n1284), .Y(new_n6408));
  AOI221xp5_ASAP7_75t_L     g06152(.A1(\b[26] ), .A2(new_n1290), .B1(\b[27] ), .B2(new_n1204), .C(new_n6408), .Y(new_n6409));
  O2A1O1Ixp33_ASAP7_75t_L   g06153(.A1(new_n1210), .A2(new_n3087), .B(new_n6409), .C(new_n1206), .Y(new_n6410));
  O2A1O1Ixp33_ASAP7_75t_L   g06154(.A1(new_n1210), .A2(new_n3087), .B(new_n6409), .C(\a[17] ), .Y(new_n6411));
  INVx1_ASAP7_75t_L         g06155(.A(new_n6411), .Y(new_n6412));
  OAI21xp33_ASAP7_75t_L     g06156(.A1(new_n1206), .A2(new_n6410), .B(new_n6412), .Y(new_n6413));
  NOR2xp33_ASAP7_75t_L      g06157(.A(new_n6212), .B(new_n6211), .Y(new_n6414));
  MAJIxp5_ASAP7_75t_L       g06158(.A(new_n6140), .B(new_n6210), .C(new_n6414), .Y(new_n6415));
  A2O1A1Ixp33_ASAP7_75t_L   g06159(.A1(new_n5961), .A2(new_n5942), .B(new_n6207), .C(new_n6206), .Y(new_n6416));
  NAND3xp33_ASAP7_75t_L     g06160(.A(new_n6166), .B(new_n6167), .C(new_n6173), .Y(new_n6417));
  NOR2xp33_ASAP7_75t_L      g06161(.A(new_n427), .B(new_n4903), .Y(new_n6418));
  AOI221xp5_ASAP7_75t_L     g06162(.A1(\b[5] ), .A2(new_n5139), .B1(\b[7] ), .B2(new_n4917), .C(new_n6418), .Y(new_n6419));
  OAI211xp5_ASAP7_75t_L     g06163(.A1(new_n4911), .A2(new_n456), .B(\a[38] ), .C(new_n6419), .Y(new_n6420));
  INVx1_ASAP7_75t_L         g06164(.A(new_n6419), .Y(new_n6421));
  A2O1A1Ixp33_ASAP7_75t_L   g06165(.A1(new_n1188), .A2(new_n4912), .B(new_n6421), .C(new_n4906), .Y(new_n6422));
  NAND2xp33_ASAP7_75t_L     g06166(.A(new_n6420), .B(new_n6422), .Y(new_n6423));
  INVx1_ASAP7_75t_L         g06167(.A(new_n6153), .Y(new_n6424));
  MAJIxp5_ASAP7_75t_L       g06168(.A(new_n6165), .B(new_n5930), .C(new_n6424), .Y(new_n6425));
  NAND2xp33_ASAP7_75t_L     g06169(.A(\b[3] ), .B(new_n5623), .Y(new_n6426));
  OAI221xp5_ASAP7_75t_L     g06170(.A1(new_n5641), .A2(new_n332), .B1(new_n289), .B2(new_n5925), .C(new_n6426), .Y(new_n6427));
  A2O1A1Ixp33_ASAP7_75t_L   g06171(.A1(new_n342), .A2(new_n5637), .B(new_n6427), .C(\a[41] ), .Y(new_n6428));
  NAND2xp33_ASAP7_75t_L     g06172(.A(\a[41] ), .B(new_n6428), .Y(new_n6429));
  NOR2xp33_ASAP7_75t_L      g06173(.A(new_n332), .B(new_n5641), .Y(new_n6430));
  AOI221xp5_ASAP7_75t_L     g06174(.A1(\b[2] ), .A2(new_n5920), .B1(\b[3] ), .B2(new_n5623), .C(new_n6430), .Y(new_n6431));
  O2A1O1Ixp33_ASAP7_75t_L   g06175(.A1(new_n5630), .A2(new_n1497), .B(new_n6431), .C(\a[41] ), .Y(new_n6432));
  INVx1_ASAP7_75t_L         g06176(.A(new_n6432), .Y(new_n6433));
  NAND2xp33_ASAP7_75t_L     g06177(.A(new_n6151), .B(new_n6150), .Y(new_n6434));
  XNOR2x2_ASAP7_75t_L       g06178(.A(\a[43] ), .B(\a[42] ), .Y(new_n6435));
  NOR2xp33_ASAP7_75t_L      g06179(.A(new_n6435), .B(new_n6434), .Y(new_n6436));
  INVx1_ASAP7_75t_L         g06180(.A(\a[43] ), .Y(new_n6437));
  NAND2xp33_ASAP7_75t_L     g06181(.A(\a[44] ), .B(new_n6437), .Y(new_n6438));
  INVx1_ASAP7_75t_L         g06182(.A(\a[44] ), .Y(new_n6439));
  NAND2xp33_ASAP7_75t_L     g06183(.A(\a[43] ), .B(new_n6439), .Y(new_n6440));
  NAND2xp33_ASAP7_75t_L     g06184(.A(new_n6440), .B(new_n6438), .Y(new_n6441));
  NOR2xp33_ASAP7_75t_L      g06185(.A(new_n6441), .B(new_n6152), .Y(new_n6442));
  NAND2xp33_ASAP7_75t_L     g06186(.A(new_n6441), .B(new_n6434), .Y(new_n6443));
  NOR2xp33_ASAP7_75t_L      g06187(.A(new_n274), .B(new_n6443), .Y(new_n6444));
  AOI221xp5_ASAP7_75t_L     g06188(.A1(\b[1] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[0] ), .C(new_n6444), .Y(new_n6445));
  NAND3xp33_ASAP7_75t_L     g06189(.A(new_n6445), .B(new_n6424), .C(\a[44] ), .Y(new_n6446));
  INVx1_ASAP7_75t_L         g06190(.A(new_n6446), .Y(new_n6447));
  A2O1A1Ixp33_ASAP7_75t_L   g06191(.A1(new_n6150), .A2(new_n6151), .B(new_n284), .C(\a[44] ), .Y(new_n6448));
  AOI22xp33_ASAP7_75t_L     g06192(.A1(new_n6436), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n6442), .Y(new_n6449));
  AOI21xp33_ASAP7_75t_L     g06193(.A1(new_n6440), .A2(new_n6438), .B(new_n6152), .Y(new_n6450));
  NAND2xp33_ASAP7_75t_L     g06194(.A(new_n275), .B(new_n6450), .Y(new_n6451));
  NAND3xp33_ASAP7_75t_L     g06195(.A(new_n6449), .B(\a[44] ), .C(new_n6451), .Y(new_n6452));
  AO21x2_ASAP7_75t_L        g06196(.A1(new_n6451), .A2(new_n6449), .B(\a[44] ), .Y(new_n6453));
  AND3x1_ASAP7_75t_L        g06197(.A(new_n6453), .B(new_n6452), .C(new_n6448), .Y(new_n6454));
  OAI211xp5_ASAP7_75t_L     g06198(.A1(new_n6447), .A2(new_n6454), .B(new_n6433), .C(new_n6429), .Y(new_n6455));
  O2A1O1Ixp33_ASAP7_75t_L   g06199(.A1(new_n5630), .A2(new_n1497), .B(new_n6431), .C(new_n5626), .Y(new_n6456));
  NOR2xp33_ASAP7_75t_L      g06200(.A(new_n5626), .B(new_n6456), .Y(new_n6457));
  O2A1O1Ixp33_ASAP7_75t_L   g06201(.A1(new_n6443), .A2(new_n274), .B(new_n6449), .C(new_n6439), .Y(new_n6458));
  A2O1A1Ixp33_ASAP7_75t_L   g06202(.A1(new_n6458), .A2(new_n6153), .B(new_n6439), .C(new_n6453), .Y(new_n6459));
  OAI211xp5_ASAP7_75t_L     g06203(.A1(new_n6432), .A2(new_n6457), .B(new_n6446), .C(new_n6459), .Y(new_n6460));
  NAND3xp33_ASAP7_75t_L     g06204(.A(new_n6425), .B(new_n6460), .C(new_n6455), .Y(new_n6461));
  NAND2xp33_ASAP7_75t_L     g06205(.A(\b[1] ), .B(new_n5920), .Y(new_n6462));
  NAND5xp2_ASAP7_75t_L      g06206(.A(new_n6161), .B(new_n6159), .C(new_n6462), .D(new_n6158), .E(\a[41] ), .Y(new_n6463));
  A2O1A1Ixp33_ASAP7_75t_L   g06207(.A1(new_n312), .A2(new_n5637), .B(new_n6160), .C(new_n5626), .Y(new_n6464));
  NAND2xp33_ASAP7_75t_L     g06208(.A(new_n6463), .B(new_n6464), .Y(new_n6465));
  MAJIxp5_ASAP7_75t_L       g06209(.A(new_n6465), .B(new_n6153), .C(new_n6156), .Y(new_n6466));
  AOI221xp5_ASAP7_75t_L     g06210(.A1(\a[41] ), .A2(new_n6428), .B1(new_n6446), .B2(new_n6459), .C(new_n6432), .Y(new_n6467));
  AOI211xp5_ASAP7_75t_L     g06211(.A1(new_n6433), .A2(new_n6429), .B(new_n6447), .C(new_n6454), .Y(new_n6468));
  OAI21xp33_ASAP7_75t_L     g06212(.A1(new_n6467), .A2(new_n6468), .B(new_n6466), .Y(new_n6469));
  NAND3xp33_ASAP7_75t_L     g06213(.A(new_n6461), .B(new_n6469), .C(new_n6423), .Y(new_n6470));
  NOR3xp33_ASAP7_75t_L      g06214(.A(new_n6468), .B(new_n6466), .C(new_n6467), .Y(new_n6471));
  AOI21xp33_ASAP7_75t_L     g06215(.A1(new_n6460), .A2(new_n6455), .B(new_n6425), .Y(new_n6472));
  NOR3xp33_ASAP7_75t_L      g06216(.A(new_n6472), .B(new_n6471), .C(new_n6423), .Y(new_n6473));
  AOI21xp33_ASAP7_75t_L     g06217(.A1(new_n6470), .A2(new_n6423), .B(new_n6473), .Y(new_n6474));
  NAND3xp33_ASAP7_75t_L     g06218(.A(new_n6474), .B(new_n6188), .C(new_n6417), .Y(new_n6475));
  A2O1A1Ixp33_ASAP7_75t_L   g06219(.A1(new_n6174), .A2(new_n6175), .B(new_n6182), .C(new_n6417), .Y(new_n6476));
  A2O1A1Ixp33_ASAP7_75t_L   g06220(.A1(new_n6470), .A2(new_n6423), .B(new_n6473), .C(new_n6476), .Y(new_n6477));
  OAI22xp33_ASAP7_75t_L     g06221(.A1(new_n4397), .A2(new_n534), .B1(new_n590), .B2(new_n4142), .Y(new_n6478));
  AOI221xp5_ASAP7_75t_L     g06222(.A1(new_n4156), .A2(\b[10] ), .B1(new_n4151), .B2(new_n690), .C(new_n6478), .Y(new_n6479));
  XNOR2x2_ASAP7_75t_L       g06223(.A(\a[35] ), .B(new_n6479), .Y(new_n6480));
  NAND3xp33_ASAP7_75t_L     g06224(.A(new_n6475), .B(new_n6477), .C(new_n6480), .Y(new_n6481));
  INVx1_ASAP7_75t_L         g06225(.A(new_n6481), .Y(new_n6482));
  AOI21xp33_ASAP7_75t_L     g06226(.A1(new_n6475), .A2(new_n6477), .B(new_n6480), .Y(new_n6483));
  OAI21xp33_ASAP7_75t_L     g06227(.A1(new_n6482), .A2(new_n6483), .B(new_n6416), .Y(new_n6484));
  A2O1A1O1Ixp25_ASAP7_75t_L g06228(.A1(new_n5960), .A2(new_n6147), .B(new_n6148), .C(new_n6205), .D(new_n6201), .Y(new_n6485));
  NAND4xp25_ASAP7_75t_L     g06229(.A(new_n6461), .B(new_n6422), .C(new_n6420), .D(new_n6469), .Y(new_n6486));
  OAI21xp33_ASAP7_75t_L     g06230(.A1(new_n6471), .A2(new_n6472), .B(new_n6423), .Y(new_n6487));
  NAND2xp33_ASAP7_75t_L     g06231(.A(new_n6487), .B(new_n6486), .Y(new_n6488));
  NOR2xp33_ASAP7_75t_L      g06232(.A(new_n6488), .B(new_n6476), .Y(new_n6489));
  A2O1A1O1Ixp25_ASAP7_75t_L g06233(.A1(new_n6175), .A2(new_n6174), .B(new_n6182), .C(new_n6417), .D(new_n6474), .Y(new_n6490));
  XNOR2x2_ASAP7_75t_L       g06234(.A(new_n4145), .B(new_n6479), .Y(new_n6491));
  OAI21xp33_ASAP7_75t_L     g06235(.A1(new_n6489), .A2(new_n6490), .B(new_n6491), .Y(new_n6492));
  NAND3xp33_ASAP7_75t_L     g06236(.A(new_n6485), .B(new_n6481), .C(new_n6492), .Y(new_n6493));
  OAI22xp33_ASAP7_75t_L     g06237(.A1(new_n3703), .A2(new_n748), .B1(new_n833), .B2(new_n3509), .Y(new_n6494));
  AOI221xp5_ASAP7_75t_L     g06238(.A1(new_n3503), .A2(\b[13] ), .B1(new_n3505), .B2(new_n1166), .C(new_n6494), .Y(new_n6495));
  XNOR2x2_ASAP7_75t_L       g06239(.A(new_n3493), .B(new_n6495), .Y(new_n6496));
  AND3x1_ASAP7_75t_L        g06240(.A(new_n6484), .B(new_n6493), .C(new_n6496), .Y(new_n6497));
  O2A1O1Ixp33_ASAP7_75t_L   g06241(.A1(new_n6195), .A2(new_n6204), .B(new_n6206), .C(new_n6483), .Y(new_n6498));
  A2O1A1O1Ixp25_ASAP7_75t_L g06242(.A1(new_n6481), .A2(new_n6498), .B(new_n6485), .C(new_n6493), .D(new_n6496), .Y(new_n6499));
  NOR3xp33_ASAP7_75t_L      g06243(.A(new_n6415), .B(new_n6497), .C(new_n6499), .Y(new_n6500));
  NAND2xp33_ASAP7_75t_L     g06244(.A(new_n6208), .B(new_n6203), .Y(new_n6501));
  MAJIxp5_ASAP7_75t_L       g06245(.A(new_n6226), .B(new_n6146), .C(new_n6501), .Y(new_n6502));
  NAND3xp33_ASAP7_75t_L     g06246(.A(new_n6484), .B(new_n6493), .C(new_n6496), .Y(new_n6503));
  AO21x2_ASAP7_75t_L        g06247(.A1(new_n6493), .A2(new_n6484), .B(new_n6496), .Y(new_n6504));
  AOI21xp33_ASAP7_75t_L     g06248(.A1(new_n6504), .A2(new_n6503), .B(new_n6502), .Y(new_n6505));
  NOR2xp33_ASAP7_75t_L      g06249(.A(new_n1043), .B(new_n2925), .Y(new_n6506));
  AOI221xp5_ASAP7_75t_L     g06250(.A1(\b[14] ), .A2(new_n3129), .B1(\b[16] ), .B2(new_n2938), .C(new_n6506), .Y(new_n6507));
  INVx1_ASAP7_75t_L         g06251(.A(new_n6507), .Y(new_n6508));
  A2O1A1Ixp33_ASAP7_75t_L   g06252(.A1(new_n1156), .A2(new_n2932), .B(new_n6508), .C(\a[29] ), .Y(new_n6509));
  INVx1_ASAP7_75t_L         g06253(.A(new_n6509), .Y(new_n6510));
  A2O1A1Ixp33_ASAP7_75t_L   g06254(.A1(new_n1156), .A2(new_n2932), .B(new_n6508), .C(new_n2928), .Y(new_n6511));
  OAI21xp33_ASAP7_75t_L     g06255(.A1(new_n2928), .A2(new_n6510), .B(new_n6511), .Y(new_n6512));
  NOR3xp33_ASAP7_75t_L      g06256(.A(new_n6512), .B(new_n6500), .C(new_n6505), .Y(new_n6513));
  NAND3xp33_ASAP7_75t_L     g06257(.A(new_n6502), .B(new_n6504), .C(new_n6503), .Y(new_n6514));
  OAI21xp33_ASAP7_75t_L     g06258(.A1(new_n6499), .A2(new_n6497), .B(new_n6415), .Y(new_n6515));
  O2A1O1Ixp33_ASAP7_75t_L   g06259(.A1(new_n2940), .A2(new_n1161), .B(new_n6507), .C(\a[29] ), .Y(new_n6516));
  AOI21xp33_ASAP7_75t_L     g06260(.A1(new_n6509), .A2(\a[29] ), .B(new_n6516), .Y(new_n6517));
  AOI21xp33_ASAP7_75t_L     g06261(.A1(new_n6514), .A2(new_n6515), .B(new_n6517), .Y(new_n6518));
  A2O1A1Ixp33_ASAP7_75t_L   g06262(.A1(new_n6224), .A2(new_n6223), .B(new_n6231), .C(new_n6233), .Y(new_n6519));
  NOR3xp33_ASAP7_75t_L      g06263(.A(new_n6519), .B(new_n6518), .C(new_n6513), .Y(new_n6520));
  NAND3xp33_ASAP7_75t_L     g06264(.A(new_n6514), .B(new_n6515), .C(new_n6517), .Y(new_n6521));
  OAI21xp33_ASAP7_75t_L     g06265(.A1(new_n6505), .A2(new_n6500), .B(new_n6512), .Y(new_n6522));
  MAJIxp5_ASAP7_75t_L       g06266(.A(new_n6139), .B(new_n6232), .C(new_n6228), .Y(new_n6523));
  AOI21xp33_ASAP7_75t_L     g06267(.A1(new_n6522), .A2(new_n6521), .B(new_n6523), .Y(new_n6524));
  NOR2xp33_ASAP7_75t_L      g06268(.A(new_n1458), .B(new_n2410), .Y(new_n6525));
  AOI221xp5_ASAP7_75t_L     g06269(.A1(\b[17] ), .A2(new_n2577), .B1(\b[19] ), .B2(new_n2423), .C(new_n6525), .Y(new_n6526));
  O2A1O1Ixp33_ASAP7_75t_L   g06270(.A1(new_n2425), .A2(new_n1628), .B(new_n6526), .C(new_n2413), .Y(new_n6527));
  O2A1O1Ixp33_ASAP7_75t_L   g06271(.A1(new_n2425), .A2(new_n1628), .B(new_n6526), .C(\a[26] ), .Y(new_n6528));
  INVx1_ASAP7_75t_L         g06272(.A(new_n6528), .Y(new_n6529));
  OAI21xp33_ASAP7_75t_L     g06273(.A1(new_n2413), .A2(new_n6527), .B(new_n6529), .Y(new_n6530));
  NOR3xp33_ASAP7_75t_L      g06274(.A(new_n6530), .B(new_n6524), .C(new_n6520), .Y(new_n6531));
  NAND3xp33_ASAP7_75t_L     g06275(.A(new_n6523), .B(new_n6522), .C(new_n6521), .Y(new_n6532));
  OAI21xp33_ASAP7_75t_L     g06276(.A1(new_n6513), .A2(new_n6518), .B(new_n6519), .Y(new_n6533));
  INVx1_ASAP7_75t_L         g06277(.A(new_n6527), .Y(new_n6534));
  AOI21xp33_ASAP7_75t_L     g06278(.A1(new_n6534), .A2(\a[26] ), .B(new_n6528), .Y(new_n6535));
  AOI21xp33_ASAP7_75t_L     g06279(.A1(new_n6532), .A2(new_n6533), .B(new_n6535), .Y(new_n6536));
  OAI21xp33_ASAP7_75t_L     g06280(.A1(new_n6249), .A2(new_n6252), .B(new_n6253), .Y(new_n6537));
  NOR3xp33_ASAP7_75t_L      g06281(.A(new_n6537), .B(new_n6536), .C(new_n6531), .Y(new_n6538));
  NOR2xp33_ASAP7_75t_L      g06282(.A(new_n6524), .B(new_n6520), .Y(new_n6539));
  NAND2xp33_ASAP7_75t_L     g06283(.A(new_n6535), .B(new_n6539), .Y(new_n6540));
  NAND2xp33_ASAP7_75t_L     g06284(.A(new_n6533), .B(new_n6532), .Y(new_n6541));
  A2O1A1Ixp33_ASAP7_75t_L   g06285(.A1(\a[26] ), .A2(new_n6534), .B(new_n6528), .C(new_n6541), .Y(new_n6542));
  A2O1A1O1Ixp25_ASAP7_75t_L g06286(.A1(new_n5990), .A2(new_n5987), .B(new_n5989), .C(new_n6254), .D(new_n6242), .Y(new_n6543));
  AOI21xp33_ASAP7_75t_L     g06287(.A1(new_n6540), .A2(new_n6542), .B(new_n6543), .Y(new_n6544));
  NOR2xp33_ASAP7_75t_L      g06288(.A(new_n1895), .B(new_n1962), .Y(new_n6545));
  AOI221xp5_ASAP7_75t_L     g06289(.A1(new_n1955), .A2(\b[22] ), .B1(new_n2093), .B2(\b[20] ), .C(new_n6545), .Y(new_n6546));
  O2A1O1Ixp33_ASAP7_75t_L   g06290(.A1(new_n1956), .A2(new_n2522), .B(new_n6546), .C(new_n1952), .Y(new_n6547));
  O2A1O1Ixp33_ASAP7_75t_L   g06291(.A1(new_n1956), .A2(new_n2522), .B(new_n6546), .C(\a[23] ), .Y(new_n6548));
  INVx1_ASAP7_75t_L         g06292(.A(new_n6548), .Y(new_n6549));
  OAI21xp33_ASAP7_75t_L     g06293(.A1(new_n1952), .A2(new_n6547), .B(new_n6549), .Y(new_n6550));
  NOR3xp33_ASAP7_75t_L      g06294(.A(new_n6544), .B(new_n6538), .C(new_n6550), .Y(new_n6551));
  NAND3xp33_ASAP7_75t_L     g06295(.A(new_n6543), .B(new_n6540), .C(new_n6542), .Y(new_n6552));
  OAI21xp33_ASAP7_75t_L     g06296(.A1(new_n6531), .A2(new_n6536), .B(new_n6537), .Y(new_n6553));
  INVx1_ASAP7_75t_L         g06297(.A(new_n6547), .Y(new_n6554));
  AOI21xp33_ASAP7_75t_L     g06298(.A1(new_n6554), .A2(\a[23] ), .B(new_n6548), .Y(new_n6555));
  AOI21xp33_ASAP7_75t_L     g06299(.A1(new_n6552), .A2(new_n6553), .B(new_n6555), .Y(new_n6556));
  NOR2xp33_ASAP7_75t_L      g06300(.A(new_n6551), .B(new_n6556), .Y(new_n6557));
  NOR3xp33_ASAP7_75t_L      g06301(.A(new_n6264), .B(new_n6265), .C(new_n6262), .Y(new_n6558));
  A2O1A1O1Ixp25_ASAP7_75t_L g06302(.A1(new_n6277), .A2(new_n6006), .B(new_n6274), .C(new_n6278), .D(new_n6558), .Y(new_n6559));
  NAND2xp33_ASAP7_75t_L     g06303(.A(new_n6557), .B(new_n6559), .Y(new_n6560));
  NAND3xp33_ASAP7_75t_L     g06304(.A(new_n6552), .B(new_n6555), .C(new_n6553), .Y(new_n6561));
  OAI21xp33_ASAP7_75t_L     g06305(.A1(new_n6538), .A2(new_n6544), .B(new_n6550), .Y(new_n6562));
  NAND2xp33_ASAP7_75t_L     g06306(.A(new_n6562), .B(new_n6561), .Y(new_n6563));
  INVx1_ASAP7_75t_L         g06307(.A(new_n6558), .Y(new_n6564));
  A2O1A1Ixp33_ASAP7_75t_L   g06308(.A1(new_n6262), .A2(new_n6263), .B(new_n6271), .C(new_n6564), .Y(new_n6565));
  NAND2xp33_ASAP7_75t_L     g06309(.A(new_n6563), .B(new_n6565), .Y(new_n6566));
  NAND2xp33_ASAP7_75t_L     g06310(.A(\b[24] ), .B(new_n1507), .Y(new_n6567));
  OAI221xp5_ASAP7_75t_L     g06311(.A1(new_n1518), .A2(new_n2377), .B1(new_n2188), .B2(new_n1654), .C(new_n6567), .Y(new_n6568));
  A2O1A1Ixp33_ASAP7_75t_L   g06312(.A1(new_n5001), .A2(new_n1513), .B(new_n6568), .C(\a[20] ), .Y(new_n6569));
  AOI211xp5_ASAP7_75t_L     g06313(.A1(new_n5001), .A2(new_n1513), .B(new_n6568), .C(new_n1501), .Y(new_n6570));
  A2O1A1O1Ixp25_ASAP7_75t_L g06314(.A1(new_n5001), .A2(new_n1513), .B(new_n6568), .C(new_n6569), .D(new_n6570), .Y(new_n6571));
  NAND3xp33_ASAP7_75t_L     g06315(.A(new_n6560), .B(new_n6566), .C(new_n6571), .Y(new_n6572));
  NOR2xp33_ASAP7_75t_L      g06316(.A(new_n6563), .B(new_n6565), .Y(new_n6573));
  O2A1O1Ixp33_ASAP7_75t_L   g06317(.A1(new_n6269), .A2(new_n6271), .B(new_n6564), .C(new_n6557), .Y(new_n6574));
  INVx1_ASAP7_75t_L         g06318(.A(new_n6571), .Y(new_n6575));
  OAI21xp33_ASAP7_75t_L     g06319(.A1(new_n6573), .A2(new_n6574), .B(new_n6575), .Y(new_n6576));
  A2O1A1O1Ixp25_ASAP7_75t_L g06320(.A1(new_n6021), .A2(new_n5894), .B(new_n6015), .C(new_n6286), .D(new_n6284), .Y(new_n6577));
  AOI21xp33_ASAP7_75t_L     g06321(.A1(new_n6576), .A2(new_n6572), .B(new_n6577), .Y(new_n6578));
  NOR3xp33_ASAP7_75t_L      g06322(.A(new_n6574), .B(new_n6575), .C(new_n6573), .Y(new_n6579));
  AOI21xp33_ASAP7_75t_L     g06323(.A1(new_n6560), .A2(new_n6566), .B(new_n6571), .Y(new_n6580));
  A2O1A1Ixp33_ASAP7_75t_L   g06324(.A1(new_n5762), .A2(new_n5764), .B(new_n6018), .C(new_n6021), .Y(new_n6581));
  A2O1A1Ixp33_ASAP7_75t_L   g06325(.A1(new_n6581), .A2(new_n6020), .B(new_n6283), .C(new_n6287), .Y(new_n6582));
  NOR3xp33_ASAP7_75t_L      g06326(.A(new_n6582), .B(new_n6580), .C(new_n6579), .Y(new_n6583));
  OAI21xp33_ASAP7_75t_L     g06327(.A1(new_n6583), .A2(new_n6578), .B(new_n6413), .Y(new_n6584));
  OAI211xp5_ASAP7_75t_L     g06328(.A1(new_n1210), .A2(new_n3087), .B(\a[17] ), .C(new_n6409), .Y(new_n6585));
  OAI21xp33_ASAP7_75t_L     g06329(.A1(new_n6579), .A2(new_n6580), .B(new_n6582), .Y(new_n6586));
  NAND3xp33_ASAP7_75t_L     g06330(.A(new_n6577), .B(new_n6576), .C(new_n6572), .Y(new_n6587));
  NAND4xp25_ASAP7_75t_L     g06331(.A(new_n6587), .B(new_n6585), .C(new_n6412), .D(new_n6586), .Y(new_n6588));
  NAND3xp33_ASAP7_75t_L     g06332(.A(new_n6407), .B(new_n6584), .C(new_n6588), .Y(new_n6589));
  MAJIxp5_ASAP7_75t_L       g06333(.A(new_n6138), .B(new_n6289), .C(new_n6303), .Y(new_n6590));
  NAND2xp33_ASAP7_75t_L     g06334(.A(new_n6584), .B(new_n6588), .Y(new_n6591));
  NAND2xp33_ASAP7_75t_L     g06335(.A(new_n6590), .B(new_n6591), .Y(new_n6592));
  NOR2xp33_ASAP7_75t_L      g06336(.A(new_n3456), .B(new_n864), .Y(new_n6593));
  AOI221xp5_ASAP7_75t_L     g06337(.A1(\b[29] ), .A2(new_n985), .B1(\b[31] ), .B2(new_n886), .C(new_n6593), .Y(new_n6594));
  O2A1O1Ixp33_ASAP7_75t_L   g06338(.A1(new_n872), .A2(new_n3681), .B(new_n6594), .C(new_n867), .Y(new_n6595));
  INVx1_ASAP7_75t_L         g06339(.A(new_n6595), .Y(new_n6596));
  O2A1O1Ixp33_ASAP7_75t_L   g06340(.A1(new_n872), .A2(new_n3681), .B(new_n6594), .C(\a[14] ), .Y(new_n6597));
  AOI21xp33_ASAP7_75t_L     g06341(.A1(new_n6596), .A2(\a[14] ), .B(new_n6597), .Y(new_n6598));
  NAND3xp33_ASAP7_75t_L     g06342(.A(new_n6589), .B(new_n6592), .C(new_n6598), .Y(new_n6599));
  O2A1O1Ixp33_ASAP7_75t_L   g06343(.A1(new_n1210), .A2(new_n2889), .B(new_n6291), .C(\a[17] ), .Y(new_n6600));
  A2O1A1Ixp33_ASAP7_75t_L   g06344(.A1(\a[17] ), .A2(new_n6293), .B(new_n6600), .C(new_n6289), .Y(new_n6601));
  A2O1A1O1Ixp25_ASAP7_75t_L g06345(.A1(new_n6304), .A2(new_n6300), .B(new_n6307), .C(new_n6601), .D(new_n6591), .Y(new_n6602));
  AOI21xp33_ASAP7_75t_L     g06346(.A1(new_n6588), .A2(new_n6584), .B(new_n6407), .Y(new_n6603));
  AO21x2_ASAP7_75t_L        g06347(.A1(\a[14] ), .A2(new_n6596), .B(new_n6597), .Y(new_n6604));
  OAI21xp33_ASAP7_75t_L     g06348(.A1(new_n6603), .A2(new_n6602), .B(new_n6604), .Y(new_n6605));
  NAND3xp33_ASAP7_75t_L     g06349(.A(new_n6406), .B(new_n6599), .C(new_n6605), .Y(new_n6606));
  A2O1A1O1Ixp25_ASAP7_75t_L g06350(.A1(new_n6053), .A2(new_n5884), .B(new_n6045), .C(new_n6324), .D(new_n6317), .Y(new_n6607));
  NOR3xp33_ASAP7_75t_L      g06351(.A(new_n6602), .B(new_n6603), .C(new_n6604), .Y(new_n6608));
  AOI21xp33_ASAP7_75t_L     g06352(.A1(new_n6589), .A2(new_n6592), .B(new_n6598), .Y(new_n6609));
  OAI21xp33_ASAP7_75t_L     g06353(.A1(new_n6609), .A2(new_n6608), .B(new_n6607), .Y(new_n6610));
  NAND2xp33_ASAP7_75t_L     g06354(.A(new_n6606), .B(new_n6610), .Y(new_n6611));
  NOR2xp33_ASAP7_75t_L      g06355(.A(new_n4101), .B(new_n1550), .Y(new_n6612));
  AOI221xp5_ASAP7_75t_L     g06356(.A1(\b[32] ), .A2(new_n713), .B1(\b[34] ), .B2(new_n640), .C(new_n6612), .Y(new_n6613));
  NAND2xp33_ASAP7_75t_L     g06357(.A(new_n718), .B(new_n5599), .Y(new_n6614));
  O2A1O1Ixp33_ASAP7_75t_L   g06358(.A1(new_n641), .A2(new_n4352), .B(new_n6613), .C(new_n637), .Y(new_n6615));
  INVx1_ASAP7_75t_L         g06359(.A(new_n6613), .Y(new_n6616));
  A2O1A1Ixp33_ASAP7_75t_L   g06360(.A1(new_n5599), .A2(new_n718), .B(new_n6616), .C(\a[11] ), .Y(new_n6617));
  NAND2xp33_ASAP7_75t_L     g06361(.A(\a[11] ), .B(new_n6617), .Y(new_n6618));
  A2O1A1Ixp33_ASAP7_75t_L   g06362(.A1(new_n6614), .A2(new_n6613), .B(new_n6615), .C(new_n6618), .Y(new_n6619));
  NOR2xp33_ASAP7_75t_L      g06363(.A(new_n6619), .B(new_n6611), .Y(new_n6620));
  NOR2xp33_ASAP7_75t_L      g06364(.A(new_n637), .B(new_n6615), .Y(new_n6621));
  A2O1A1O1Ixp25_ASAP7_75t_L g06365(.A1(new_n5599), .A2(new_n718), .B(new_n6616), .C(new_n6617), .D(new_n6621), .Y(new_n6622));
  AOI21xp33_ASAP7_75t_L     g06366(.A1(new_n6606), .A2(new_n6610), .B(new_n6622), .Y(new_n6623));
  NAND2xp33_ASAP7_75t_L     g06367(.A(new_n6335), .B(new_n6334), .Y(new_n6624));
  MAJIxp5_ASAP7_75t_L       g06368(.A(new_n6136), .B(new_n6336), .C(new_n6624), .Y(new_n6625));
  NOR3xp33_ASAP7_75t_L      g06369(.A(new_n6620), .B(new_n6625), .C(new_n6623), .Y(new_n6626));
  NOR2xp33_ASAP7_75t_L      g06370(.A(new_n6622), .B(new_n6611), .Y(new_n6627));
  NAND3xp33_ASAP7_75t_L     g06371(.A(new_n6622), .B(new_n6610), .C(new_n6606), .Y(new_n6628));
  NOR2xp33_ASAP7_75t_L      g06372(.A(new_n6322), .B(new_n6325), .Y(new_n6629));
  MAJIxp5_ASAP7_75t_L       g06373(.A(new_n6339), .B(new_n6629), .C(new_n6331), .Y(new_n6630));
  O2A1O1Ixp33_ASAP7_75t_L   g06374(.A1(new_n6622), .A2(new_n6627), .B(new_n6628), .C(new_n6630), .Y(new_n6631));
  NOR2xp33_ASAP7_75t_L      g06375(.A(new_n4581), .B(new_n506), .Y(new_n6632));
  AOI221xp5_ASAP7_75t_L     g06376(.A1(\b[37] ), .A2(new_n475), .B1(new_n470), .B2(\b[36] ), .C(new_n6632), .Y(new_n6633));
  O2A1O1Ixp33_ASAP7_75t_L   g06377(.A1(new_n477), .A2(new_n5083), .B(new_n6633), .C(new_n466), .Y(new_n6634));
  OAI21xp33_ASAP7_75t_L     g06378(.A1(new_n477), .A2(new_n5083), .B(new_n6633), .Y(new_n6635));
  NAND2xp33_ASAP7_75t_L     g06379(.A(new_n466), .B(new_n6635), .Y(new_n6636));
  OAI21xp33_ASAP7_75t_L     g06380(.A1(new_n466), .A2(new_n6634), .B(new_n6636), .Y(new_n6637));
  INVx1_ASAP7_75t_L         g06381(.A(new_n6637), .Y(new_n6638));
  NOR3xp33_ASAP7_75t_L      g06382(.A(new_n6631), .B(new_n6638), .C(new_n6626), .Y(new_n6639));
  OAI211xp5_ASAP7_75t_L     g06383(.A1(new_n6622), .A2(new_n6627), .B(new_n6628), .C(new_n6630), .Y(new_n6640));
  OAI21xp33_ASAP7_75t_L     g06384(.A1(new_n6623), .A2(new_n6620), .B(new_n6625), .Y(new_n6641));
  AOI21xp33_ASAP7_75t_L     g06385(.A1(new_n6640), .A2(new_n6641), .B(new_n6637), .Y(new_n6642));
  OAI22xp33_ASAP7_75t_L     g06386(.A1(new_n6366), .A2(new_n6355), .B1(new_n6642), .B2(new_n6639), .Y(new_n6643));
  A2O1A1O1Ixp25_ASAP7_75t_L g06387(.A1(new_n6092), .A2(new_n6095), .B(new_n6097), .C(new_n6359), .D(new_n6355), .Y(new_n6644));
  NAND3xp33_ASAP7_75t_L     g06388(.A(new_n6640), .B(new_n6641), .C(new_n6637), .Y(new_n6645));
  OAI21xp33_ASAP7_75t_L     g06389(.A1(new_n6626), .A2(new_n6631), .B(new_n6638), .Y(new_n6646));
  NAND3xp33_ASAP7_75t_L     g06390(.A(new_n6644), .B(new_n6645), .C(new_n6646), .Y(new_n6647));
  NOR2xp33_ASAP7_75t_L      g06391(.A(new_n5311), .B(new_n375), .Y(new_n6648));
  AOI221xp5_ASAP7_75t_L     g06392(.A1(\b[40] ), .A2(new_n361), .B1(new_n349), .B2(\b[39] ), .C(new_n6648), .Y(new_n6649));
  O2A1O1Ixp33_ASAP7_75t_L   g06393(.A1(new_n356), .A2(new_n5862), .B(new_n6649), .C(new_n346), .Y(new_n6650));
  INVx1_ASAP7_75t_L         g06394(.A(new_n5862), .Y(new_n6651));
  INVx1_ASAP7_75t_L         g06395(.A(new_n6649), .Y(new_n6652));
  A2O1A1Ixp33_ASAP7_75t_L   g06396(.A1(new_n6651), .A2(new_n359), .B(new_n6652), .C(new_n346), .Y(new_n6653));
  OAI21xp33_ASAP7_75t_L     g06397(.A1(new_n346), .A2(new_n6650), .B(new_n6653), .Y(new_n6654));
  INVx1_ASAP7_75t_L         g06398(.A(new_n6654), .Y(new_n6655));
  NAND3xp33_ASAP7_75t_L     g06399(.A(new_n6647), .B(new_n6643), .C(new_n6655), .Y(new_n6656));
  AOI21xp33_ASAP7_75t_L     g06400(.A1(new_n6646), .A2(new_n6645), .B(new_n6644), .Y(new_n6657));
  OAI21xp33_ASAP7_75t_L     g06401(.A1(new_n6074), .A2(new_n6076), .B(new_n6078), .Y(new_n6658));
  A2O1A1O1Ixp25_ASAP7_75t_L g06402(.A1(new_n6359), .A2(new_n6658), .B(new_n6355), .C(new_n6646), .D(new_n6639), .Y(new_n6659));
  A2O1A1Ixp33_ASAP7_75t_L   g06403(.A1(new_n6659), .A2(new_n6646), .B(new_n6657), .C(new_n6654), .Y(new_n6660));
  NAND3xp33_ASAP7_75t_L     g06404(.A(new_n6405), .B(new_n6656), .C(new_n6660), .Y(new_n6661));
  NOR2xp33_ASAP7_75t_L      g06405(.A(new_n6367), .B(new_n6366), .Y(new_n6662));
  A2O1A1Ixp33_ASAP7_75t_L   g06406(.A1(new_n6133), .A2(\a[5] ), .B(new_n6134), .C(new_n6662), .Y(new_n6663));
  NOR2xp33_ASAP7_75t_L      g06407(.A(new_n6363), .B(new_n6368), .Y(new_n6664));
  AOI211xp5_ASAP7_75t_L     g06408(.A1(new_n6659), .A2(new_n6646), .B(new_n6654), .C(new_n6657), .Y(new_n6665));
  AOI21xp33_ASAP7_75t_L     g06409(.A1(new_n6647), .A2(new_n6643), .B(new_n6655), .Y(new_n6666));
  OAI221xp5_ASAP7_75t_L     g06410(.A1(new_n6664), .A2(new_n6129), .B1(new_n6666), .B2(new_n6665), .C(new_n6663), .Y(new_n6667));
  NOR2xp33_ASAP7_75t_L      g06411(.A(new_n6110), .B(new_n287), .Y(new_n6668));
  AOI221xp5_ASAP7_75t_L     g06412(.A1(\b[42] ), .A2(new_n264), .B1(\b[43] ), .B2(new_n283), .C(new_n6668), .Y(new_n6669));
  NOR2xp33_ASAP7_75t_L      g06413(.A(\b[42] ), .B(\b[43] ), .Y(new_n6670));
  INVx1_ASAP7_75t_L         g06414(.A(\b[43] ), .Y(new_n6671));
  NOR2xp33_ASAP7_75t_L      g06415(.A(new_n6378), .B(new_n6671), .Y(new_n6672));
  NOR2xp33_ASAP7_75t_L      g06416(.A(new_n6670), .B(new_n6672), .Y(new_n6673));
  A2O1A1Ixp33_ASAP7_75t_L   g06417(.A1(\b[42] ), .A2(\b[41] ), .B(new_n6382), .C(new_n6673), .Y(new_n6674));
  O2A1O1Ixp33_ASAP7_75t_L   g06418(.A1(new_n5570), .A2(new_n5855), .B(new_n5858), .C(new_n6115), .Y(new_n6675));
  O2A1O1Ixp33_ASAP7_75t_L   g06419(.A1(new_n6111), .A2(new_n6675), .B(new_n6380), .C(new_n6379), .Y(new_n6676));
  INVx1_ASAP7_75t_L         g06420(.A(new_n6673), .Y(new_n6677));
  NAND2xp33_ASAP7_75t_L     g06421(.A(new_n6677), .B(new_n6676), .Y(new_n6678));
  NAND2xp33_ASAP7_75t_L     g06422(.A(new_n6674), .B(new_n6678), .Y(new_n6679));
  O2A1O1Ixp33_ASAP7_75t_L   g06423(.A1(new_n279), .A2(new_n6679), .B(new_n6669), .C(new_n257), .Y(new_n6680));
  INVx1_ASAP7_75t_L         g06424(.A(new_n6669), .Y(new_n6681));
  INVx1_ASAP7_75t_L         g06425(.A(new_n6679), .Y(new_n6682));
  A2O1A1Ixp33_ASAP7_75t_L   g06426(.A1(new_n6682), .A2(new_n273), .B(new_n6681), .C(new_n257), .Y(new_n6683));
  OAI21xp33_ASAP7_75t_L     g06427(.A1(new_n257), .A2(new_n6680), .B(new_n6683), .Y(new_n6684));
  NAND3xp33_ASAP7_75t_L     g06428(.A(new_n6661), .B(new_n6667), .C(new_n6684), .Y(new_n6685));
  INVx1_ASAP7_75t_L         g06429(.A(new_n6684), .Y(new_n6686));
  AOI21xp33_ASAP7_75t_L     g06430(.A1(new_n6661), .A2(new_n6667), .B(new_n6686), .Y(new_n6687));
  AOI31xp33_ASAP7_75t_L     g06431(.A1(new_n6685), .A2(new_n6661), .A3(new_n6667), .B(new_n6687), .Y(new_n6688));
  O2A1O1Ixp33_ASAP7_75t_L   g06432(.A1(new_n6129), .A2(new_n6394), .B(new_n6396), .C(new_n6392), .Y(new_n6689));
  AOI21xp33_ASAP7_75t_L     g06433(.A1(new_n6401), .A2(new_n6398), .B(new_n6689), .Y(new_n6690));
  XOR2x2_ASAP7_75t_L        g06434(.A(new_n6688), .B(new_n6690), .Y(\f[43] ));
  NOR2xp33_ASAP7_75t_L      g06435(.A(new_n5570), .B(new_n375), .Y(new_n6692));
  AOI221xp5_ASAP7_75t_L     g06436(.A1(\b[41] ), .A2(new_n361), .B1(new_n349), .B2(\b[40] ), .C(new_n6692), .Y(new_n6693));
  O2A1O1Ixp33_ASAP7_75t_L   g06437(.A1(new_n356), .A2(new_n6117), .B(new_n6693), .C(new_n346), .Y(new_n6694));
  INVx1_ASAP7_75t_L         g06438(.A(new_n6693), .Y(new_n6695));
  A2O1A1Ixp33_ASAP7_75t_L   g06439(.A1(new_n6118), .A2(new_n359), .B(new_n6695), .C(new_n346), .Y(new_n6696));
  OAI21xp33_ASAP7_75t_L     g06440(.A1(new_n346), .A2(new_n6694), .B(new_n6696), .Y(new_n6697));
  A2O1A1Ixp33_ASAP7_75t_L   g06441(.A1(new_n6658), .A2(new_n6356), .B(new_n6355), .C(new_n6646), .Y(new_n6698));
  A2O1A1O1Ixp25_ASAP7_75t_L g06442(.A1(new_n6324), .A2(new_n6333), .B(new_n6317), .C(new_n6599), .D(new_n6609), .Y(new_n6699));
  NOR2xp33_ASAP7_75t_L      g06443(.A(new_n3674), .B(new_n864), .Y(new_n6700));
  AOI221xp5_ASAP7_75t_L     g06444(.A1(\b[30] ), .A2(new_n985), .B1(\b[32] ), .B2(new_n886), .C(new_n6700), .Y(new_n6701));
  O2A1O1Ixp33_ASAP7_75t_L   g06445(.A1(new_n872), .A2(new_n3897), .B(new_n6701), .C(new_n867), .Y(new_n6702));
  INVx1_ASAP7_75t_L         g06446(.A(new_n6701), .Y(new_n6703));
  A2O1A1Ixp33_ASAP7_75t_L   g06447(.A1(new_n3900), .A2(new_n873), .B(new_n6703), .C(new_n867), .Y(new_n6704));
  OAI21xp33_ASAP7_75t_L     g06448(.A1(new_n867), .A2(new_n6702), .B(new_n6704), .Y(new_n6705));
  NAND2xp33_ASAP7_75t_L     g06449(.A(new_n6586), .B(new_n6587), .Y(new_n6706));
  NOR2xp33_ASAP7_75t_L      g06450(.A(new_n6583), .B(new_n6578), .Y(new_n6707));
  NAND2xp33_ASAP7_75t_L     g06451(.A(new_n6413), .B(new_n6707), .Y(new_n6708));
  A2O1A1Ixp33_ASAP7_75t_L   g06452(.A1(new_n6584), .A2(new_n6706), .B(new_n6590), .C(new_n6708), .Y(new_n6709));
  OAI22xp33_ASAP7_75t_L     g06453(.A1(new_n1285), .A2(new_n2879), .B1(new_n3079), .B2(new_n2118), .Y(new_n6710));
  AOI221xp5_ASAP7_75t_L     g06454(.A1(new_n1209), .A2(\b[29] ), .B1(new_n1216), .B2(new_n3873), .C(new_n6710), .Y(new_n6711));
  XNOR2x2_ASAP7_75t_L       g06455(.A(new_n1206), .B(new_n6711), .Y(new_n6712));
  NOR2xp33_ASAP7_75t_L      g06456(.A(new_n6573), .B(new_n6574), .Y(new_n6713));
  MAJIxp5_ASAP7_75t_L       g06457(.A(new_n6582), .B(new_n6575), .C(new_n6713), .Y(new_n6714));
  NAND2xp33_ASAP7_75t_L     g06458(.A(new_n6515), .B(new_n6514), .Y(new_n6715));
  O2A1O1Ixp33_ASAP7_75t_L   g06459(.A1(new_n6510), .A2(new_n2928), .B(new_n6511), .C(new_n6715), .Y(new_n6716));
  NAND2xp33_ASAP7_75t_L     g06460(.A(new_n6521), .B(new_n6522), .Y(new_n6717));
  NAND2xp33_ASAP7_75t_L     g06461(.A(\b[16] ), .B(new_n2936), .Y(new_n6718));
  OAI221xp5_ASAP7_75t_L     g06462(.A1(new_n2930), .A2(new_n1349), .B1(new_n1043), .B2(new_n3133), .C(new_n6718), .Y(new_n6719));
  AOI211xp5_ASAP7_75t_L     g06463(.A1(new_n1633), .A2(new_n2932), .B(new_n6719), .C(new_n2928), .Y(new_n6720));
  INVx1_ASAP7_75t_L         g06464(.A(new_n6720), .Y(new_n6721));
  A2O1A1Ixp33_ASAP7_75t_L   g06465(.A1(new_n1633), .A2(new_n2932), .B(new_n6719), .C(new_n2928), .Y(new_n6722));
  NAND2xp33_ASAP7_75t_L     g06466(.A(new_n6722), .B(new_n6721), .Y(new_n6723));
  NAND2xp33_ASAP7_75t_L     g06467(.A(new_n6210), .B(new_n6414), .Y(new_n6724));
  A2O1A1Ixp33_ASAP7_75t_L   g06468(.A1(new_n6214), .A2(new_n6724), .B(new_n6497), .C(new_n6504), .Y(new_n6725));
  NOR2xp33_ASAP7_75t_L      g06469(.A(new_n936), .B(new_n3509), .Y(new_n6726));
  AOI221xp5_ASAP7_75t_L     g06470(.A1(\b[12] ), .A2(new_n3708), .B1(\b[14] ), .B2(new_n3503), .C(new_n6726), .Y(new_n6727));
  INVx1_ASAP7_75t_L         g06471(.A(new_n6727), .Y(new_n6728));
  A2O1A1Ixp33_ASAP7_75t_L   g06472(.A1(new_n971), .A2(new_n3505), .B(new_n6728), .C(\a[32] ), .Y(new_n6729));
  O2A1O1Ixp33_ASAP7_75t_L   g06473(.A1(new_n3513), .A2(new_n1268), .B(new_n6727), .C(\a[32] ), .Y(new_n6730));
  AOI21xp33_ASAP7_75t_L     g06474(.A1(new_n6729), .A2(\a[32] ), .B(new_n6730), .Y(new_n6731));
  OAI21xp33_ASAP7_75t_L     g06475(.A1(new_n5946), .A2(new_n5948), .B(new_n5942), .Y(new_n6732));
  A2O1A1Ixp33_ASAP7_75t_L   g06476(.A1(new_n6732), .A2(new_n6205), .B(new_n6201), .C(new_n6492), .Y(new_n6733));
  NOR2xp33_ASAP7_75t_L      g06477(.A(new_n448), .B(new_n4903), .Y(new_n6734));
  AOI221xp5_ASAP7_75t_L     g06478(.A1(\b[6] ), .A2(new_n5139), .B1(\b[8] ), .B2(new_n4917), .C(new_n6734), .Y(new_n6735));
  O2A1O1Ixp33_ASAP7_75t_L   g06479(.A1(new_n4911), .A2(new_n540), .B(new_n6735), .C(new_n4906), .Y(new_n6736));
  O2A1O1Ixp33_ASAP7_75t_L   g06480(.A1(new_n4911), .A2(new_n540), .B(new_n6735), .C(\a[38] ), .Y(new_n6737));
  INVx1_ASAP7_75t_L         g06481(.A(new_n6737), .Y(new_n6738));
  OAI21xp33_ASAP7_75t_L     g06482(.A1(new_n4906), .A2(new_n6736), .B(new_n6738), .Y(new_n6739));
  NAND2xp33_ASAP7_75t_L     g06483(.A(\b[2] ), .B(new_n6442), .Y(new_n6740));
  NAND3xp33_ASAP7_75t_L     g06484(.A(new_n6152), .B(new_n6435), .C(new_n6441), .Y(new_n6741));
  INVx1_ASAP7_75t_L         g06485(.A(new_n6741), .Y(new_n6742));
  NAND2xp33_ASAP7_75t_L     g06486(.A(\b[0] ), .B(new_n6742), .Y(new_n6743));
  NAND2xp33_ASAP7_75t_L     g06487(.A(\b[1] ), .B(new_n6436), .Y(new_n6744));
  NOR2xp33_ASAP7_75t_L      g06488(.A(new_n6443), .B(new_n509), .Y(new_n6745));
  INVx1_ASAP7_75t_L         g06489(.A(new_n6745), .Y(new_n6746));
  NAND5xp2_ASAP7_75t_L      g06490(.A(\a[44] ), .B(new_n6743), .C(new_n6746), .D(new_n6744), .E(new_n6740), .Y(new_n6747));
  OAI211xp5_ASAP7_75t_L     g06491(.A1(new_n284), .A2(new_n6741), .B(new_n6740), .C(new_n6744), .Y(new_n6748));
  A2O1A1Ixp33_ASAP7_75t_L   g06492(.A1(new_n294), .A2(new_n6450), .B(new_n6748), .C(new_n6439), .Y(new_n6749));
  NAND3xp33_ASAP7_75t_L     g06493(.A(new_n6749), .B(new_n6747), .C(new_n6446), .Y(new_n6750));
  NOR2xp33_ASAP7_75t_L      g06494(.A(new_n284), .B(new_n6741), .Y(new_n6751));
  AOI221xp5_ASAP7_75t_L     g06495(.A1(\b[2] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[1] ), .C(new_n6751), .Y(new_n6752));
  NAND5xp2_ASAP7_75t_L      g06496(.A(\a[44] ), .B(new_n6752), .C(new_n6746), .D(new_n6445), .E(new_n6424), .Y(new_n6753));
  NOR2xp33_ASAP7_75t_L      g06497(.A(new_n384), .B(new_n5641), .Y(new_n6754));
  AOI221xp5_ASAP7_75t_L     g06498(.A1(\b[3] ), .A2(new_n5920), .B1(\b[4] ), .B2(new_n5623), .C(new_n6754), .Y(new_n6755));
  OAI211xp5_ASAP7_75t_L     g06499(.A1(new_n5630), .A2(new_n728), .B(\a[41] ), .C(new_n6755), .Y(new_n6756));
  OAI21xp33_ASAP7_75t_L     g06500(.A1(new_n5630), .A2(new_n728), .B(new_n6755), .Y(new_n6757));
  NAND2xp33_ASAP7_75t_L     g06501(.A(new_n5626), .B(new_n6757), .Y(new_n6758));
  AND4x1_ASAP7_75t_L        g06502(.A(new_n6750), .B(new_n6758), .C(new_n6753), .D(new_n6756), .Y(new_n6759));
  AOI22xp33_ASAP7_75t_L     g06503(.A1(new_n6756), .A2(new_n6758), .B1(new_n6753), .B2(new_n6750), .Y(new_n6760));
  NOR2xp33_ASAP7_75t_L      g06504(.A(new_n6760), .B(new_n6759), .Y(new_n6761));
  O2A1O1Ixp33_ASAP7_75t_L   g06505(.A1(new_n6466), .A2(new_n6467), .B(new_n6460), .C(new_n6761), .Y(new_n6762));
  OAI21xp33_ASAP7_75t_L     g06506(.A1(new_n6467), .A2(new_n6466), .B(new_n6460), .Y(new_n6763));
  NOR3xp33_ASAP7_75t_L      g06507(.A(new_n6763), .B(new_n6759), .C(new_n6760), .Y(new_n6764));
  OAI21xp33_ASAP7_75t_L     g06508(.A1(new_n6764), .A2(new_n6762), .B(new_n6739), .Y(new_n6765));
  INVx1_ASAP7_75t_L         g06509(.A(new_n6736), .Y(new_n6766));
  AOI21xp33_ASAP7_75t_L     g06510(.A1(new_n6766), .A2(\a[38] ), .B(new_n6737), .Y(new_n6767));
  OAI21xp33_ASAP7_75t_L     g06511(.A1(new_n6759), .A2(new_n6760), .B(new_n6763), .Y(new_n6768));
  AOI21xp33_ASAP7_75t_L     g06512(.A1(new_n6425), .A2(new_n6455), .B(new_n6468), .Y(new_n6769));
  NAND2xp33_ASAP7_75t_L     g06513(.A(new_n6761), .B(new_n6769), .Y(new_n6770));
  NAND3xp33_ASAP7_75t_L     g06514(.A(new_n6770), .B(new_n6767), .C(new_n6768), .Y(new_n6771));
  NAND2xp33_ASAP7_75t_L     g06515(.A(new_n6771), .B(new_n6765), .Y(new_n6772));
  A2O1A1O1Ixp25_ASAP7_75t_L g06516(.A1(new_n6188), .A2(new_n6417), .B(new_n6474), .C(new_n6470), .D(new_n6772), .Y(new_n6773));
  A2O1A1Ixp33_ASAP7_75t_L   g06517(.A1(new_n6188), .A2(new_n6417), .B(new_n6474), .C(new_n6470), .Y(new_n6774));
  AOI21xp33_ASAP7_75t_L     g06518(.A1(new_n6770), .A2(new_n6768), .B(new_n6767), .Y(new_n6775));
  NOR3xp33_ASAP7_75t_L      g06519(.A(new_n6762), .B(new_n6764), .C(new_n6739), .Y(new_n6776));
  NOR2xp33_ASAP7_75t_L      g06520(.A(new_n6775), .B(new_n6776), .Y(new_n6777));
  NOR2xp33_ASAP7_75t_L      g06521(.A(new_n6777), .B(new_n6774), .Y(new_n6778));
  NOR2xp33_ASAP7_75t_L      g06522(.A(new_n680), .B(new_n4142), .Y(new_n6779));
  AOI221xp5_ASAP7_75t_L     g06523(.A1(\b[9] ), .A2(new_n4402), .B1(\b[11] ), .B2(new_n4156), .C(new_n6779), .Y(new_n6780));
  O2A1O1Ixp33_ASAP7_75t_L   g06524(.A1(new_n4150), .A2(new_n754), .B(new_n6780), .C(new_n4145), .Y(new_n6781));
  INVx1_ASAP7_75t_L         g06525(.A(new_n6781), .Y(new_n6782));
  O2A1O1Ixp33_ASAP7_75t_L   g06526(.A1(new_n4150), .A2(new_n754), .B(new_n6780), .C(\a[35] ), .Y(new_n6783));
  AOI21xp33_ASAP7_75t_L     g06527(.A1(new_n6782), .A2(\a[35] ), .B(new_n6783), .Y(new_n6784));
  INVx1_ASAP7_75t_L         g06528(.A(new_n6784), .Y(new_n6785));
  NOR3xp33_ASAP7_75t_L      g06529(.A(new_n6785), .B(new_n6773), .C(new_n6778), .Y(new_n6786));
  INVx1_ASAP7_75t_L         g06530(.A(new_n6470), .Y(new_n6787));
  AOI21xp33_ASAP7_75t_L     g06531(.A1(new_n6476), .A2(new_n6488), .B(new_n6787), .Y(new_n6788));
  NOR2xp33_ASAP7_75t_L      g06532(.A(new_n6777), .B(new_n6788), .Y(new_n6789));
  NAND2xp33_ASAP7_75t_L     g06533(.A(new_n6772), .B(new_n6788), .Y(new_n6790));
  O2A1O1Ixp33_ASAP7_75t_L   g06534(.A1(new_n6788), .A2(new_n6789), .B(new_n6790), .C(new_n6784), .Y(new_n6791));
  AOI211xp5_ASAP7_75t_L     g06535(.A1(new_n6733), .A2(new_n6481), .B(new_n6786), .C(new_n6791), .Y(new_n6792));
  A2O1A1Ixp33_ASAP7_75t_L   g06536(.A1(new_n6488), .A2(new_n6476), .B(new_n6787), .C(new_n6777), .Y(new_n6793));
  NAND3xp33_ASAP7_75t_L     g06537(.A(new_n6793), .B(new_n6790), .C(new_n6784), .Y(new_n6794));
  OAI21xp33_ASAP7_75t_L     g06538(.A1(new_n6778), .A2(new_n6773), .B(new_n6785), .Y(new_n6795));
  AOI211xp5_ASAP7_75t_L     g06539(.A1(new_n6795), .A2(new_n6794), .B(new_n6482), .C(new_n6498), .Y(new_n6796));
  OAI21xp33_ASAP7_75t_L     g06540(.A1(new_n6796), .A2(new_n6792), .B(new_n6731), .Y(new_n6797));
  NOR3xp33_ASAP7_75t_L      g06541(.A(new_n6792), .B(new_n6796), .C(new_n6731), .Y(new_n6798));
  INVx1_ASAP7_75t_L         g06542(.A(new_n6798), .Y(new_n6799));
  NAND3xp33_ASAP7_75t_L     g06543(.A(new_n6725), .B(new_n6799), .C(new_n6797), .Y(new_n6800));
  O2A1O1Ixp33_ASAP7_75t_L   g06544(.A1(new_n3493), .A2(new_n6143), .B(new_n6145), .C(new_n6501), .Y(new_n6801));
  NAND2xp33_ASAP7_75t_L     g06545(.A(new_n6216), .B(new_n6215), .Y(new_n6802));
  A2O1A1O1Ixp25_ASAP7_75t_L g06546(.A1(new_n6140), .A2(new_n6802), .B(new_n6801), .C(new_n6503), .D(new_n6499), .Y(new_n6803));
  INVx1_ASAP7_75t_L         g06547(.A(new_n6797), .Y(new_n6804));
  OAI21xp33_ASAP7_75t_L     g06548(.A1(new_n6798), .A2(new_n6804), .B(new_n6803), .Y(new_n6805));
  AOI21xp33_ASAP7_75t_L     g06549(.A1(new_n6800), .A2(new_n6805), .B(new_n6723), .Y(new_n6806));
  A2O1A1Ixp33_ASAP7_75t_L   g06550(.A1(new_n1633), .A2(new_n2932), .B(new_n6719), .C(\a[29] ), .Y(new_n6807));
  A2O1A1O1Ixp25_ASAP7_75t_L g06551(.A1(new_n2932), .A2(new_n1633), .B(new_n6719), .C(new_n6807), .D(new_n6720), .Y(new_n6808));
  NOR3xp33_ASAP7_75t_L      g06552(.A(new_n6803), .B(new_n6804), .C(new_n6798), .Y(new_n6809));
  AOI21xp33_ASAP7_75t_L     g06553(.A1(new_n6799), .A2(new_n6797), .B(new_n6725), .Y(new_n6810));
  NOR3xp33_ASAP7_75t_L      g06554(.A(new_n6809), .B(new_n6810), .C(new_n6808), .Y(new_n6811));
  NOR2xp33_ASAP7_75t_L      g06555(.A(new_n6806), .B(new_n6811), .Y(new_n6812));
  A2O1A1Ixp33_ASAP7_75t_L   g06556(.A1(new_n6717), .A2(new_n6519), .B(new_n6716), .C(new_n6812), .Y(new_n6813));
  O2A1O1Ixp33_ASAP7_75t_L   g06557(.A1(new_n6513), .A2(new_n6512), .B(new_n6519), .C(new_n6716), .Y(new_n6814));
  OAI21xp33_ASAP7_75t_L     g06558(.A1(new_n6810), .A2(new_n6809), .B(new_n6808), .Y(new_n6815));
  NAND3xp33_ASAP7_75t_L     g06559(.A(new_n6800), .B(new_n6805), .C(new_n6723), .Y(new_n6816));
  NAND2xp33_ASAP7_75t_L     g06560(.A(new_n6816), .B(new_n6815), .Y(new_n6817));
  NAND2xp33_ASAP7_75t_L     g06561(.A(new_n6814), .B(new_n6817), .Y(new_n6818));
  NOR2xp33_ASAP7_75t_L      g06562(.A(new_n1745), .B(new_n2415), .Y(new_n6819));
  AOI221xp5_ASAP7_75t_L     g06563(.A1(\b[18] ), .A2(new_n2577), .B1(\b[19] ), .B2(new_n2421), .C(new_n6819), .Y(new_n6820));
  O2A1O1Ixp33_ASAP7_75t_L   g06564(.A1(new_n2425), .A2(new_n1754), .B(new_n6820), .C(new_n2413), .Y(new_n6821));
  OAI21xp33_ASAP7_75t_L     g06565(.A1(new_n2425), .A2(new_n1754), .B(new_n6820), .Y(new_n6822));
  NAND2xp33_ASAP7_75t_L     g06566(.A(new_n2413), .B(new_n6822), .Y(new_n6823));
  OAI21xp33_ASAP7_75t_L     g06567(.A1(new_n2413), .A2(new_n6821), .B(new_n6823), .Y(new_n6824));
  INVx1_ASAP7_75t_L         g06568(.A(new_n6824), .Y(new_n6825));
  NAND3xp33_ASAP7_75t_L     g06569(.A(new_n6825), .B(new_n6813), .C(new_n6818), .Y(new_n6826));
  O2A1O1Ixp33_ASAP7_75t_L   g06570(.A1(new_n6715), .A2(new_n6517), .B(new_n6533), .C(new_n6817), .Y(new_n6827));
  MAJIxp5_ASAP7_75t_L       g06571(.A(new_n6523), .B(new_n6715), .C(new_n6517), .Y(new_n6828));
  NOR2xp33_ASAP7_75t_L      g06572(.A(new_n6828), .B(new_n6812), .Y(new_n6829));
  OAI21xp33_ASAP7_75t_L     g06573(.A1(new_n6829), .A2(new_n6827), .B(new_n6824), .Y(new_n6830));
  MAJIxp5_ASAP7_75t_L       g06574(.A(new_n6537), .B(new_n6539), .C(new_n6530), .Y(new_n6831));
  AND3x1_ASAP7_75t_L        g06575(.A(new_n6831), .B(new_n6830), .C(new_n6826), .Y(new_n6832));
  AOI21xp33_ASAP7_75t_L     g06576(.A1(new_n6830), .A2(new_n6826), .B(new_n6831), .Y(new_n6833));
  NOR2xp33_ASAP7_75t_L      g06577(.A(new_n2045), .B(new_n1962), .Y(new_n6834));
  AOI221xp5_ASAP7_75t_L     g06578(.A1(new_n1955), .A2(\b[23] ), .B1(new_n2093), .B2(\b[21] ), .C(new_n6834), .Y(new_n6835));
  O2A1O1Ixp33_ASAP7_75t_L   g06579(.A1(new_n1956), .A2(new_n2194), .B(new_n6835), .C(new_n1952), .Y(new_n6836));
  INVx1_ASAP7_75t_L         g06580(.A(new_n6836), .Y(new_n6837));
  O2A1O1Ixp33_ASAP7_75t_L   g06581(.A1(new_n1956), .A2(new_n2194), .B(new_n6835), .C(\a[23] ), .Y(new_n6838));
  AOI21xp33_ASAP7_75t_L     g06582(.A1(new_n6837), .A2(\a[23] ), .B(new_n6838), .Y(new_n6839));
  OAI21xp33_ASAP7_75t_L     g06583(.A1(new_n6833), .A2(new_n6832), .B(new_n6839), .Y(new_n6840));
  NAND2xp33_ASAP7_75t_L     g06584(.A(new_n6553), .B(new_n6552), .Y(new_n6841));
  O2A1O1Ixp33_ASAP7_75t_L   g06585(.A1(new_n6547), .A2(new_n1952), .B(new_n6549), .C(new_n6841), .Y(new_n6842));
  O2A1O1Ixp33_ASAP7_75t_L   g06586(.A1(new_n6551), .A2(new_n6550), .B(new_n6565), .C(new_n6842), .Y(new_n6843));
  NOR3xp33_ASAP7_75t_L      g06587(.A(new_n6832), .B(new_n6839), .C(new_n6833), .Y(new_n6844));
  INVx1_ASAP7_75t_L         g06588(.A(new_n6844), .Y(new_n6845));
  AOI21xp33_ASAP7_75t_L     g06589(.A1(new_n6840), .A2(new_n6845), .B(new_n6843), .Y(new_n6846));
  A2O1A1O1Ixp25_ASAP7_75t_L g06590(.A1(new_n6563), .A2(new_n6565), .B(new_n6842), .C(new_n6840), .D(new_n6844), .Y(new_n6847));
  NAND2xp33_ASAP7_75t_L     g06591(.A(\b[25] ), .B(new_n1507), .Y(new_n6848));
  OAI221xp5_ASAP7_75t_L     g06592(.A1(new_n1518), .A2(new_n2703), .B1(new_n2205), .B2(new_n1654), .C(new_n6848), .Y(new_n6849));
  A2O1A1Ixp33_ASAP7_75t_L   g06593(.A1(new_n2709), .A2(new_n1513), .B(new_n6849), .C(\a[20] ), .Y(new_n6850));
  AOI211xp5_ASAP7_75t_L     g06594(.A1(new_n2709), .A2(new_n1513), .B(new_n6849), .C(new_n1501), .Y(new_n6851));
  A2O1A1O1Ixp25_ASAP7_75t_L g06595(.A1(new_n2709), .A2(new_n1513), .B(new_n6849), .C(new_n6850), .D(new_n6851), .Y(new_n6852));
  INVx1_ASAP7_75t_L         g06596(.A(new_n6852), .Y(new_n6853));
  AOI211xp5_ASAP7_75t_L     g06597(.A1(new_n6847), .A2(new_n6840), .B(new_n6846), .C(new_n6853), .Y(new_n6854));
  NOR2xp33_ASAP7_75t_L      g06598(.A(new_n6538), .B(new_n6544), .Y(new_n6855));
  A2O1A1Ixp33_ASAP7_75t_L   g06599(.A1(\a[23] ), .A2(new_n6554), .B(new_n6548), .C(new_n6855), .Y(new_n6856));
  OA21x2_ASAP7_75t_L        g06600(.A1(new_n6833), .A2(new_n6832), .B(new_n6839), .Y(new_n6857));
  O2A1O1Ixp33_ASAP7_75t_L   g06601(.A1(new_n6557), .A2(new_n6559), .B(new_n6856), .C(new_n6857), .Y(new_n6858));
  NAND4xp25_ASAP7_75t_L     g06602(.A(new_n6845), .B(new_n6566), .C(new_n6856), .D(new_n6840), .Y(new_n6859));
  A2O1A1O1Ixp25_ASAP7_75t_L g06603(.A1(new_n6845), .A2(new_n6858), .B(new_n6843), .C(new_n6859), .D(new_n6852), .Y(new_n6860));
  NOR3xp33_ASAP7_75t_L      g06604(.A(new_n6714), .B(new_n6854), .C(new_n6860), .Y(new_n6861));
  NAND2xp33_ASAP7_75t_L     g06605(.A(new_n6566), .B(new_n6560), .Y(new_n6862));
  NOR2xp33_ASAP7_75t_L      g06606(.A(new_n6571), .B(new_n6862), .Y(new_n6863));
  NAND2xp33_ASAP7_75t_L     g06607(.A(new_n6572), .B(new_n6576), .Y(new_n6864));
  A2O1A1Ixp33_ASAP7_75t_L   g06608(.A1(new_n6279), .A2(new_n6564), .B(new_n6557), .C(new_n6856), .Y(new_n6865));
  OAI21xp33_ASAP7_75t_L     g06609(.A1(new_n6844), .A2(new_n6857), .B(new_n6865), .Y(new_n6866));
  NAND3xp33_ASAP7_75t_L     g06610(.A(new_n6866), .B(new_n6859), .C(new_n6852), .Y(new_n6867));
  A2O1A1Ixp33_ASAP7_75t_L   g06611(.A1(new_n6847), .A2(new_n6840), .B(new_n6846), .C(new_n6853), .Y(new_n6868));
  AOI221xp5_ASAP7_75t_L     g06612(.A1(new_n6582), .A2(new_n6864), .B1(new_n6867), .B2(new_n6868), .C(new_n6863), .Y(new_n6869));
  OAI21xp33_ASAP7_75t_L     g06613(.A1(new_n6869), .A2(new_n6861), .B(new_n6712), .Y(new_n6870));
  XNOR2x2_ASAP7_75t_L       g06614(.A(\a[17] ), .B(new_n6711), .Y(new_n6871));
  MAJIxp5_ASAP7_75t_L       g06615(.A(new_n6577), .B(new_n6862), .C(new_n6571), .Y(new_n6872));
  NAND3xp33_ASAP7_75t_L     g06616(.A(new_n6872), .B(new_n6867), .C(new_n6868), .Y(new_n6873));
  OAI21xp33_ASAP7_75t_L     g06617(.A1(new_n6854), .A2(new_n6860), .B(new_n6714), .Y(new_n6874));
  NAND3xp33_ASAP7_75t_L     g06618(.A(new_n6873), .B(new_n6871), .C(new_n6874), .Y(new_n6875));
  NAND3xp33_ASAP7_75t_L     g06619(.A(new_n6709), .B(new_n6870), .C(new_n6875), .Y(new_n6876));
  MAJIxp5_ASAP7_75t_L       g06620(.A(new_n6407), .B(new_n6413), .C(new_n6707), .Y(new_n6877));
  NAND2xp33_ASAP7_75t_L     g06621(.A(new_n6870), .B(new_n6875), .Y(new_n6878));
  NAND2xp33_ASAP7_75t_L     g06622(.A(new_n6877), .B(new_n6878), .Y(new_n6879));
  AOI21xp33_ASAP7_75t_L     g06623(.A1(new_n6876), .A2(new_n6879), .B(new_n6705), .Y(new_n6880));
  INVx1_ASAP7_75t_L         g06624(.A(new_n6705), .Y(new_n6881));
  NOR2xp33_ASAP7_75t_L      g06625(.A(new_n6877), .B(new_n6878), .Y(new_n6882));
  O2A1O1Ixp33_ASAP7_75t_L   g06626(.A1(new_n1206), .A2(new_n6410), .B(new_n6412), .C(new_n6706), .Y(new_n6883));
  AOI221xp5_ASAP7_75t_L     g06627(.A1(new_n6407), .A2(new_n6591), .B1(new_n6870), .B2(new_n6875), .C(new_n6883), .Y(new_n6884));
  NOR3xp33_ASAP7_75t_L      g06628(.A(new_n6882), .B(new_n6884), .C(new_n6881), .Y(new_n6885));
  NOR3xp33_ASAP7_75t_L      g06629(.A(new_n6699), .B(new_n6880), .C(new_n6885), .Y(new_n6886));
  OAI21xp33_ASAP7_75t_L     g06630(.A1(new_n6884), .A2(new_n6882), .B(new_n6881), .Y(new_n6887));
  NAND3xp33_ASAP7_75t_L     g06631(.A(new_n6876), .B(new_n6879), .C(new_n6705), .Y(new_n6888));
  AOI221xp5_ASAP7_75t_L     g06632(.A1(new_n6406), .A2(new_n6599), .B1(new_n6888), .B2(new_n6887), .C(new_n6609), .Y(new_n6889));
  NOR2xp33_ASAP7_75t_L      g06633(.A(new_n4344), .B(new_n1550), .Y(new_n6890));
  AOI221xp5_ASAP7_75t_L     g06634(.A1(\b[33] ), .A2(new_n713), .B1(\b[35] ), .B2(new_n640), .C(new_n6890), .Y(new_n6891));
  O2A1O1Ixp33_ASAP7_75t_L   g06635(.A1(new_n641), .A2(new_n4589), .B(new_n6891), .C(new_n637), .Y(new_n6892));
  INVx1_ASAP7_75t_L         g06636(.A(new_n6892), .Y(new_n6893));
  O2A1O1Ixp33_ASAP7_75t_L   g06637(.A1(new_n641), .A2(new_n4589), .B(new_n6891), .C(\a[11] ), .Y(new_n6894));
  AOI21xp33_ASAP7_75t_L     g06638(.A1(new_n6893), .A2(\a[11] ), .B(new_n6894), .Y(new_n6895));
  INVx1_ASAP7_75t_L         g06639(.A(new_n6895), .Y(new_n6896));
  NOR3xp33_ASAP7_75t_L      g06640(.A(new_n6896), .B(new_n6889), .C(new_n6886), .Y(new_n6897));
  OAI21xp33_ASAP7_75t_L     g06641(.A1(new_n6608), .A2(new_n6607), .B(new_n6605), .Y(new_n6898));
  NAND3xp33_ASAP7_75t_L     g06642(.A(new_n6898), .B(new_n6887), .C(new_n6888), .Y(new_n6899));
  OAI21xp33_ASAP7_75t_L     g06643(.A1(new_n6885), .A2(new_n6880), .B(new_n6699), .Y(new_n6900));
  AOI21xp33_ASAP7_75t_L     g06644(.A1(new_n6899), .A2(new_n6900), .B(new_n6895), .Y(new_n6901));
  NOR2xp33_ASAP7_75t_L      g06645(.A(new_n6901), .B(new_n6897), .Y(new_n6902));
  AND2x2_ASAP7_75t_L        g06646(.A(new_n6606), .B(new_n6610), .Y(new_n6903));
  MAJIxp5_ASAP7_75t_L       g06647(.A(new_n6625), .B(new_n6619), .C(new_n6903), .Y(new_n6904));
  NAND2xp33_ASAP7_75t_L     g06648(.A(new_n6904), .B(new_n6902), .Y(new_n6905));
  MAJIxp5_ASAP7_75t_L       g06649(.A(new_n6630), .B(new_n6611), .C(new_n6622), .Y(new_n6906));
  OAI21xp33_ASAP7_75t_L     g06650(.A1(new_n6897), .A2(new_n6901), .B(new_n6906), .Y(new_n6907));
  NOR2xp33_ASAP7_75t_L      g06651(.A(new_n5074), .B(new_n513), .Y(new_n6908));
  AOI221xp5_ASAP7_75t_L     g06652(.A1(\b[36] ), .A2(new_n560), .B1(\b[38] ), .B2(new_n475), .C(new_n6908), .Y(new_n6909));
  O2A1O1Ixp33_ASAP7_75t_L   g06653(.A1(new_n477), .A2(new_n5318), .B(new_n6909), .C(new_n466), .Y(new_n6910));
  INVx1_ASAP7_75t_L         g06654(.A(new_n6910), .Y(new_n6911));
  O2A1O1Ixp33_ASAP7_75t_L   g06655(.A1(new_n477), .A2(new_n5318), .B(new_n6909), .C(\a[8] ), .Y(new_n6912));
  AOI21xp33_ASAP7_75t_L     g06656(.A1(new_n6911), .A2(\a[8] ), .B(new_n6912), .Y(new_n6913));
  NAND3xp33_ASAP7_75t_L     g06657(.A(new_n6905), .B(new_n6907), .C(new_n6913), .Y(new_n6914));
  NAND3xp33_ASAP7_75t_L     g06658(.A(new_n6899), .B(new_n6900), .C(new_n6895), .Y(new_n6915));
  OAI21xp33_ASAP7_75t_L     g06659(.A1(new_n6886), .A2(new_n6889), .B(new_n6896), .Y(new_n6916));
  NAND2xp33_ASAP7_75t_L     g06660(.A(new_n6916), .B(new_n6915), .Y(new_n6917));
  NOR2xp33_ASAP7_75t_L      g06661(.A(new_n6906), .B(new_n6917), .Y(new_n6918));
  AOI21xp33_ASAP7_75t_L     g06662(.A1(new_n6916), .A2(new_n6915), .B(new_n6904), .Y(new_n6919));
  INVx1_ASAP7_75t_L         g06663(.A(new_n6912), .Y(new_n6920));
  OAI21xp33_ASAP7_75t_L     g06664(.A1(new_n466), .A2(new_n6910), .B(new_n6920), .Y(new_n6921));
  OAI21xp33_ASAP7_75t_L     g06665(.A1(new_n6919), .A2(new_n6918), .B(new_n6921), .Y(new_n6922));
  AOI22xp33_ASAP7_75t_L     g06666(.A1(new_n6914), .A2(new_n6922), .B1(new_n6645), .B2(new_n6698), .Y(new_n6923));
  A2O1A1O1Ixp25_ASAP7_75t_L g06667(.A1(new_n5829), .A2(new_n5875), .B(new_n5828), .C(new_n6092), .D(new_n6097), .Y(new_n6924));
  O2A1O1Ixp33_ASAP7_75t_L   g06668(.A1(new_n6361), .A2(new_n6924), .B(new_n6360), .C(new_n6642), .Y(new_n6925));
  NOR3xp33_ASAP7_75t_L      g06669(.A(new_n6918), .B(new_n6919), .C(new_n6921), .Y(new_n6926));
  AOI21xp33_ASAP7_75t_L     g06670(.A1(new_n6905), .A2(new_n6907), .B(new_n6913), .Y(new_n6927));
  NOR4xp25_ASAP7_75t_L      g06671(.A(new_n6925), .B(new_n6927), .C(new_n6639), .D(new_n6926), .Y(new_n6928));
  OAI21xp33_ASAP7_75t_L     g06672(.A1(new_n6923), .A2(new_n6928), .B(new_n6697), .Y(new_n6929));
  INVx1_ASAP7_75t_L         g06673(.A(new_n6697), .Y(new_n6930));
  OAI22xp33_ASAP7_75t_L     g06674(.A1(new_n6925), .A2(new_n6639), .B1(new_n6927), .B2(new_n6926), .Y(new_n6931));
  NAND3xp33_ASAP7_75t_L     g06675(.A(new_n6659), .B(new_n6914), .C(new_n6922), .Y(new_n6932));
  NAND3xp33_ASAP7_75t_L     g06676(.A(new_n6930), .B(new_n6932), .C(new_n6931), .Y(new_n6933));
  NAND2xp33_ASAP7_75t_L     g06677(.A(new_n6933), .B(new_n6929), .Y(new_n6934));
  NOR2xp33_ASAP7_75t_L      g06678(.A(new_n6666), .B(new_n6665), .Y(new_n6935));
  A2O1A1Ixp33_ASAP7_75t_L   g06679(.A1(new_n6935), .A2(new_n6405), .B(new_n6666), .C(new_n6934), .Y(new_n6936));
  A2O1A1O1Ixp25_ASAP7_75t_L g06680(.A1(new_n6641), .A2(new_n6640), .B(new_n6637), .C(new_n6659), .D(new_n6657), .Y(new_n6937));
  O2A1O1Ixp33_ASAP7_75t_L   g06681(.A1(new_n6937), .A2(new_n6655), .B(new_n6661), .C(new_n6934), .Y(new_n6938));
  NOR2xp33_ASAP7_75t_L      g06682(.A(new_n6378), .B(new_n287), .Y(new_n6939));
  AOI221xp5_ASAP7_75t_L     g06683(.A1(\b[43] ), .A2(new_n264), .B1(\b[44] ), .B2(new_n283), .C(new_n6939), .Y(new_n6940));
  INVx1_ASAP7_75t_L         g06684(.A(new_n6379), .Y(new_n6941));
  A2O1A1Ixp33_ASAP7_75t_L   g06685(.A1(new_n6113), .A2(new_n6376), .B(new_n6377), .C(new_n6941), .Y(new_n6942));
  NOR2xp33_ASAP7_75t_L      g06686(.A(\b[43] ), .B(\b[44] ), .Y(new_n6943));
  INVx1_ASAP7_75t_L         g06687(.A(\b[44] ), .Y(new_n6944));
  NOR2xp33_ASAP7_75t_L      g06688(.A(new_n6671), .B(new_n6944), .Y(new_n6945));
  NOR2xp33_ASAP7_75t_L      g06689(.A(new_n6943), .B(new_n6945), .Y(new_n6946));
  A2O1A1Ixp33_ASAP7_75t_L   g06690(.A1(new_n6942), .A2(new_n6673), .B(new_n6672), .C(new_n6946), .Y(new_n6947));
  O2A1O1Ixp33_ASAP7_75t_L   g06691(.A1(new_n6379), .A2(new_n6382), .B(new_n6673), .C(new_n6672), .Y(new_n6948));
  INVx1_ASAP7_75t_L         g06692(.A(new_n6946), .Y(new_n6949));
  NAND2xp33_ASAP7_75t_L     g06693(.A(new_n6949), .B(new_n6948), .Y(new_n6950));
  NAND2xp33_ASAP7_75t_L     g06694(.A(new_n6950), .B(new_n6947), .Y(new_n6951));
  O2A1O1Ixp33_ASAP7_75t_L   g06695(.A1(new_n279), .A2(new_n6951), .B(new_n6940), .C(new_n257), .Y(new_n6952));
  O2A1O1Ixp33_ASAP7_75t_L   g06696(.A1(new_n279), .A2(new_n6951), .B(new_n6940), .C(\a[2] ), .Y(new_n6953));
  INVx1_ASAP7_75t_L         g06697(.A(new_n6953), .Y(new_n6954));
  OAI21xp33_ASAP7_75t_L     g06698(.A1(new_n257), .A2(new_n6952), .B(new_n6954), .Y(new_n6955));
  INVx1_ASAP7_75t_L         g06699(.A(new_n6955), .Y(new_n6956));
  A2O1A1Ixp33_ASAP7_75t_L   g06700(.A1(new_n6936), .A2(new_n6934), .B(new_n6938), .C(new_n6956), .Y(new_n6957));
  AO21x2_ASAP7_75t_L        g06701(.A1(new_n6660), .A2(new_n6661), .B(new_n6934), .Y(new_n6958));
  AOI21xp33_ASAP7_75t_L     g06702(.A1(new_n6405), .A2(new_n6656), .B(new_n6666), .Y(new_n6959));
  NAND2xp33_ASAP7_75t_L     g06703(.A(new_n6934), .B(new_n6959), .Y(new_n6960));
  NAND3xp33_ASAP7_75t_L     g06704(.A(new_n6958), .B(new_n6960), .C(new_n6955), .Y(new_n6961));
  NAND2xp33_ASAP7_75t_L     g06705(.A(new_n6961), .B(new_n6957), .Y(new_n6962));
  INVx1_ASAP7_75t_L         g06706(.A(new_n6962), .Y(new_n6963));
  O2A1O1Ixp33_ASAP7_75t_L   g06707(.A1(new_n6688), .A2(new_n6690), .B(new_n6685), .C(new_n6963), .Y(new_n6964));
  OAI21xp33_ASAP7_75t_L     g06708(.A1(new_n6688), .A2(new_n6690), .B(new_n6685), .Y(new_n6965));
  NOR2xp33_ASAP7_75t_L      g06709(.A(new_n6962), .B(new_n6965), .Y(new_n6966));
  NOR2xp33_ASAP7_75t_L      g06710(.A(new_n6966), .B(new_n6964), .Y(\f[44] ));
  INVx1_ASAP7_75t_L         g06711(.A(new_n6957), .Y(new_n6968));
  INVx1_ASAP7_75t_L         g06712(.A(new_n6961), .Y(new_n6969));
  INVx1_ASAP7_75t_L         g06713(.A(new_n6936), .Y(new_n6970));
  O2A1O1Ixp33_ASAP7_75t_L   g06714(.A1(new_n6959), .A2(new_n6970), .B(new_n6960), .C(new_n6956), .Y(new_n6971));
  O2A1O1Ixp33_ASAP7_75t_L   g06715(.A1(new_n6968), .A2(new_n6969), .B(new_n6965), .C(new_n6971), .Y(new_n6972));
  NOR2xp33_ASAP7_75t_L      g06716(.A(new_n6919), .B(new_n6918), .Y(new_n6973));
  A2O1A1Ixp33_ASAP7_75t_L   g06717(.A1(\a[8] ), .A2(new_n6911), .B(new_n6912), .C(new_n6973), .Y(new_n6974));
  NOR2xp33_ASAP7_75t_L      g06718(.A(new_n6886), .B(new_n6889), .Y(new_n6975));
  A2O1A1Ixp33_ASAP7_75t_L   g06719(.A1(\a[11] ), .A2(new_n6893), .B(new_n6894), .C(new_n6975), .Y(new_n6976));
  OAI21xp33_ASAP7_75t_L     g06720(.A1(new_n6880), .A2(new_n6699), .B(new_n6888), .Y(new_n6977));
  NOR3xp33_ASAP7_75t_L      g06721(.A(new_n6712), .B(new_n6861), .C(new_n6869), .Y(new_n6978));
  NAND2xp33_ASAP7_75t_L     g06722(.A(new_n6575), .B(new_n6713), .Y(new_n6979));
  A2O1A1Ixp33_ASAP7_75t_L   g06723(.A1(new_n6586), .A2(new_n6979), .B(new_n6854), .C(new_n6868), .Y(new_n6980));
  INVx1_ASAP7_75t_L         g06724(.A(new_n6716), .Y(new_n6981));
  A2O1A1Ixp33_ASAP7_75t_L   g06725(.A1(new_n6533), .A2(new_n6981), .B(new_n6806), .C(new_n6816), .Y(new_n6982));
  A2O1A1O1Ixp25_ASAP7_75t_L g06726(.A1(new_n6503), .A2(new_n6502), .B(new_n6499), .C(new_n6797), .D(new_n6798), .Y(new_n6983));
  A2O1A1Ixp33_ASAP7_75t_L   g06727(.A1(new_n6733), .A2(new_n6481), .B(new_n6786), .C(new_n6795), .Y(new_n6984));
  NOR2xp33_ASAP7_75t_L      g06728(.A(new_n833), .B(new_n4147), .Y(new_n6985));
  AOI221xp5_ASAP7_75t_L     g06729(.A1(\b[10] ), .A2(new_n4402), .B1(\b[11] ), .B2(new_n4155), .C(new_n6985), .Y(new_n6986));
  O2A1O1Ixp33_ASAP7_75t_L   g06730(.A1(new_n4150), .A2(new_n841), .B(new_n6986), .C(new_n4145), .Y(new_n6987));
  OAI21xp33_ASAP7_75t_L     g06731(.A1(new_n4150), .A2(new_n841), .B(new_n6986), .Y(new_n6988));
  NAND2xp33_ASAP7_75t_L     g06732(.A(new_n4145), .B(new_n6988), .Y(new_n6989));
  OAI21xp33_ASAP7_75t_L     g06733(.A1(new_n4145), .A2(new_n6987), .B(new_n6989), .Y(new_n6990));
  NOR2xp33_ASAP7_75t_L      g06734(.A(new_n6764), .B(new_n6762), .Y(new_n6991));
  A2O1A1Ixp33_ASAP7_75t_L   g06735(.A1(new_n6766), .A2(\a[38] ), .B(new_n6737), .C(new_n6991), .Y(new_n6992));
  NAND2xp33_ASAP7_75t_L     g06736(.A(new_n6753), .B(new_n6750), .Y(new_n6993));
  O2A1O1Ixp33_ASAP7_75t_L   g06737(.A1(new_n5630), .A2(new_n728), .B(new_n6755), .C(new_n5626), .Y(new_n6994));
  O2A1O1Ixp33_ASAP7_75t_L   g06738(.A1(new_n6994), .A2(new_n5626), .B(new_n6758), .C(new_n6993), .Y(new_n6995));
  INVx1_ASAP7_75t_L         g06739(.A(new_n6995), .Y(new_n6996));
  INVx1_ASAP7_75t_L         g06740(.A(\a[45] ), .Y(new_n6997));
  NAND2xp33_ASAP7_75t_L     g06741(.A(\a[44] ), .B(new_n6997), .Y(new_n6998));
  NAND2xp33_ASAP7_75t_L     g06742(.A(\a[45] ), .B(new_n6439), .Y(new_n6999));
  AND2x2_ASAP7_75t_L        g06743(.A(new_n6998), .B(new_n6999), .Y(new_n7000));
  NOR2xp33_ASAP7_75t_L      g06744(.A(new_n284), .B(new_n7000), .Y(new_n7001));
  A2O1A1Ixp33_ASAP7_75t_L   g06745(.A1(new_n6749), .A2(new_n6747), .B(new_n6446), .C(new_n7001), .Y(new_n7002));
  NAND2xp33_ASAP7_75t_L     g06746(.A(new_n6451), .B(new_n6449), .Y(new_n7003));
  NOR5xp2_ASAP7_75t_L       g06747(.A(new_n7003), .B(new_n6748), .C(new_n6745), .D(new_n6153), .E(new_n6439), .Y(new_n7004));
  A2O1A1Ixp33_ASAP7_75t_L   g06748(.A1(new_n6998), .A2(new_n6999), .B(new_n284), .C(new_n7004), .Y(new_n7005));
  NAND2xp33_ASAP7_75t_L     g06749(.A(\b[3] ), .B(new_n6442), .Y(new_n7006));
  NAND2xp33_ASAP7_75t_L     g06750(.A(\b[1] ), .B(new_n6742), .Y(new_n7007));
  NAND2xp33_ASAP7_75t_L     g06751(.A(\b[2] ), .B(new_n6436), .Y(new_n7008));
  NAND2xp33_ASAP7_75t_L     g06752(.A(new_n6450), .B(new_n312), .Y(new_n7009));
  NAND5xp2_ASAP7_75t_L      g06753(.A(new_n7009), .B(new_n7008), .C(new_n7007), .D(new_n7006), .E(\a[44] ), .Y(new_n7010));
  OAI211xp5_ASAP7_75t_L     g06754(.A1(new_n6741), .A2(new_n262), .B(new_n7006), .C(new_n7008), .Y(new_n7011));
  A2O1A1Ixp33_ASAP7_75t_L   g06755(.A1(new_n312), .A2(new_n6450), .B(new_n7011), .C(new_n6439), .Y(new_n7012));
  AND2x2_ASAP7_75t_L        g06756(.A(new_n7010), .B(new_n7012), .Y(new_n7013));
  AO21x2_ASAP7_75t_L        g06757(.A1(new_n7002), .A2(new_n7005), .B(new_n7013), .Y(new_n7014));
  NAND3xp33_ASAP7_75t_L     g06758(.A(new_n7005), .B(new_n7002), .C(new_n7013), .Y(new_n7015));
  NAND2xp33_ASAP7_75t_L     g06759(.A(\b[5] ), .B(new_n5623), .Y(new_n7016));
  OAI221xp5_ASAP7_75t_L     g06760(.A1(new_n5641), .A2(new_n427), .B1(new_n332), .B2(new_n5925), .C(new_n7016), .Y(new_n7017));
  A2O1A1Ixp33_ASAP7_75t_L   g06761(.A1(new_n5363), .A2(new_n5637), .B(new_n7017), .C(\a[41] ), .Y(new_n7018));
  NAND2xp33_ASAP7_75t_L     g06762(.A(\a[41] ), .B(new_n7018), .Y(new_n7019));
  A2O1A1Ixp33_ASAP7_75t_L   g06763(.A1(new_n5363), .A2(new_n5637), .B(new_n7017), .C(new_n5626), .Y(new_n7020));
  NAND4xp25_ASAP7_75t_L     g06764(.A(new_n7014), .B(new_n7020), .C(new_n7019), .D(new_n7015), .Y(new_n7021));
  AOI21xp33_ASAP7_75t_L     g06765(.A1(new_n7005), .A2(new_n7002), .B(new_n7013), .Y(new_n7022));
  AND3x1_ASAP7_75t_L        g06766(.A(new_n7005), .B(new_n7013), .C(new_n7002), .Y(new_n7023));
  NAND2xp33_ASAP7_75t_L     g06767(.A(new_n7020), .B(new_n7019), .Y(new_n7024));
  OAI21xp33_ASAP7_75t_L     g06768(.A1(new_n7022), .A2(new_n7023), .B(new_n7024), .Y(new_n7025));
  AND4x1_ASAP7_75t_L        g06769(.A(new_n6768), .B(new_n6996), .C(new_n7025), .D(new_n7021), .Y(new_n7026));
  O2A1O1Ixp33_ASAP7_75t_L   g06770(.A1(new_n6759), .A2(new_n6760), .B(new_n6763), .C(new_n6995), .Y(new_n7027));
  AOI21xp33_ASAP7_75t_L     g06771(.A1(new_n7025), .A2(new_n7021), .B(new_n7027), .Y(new_n7028));
  NOR2xp33_ASAP7_75t_L      g06772(.A(new_n590), .B(new_n4908), .Y(new_n7029));
  AOI221xp5_ASAP7_75t_L     g06773(.A1(\b[7] ), .A2(new_n5139), .B1(\b[8] ), .B2(new_n4916), .C(new_n7029), .Y(new_n7030));
  OAI21xp33_ASAP7_75t_L     g06774(.A1(new_n4911), .A2(new_n1066), .B(new_n7030), .Y(new_n7031));
  NOR2xp33_ASAP7_75t_L      g06775(.A(new_n4906), .B(new_n7031), .Y(new_n7032));
  O2A1O1Ixp33_ASAP7_75t_L   g06776(.A1(new_n4911), .A2(new_n1066), .B(new_n7030), .C(\a[38] ), .Y(new_n7033));
  NOR2xp33_ASAP7_75t_L      g06777(.A(new_n7033), .B(new_n7032), .Y(new_n7034));
  OAI21xp33_ASAP7_75t_L     g06778(.A1(new_n7028), .A2(new_n7026), .B(new_n7034), .Y(new_n7035));
  NAND3xp33_ASAP7_75t_L     g06779(.A(new_n7027), .B(new_n7025), .C(new_n7021), .Y(new_n7036));
  AO22x1_ASAP7_75t_L        g06780(.A1(new_n7025), .A2(new_n7021), .B1(new_n6996), .B2(new_n6768), .Y(new_n7037));
  O2A1O1Ixp33_ASAP7_75t_L   g06781(.A1(new_n4911), .A2(new_n1066), .B(new_n7030), .C(new_n4906), .Y(new_n7038));
  INVx1_ASAP7_75t_L         g06782(.A(new_n7033), .Y(new_n7039));
  OAI21xp33_ASAP7_75t_L     g06783(.A1(new_n4906), .A2(new_n7038), .B(new_n7039), .Y(new_n7040));
  NAND3xp33_ASAP7_75t_L     g06784(.A(new_n7037), .B(new_n7040), .C(new_n7036), .Y(new_n7041));
  NAND2xp33_ASAP7_75t_L     g06785(.A(new_n7035), .B(new_n7041), .Y(new_n7042));
  O2A1O1Ixp33_ASAP7_75t_L   g06786(.A1(new_n6788), .A2(new_n6777), .B(new_n6992), .C(new_n7042), .Y(new_n7043));
  NAND2xp33_ASAP7_75t_L     g06787(.A(new_n6768), .B(new_n6770), .Y(new_n7044));
  O2A1O1Ixp33_ASAP7_75t_L   g06788(.A1(new_n4906), .A2(new_n6736), .B(new_n6738), .C(new_n7044), .Y(new_n7045));
  AOI221xp5_ASAP7_75t_L     g06789(.A1(new_n7041), .A2(new_n7035), .B1(new_n6772), .B2(new_n6774), .C(new_n7045), .Y(new_n7046));
  OAI21xp33_ASAP7_75t_L     g06790(.A1(new_n7046), .A2(new_n7043), .B(new_n6990), .Y(new_n7047));
  OA21x2_ASAP7_75t_L        g06791(.A1(new_n4145), .A2(new_n6987), .B(new_n6989), .Y(new_n7048));
  OAI21xp33_ASAP7_75t_L     g06792(.A1(new_n6777), .A2(new_n6788), .B(new_n6992), .Y(new_n7049));
  AOI21xp33_ASAP7_75t_L     g06793(.A1(new_n7037), .A2(new_n7036), .B(new_n7040), .Y(new_n7050));
  NOR3xp33_ASAP7_75t_L      g06794(.A(new_n7026), .B(new_n7034), .C(new_n7028), .Y(new_n7051));
  NOR2xp33_ASAP7_75t_L      g06795(.A(new_n7051), .B(new_n7050), .Y(new_n7052));
  NAND2xp33_ASAP7_75t_L     g06796(.A(new_n7052), .B(new_n7049), .Y(new_n7053));
  OAI221xp5_ASAP7_75t_L     g06797(.A1(new_n6788), .A2(new_n6777), .B1(new_n7050), .B2(new_n7051), .C(new_n6992), .Y(new_n7054));
  NAND3xp33_ASAP7_75t_L     g06798(.A(new_n7053), .B(new_n7048), .C(new_n7054), .Y(new_n7055));
  NAND3xp33_ASAP7_75t_L     g06799(.A(new_n6984), .B(new_n7047), .C(new_n7055), .Y(new_n7056));
  A2O1A1O1Ixp25_ASAP7_75t_L g06800(.A1(new_n6492), .A2(new_n6416), .B(new_n6482), .C(new_n6794), .D(new_n6791), .Y(new_n7057));
  NAND2xp33_ASAP7_75t_L     g06801(.A(new_n7055), .B(new_n7047), .Y(new_n7058));
  NAND2xp33_ASAP7_75t_L     g06802(.A(new_n7057), .B(new_n7058), .Y(new_n7059));
  NOR2xp33_ASAP7_75t_L      g06803(.A(new_n960), .B(new_n3509), .Y(new_n7060));
  AOI221xp5_ASAP7_75t_L     g06804(.A1(\b[13] ), .A2(new_n3708), .B1(\b[15] ), .B2(new_n3503), .C(new_n7060), .Y(new_n7061));
  INVx1_ASAP7_75t_L         g06805(.A(new_n7061), .Y(new_n7062));
  A2O1A1Ixp33_ASAP7_75t_L   g06806(.A1(new_n1052), .A2(new_n3505), .B(new_n7062), .C(\a[32] ), .Y(new_n7063));
  O2A1O1Ixp33_ASAP7_75t_L   g06807(.A1(new_n3513), .A2(new_n1774), .B(new_n7061), .C(\a[32] ), .Y(new_n7064));
  AO21x2_ASAP7_75t_L        g06808(.A1(\a[32] ), .A2(new_n7063), .B(new_n7064), .Y(new_n7065));
  AOI21xp33_ASAP7_75t_L     g06809(.A1(new_n7059), .A2(new_n7056), .B(new_n7065), .Y(new_n7066));
  AOI21xp33_ASAP7_75t_L     g06810(.A1(new_n7053), .A2(new_n7054), .B(new_n7048), .Y(new_n7067));
  NOR3xp33_ASAP7_75t_L      g06811(.A(new_n7043), .B(new_n7046), .C(new_n6990), .Y(new_n7068));
  OAI21xp33_ASAP7_75t_L     g06812(.A1(new_n7067), .A2(new_n7068), .B(new_n6984), .Y(new_n7069));
  AOI21xp33_ASAP7_75t_L     g06813(.A1(new_n7055), .A2(new_n7047), .B(new_n6984), .Y(new_n7070));
  AOI21xp33_ASAP7_75t_L     g06814(.A1(new_n7063), .A2(\a[32] ), .B(new_n7064), .Y(new_n7071));
  AOI211xp5_ASAP7_75t_L     g06815(.A1(new_n7069), .A2(new_n6984), .B(new_n7070), .C(new_n7071), .Y(new_n7072));
  OR3x1_ASAP7_75t_L         g06816(.A(new_n6983), .B(new_n7066), .C(new_n7072), .Y(new_n7073));
  A2O1A1Ixp33_ASAP7_75t_L   g06817(.A1(new_n7069), .A2(new_n6984), .B(new_n7070), .C(new_n7065), .Y(new_n7074));
  A2O1A1Ixp33_ASAP7_75t_L   g06818(.A1(new_n7065), .A2(new_n7074), .B(new_n7066), .C(new_n6983), .Y(new_n7075));
  NOR2xp33_ASAP7_75t_L      g06819(.A(new_n1349), .B(new_n2925), .Y(new_n7076));
  AOI221xp5_ASAP7_75t_L     g06820(.A1(\b[16] ), .A2(new_n3129), .B1(\b[18] ), .B2(new_n2938), .C(new_n7076), .Y(new_n7077));
  O2A1O1Ixp33_ASAP7_75t_L   g06821(.A1(new_n2940), .A2(new_n1464), .B(new_n7077), .C(new_n2928), .Y(new_n7078));
  INVx1_ASAP7_75t_L         g06822(.A(new_n7077), .Y(new_n7079));
  A2O1A1Ixp33_ASAP7_75t_L   g06823(.A1(new_n2329), .A2(new_n2932), .B(new_n7079), .C(new_n2928), .Y(new_n7080));
  OA21x2_ASAP7_75t_L        g06824(.A1(new_n2928), .A2(new_n7078), .B(new_n7080), .Y(new_n7081));
  AOI21xp33_ASAP7_75t_L     g06825(.A1(new_n7073), .A2(new_n7075), .B(new_n7081), .Y(new_n7082));
  NOR3xp33_ASAP7_75t_L      g06826(.A(new_n6983), .B(new_n7066), .C(new_n7072), .Y(new_n7083));
  A2O1A1Ixp33_ASAP7_75t_L   g06827(.A1(new_n7069), .A2(new_n6984), .B(new_n7070), .C(new_n7071), .Y(new_n7084));
  NAND3xp33_ASAP7_75t_L     g06828(.A(new_n7059), .B(new_n7056), .C(new_n7065), .Y(new_n7085));
  AOI221xp5_ASAP7_75t_L     g06829(.A1(new_n6725), .A2(new_n6797), .B1(new_n7084), .B2(new_n7085), .C(new_n6798), .Y(new_n7086));
  OAI21xp33_ASAP7_75t_L     g06830(.A1(new_n2928), .A2(new_n7078), .B(new_n7080), .Y(new_n7087));
  NOR3xp33_ASAP7_75t_L      g06831(.A(new_n7086), .B(new_n7083), .C(new_n7087), .Y(new_n7088));
  NOR2xp33_ASAP7_75t_L      g06832(.A(new_n7088), .B(new_n7082), .Y(new_n7089));
  NAND2xp33_ASAP7_75t_L     g06833(.A(new_n6982), .B(new_n7089), .Y(new_n7090));
  A2O1A1O1Ixp25_ASAP7_75t_L g06834(.A1(new_n6519), .A2(new_n6717), .B(new_n6716), .C(new_n6815), .D(new_n6811), .Y(new_n7091));
  OAI21xp33_ASAP7_75t_L     g06835(.A1(new_n7082), .A2(new_n7088), .B(new_n7091), .Y(new_n7092));
  NOR2xp33_ASAP7_75t_L      g06836(.A(new_n1745), .B(new_n2410), .Y(new_n7093));
  AOI221xp5_ASAP7_75t_L     g06837(.A1(\b[19] ), .A2(new_n2577), .B1(\b[21] ), .B2(new_n2423), .C(new_n7093), .Y(new_n7094));
  O2A1O1Ixp33_ASAP7_75t_L   g06838(.A1(new_n2425), .A2(new_n1901), .B(new_n7094), .C(new_n2413), .Y(new_n7095));
  INVx1_ASAP7_75t_L         g06839(.A(new_n7095), .Y(new_n7096));
  O2A1O1Ixp33_ASAP7_75t_L   g06840(.A1(new_n2425), .A2(new_n1901), .B(new_n7094), .C(\a[26] ), .Y(new_n7097));
  AOI21xp33_ASAP7_75t_L     g06841(.A1(new_n7096), .A2(\a[26] ), .B(new_n7097), .Y(new_n7098));
  NAND3xp33_ASAP7_75t_L     g06842(.A(new_n7090), .B(new_n7092), .C(new_n7098), .Y(new_n7099));
  NOR3xp33_ASAP7_75t_L      g06843(.A(new_n7091), .B(new_n7082), .C(new_n7088), .Y(new_n7100));
  OAI21xp33_ASAP7_75t_L     g06844(.A1(new_n7083), .A2(new_n7086), .B(new_n7087), .Y(new_n7101));
  NAND3xp33_ASAP7_75t_L     g06845(.A(new_n7073), .B(new_n7075), .C(new_n7081), .Y(new_n7102));
  AOI221xp5_ASAP7_75t_L     g06846(.A1(new_n6828), .A2(new_n6815), .B1(new_n7101), .B2(new_n7102), .C(new_n6811), .Y(new_n7103));
  INVx1_ASAP7_75t_L         g06847(.A(new_n7097), .Y(new_n7104));
  OAI21xp33_ASAP7_75t_L     g06848(.A1(new_n2413), .A2(new_n7095), .B(new_n7104), .Y(new_n7105));
  OAI21xp33_ASAP7_75t_L     g06849(.A1(new_n7103), .A2(new_n7100), .B(new_n7105), .Y(new_n7106));
  NAND2xp33_ASAP7_75t_L     g06850(.A(new_n7106), .B(new_n7099), .Y(new_n7107));
  XNOR2x2_ASAP7_75t_L       g06851(.A(new_n6814), .B(new_n6817), .Y(new_n7108));
  MAJIxp5_ASAP7_75t_L       g06852(.A(new_n6831), .B(new_n7108), .C(new_n6825), .Y(new_n7109));
  NOR2xp33_ASAP7_75t_L      g06853(.A(new_n7109), .B(new_n7107), .Y(new_n7110));
  NAND2xp33_ASAP7_75t_L     g06854(.A(new_n7092), .B(new_n7090), .Y(new_n7111));
  O2A1O1Ixp33_ASAP7_75t_L   g06855(.A1(new_n7095), .A2(new_n2413), .B(new_n7104), .C(new_n7111), .Y(new_n7112));
  NOR2xp33_ASAP7_75t_L      g06856(.A(new_n6829), .B(new_n6827), .Y(new_n7113));
  MAJIxp5_ASAP7_75t_L       g06857(.A(new_n6543), .B(new_n6541), .C(new_n6535), .Y(new_n7114));
  MAJIxp5_ASAP7_75t_L       g06858(.A(new_n7114), .B(new_n7113), .C(new_n6824), .Y(new_n7115));
  O2A1O1Ixp33_ASAP7_75t_L   g06859(.A1(new_n7111), .A2(new_n7112), .B(new_n7106), .C(new_n7115), .Y(new_n7116));
  OAI22xp33_ASAP7_75t_L     g06860(.A1(new_n2089), .A2(new_n2045), .B1(new_n2188), .B2(new_n1962), .Y(new_n7117));
  AOI221xp5_ASAP7_75t_L     g06861(.A1(new_n1955), .A2(\b[24] ), .B1(new_n1964), .B2(new_n2216), .C(new_n7117), .Y(new_n7118));
  XNOR2x2_ASAP7_75t_L       g06862(.A(new_n1952), .B(new_n7118), .Y(new_n7119));
  OAI21xp33_ASAP7_75t_L     g06863(.A1(new_n7110), .A2(new_n7116), .B(new_n7119), .Y(new_n7120));
  NOR3xp33_ASAP7_75t_L      g06864(.A(new_n7100), .B(new_n7105), .C(new_n7103), .Y(new_n7121));
  AOI21xp33_ASAP7_75t_L     g06865(.A1(new_n7090), .A2(new_n7092), .B(new_n7098), .Y(new_n7122));
  NOR2xp33_ASAP7_75t_L      g06866(.A(new_n7121), .B(new_n7122), .Y(new_n7123));
  NAND2xp33_ASAP7_75t_L     g06867(.A(new_n7123), .B(new_n7115), .Y(new_n7124));
  OAI21xp33_ASAP7_75t_L     g06868(.A1(new_n7121), .A2(new_n7122), .B(new_n7109), .Y(new_n7125));
  XNOR2x2_ASAP7_75t_L       g06869(.A(\a[23] ), .B(new_n7118), .Y(new_n7126));
  NAND3xp33_ASAP7_75t_L     g06870(.A(new_n7124), .B(new_n7126), .C(new_n7125), .Y(new_n7127));
  OAI211xp5_ASAP7_75t_L     g06871(.A1(new_n6844), .A2(new_n6858), .B(new_n7120), .C(new_n7127), .Y(new_n7128));
  AOI21xp33_ASAP7_75t_L     g06872(.A1(new_n7124), .A2(new_n7125), .B(new_n7126), .Y(new_n7129));
  NOR3xp33_ASAP7_75t_L      g06873(.A(new_n7116), .B(new_n7119), .C(new_n7110), .Y(new_n7130));
  OAI21xp33_ASAP7_75t_L     g06874(.A1(new_n7129), .A2(new_n7130), .B(new_n6847), .Y(new_n7131));
  NOR2xp33_ASAP7_75t_L      g06875(.A(new_n2703), .B(new_n1517), .Y(new_n7132));
  AOI221xp5_ASAP7_75t_L     g06876(.A1(\b[25] ), .A2(new_n1659), .B1(\b[27] ), .B2(new_n1511), .C(new_n7132), .Y(new_n7133));
  O2A1O1Ixp33_ASAP7_75t_L   g06877(.A1(new_n1521), .A2(new_n2889), .B(new_n7133), .C(new_n1501), .Y(new_n7134));
  INVx1_ASAP7_75t_L         g06878(.A(new_n7134), .Y(new_n7135));
  O2A1O1Ixp33_ASAP7_75t_L   g06879(.A1(new_n1521), .A2(new_n2889), .B(new_n7133), .C(\a[20] ), .Y(new_n7136));
  AOI21xp33_ASAP7_75t_L     g06880(.A1(new_n7135), .A2(\a[20] ), .B(new_n7136), .Y(new_n7137));
  NAND3xp33_ASAP7_75t_L     g06881(.A(new_n7128), .B(new_n7131), .C(new_n7137), .Y(new_n7138));
  NOR3xp33_ASAP7_75t_L      g06882(.A(new_n6847), .B(new_n7130), .C(new_n7129), .Y(new_n7139));
  AOI211xp5_ASAP7_75t_L     g06883(.A1(new_n7120), .A2(new_n7127), .B(new_n6858), .C(new_n6844), .Y(new_n7140));
  AO21x2_ASAP7_75t_L        g06884(.A1(\a[20] ), .A2(new_n7135), .B(new_n7136), .Y(new_n7141));
  OAI21xp33_ASAP7_75t_L     g06885(.A1(new_n7139), .A2(new_n7140), .B(new_n7141), .Y(new_n7142));
  NAND3xp33_ASAP7_75t_L     g06886(.A(new_n6980), .B(new_n7138), .C(new_n7142), .Y(new_n7143));
  A2O1A1O1Ixp25_ASAP7_75t_L g06887(.A1(new_n6582), .A2(new_n6864), .B(new_n6863), .C(new_n6867), .D(new_n6860), .Y(new_n7144));
  INVx1_ASAP7_75t_L         g06888(.A(new_n7138), .Y(new_n7145));
  AOI21xp33_ASAP7_75t_L     g06889(.A1(new_n7128), .A2(new_n7131), .B(new_n7137), .Y(new_n7146));
  OAI21xp33_ASAP7_75t_L     g06890(.A1(new_n7146), .A2(new_n7145), .B(new_n7144), .Y(new_n7147));
  NOR2xp33_ASAP7_75t_L      g06891(.A(new_n3098), .B(new_n2118), .Y(new_n7148));
  AOI221xp5_ASAP7_75t_L     g06892(.A1(\b[28] ), .A2(new_n1290), .B1(\b[30] ), .B2(new_n1209), .C(new_n7148), .Y(new_n7149));
  O2A1O1Ixp33_ASAP7_75t_L   g06893(.A1(new_n1210), .A2(new_n3464), .B(new_n7149), .C(new_n1206), .Y(new_n7150));
  INVx1_ASAP7_75t_L         g06894(.A(new_n7150), .Y(new_n7151));
  O2A1O1Ixp33_ASAP7_75t_L   g06895(.A1(new_n1210), .A2(new_n3464), .B(new_n7149), .C(\a[17] ), .Y(new_n7152));
  AOI21xp33_ASAP7_75t_L     g06896(.A1(new_n7151), .A2(\a[17] ), .B(new_n7152), .Y(new_n7153));
  AOI21xp33_ASAP7_75t_L     g06897(.A1(new_n7147), .A2(new_n7143), .B(new_n7153), .Y(new_n7154));
  NOR3xp33_ASAP7_75t_L      g06898(.A(new_n7144), .B(new_n7145), .C(new_n7146), .Y(new_n7155));
  AOI21xp33_ASAP7_75t_L     g06899(.A1(new_n7142), .A2(new_n7138), .B(new_n6980), .Y(new_n7156));
  AO21x2_ASAP7_75t_L        g06900(.A1(\a[17] ), .A2(new_n7151), .B(new_n7152), .Y(new_n7157));
  NOR3xp33_ASAP7_75t_L      g06901(.A(new_n7155), .B(new_n7156), .C(new_n7157), .Y(new_n7158));
  NOR2xp33_ASAP7_75t_L      g06902(.A(new_n7154), .B(new_n7158), .Y(new_n7159));
  A2O1A1Ixp33_ASAP7_75t_L   g06903(.A1(new_n6870), .A2(new_n6709), .B(new_n6978), .C(new_n7159), .Y(new_n7160));
  A2O1A1O1Ixp25_ASAP7_75t_L g06904(.A1(new_n6407), .A2(new_n6591), .B(new_n6883), .C(new_n6870), .D(new_n6978), .Y(new_n7161));
  OAI21xp33_ASAP7_75t_L     g06905(.A1(new_n7156), .A2(new_n7155), .B(new_n7157), .Y(new_n7162));
  NAND3xp33_ASAP7_75t_L     g06906(.A(new_n7147), .B(new_n7143), .C(new_n7153), .Y(new_n7163));
  NAND2xp33_ASAP7_75t_L     g06907(.A(new_n7163), .B(new_n7162), .Y(new_n7164));
  NAND2xp33_ASAP7_75t_L     g06908(.A(new_n7161), .B(new_n7164), .Y(new_n7165));
  NOR2xp33_ASAP7_75t_L      g06909(.A(new_n3891), .B(new_n864), .Y(new_n7166));
  AOI221xp5_ASAP7_75t_L     g06910(.A1(\b[31] ), .A2(new_n985), .B1(\b[33] ), .B2(new_n886), .C(new_n7166), .Y(new_n7167));
  O2A1O1Ixp33_ASAP7_75t_L   g06911(.A1(new_n872), .A2(new_n4108), .B(new_n7167), .C(new_n867), .Y(new_n7168));
  INVx1_ASAP7_75t_L         g06912(.A(new_n7168), .Y(new_n7169));
  O2A1O1Ixp33_ASAP7_75t_L   g06913(.A1(new_n872), .A2(new_n4108), .B(new_n7167), .C(\a[14] ), .Y(new_n7170));
  AOI21xp33_ASAP7_75t_L     g06914(.A1(new_n7169), .A2(\a[14] ), .B(new_n7170), .Y(new_n7171));
  NAND3xp33_ASAP7_75t_L     g06915(.A(new_n7160), .B(new_n7165), .C(new_n7171), .Y(new_n7172));
  NOR2xp33_ASAP7_75t_L      g06916(.A(new_n7161), .B(new_n7164), .Y(new_n7173));
  AOI221xp5_ASAP7_75t_L     g06917(.A1(new_n6709), .A2(new_n6870), .B1(new_n7162), .B2(new_n7163), .C(new_n6978), .Y(new_n7174));
  INVx1_ASAP7_75t_L         g06918(.A(new_n7171), .Y(new_n7175));
  OAI21xp33_ASAP7_75t_L     g06919(.A1(new_n7174), .A2(new_n7173), .B(new_n7175), .Y(new_n7176));
  NAND3xp33_ASAP7_75t_L     g06920(.A(new_n6977), .B(new_n7172), .C(new_n7176), .Y(new_n7177));
  A2O1A1O1Ixp25_ASAP7_75t_L g06921(.A1(new_n6599), .A2(new_n6406), .B(new_n6609), .C(new_n6887), .D(new_n6885), .Y(new_n7178));
  NOR3xp33_ASAP7_75t_L      g06922(.A(new_n7175), .B(new_n7173), .C(new_n7174), .Y(new_n7179));
  AOI21xp33_ASAP7_75t_L     g06923(.A1(new_n7160), .A2(new_n7165), .B(new_n7171), .Y(new_n7180));
  OAI21xp33_ASAP7_75t_L     g06924(.A1(new_n7179), .A2(new_n7180), .B(new_n7178), .Y(new_n7181));
  NOR2xp33_ASAP7_75t_L      g06925(.A(new_n4581), .B(new_n1550), .Y(new_n7182));
  AOI221xp5_ASAP7_75t_L     g06926(.A1(\b[34] ), .A2(new_n713), .B1(\b[36] ), .B2(new_n640), .C(new_n7182), .Y(new_n7183));
  INVx1_ASAP7_75t_L         g06927(.A(new_n7183), .Y(new_n7184));
  A2O1A1Ixp33_ASAP7_75t_L   g06928(.A1(new_n4621), .A2(new_n718), .B(new_n7184), .C(\a[11] ), .Y(new_n7185));
  A2O1A1Ixp33_ASAP7_75t_L   g06929(.A1(new_n4621), .A2(new_n718), .B(new_n7184), .C(new_n637), .Y(new_n7186));
  INVx1_ASAP7_75t_L         g06930(.A(new_n7186), .Y(new_n7187));
  AOI21xp33_ASAP7_75t_L     g06931(.A1(new_n7185), .A2(\a[11] ), .B(new_n7187), .Y(new_n7188));
  AOI21xp33_ASAP7_75t_L     g06932(.A1(new_n7177), .A2(new_n7181), .B(new_n7188), .Y(new_n7189));
  NOR3xp33_ASAP7_75t_L      g06933(.A(new_n7178), .B(new_n7179), .C(new_n7180), .Y(new_n7190));
  AOI21xp33_ASAP7_75t_L     g06934(.A1(new_n7176), .A2(new_n7172), .B(new_n6977), .Y(new_n7191));
  AO21x2_ASAP7_75t_L        g06935(.A1(\a[11] ), .A2(new_n7185), .B(new_n7187), .Y(new_n7192));
  NOR3xp33_ASAP7_75t_L      g06936(.A(new_n7190), .B(new_n7191), .C(new_n7192), .Y(new_n7193));
  OAI221xp5_ASAP7_75t_L     g06937(.A1(new_n7193), .A2(new_n7189), .B1(new_n6902), .B2(new_n6904), .C(new_n6976), .Y(new_n7194));
  NAND2xp33_ASAP7_75t_L     g06938(.A(new_n6900), .B(new_n6899), .Y(new_n7195));
  INVx1_ASAP7_75t_L         g06939(.A(new_n6894), .Y(new_n7196));
  O2A1O1Ixp33_ASAP7_75t_L   g06940(.A1(new_n6892), .A2(new_n637), .B(new_n7196), .C(new_n7195), .Y(new_n7197));
  NOR2xp33_ASAP7_75t_L      g06941(.A(new_n7189), .B(new_n7193), .Y(new_n7198));
  OAI21xp33_ASAP7_75t_L     g06942(.A1(new_n7197), .A2(new_n6919), .B(new_n7198), .Y(new_n7199));
  NOR2xp33_ASAP7_75t_L      g06943(.A(new_n5311), .B(new_n513), .Y(new_n7200));
  AOI221xp5_ASAP7_75t_L     g06944(.A1(\b[37] ), .A2(new_n560), .B1(\b[39] ), .B2(new_n475), .C(new_n7200), .Y(new_n7201));
  O2A1O1Ixp33_ASAP7_75t_L   g06945(.A1(new_n477), .A2(new_n5578), .B(new_n7201), .C(new_n466), .Y(new_n7202));
  INVx1_ASAP7_75t_L         g06946(.A(new_n7202), .Y(new_n7203));
  O2A1O1Ixp33_ASAP7_75t_L   g06947(.A1(new_n477), .A2(new_n5578), .B(new_n7201), .C(\a[8] ), .Y(new_n7204));
  AOI21xp33_ASAP7_75t_L     g06948(.A1(new_n7203), .A2(\a[8] ), .B(new_n7204), .Y(new_n7205));
  NAND3xp33_ASAP7_75t_L     g06949(.A(new_n7199), .B(new_n7194), .C(new_n7205), .Y(new_n7206));
  OAI21xp33_ASAP7_75t_L     g06950(.A1(new_n7191), .A2(new_n7190), .B(new_n7192), .Y(new_n7207));
  NAND3xp33_ASAP7_75t_L     g06951(.A(new_n7177), .B(new_n7181), .C(new_n7188), .Y(new_n7208));
  AOI221xp5_ASAP7_75t_L     g06952(.A1(new_n7207), .A2(new_n7208), .B1(new_n6906), .B2(new_n6917), .C(new_n7197), .Y(new_n7209));
  NAND2xp33_ASAP7_75t_L     g06953(.A(new_n7208), .B(new_n7207), .Y(new_n7210));
  AOI21xp33_ASAP7_75t_L     g06954(.A1(new_n6907), .A2(new_n6976), .B(new_n7210), .Y(new_n7211));
  INVx1_ASAP7_75t_L         g06955(.A(new_n7204), .Y(new_n7212));
  OAI21xp33_ASAP7_75t_L     g06956(.A1(new_n466), .A2(new_n7202), .B(new_n7212), .Y(new_n7213));
  OAI21xp33_ASAP7_75t_L     g06957(.A1(new_n7209), .A2(new_n7211), .B(new_n7213), .Y(new_n7214));
  NAND4xp25_ASAP7_75t_L     g06958(.A(new_n6931), .B(new_n7206), .C(new_n7214), .D(new_n6974), .Y(new_n7215));
  NAND2xp33_ASAP7_75t_L     g06959(.A(new_n7206), .B(new_n7214), .Y(new_n7216));
  NAND2xp33_ASAP7_75t_L     g06960(.A(new_n6907), .B(new_n6905), .Y(new_n7217));
  MAJIxp5_ASAP7_75t_L       g06961(.A(new_n6659), .B(new_n6913), .C(new_n7217), .Y(new_n7218));
  NAND2xp33_ASAP7_75t_L     g06962(.A(new_n7218), .B(new_n7216), .Y(new_n7219));
  NOR2xp33_ASAP7_75t_L      g06963(.A(new_n5855), .B(new_n375), .Y(new_n7220));
  AOI221xp5_ASAP7_75t_L     g06964(.A1(\b[42] ), .A2(new_n361), .B1(new_n349), .B2(\b[41] ), .C(new_n7220), .Y(new_n7221));
  O2A1O1Ixp33_ASAP7_75t_L   g06965(.A1(new_n356), .A2(new_n6386), .B(new_n7221), .C(new_n346), .Y(new_n7222));
  O2A1O1Ixp33_ASAP7_75t_L   g06966(.A1(new_n356), .A2(new_n6386), .B(new_n7221), .C(\a[5] ), .Y(new_n7223));
  INVx1_ASAP7_75t_L         g06967(.A(new_n7223), .Y(new_n7224));
  OA21x2_ASAP7_75t_L        g06968(.A1(new_n346), .A2(new_n7222), .B(new_n7224), .Y(new_n7225));
  NAND3xp33_ASAP7_75t_L     g06969(.A(new_n7219), .B(new_n7215), .C(new_n7225), .Y(new_n7226));
  O2A1O1Ixp33_ASAP7_75t_L   g06970(.A1(new_n6910), .A2(new_n466), .B(new_n6920), .C(new_n7217), .Y(new_n7227));
  NOR3xp33_ASAP7_75t_L      g06971(.A(new_n7211), .B(new_n7213), .C(new_n7209), .Y(new_n7228));
  AOI21xp33_ASAP7_75t_L     g06972(.A1(new_n7199), .A2(new_n7194), .B(new_n7205), .Y(new_n7229));
  NOR4xp25_ASAP7_75t_L      g06973(.A(new_n6923), .B(new_n7229), .C(new_n7227), .D(new_n7228), .Y(new_n7230));
  AOI22xp33_ASAP7_75t_L     g06974(.A1(new_n7206), .A2(new_n7214), .B1(new_n6974), .B2(new_n6931), .Y(new_n7231));
  OAI21xp33_ASAP7_75t_L     g06975(.A1(new_n346), .A2(new_n7222), .B(new_n7224), .Y(new_n7232));
  OAI21xp33_ASAP7_75t_L     g06976(.A1(new_n7230), .A2(new_n7231), .B(new_n7232), .Y(new_n7233));
  NAND2xp33_ASAP7_75t_L     g06977(.A(new_n7233), .B(new_n7226), .Y(new_n7234));
  NAND2xp33_ASAP7_75t_L     g06978(.A(new_n6931), .B(new_n6932), .Y(new_n7235));
  MAJIxp5_ASAP7_75t_L       g06979(.A(new_n6959), .B(new_n6930), .C(new_n7235), .Y(new_n7236));
  NOR2xp33_ASAP7_75t_L      g06980(.A(new_n7234), .B(new_n7236), .Y(new_n7237));
  NAND3xp33_ASAP7_75t_L     g06981(.A(new_n7219), .B(new_n7215), .C(new_n7232), .Y(new_n7238));
  INVx1_ASAP7_75t_L         g06982(.A(new_n7238), .Y(new_n7239));
  O2A1O1Ixp33_ASAP7_75t_L   g06983(.A1(new_n346), .A2(new_n6694), .B(new_n6696), .C(new_n7235), .Y(new_n7240));
  A2O1A1O1Ixp25_ASAP7_75t_L g06984(.A1(new_n6405), .A2(new_n6935), .B(new_n6666), .C(new_n6934), .D(new_n7240), .Y(new_n7241));
  O2A1O1Ixp33_ASAP7_75t_L   g06985(.A1(new_n7225), .A2(new_n7239), .B(new_n7226), .C(new_n7241), .Y(new_n7242));
  NOR2xp33_ASAP7_75t_L      g06986(.A(new_n6671), .B(new_n287), .Y(new_n7243));
  AOI221xp5_ASAP7_75t_L     g06987(.A1(\b[44] ), .A2(new_n264), .B1(\b[45] ), .B2(new_n283), .C(new_n7243), .Y(new_n7244));
  INVx1_ASAP7_75t_L         g06988(.A(new_n7244), .Y(new_n7245));
  INVx1_ASAP7_75t_L         g06989(.A(new_n6672), .Y(new_n7246));
  A2O1A1O1Ixp25_ASAP7_75t_L g06990(.A1(new_n6941), .A2(new_n6383), .B(new_n6670), .C(new_n7246), .D(new_n6949), .Y(new_n7247));
  NOR2xp33_ASAP7_75t_L      g06991(.A(\b[44] ), .B(\b[45] ), .Y(new_n7248));
  INVx1_ASAP7_75t_L         g06992(.A(\b[45] ), .Y(new_n7249));
  NOR2xp33_ASAP7_75t_L      g06993(.A(new_n6944), .B(new_n7249), .Y(new_n7250));
  NOR2xp33_ASAP7_75t_L      g06994(.A(new_n7248), .B(new_n7250), .Y(new_n7251));
  A2O1A1Ixp33_ASAP7_75t_L   g06995(.A1(\b[44] ), .A2(\b[43] ), .B(new_n7247), .C(new_n7251), .Y(new_n7252));
  INVx1_ASAP7_75t_L         g06996(.A(new_n6945), .Y(new_n7253));
  OAI211xp5_ASAP7_75t_L     g06997(.A1(new_n7248), .A2(new_n7250), .B(new_n6947), .C(new_n7253), .Y(new_n7254));
  NAND2xp33_ASAP7_75t_L     g06998(.A(new_n7252), .B(new_n7254), .Y(new_n7255));
  INVx1_ASAP7_75t_L         g06999(.A(new_n7255), .Y(new_n7256));
  A2O1A1Ixp33_ASAP7_75t_L   g07000(.A1(new_n7256), .A2(new_n273), .B(new_n7245), .C(\a[2] ), .Y(new_n7257));
  O2A1O1Ixp33_ASAP7_75t_L   g07001(.A1(new_n279), .A2(new_n7255), .B(new_n7244), .C(new_n257), .Y(new_n7258));
  NOR2xp33_ASAP7_75t_L      g07002(.A(new_n257), .B(new_n7258), .Y(new_n7259));
  A2O1A1O1Ixp25_ASAP7_75t_L g07003(.A1(new_n273), .A2(new_n7256), .B(new_n7245), .C(new_n7257), .D(new_n7259), .Y(new_n7260));
  OAI21xp33_ASAP7_75t_L     g07004(.A1(new_n7237), .A2(new_n7242), .B(new_n7260), .Y(new_n7261));
  NOR3xp33_ASAP7_75t_L      g07005(.A(new_n7242), .B(new_n7237), .C(new_n7260), .Y(new_n7262));
  INVx1_ASAP7_75t_L         g07006(.A(new_n7262), .Y(new_n7263));
  NAND2xp33_ASAP7_75t_L     g07007(.A(new_n7261), .B(new_n7263), .Y(new_n7264));
  XOR2x2_ASAP7_75t_L        g07008(.A(new_n6972), .B(new_n7264), .Y(\f[45] ));
  NOR2xp33_ASAP7_75t_L      g07009(.A(new_n6944), .B(new_n287), .Y(new_n7266));
  AOI221xp5_ASAP7_75t_L     g07010(.A1(\b[45] ), .A2(new_n264), .B1(\b[46] ), .B2(new_n283), .C(new_n7266), .Y(new_n7267));
  A2O1A1Ixp33_ASAP7_75t_L   g07011(.A1(new_n6674), .A2(new_n7246), .B(new_n6949), .C(new_n7253), .Y(new_n7268));
  NOR2xp33_ASAP7_75t_L      g07012(.A(\b[45] ), .B(\b[46] ), .Y(new_n7269));
  INVx1_ASAP7_75t_L         g07013(.A(\b[46] ), .Y(new_n7270));
  NOR2xp33_ASAP7_75t_L      g07014(.A(new_n7249), .B(new_n7270), .Y(new_n7271));
  NOR2xp33_ASAP7_75t_L      g07015(.A(new_n7269), .B(new_n7271), .Y(new_n7272));
  A2O1A1Ixp33_ASAP7_75t_L   g07016(.A1(new_n7268), .A2(new_n7251), .B(new_n7250), .C(new_n7272), .Y(new_n7273));
  INVx1_ASAP7_75t_L         g07017(.A(new_n7273), .Y(new_n7274));
  INVx1_ASAP7_75t_L         g07018(.A(new_n7250), .Y(new_n7275));
  A2O1A1Ixp33_ASAP7_75t_L   g07019(.A1(new_n6947), .A2(new_n7253), .B(new_n7248), .C(new_n7275), .Y(new_n7276));
  NOR2xp33_ASAP7_75t_L      g07020(.A(new_n7272), .B(new_n7276), .Y(new_n7277));
  NOR2xp33_ASAP7_75t_L      g07021(.A(new_n7274), .B(new_n7277), .Y(new_n7278));
  INVx1_ASAP7_75t_L         g07022(.A(new_n7278), .Y(new_n7279));
  O2A1O1Ixp33_ASAP7_75t_L   g07023(.A1(new_n279), .A2(new_n7279), .B(new_n7267), .C(new_n257), .Y(new_n7280));
  INVx1_ASAP7_75t_L         g07024(.A(new_n7280), .Y(new_n7281));
  O2A1O1Ixp33_ASAP7_75t_L   g07025(.A1(new_n279), .A2(new_n7279), .B(new_n7267), .C(\a[2] ), .Y(new_n7282));
  OAI21xp33_ASAP7_75t_L     g07026(.A1(new_n7158), .A2(new_n7161), .B(new_n7162), .Y(new_n7283));
  NAND2xp33_ASAP7_75t_L     g07027(.A(new_n7131), .B(new_n7128), .Y(new_n7284));
  MAJIxp5_ASAP7_75t_L       g07028(.A(new_n7144), .B(new_n7284), .C(new_n7137), .Y(new_n7285));
  NOR2xp33_ASAP7_75t_L      g07029(.A(new_n2879), .B(new_n1517), .Y(new_n7286));
  AOI221xp5_ASAP7_75t_L     g07030(.A1(\b[26] ), .A2(new_n1659), .B1(\b[28] ), .B2(new_n1511), .C(new_n7286), .Y(new_n7287));
  INVx1_ASAP7_75t_L         g07031(.A(new_n7287), .Y(new_n7288));
  A2O1A1Ixp33_ASAP7_75t_L   g07032(.A1(new_n3085), .A2(new_n1513), .B(new_n7288), .C(\a[20] ), .Y(new_n7289));
  O2A1O1Ixp33_ASAP7_75t_L   g07033(.A1(new_n1521), .A2(new_n3087), .B(new_n7287), .C(\a[20] ), .Y(new_n7290));
  AOI21xp33_ASAP7_75t_L     g07034(.A1(new_n7289), .A2(\a[20] ), .B(new_n7290), .Y(new_n7291));
  INVx1_ASAP7_75t_L         g07035(.A(new_n7291), .Y(new_n7292));
  NOR2xp33_ASAP7_75t_L      g07036(.A(new_n1895), .B(new_n2410), .Y(new_n7293));
  AOI221xp5_ASAP7_75t_L     g07037(.A1(\b[20] ), .A2(new_n2577), .B1(\b[22] ), .B2(new_n2423), .C(new_n7293), .Y(new_n7294));
  O2A1O1Ixp33_ASAP7_75t_L   g07038(.A1(new_n2425), .A2(new_n2522), .B(new_n7294), .C(new_n2413), .Y(new_n7295));
  O2A1O1Ixp33_ASAP7_75t_L   g07039(.A1(new_n2425), .A2(new_n2522), .B(new_n7294), .C(\a[26] ), .Y(new_n7296));
  INVx1_ASAP7_75t_L         g07040(.A(new_n7296), .Y(new_n7297));
  OAI21xp33_ASAP7_75t_L     g07041(.A1(new_n2413), .A2(new_n7295), .B(new_n7297), .Y(new_n7298));
  NAND2xp33_ASAP7_75t_L     g07042(.A(new_n7054), .B(new_n7053), .Y(new_n7299));
  MAJIxp5_ASAP7_75t_L       g07043(.A(new_n7057), .B(new_n7048), .C(new_n7299), .Y(new_n7300));
  A2O1A1O1Ixp25_ASAP7_75t_L g07044(.A1(new_n6772), .A2(new_n6774), .B(new_n7045), .C(new_n7035), .D(new_n7051), .Y(new_n7301));
  INVx1_ASAP7_75t_L         g07045(.A(new_n7001), .Y(new_n7302));
  MAJIxp5_ASAP7_75t_L       g07046(.A(new_n7013), .B(new_n6753), .C(new_n7302), .Y(new_n7303));
  OR2x4_ASAP7_75t_L         g07047(.A(new_n6435), .B(new_n6434), .Y(new_n7304));
  NAND2xp33_ASAP7_75t_L     g07048(.A(\b[4] ), .B(new_n6442), .Y(new_n7305));
  OAI221xp5_ASAP7_75t_L     g07049(.A1(new_n7304), .A2(new_n301), .B1(new_n289), .B2(new_n6741), .C(new_n7305), .Y(new_n7306));
  A2O1A1Ixp33_ASAP7_75t_L   g07050(.A1(new_n342), .A2(new_n6450), .B(new_n7306), .C(\a[44] ), .Y(new_n7307));
  AOI211xp5_ASAP7_75t_L     g07051(.A1(new_n342), .A2(new_n6450), .B(new_n6439), .C(new_n7306), .Y(new_n7308));
  A2O1A1O1Ixp25_ASAP7_75t_L g07052(.A1(new_n6450), .A2(new_n342), .B(new_n7306), .C(new_n7307), .D(new_n7308), .Y(new_n7309));
  XNOR2x2_ASAP7_75t_L       g07053(.A(\a[46] ), .B(\a[45] ), .Y(new_n7310));
  INVx1_ASAP7_75t_L         g07054(.A(new_n7310), .Y(new_n7311));
  NAND2xp33_ASAP7_75t_L     g07055(.A(new_n7311), .B(new_n7000), .Y(new_n7312));
  NAND2xp33_ASAP7_75t_L     g07056(.A(new_n6999), .B(new_n6998), .Y(new_n7313));
  INVx1_ASAP7_75t_L         g07057(.A(\a[46] ), .Y(new_n7314));
  NAND2xp33_ASAP7_75t_L     g07058(.A(\a[47] ), .B(new_n7314), .Y(new_n7315));
  INVx1_ASAP7_75t_L         g07059(.A(\a[47] ), .Y(new_n7316));
  NAND2xp33_ASAP7_75t_L     g07060(.A(\a[46] ), .B(new_n7316), .Y(new_n7317));
  NAND3xp33_ASAP7_75t_L     g07061(.A(new_n7313), .B(new_n7315), .C(new_n7317), .Y(new_n7318));
  OAI22xp33_ASAP7_75t_L     g07062(.A1(new_n7312), .A2(new_n284), .B1(new_n262), .B2(new_n7318), .Y(new_n7319));
  NAND2xp33_ASAP7_75t_L     g07063(.A(new_n7317), .B(new_n7315), .Y(new_n7320));
  NAND2xp33_ASAP7_75t_L     g07064(.A(new_n7320), .B(new_n7313), .Y(new_n7321));
  INVx1_ASAP7_75t_L         g07065(.A(new_n7321), .Y(new_n7322));
  AOI21xp33_ASAP7_75t_L     g07066(.A1(new_n275), .A2(new_n7322), .B(new_n7319), .Y(new_n7323));
  NAND3xp33_ASAP7_75t_L     g07067(.A(new_n7323), .B(new_n7302), .C(\a[47] ), .Y(new_n7324));
  INVx1_ASAP7_75t_L         g07068(.A(new_n7324), .Y(new_n7325));
  A2O1A1Ixp33_ASAP7_75t_L   g07069(.A1(new_n7322), .A2(new_n275), .B(new_n7319), .C(\a[47] ), .Y(new_n7326));
  A2O1A1Ixp33_ASAP7_75t_L   g07070(.A1(new_n7322), .A2(new_n275), .B(new_n7319), .C(new_n7316), .Y(new_n7327));
  INVx1_ASAP7_75t_L         g07071(.A(new_n7327), .Y(new_n7328));
  O2A1O1Ixp33_ASAP7_75t_L   g07072(.A1(new_n7302), .A2(new_n7326), .B(\a[47] ), .C(new_n7328), .Y(new_n7329));
  OAI21xp33_ASAP7_75t_L     g07073(.A1(new_n7325), .A2(new_n7329), .B(new_n7309), .Y(new_n7330));
  A2O1A1Ixp33_ASAP7_75t_L   g07074(.A1(new_n342), .A2(new_n6450), .B(new_n7306), .C(new_n6439), .Y(new_n7331));
  INVx1_ASAP7_75t_L         g07075(.A(new_n7331), .Y(new_n7332));
  NOR2xp33_ASAP7_75t_L      g07076(.A(new_n7310), .B(new_n7313), .Y(new_n7333));
  NOR2xp33_ASAP7_75t_L      g07077(.A(new_n7320), .B(new_n7000), .Y(new_n7334));
  AOI22xp33_ASAP7_75t_L     g07078(.A1(new_n7333), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n7334), .Y(new_n7335));
  O2A1O1Ixp33_ASAP7_75t_L   g07079(.A1(new_n7321), .A2(new_n274), .B(new_n7335), .C(new_n7316), .Y(new_n7336));
  A2O1A1Ixp33_ASAP7_75t_L   g07080(.A1(new_n7336), .A2(new_n7001), .B(new_n7316), .C(new_n7327), .Y(new_n7337));
  OAI211xp5_ASAP7_75t_L     g07081(.A1(new_n7308), .A2(new_n7332), .B(new_n7337), .C(new_n7324), .Y(new_n7338));
  NAND3xp33_ASAP7_75t_L     g07082(.A(new_n7303), .B(new_n7330), .C(new_n7338), .Y(new_n7339));
  NAND2xp33_ASAP7_75t_L     g07083(.A(new_n7010), .B(new_n7012), .Y(new_n7340));
  MAJIxp5_ASAP7_75t_L       g07084(.A(new_n7340), .B(new_n7001), .C(new_n7004), .Y(new_n7341));
  AOI211xp5_ASAP7_75t_L     g07085(.A1(new_n7337), .A2(new_n7324), .B(new_n7308), .C(new_n7332), .Y(new_n7342));
  INVx1_ASAP7_75t_L         g07086(.A(new_n7306), .Y(new_n7343));
  OAI211xp5_ASAP7_75t_L     g07087(.A1(new_n1497), .A2(new_n6443), .B(new_n7343), .C(\a[44] ), .Y(new_n7344));
  AOI211xp5_ASAP7_75t_L     g07088(.A1(new_n7344), .A2(new_n7331), .B(new_n7325), .C(new_n7329), .Y(new_n7345));
  OAI21xp33_ASAP7_75t_L     g07089(.A1(new_n7342), .A2(new_n7345), .B(new_n7341), .Y(new_n7346));
  NOR2xp33_ASAP7_75t_L      g07090(.A(new_n427), .B(new_n5640), .Y(new_n7347));
  AOI221xp5_ASAP7_75t_L     g07091(.A1(\b[5] ), .A2(new_n5920), .B1(\b[7] ), .B2(new_n5629), .C(new_n7347), .Y(new_n7348));
  OAI211xp5_ASAP7_75t_L     g07092(.A1(new_n5630), .A2(new_n456), .B(\a[41] ), .C(new_n7348), .Y(new_n7349));
  INVx1_ASAP7_75t_L         g07093(.A(new_n7348), .Y(new_n7350));
  A2O1A1Ixp33_ASAP7_75t_L   g07094(.A1(new_n1188), .A2(new_n5637), .B(new_n7350), .C(new_n5626), .Y(new_n7351));
  NAND4xp25_ASAP7_75t_L     g07095(.A(new_n7339), .B(new_n7351), .C(new_n7346), .D(new_n7349), .Y(new_n7352));
  NOR3xp33_ASAP7_75t_L      g07096(.A(new_n7345), .B(new_n7341), .C(new_n7342), .Y(new_n7353));
  AOI21xp33_ASAP7_75t_L     g07097(.A1(new_n7338), .A2(new_n7330), .B(new_n7303), .Y(new_n7354));
  NAND2xp33_ASAP7_75t_L     g07098(.A(new_n7349), .B(new_n7351), .Y(new_n7355));
  OAI21xp33_ASAP7_75t_L     g07099(.A1(new_n7353), .A2(new_n7354), .B(new_n7355), .Y(new_n7356));
  NAND2xp33_ASAP7_75t_L     g07100(.A(new_n7356), .B(new_n7352), .Y(new_n7357));
  NAND3xp33_ASAP7_75t_L     g07101(.A(new_n7014), .B(new_n7024), .C(new_n7015), .Y(new_n7358));
  A2O1A1Ixp33_ASAP7_75t_L   g07102(.A1(new_n7021), .A2(new_n7025), .B(new_n7027), .C(new_n7358), .Y(new_n7359));
  NOR2xp33_ASAP7_75t_L      g07103(.A(new_n7357), .B(new_n7359), .Y(new_n7360));
  AOI22xp33_ASAP7_75t_L     g07104(.A1(new_n7352), .A2(new_n7356), .B1(new_n7358), .B2(new_n7037), .Y(new_n7361));
  OAI22xp33_ASAP7_75t_L     g07105(.A1(new_n5144), .A2(new_n534), .B1(new_n590), .B2(new_n4903), .Y(new_n7362));
  AOI221xp5_ASAP7_75t_L     g07106(.A1(new_n4917), .A2(\b[10] ), .B1(new_n4912), .B2(new_n690), .C(new_n7362), .Y(new_n7363));
  XNOR2x2_ASAP7_75t_L       g07107(.A(new_n4906), .B(new_n7363), .Y(new_n7364));
  OR3x1_ASAP7_75t_L         g07108(.A(new_n7361), .B(new_n7360), .C(new_n7364), .Y(new_n7365));
  OAI21xp33_ASAP7_75t_L     g07109(.A1(new_n7360), .A2(new_n7361), .B(new_n7364), .Y(new_n7366));
  AO21x2_ASAP7_75t_L        g07110(.A1(new_n7366), .A2(new_n7365), .B(new_n7301), .Y(new_n7367));
  NAND3xp33_ASAP7_75t_L     g07111(.A(new_n7301), .B(new_n7365), .C(new_n7366), .Y(new_n7368));
  NAND2xp33_ASAP7_75t_L     g07112(.A(\b[12] ), .B(new_n4155), .Y(new_n7369));
  OAI221xp5_ASAP7_75t_L     g07113(.A1(new_n4147), .A2(new_n936), .B1(new_n748), .B2(new_n4397), .C(new_n7369), .Y(new_n7370));
  A2O1A1Ixp33_ASAP7_75t_L   g07114(.A1(new_n1166), .A2(new_n4151), .B(new_n7370), .C(\a[35] ), .Y(new_n7371));
  AOI211xp5_ASAP7_75t_L     g07115(.A1(new_n1166), .A2(new_n4151), .B(new_n7370), .C(new_n4145), .Y(new_n7372));
  A2O1A1O1Ixp25_ASAP7_75t_L g07116(.A1(new_n4151), .A2(new_n1166), .B(new_n7370), .C(new_n7371), .D(new_n7372), .Y(new_n7373));
  NAND3xp33_ASAP7_75t_L     g07117(.A(new_n7367), .B(new_n7368), .C(new_n7373), .Y(new_n7374));
  AOI21xp33_ASAP7_75t_L     g07118(.A1(new_n7365), .A2(new_n7366), .B(new_n7301), .Y(new_n7375));
  NOR3xp33_ASAP7_75t_L      g07119(.A(new_n7361), .B(new_n7364), .C(new_n7360), .Y(new_n7376));
  A2O1A1O1Ixp25_ASAP7_75t_L g07120(.A1(new_n7035), .A2(new_n7049), .B(new_n7051), .C(new_n7366), .D(new_n7376), .Y(new_n7377));
  INVx1_ASAP7_75t_L         g07121(.A(new_n7372), .Y(new_n7378));
  A2O1A1Ixp33_ASAP7_75t_L   g07122(.A1(new_n1166), .A2(new_n4151), .B(new_n7370), .C(new_n4145), .Y(new_n7379));
  NAND2xp33_ASAP7_75t_L     g07123(.A(new_n7379), .B(new_n7378), .Y(new_n7380));
  A2O1A1Ixp33_ASAP7_75t_L   g07124(.A1(new_n7377), .A2(new_n7366), .B(new_n7375), .C(new_n7380), .Y(new_n7381));
  NAND3xp33_ASAP7_75t_L     g07125(.A(new_n7300), .B(new_n7374), .C(new_n7381), .Y(new_n7382));
  NOR2xp33_ASAP7_75t_L      g07126(.A(new_n7046), .B(new_n7043), .Y(new_n7383));
  MAJIxp5_ASAP7_75t_L       g07127(.A(new_n6984), .B(new_n6990), .C(new_n7383), .Y(new_n7384));
  NAND2xp33_ASAP7_75t_L     g07128(.A(new_n7381), .B(new_n7374), .Y(new_n7385));
  NAND2xp33_ASAP7_75t_L     g07129(.A(new_n7384), .B(new_n7385), .Y(new_n7386));
  NAND2xp33_ASAP7_75t_L     g07130(.A(\b[15] ), .B(new_n3499), .Y(new_n7387));
  OAI221xp5_ASAP7_75t_L     g07131(.A1(new_n3510), .A2(new_n1150), .B1(new_n960), .B2(new_n3703), .C(new_n7387), .Y(new_n7388));
  A2O1A1Ixp33_ASAP7_75t_L   g07132(.A1(new_n1156), .A2(new_n3505), .B(new_n7388), .C(\a[32] ), .Y(new_n7389));
  AOI211xp5_ASAP7_75t_L     g07133(.A1(new_n1156), .A2(new_n3505), .B(new_n7388), .C(new_n3493), .Y(new_n7390));
  A2O1A1O1Ixp25_ASAP7_75t_L g07134(.A1(new_n3505), .A2(new_n1156), .B(new_n7388), .C(new_n7389), .D(new_n7390), .Y(new_n7391));
  NAND3xp33_ASAP7_75t_L     g07135(.A(new_n7382), .B(new_n7386), .C(new_n7391), .Y(new_n7392));
  NOR2xp33_ASAP7_75t_L      g07136(.A(new_n7384), .B(new_n7385), .Y(new_n7393));
  AOI21xp33_ASAP7_75t_L     g07137(.A1(new_n7381), .A2(new_n7374), .B(new_n7300), .Y(new_n7394));
  INVx1_ASAP7_75t_L         g07138(.A(new_n7390), .Y(new_n7395));
  A2O1A1Ixp33_ASAP7_75t_L   g07139(.A1(new_n1156), .A2(new_n3505), .B(new_n7388), .C(new_n3493), .Y(new_n7396));
  NAND2xp33_ASAP7_75t_L     g07140(.A(new_n7396), .B(new_n7395), .Y(new_n7397));
  OAI21xp33_ASAP7_75t_L     g07141(.A1(new_n7394), .A2(new_n7393), .B(new_n7397), .Y(new_n7398));
  AO21x2_ASAP7_75t_L        g07142(.A1(new_n7085), .A2(new_n7084), .B(new_n6983), .Y(new_n7399));
  NAND4xp25_ASAP7_75t_L     g07143(.A(new_n7399), .B(new_n7398), .C(new_n7074), .D(new_n7392), .Y(new_n7400));
  NOR3xp33_ASAP7_75t_L      g07144(.A(new_n7393), .B(new_n7394), .C(new_n7397), .Y(new_n7401));
  AOI21xp33_ASAP7_75t_L     g07145(.A1(new_n7382), .A2(new_n7386), .B(new_n7391), .Y(new_n7402));
  A2O1A1Ixp33_ASAP7_75t_L   g07146(.A1(new_n7084), .A2(new_n7071), .B(new_n6983), .C(new_n7074), .Y(new_n7403));
  OAI21xp33_ASAP7_75t_L     g07147(.A1(new_n7402), .A2(new_n7401), .B(new_n7403), .Y(new_n7404));
  NOR2xp33_ASAP7_75t_L      g07148(.A(new_n1458), .B(new_n2925), .Y(new_n7405));
  AOI221xp5_ASAP7_75t_L     g07149(.A1(\b[17] ), .A2(new_n3129), .B1(\b[19] ), .B2(new_n2938), .C(new_n7405), .Y(new_n7406));
  INVx1_ASAP7_75t_L         g07150(.A(new_n7406), .Y(new_n7407));
  A2O1A1Ixp33_ASAP7_75t_L   g07151(.A1(new_n1607), .A2(new_n2932), .B(new_n7407), .C(\a[29] ), .Y(new_n7408));
  O2A1O1Ixp33_ASAP7_75t_L   g07152(.A1(new_n2940), .A2(new_n1628), .B(new_n7406), .C(\a[29] ), .Y(new_n7409));
  AOI21xp33_ASAP7_75t_L     g07153(.A1(new_n7408), .A2(\a[29] ), .B(new_n7409), .Y(new_n7410));
  NAND3xp33_ASAP7_75t_L     g07154(.A(new_n7400), .B(new_n7404), .C(new_n7410), .Y(new_n7411));
  NOR3xp33_ASAP7_75t_L      g07155(.A(new_n7403), .B(new_n7402), .C(new_n7401), .Y(new_n7412));
  AOI22xp33_ASAP7_75t_L     g07156(.A1(new_n7398), .A2(new_n7392), .B1(new_n7074), .B2(new_n7399), .Y(new_n7413));
  INVx1_ASAP7_75t_L         g07157(.A(new_n7410), .Y(new_n7414));
  OAI21xp33_ASAP7_75t_L     g07158(.A1(new_n7412), .A2(new_n7413), .B(new_n7414), .Y(new_n7415));
  A2O1A1O1Ixp25_ASAP7_75t_L g07159(.A1(new_n6815), .A2(new_n6828), .B(new_n6811), .C(new_n7102), .D(new_n7082), .Y(new_n7416));
  NAND3xp33_ASAP7_75t_L     g07160(.A(new_n7416), .B(new_n7415), .C(new_n7411), .Y(new_n7417));
  AO21x2_ASAP7_75t_L        g07161(.A1(new_n7411), .A2(new_n7415), .B(new_n7416), .Y(new_n7418));
  NAND3xp33_ASAP7_75t_L     g07162(.A(new_n7418), .B(new_n7298), .C(new_n7417), .Y(new_n7419));
  AND3x1_ASAP7_75t_L        g07163(.A(new_n7416), .B(new_n7415), .C(new_n7411), .Y(new_n7420));
  AOI21xp33_ASAP7_75t_L     g07164(.A1(new_n7415), .A2(new_n7411), .B(new_n7416), .Y(new_n7421));
  NOR3xp33_ASAP7_75t_L      g07165(.A(new_n7420), .B(new_n7421), .C(new_n7298), .Y(new_n7422));
  AOI21xp33_ASAP7_75t_L     g07166(.A1(new_n7419), .A2(new_n7298), .B(new_n7422), .Y(new_n7423));
  AOI21xp33_ASAP7_75t_L     g07167(.A1(new_n7107), .A2(new_n7109), .B(new_n7112), .Y(new_n7424));
  NAND2xp33_ASAP7_75t_L     g07168(.A(new_n7423), .B(new_n7424), .Y(new_n7425));
  INVx1_ASAP7_75t_L         g07169(.A(new_n7294), .Y(new_n7426));
  A2O1A1Ixp33_ASAP7_75t_L   g07170(.A1(new_n2056), .A2(new_n2417), .B(new_n7426), .C(\a[26] ), .Y(new_n7427));
  AOI21xp33_ASAP7_75t_L     g07171(.A1(new_n7427), .A2(\a[26] ), .B(new_n7296), .Y(new_n7428));
  NAND3xp33_ASAP7_75t_L     g07172(.A(new_n7418), .B(new_n7417), .C(new_n7428), .Y(new_n7429));
  OAI21xp33_ASAP7_75t_L     g07173(.A1(new_n7421), .A2(new_n7420), .B(new_n7298), .Y(new_n7430));
  NAND2xp33_ASAP7_75t_L     g07174(.A(new_n7429), .B(new_n7430), .Y(new_n7431));
  A2O1A1Ixp33_ASAP7_75t_L   g07175(.A1(new_n7107), .A2(new_n7109), .B(new_n7112), .C(new_n7431), .Y(new_n7432));
  NAND2xp33_ASAP7_75t_L     g07176(.A(\b[25] ), .B(new_n1955), .Y(new_n7433));
  OAI221xp5_ASAP7_75t_L     g07177(.A1(new_n1962), .A2(new_n2205), .B1(new_n2188), .B2(new_n2089), .C(new_n7433), .Y(new_n7434));
  A2O1A1Ixp33_ASAP7_75t_L   g07178(.A1(new_n5001), .A2(new_n1964), .B(new_n7434), .C(\a[23] ), .Y(new_n7435));
  AOI211xp5_ASAP7_75t_L     g07179(.A1(new_n5001), .A2(new_n1964), .B(new_n7434), .C(new_n1952), .Y(new_n7436));
  A2O1A1O1Ixp25_ASAP7_75t_L g07180(.A1(new_n5001), .A2(new_n1964), .B(new_n7434), .C(new_n7435), .D(new_n7436), .Y(new_n7437));
  NAND3xp33_ASAP7_75t_L     g07181(.A(new_n7425), .B(new_n7432), .C(new_n7437), .Y(new_n7438));
  AOI211xp5_ASAP7_75t_L     g07182(.A1(new_n7107), .A2(new_n7109), .B(new_n7112), .C(new_n7431), .Y(new_n7439));
  NOR2xp33_ASAP7_75t_L      g07183(.A(new_n7103), .B(new_n7100), .Y(new_n7440));
  A2O1A1Ixp33_ASAP7_75t_L   g07184(.A1(\a[26] ), .A2(new_n7096), .B(new_n7097), .C(new_n7440), .Y(new_n7441));
  AOI21xp33_ASAP7_75t_L     g07185(.A1(new_n7125), .A2(new_n7441), .B(new_n7423), .Y(new_n7442));
  INVx1_ASAP7_75t_L         g07186(.A(new_n7437), .Y(new_n7443));
  OAI21xp33_ASAP7_75t_L     g07187(.A1(new_n7442), .A2(new_n7439), .B(new_n7443), .Y(new_n7444));
  A2O1A1O1Ixp25_ASAP7_75t_L g07188(.A1(new_n6840), .A2(new_n6865), .B(new_n6844), .C(new_n7120), .D(new_n7130), .Y(new_n7445));
  AOI21xp33_ASAP7_75t_L     g07189(.A1(new_n7444), .A2(new_n7438), .B(new_n7445), .Y(new_n7446));
  NOR3xp33_ASAP7_75t_L      g07190(.A(new_n7443), .B(new_n7439), .C(new_n7442), .Y(new_n7447));
  AOI21xp33_ASAP7_75t_L     g07191(.A1(new_n7425), .A2(new_n7432), .B(new_n7437), .Y(new_n7448));
  A2O1A1Ixp33_ASAP7_75t_L   g07192(.A1(new_n6565), .A2(new_n6563), .B(new_n6842), .C(new_n6840), .Y(new_n7449));
  A2O1A1Ixp33_ASAP7_75t_L   g07193(.A1(new_n7449), .A2(new_n6845), .B(new_n7129), .C(new_n7127), .Y(new_n7450));
  NOR3xp33_ASAP7_75t_L      g07194(.A(new_n7450), .B(new_n7448), .C(new_n7447), .Y(new_n7451));
  OAI21xp33_ASAP7_75t_L     g07195(.A1(new_n7451), .A2(new_n7446), .B(new_n7292), .Y(new_n7452));
  NOR2xp33_ASAP7_75t_L      g07196(.A(new_n7442), .B(new_n7439), .Y(new_n7453));
  NAND3xp33_ASAP7_75t_L     g07197(.A(new_n7443), .B(new_n7425), .C(new_n7432), .Y(new_n7454));
  A2O1A1Ixp33_ASAP7_75t_L   g07198(.A1(new_n7454), .A2(new_n7453), .B(new_n7448), .C(new_n7450), .Y(new_n7455));
  NAND3xp33_ASAP7_75t_L     g07199(.A(new_n7445), .B(new_n7444), .C(new_n7438), .Y(new_n7456));
  NAND3xp33_ASAP7_75t_L     g07200(.A(new_n7456), .B(new_n7455), .C(new_n7291), .Y(new_n7457));
  NAND3xp33_ASAP7_75t_L     g07201(.A(new_n7285), .B(new_n7452), .C(new_n7457), .Y(new_n7458));
  NOR2xp33_ASAP7_75t_L      g07202(.A(new_n7139), .B(new_n7140), .Y(new_n7459));
  MAJIxp5_ASAP7_75t_L       g07203(.A(new_n6980), .B(new_n7459), .C(new_n7141), .Y(new_n7460));
  NAND2xp33_ASAP7_75t_L     g07204(.A(new_n7457), .B(new_n7452), .Y(new_n7461));
  NAND2xp33_ASAP7_75t_L     g07205(.A(new_n7461), .B(new_n7460), .Y(new_n7462));
  NOR2xp33_ASAP7_75t_L      g07206(.A(new_n3456), .B(new_n2118), .Y(new_n7463));
  AOI221xp5_ASAP7_75t_L     g07207(.A1(\b[29] ), .A2(new_n1290), .B1(\b[31] ), .B2(new_n1209), .C(new_n7463), .Y(new_n7464));
  O2A1O1Ixp33_ASAP7_75t_L   g07208(.A1(new_n1210), .A2(new_n3681), .B(new_n7464), .C(new_n1206), .Y(new_n7465));
  INVx1_ASAP7_75t_L         g07209(.A(new_n7465), .Y(new_n7466));
  O2A1O1Ixp33_ASAP7_75t_L   g07210(.A1(new_n1210), .A2(new_n3681), .B(new_n7464), .C(\a[17] ), .Y(new_n7467));
  AOI21xp33_ASAP7_75t_L     g07211(.A1(new_n7466), .A2(\a[17] ), .B(new_n7467), .Y(new_n7468));
  NAND3xp33_ASAP7_75t_L     g07212(.A(new_n7458), .B(new_n7462), .C(new_n7468), .Y(new_n7469));
  NAND2xp33_ASAP7_75t_L     g07213(.A(new_n7461), .B(new_n7285), .Y(new_n7470));
  NAND2xp33_ASAP7_75t_L     g07214(.A(new_n7455), .B(new_n7456), .Y(new_n7471));
  NOR2xp33_ASAP7_75t_L      g07215(.A(new_n7291), .B(new_n7471), .Y(new_n7472));
  O2A1O1Ixp33_ASAP7_75t_L   g07216(.A1(new_n7291), .A2(new_n7472), .B(new_n7457), .C(new_n7285), .Y(new_n7473));
  AO21x2_ASAP7_75t_L        g07217(.A1(\a[17] ), .A2(new_n7466), .B(new_n7467), .Y(new_n7474));
  A2O1A1Ixp33_ASAP7_75t_L   g07218(.A1(new_n7470), .A2(new_n7285), .B(new_n7473), .C(new_n7474), .Y(new_n7475));
  NAND3xp33_ASAP7_75t_L     g07219(.A(new_n7283), .B(new_n7469), .C(new_n7475), .Y(new_n7476));
  A2O1A1O1Ixp25_ASAP7_75t_L g07220(.A1(new_n6870), .A2(new_n6709), .B(new_n6978), .C(new_n7163), .D(new_n7154), .Y(new_n7477));
  NAND2xp33_ASAP7_75t_L     g07221(.A(new_n7469), .B(new_n7475), .Y(new_n7478));
  NAND2xp33_ASAP7_75t_L     g07222(.A(new_n7477), .B(new_n7478), .Y(new_n7479));
  OAI22xp33_ASAP7_75t_L     g07223(.A1(new_n980), .A2(new_n3891), .B1(new_n4101), .B2(new_n864), .Y(new_n7480));
  AOI221xp5_ASAP7_75t_L     g07224(.A1(new_n886), .A2(\b[34] ), .B1(new_n873), .B2(new_n5599), .C(new_n7480), .Y(new_n7481));
  XNOR2x2_ASAP7_75t_L       g07225(.A(new_n867), .B(new_n7481), .Y(new_n7482));
  NAND3xp33_ASAP7_75t_L     g07226(.A(new_n7479), .B(new_n7476), .C(new_n7482), .Y(new_n7483));
  NOR2xp33_ASAP7_75t_L      g07227(.A(new_n7477), .B(new_n7478), .Y(new_n7484));
  AOI21xp33_ASAP7_75t_L     g07228(.A1(new_n7475), .A2(new_n7469), .B(new_n7283), .Y(new_n7485));
  XNOR2x2_ASAP7_75t_L       g07229(.A(\a[14] ), .B(new_n7481), .Y(new_n7486));
  OAI21xp33_ASAP7_75t_L     g07230(.A1(new_n7485), .A2(new_n7484), .B(new_n7486), .Y(new_n7487));
  NOR2xp33_ASAP7_75t_L      g07231(.A(new_n7174), .B(new_n7173), .Y(new_n7488));
  MAJIxp5_ASAP7_75t_L       g07232(.A(new_n6977), .B(new_n7175), .C(new_n7488), .Y(new_n7489));
  NAND3xp33_ASAP7_75t_L     g07233(.A(new_n7489), .B(new_n7487), .C(new_n7483), .Y(new_n7490));
  NOR3xp33_ASAP7_75t_L      g07234(.A(new_n7484), .B(new_n7485), .C(new_n7486), .Y(new_n7491));
  AOI21xp33_ASAP7_75t_L     g07235(.A1(new_n7479), .A2(new_n7476), .B(new_n7482), .Y(new_n7492));
  NAND2xp33_ASAP7_75t_L     g07236(.A(new_n7165), .B(new_n7160), .Y(new_n7493));
  MAJIxp5_ASAP7_75t_L       g07237(.A(new_n7178), .B(new_n7171), .C(new_n7493), .Y(new_n7494));
  OAI21xp33_ASAP7_75t_L     g07238(.A1(new_n7491), .A2(new_n7492), .B(new_n7494), .Y(new_n7495));
  NOR2xp33_ASAP7_75t_L      g07239(.A(new_n5074), .B(new_n710), .Y(new_n7496));
  AOI221xp5_ASAP7_75t_L     g07240(.A1(\b[36] ), .A2(new_n635), .B1(\b[35] ), .B2(new_n713), .C(new_n7496), .Y(new_n7497));
  O2A1O1Ixp33_ASAP7_75t_L   g07241(.A1(new_n641), .A2(new_n5083), .B(new_n7497), .C(new_n637), .Y(new_n7498));
  OAI21xp33_ASAP7_75t_L     g07242(.A1(new_n641), .A2(new_n5083), .B(new_n7497), .Y(new_n7499));
  NAND2xp33_ASAP7_75t_L     g07243(.A(new_n637), .B(new_n7499), .Y(new_n7500));
  OA21x2_ASAP7_75t_L        g07244(.A1(new_n637), .A2(new_n7498), .B(new_n7500), .Y(new_n7501));
  NAND3xp33_ASAP7_75t_L     g07245(.A(new_n7495), .B(new_n7490), .C(new_n7501), .Y(new_n7502));
  AO21x2_ASAP7_75t_L        g07246(.A1(new_n7490), .A2(new_n7495), .B(new_n7501), .Y(new_n7503));
  A2O1A1O1Ixp25_ASAP7_75t_L g07247(.A1(new_n6906), .A2(new_n6917), .B(new_n7197), .C(new_n7208), .D(new_n7189), .Y(new_n7504));
  AND3x1_ASAP7_75t_L        g07248(.A(new_n7504), .B(new_n7503), .C(new_n7502), .Y(new_n7505));
  AOI21xp33_ASAP7_75t_L     g07249(.A1(new_n7503), .A2(new_n7502), .B(new_n7504), .Y(new_n7506));
  NOR2xp33_ASAP7_75t_L      g07250(.A(new_n5570), .B(new_n513), .Y(new_n7507));
  AOI221xp5_ASAP7_75t_L     g07251(.A1(\b[38] ), .A2(new_n560), .B1(\b[40] ), .B2(new_n475), .C(new_n7507), .Y(new_n7508));
  O2A1O1Ixp33_ASAP7_75t_L   g07252(.A1(new_n477), .A2(new_n5862), .B(new_n7508), .C(new_n466), .Y(new_n7509));
  INVx1_ASAP7_75t_L         g07253(.A(new_n7508), .Y(new_n7510));
  A2O1A1Ixp33_ASAP7_75t_L   g07254(.A1(new_n6651), .A2(new_n483), .B(new_n7510), .C(new_n466), .Y(new_n7511));
  OAI21xp33_ASAP7_75t_L     g07255(.A1(new_n466), .A2(new_n7509), .B(new_n7511), .Y(new_n7512));
  INVx1_ASAP7_75t_L         g07256(.A(new_n7512), .Y(new_n7513));
  OAI21xp33_ASAP7_75t_L     g07257(.A1(new_n7506), .A2(new_n7505), .B(new_n7513), .Y(new_n7514));
  NOR3xp33_ASAP7_75t_L      g07258(.A(new_n7211), .B(new_n7205), .C(new_n7209), .Y(new_n7515));
  O2A1O1Ixp33_ASAP7_75t_L   g07259(.A1(new_n7228), .A2(new_n7213), .B(new_n7218), .C(new_n7515), .Y(new_n7516));
  NOR3xp33_ASAP7_75t_L      g07260(.A(new_n7505), .B(new_n7506), .C(new_n7513), .Y(new_n7517));
  INVx1_ASAP7_75t_L         g07261(.A(new_n7517), .Y(new_n7518));
  AOI21xp33_ASAP7_75t_L     g07262(.A1(new_n7514), .A2(new_n7518), .B(new_n7516), .Y(new_n7519));
  A2O1A1O1Ixp25_ASAP7_75t_L g07263(.A1(new_n7218), .A2(new_n7216), .B(new_n7515), .C(new_n7514), .D(new_n7517), .Y(new_n7520));
  NOR2xp33_ASAP7_75t_L      g07264(.A(new_n6110), .B(new_n375), .Y(new_n7521));
  AOI221xp5_ASAP7_75t_L     g07265(.A1(\b[43] ), .A2(new_n361), .B1(new_n349), .B2(\b[42] ), .C(new_n7521), .Y(new_n7522));
  O2A1O1Ixp33_ASAP7_75t_L   g07266(.A1(new_n356), .A2(new_n6679), .B(new_n7522), .C(new_n346), .Y(new_n7523));
  INVx1_ASAP7_75t_L         g07267(.A(new_n7522), .Y(new_n7524));
  A2O1A1Ixp33_ASAP7_75t_L   g07268(.A1(new_n6682), .A2(new_n359), .B(new_n7524), .C(new_n346), .Y(new_n7525));
  OAI21xp33_ASAP7_75t_L     g07269(.A1(new_n346), .A2(new_n7523), .B(new_n7525), .Y(new_n7526));
  INVx1_ASAP7_75t_L         g07270(.A(new_n7526), .Y(new_n7527));
  A2O1A1Ixp33_ASAP7_75t_L   g07271(.A1(new_n7520), .A2(new_n7514), .B(new_n7519), .C(new_n7527), .Y(new_n7528));
  INVx1_ASAP7_75t_L         g07272(.A(new_n7515), .Y(new_n7529));
  NOR2xp33_ASAP7_75t_L      g07273(.A(new_n7229), .B(new_n7228), .Y(new_n7530));
  A2O1A1Ixp33_ASAP7_75t_L   g07274(.A1(new_n6974), .A2(new_n6931), .B(new_n7530), .C(new_n7529), .Y(new_n7531));
  NAND3xp33_ASAP7_75t_L     g07275(.A(new_n7504), .B(new_n7503), .C(new_n7502), .Y(new_n7532));
  AO21x2_ASAP7_75t_L        g07276(.A1(new_n7502), .A2(new_n7503), .B(new_n7504), .Y(new_n7533));
  AOI21xp33_ASAP7_75t_L     g07277(.A1(new_n7533), .A2(new_n7532), .B(new_n7512), .Y(new_n7534));
  OAI21xp33_ASAP7_75t_L     g07278(.A1(new_n7517), .A2(new_n7534), .B(new_n7531), .Y(new_n7535));
  NAND3xp33_ASAP7_75t_L     g07279(.A(new_n7516), .B(new_n7518), .C(new_n7514), .Y(new_n7536));
  NAND3xp33_ASAP7_75t_L     g07280(.A(new_n7535), .B(new_n7536), .C(new_n7526), .Y(new_n7537));
  NAND2xp33_ASAP7_75t_L     g07281(.A(new_n7528), .B(new_n7537), .Y(new_n7538));
  AOI21xp33_ASAP7_75t_L     g07282(.A1(new_n7236), .A2(new_n7234), .B(new_n7239), .Y(new_n7539));
  XOR2x2_ASAP7_75t_L        g07283(.A(new_n7539), .B(new_n7538), .Y(new_n7540));
  INVx1_ASAP7_75t_L         g07284(.A(new_n7282), .Y(new_n7541));
  O2A1O1Ixp33_ASAP7_75t_L   g07285(.A1(new_n7280), .A2(new_n257), .B(new_n7541), .C(new_n7540), .Y(new_n7542));
  INVx1_ASAP7_75t_L         g07286(.A(new_n7542), .Y(new_n7543));
  NOR2xp33_ASAP7_75t_L      g07287(.A(new_n7540), .B(new_n7542), .Y(new_n7544));
  A2O1A1O1Ixp25_ASAP7_75t_L g07288(.A1(new_n7281), .A2(\a[2] ), .B(new_n7282), .C(new_n7543), .D(new_n7544), .Y(new_n7545));
  A2O1A1O1Ixp25_ASAP7_75t_L g07289(.A1(new_n6962), .A2(new_n6965), .B(new_n6971), .C(new_n7261), .D(new_n7262), .Y(new_n7546));
  INVx1_ASAP7_75t_L         g07290(.A(new_n7546), .Y(new_n7547));
  XNOR2x2_ASAP7_75t_L       g07291(.A(new_n7547), .B(new_n7545), .Y(\f[46] ));
  NOR2xp33_ASAP7_75t_L      g07292(.A(new_n7249), .B(new_n287), .Y(new_n7549));
  AOI221xp5_ASAP7_75t_L     g07293(.A1(\b[46] ), .A2(new_n264), .B1(\b[47] ), .B2(new_n283), .C(new_n7549), .Y(new_n7550));
  NOR2xp33_ASAP7_75t_L      g07294(.A(\b[46] ), .B(\b[47] ), .Y(new_n7551));
  INVx1_ASAP7_75t_L         g07295(.A(\b[47] ), .Y(new_n7552));
  NOR2xp33_ASAP7_75t_L      g07296(.A(new_n7270), .B(new_n7552), .Y(new_n7553));
  NOR2xp33_ASAP7_75t_L      g07297(.A(new_n7551), .B(new_n7553), .Y(new_n7554));
  INVx1_ASAP7_75t_L         g07298(.A(new_n7554), .Y(new_n7555));
  O2A1O1Ixp33_ASAP7_75t_L   g07299(.A1(new_n7249), .A2(new_n7270), .B(new_n7273), .C(new_n7555), .Y(new_n7556));
  INVx1_ASAP7_75t_L         g07300(.A(new_n7556), .Y(new_n7557));
  A2O1A1O1Ixp25_ASAP7_75t_L g07301(.A1(new_n7251), .A2(new_n7268), .B(new_n7250), .C(new_n7272), .D(new_n7271), .Y(new_n7558));
  NAND2xp33_ASAP7_75t_L     g07302(.A(new_n7555), .B(new_n7558), .Y(new_n7559));
  NAND2xp33_ASAP7_75t_L     g07303(.A(new_n7559), .B(new_n7557), .Y(new_n7560));
  O2A1O1Ixp33_ASAP7_75t_L   g07304(.A1(new_n279), .A2(new_n7560), .B(new_n7550), .C(new_n257), .Y(new_n7561));
  INVx1_ASAP7_75t_L         g07305(.A(new_n7561), .Y(new_n7562));
  O2A1O1Ixp33_ASAP7_75t_L   g07306(.A1(new_n279), .A2(new_n7560), .B(new_n7550), .C(\a[2] ), .Y(new_n7563));
  AOI21xp33_ASAP7_75t_L     g07307(.A1(new_n7562), .A2(\a[2] ), .B(new_n7563), .Y(new_n7564));
  A2O1A1Ixp33_ASAP7_75t_L   g07308(.A1(new_n7520), .A2(new_n7514), .B(new_n7519), .C(new_n7526), .Y(new_n7565));
  A2O1A1O1Ixp25_ASAP7_75t_L g07309(.A1(new_n6931), .A2(new_n6974), .B(new_n7530), .C(new_n7529), .D(new_n7534), .Y(new_n7566));
  A2O1A1O1Ixp25_ASAP7_75t_L g07310(.A1(new_n7518), .A2(new_n7566), .B(new_n7516), .C(new_n7536), .D(new_n7526), .Y(new_n7567));
  AOI21xp33_ASAP7_75t_L     g07311(.A1(new_n7565), .A2(new_n7526), .B(new_n7567), .Y(new_n7568));
  A2O1A1Ixp33_ASAP7_75t_L   g07312(.A1(\a[20] ), .A2(new_n7135), .B(new_n7136), .C(new_n7459), .Y(new_n7569));
  A2O1A1O1Ixp25_ASAP7_75t_L g07313(.A1(new_n7142), .A2(new_n7284), .B(new_n7144), .C(new_n7569), .D(new_n7461), .Y(new_n7570));
  NOR3xp33_ASAP7_75t_L      g07314(.A(new_n7570), .B(new_n7473), .C(new_n7474), .Y(new_n7571));
  OAI21xp33_ASAP7_75t_L     g07315(.A1(new_n7571), .A2(new_n7477), .B(new_n7475), .Y(new_n7572));
  NOR2xp33_ASAP7_75t_L      g07316(.A(new_n3674), .B(new_n2118), .Y(new_n7573));
  AOI221xp5_ASAP7_75t_L     g07317(.A1(\b[30] ), .A2(new_n1290), .B1(\b[32] ), .B2(new_n1209), .C(new_n7573), .Y(new_n7574));
  O2A1O1Ixp33_ASAP7_75t_L   g07318(.A1(new_n1210), .A2(new_n3897), .B(new_n7574), .C(new_n1206), .Y(new_n7575));
  INVx1_ASAP7_75t_L         g07319(.A(new_n7574), .Y(new_n7576));
  A2O1A1Ixp33_ASAP7_75t_L   g07320(.A1(new_n3900), .A2(new_n1216), .B(new_n7576), .C(new_n1206), .Y(new_n7577));
  OAI21xp33_ASAP7_75t_L     g07321(.A1(new_n1206), .A2(new_n7575), .B(new_n7577), .Y(new_n7578));
  INVx1_ASAP7_75t_L         g07322(.A(new_n7578), .Y(new_n7579));
  NOR2xp33_ASAP7_75t_L      g07323(.A(new_n7292), .B(new_n7471), .Y(new_n7580));
  O2A1O1Ixp33_ASAP7_75t_L   g07324(.A1(new_n7292), .A2(new_n7580), .B(new_n7285), .C(new_n7472), .Y(new_n7581));
  OAI22xp33_ASAP7_75t_L     g07325(.A1(new_n1654), .A2(new_n2879), .B1(new_n3079), .B2(new_n1517), .Y(new_n7582));
  AOI221xp5_ASAP7_75t_L     g07326(.A1(new_n1511), .A2(\b[29] ), .B1(new_n1513), .B2(new_n3873), .C(new_n7582), .Y(new_n7583));
  XNOR2x2_ASAP7_75t_L       g07327(.A(new_n1501), .B(new_n7583), .Y(new_n7584));
  MAJIxp5_ASAP7_75t_L       g07328(.A(new_n7450), .B(new_n7443), .C(new_n7453), .Y(new_n7585));
  NOR3xp33_ASAP7_75t_L      g07329(.A(new_n7393), .B(new_n7394), .C(new_n7391), .Y(new_n7586));
  O2A1O1Ixp33_ASAP7_75t_L   g07330(.A1(new_n7397), .A2(new_n7401), .B(new_n7403), .C(new_n7586), .Y(new_n7587));
  OAI22xp33_ASAP7_75t_L     g07331(.A1(new_n3703), .A2(new_n1043), .B1(new_n1150), .B2(new_n3509), .Y(new_n7588));
  AOI221xp5_ASAP7_75t_L     g07332(.A1(new_n3503), .A2(\b[17] ), .B1(new_n3505), .B2(new_n1633), .C(new_n7588), .Y(new_n7589));
  XNOR2x2_ASAP7_75t_L       g07333(.A(\a[32] ), .B(new_n7589), .Y(new_n7590));
  O2A1O1Ixp33_ASAP7_75t_L   g07334(.A1(new_n4145), .A2(new_n6987), .B(new_n6989), .C(new_n7299), .Y(new_n7591));
  XNOR2x2_ASAP7_75t_L       g07335(.A(new_n7357), .B(new_n7359), .Y(new_n7592));
  MAJIxp5_ASAP7_75t_L       g07336(.A(new_n7301), .B(new_n7592), .C(new_n7364), .Y(new_n7593));
  A2O1A1O1Ixp25_ASAP7_75t_L g07337(.A1(new_n7364), .A2(new_n7592), .B(new_n7593), .C(new_n7367), .D(new_n7373), .Y(new_n7594));
  A2O1A1O1Ixp25_ASAP7_75t_L g07338(.A1(new_n6984), .A2(new_n7058), .B(new_n7591), .C(new_n7374), .D(new_n7594), .Y(new_n7595));
  NAND2xp33_ASAP7_75t_L     g07339(.A(new_n7346), .B(new_n7339), .Y(new_n7596));
  O2A1O1Ixp33_ASAP7_75t_L   g07340(.A1(new_n5630), .A2(new_n456), .B(new_n7348), .C(new_n5626), .Y(new_n7597));
  O2A1O1Ixp33_ASAP7_75t_L   g07341(.A1(new_n7597), .A2(new_n5626), .B(new_n7351), .C(new_n7596), .Y(new_n7598));
  AOI21xp33_ASAP7_75t_L     g07342(.A1(new_n7359), .A2(new_n7357), .B(new_n7598), .Y(new_n7599));
  NOR2xp33_ASAP7_75t_L      g07343(.A(new_n448), .B(new_n5640), .Y(new_n7600));
  AOI221xp5_ASAP7_75t_L     g07344(.A1(\b[6] ), .A2(new_n5920), .B1(\b[8] ), .B2(new_n5629), .C(new_n7600), .Y(new_n7601));
  O2A1O1Ixp33_ASAP7_75t_L   g07345(.A1(new_n5630), .A2(new_n540), .B(new_n7601), .C(new_n5626), .Y(new_n7602));
  INVx1_ASAP7_75t_L         g07346(.A(new_n7602), .Y(new_n7603));
  O2A1O1Ixp33_ASAP7_75t_L   g07347(.A1(new_n5630), .A2(new_n540), .B(new_n7601), .C(\a[41] ), .Y(new_n7604));
  AOI21xp33_ASAP7_75t_L     g07348(.A1(new_n7603), .A2(\a[41] ), .B(new_n7604), .Y(new_n7605));
  INVx1_ASAP7_75t_L         g07349(.A(new_n7604), .Y(new_n7606));
  OAI21xp33_ASAP7_75t_L     g07350(.A1(new_n7342), .A2(new_n7341), .B(new_n7338), .Y(new_n7607));
  NOR2xp33_ASAP7_75t_L      g07351(.A(new_n289), .B(new_n7318), .Y(new_n7608));
  AOI211xp5_ASAP7_75t_L     g07352(.A1(new_n7315), .A2(new_n7317), .B(new_n7311), .C(new_n7313), .Y(new_n7609));
  AOI221xp5_ASAP7_75t_L     g07353(.A1(new_n7333), .A2(\b[1] ), .B1(new_n7609), .B2(\b[0] ), .C(new_n7608), .Y(new_n7610));
  NOR2xp33_ASAP7_75t_L      g07354(.A(new_n7321), .B(new_n509), .Y(new_n7611));
  INVx1_ASAP7_75t_L         g07355(.A(new_n7611), .Y(new_n7612));
  NAND3xp33_ASAP7_75t_L     g07356(.A(new_n7610), .B(\a[47] ), .C(new_n7612), .Y(new_n7613));
  INVx1_ASAP7_75t_L         g07357(.A(new_n7609), .Y(new_n7614));
  NAND2xp33_ASAP7_75t_L     g07358(.A(\b[1] ), .B(new_n7333), .Y(new_n7615));
  OAI221xp5_ASAP7_75t_L     g07359(.A1(new_n7318), .A2(new_n289), .B1(new_n284), .B2(new_n7614), .C(new_n7615), .Y(new_n7616));
  A2O1A1Ixp33_ASAP7_75t_L   g07360(.A1(new_n294), .A2(new_n7322), .B(new_n7616), .C(new_n7316), .Y(new_n7617));
  NAND3xp33_ASAP7_75t_L     g07361(.A(new_n7617), .B(new_n7324), .C(new_n7613), .Y(new_n7618));
  NAND5xp2_ASAP7_75t_L      g07362(.A(\a[47] ), .B(new_n7323), .C(new_n7612), .D(new_n7610), .E(new_n7302), .Y(new_n7619));
  NOR2xp33_ASAP7_75t_L      g07363(.A(new_n301), .B(new_n6741), .Y(new_n7620));
  AOI221xp5_ASAP7_75t_L     g07364(.A1(\b[5] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[4] ), .C(new_n7620), .Y(new_n7621));
  NAND2xp33_ASAP7_75t_L     g07365(.A(new_n6450), .B(new_n394), .Y(new_n7622));
  NAND3xp33_ASAP7_75t_L     g07366(.A(new_n7622), .B(new_n7621), .C(\a[44] ), .Y(new_n7623));
  OAI21xp33_ASAP7_75t_L     g07367(.A1(new_n728), .A2(new_n6443), .B(new_n7621), .Y(new_n7624));
  NAND2xp33_ASAP7_75t_L     g07368(.A(new_n6439), .B(new_n7624), .Y(new_n7625));
  AND4x1_ASAP7_75t_L        g07369(.A(new_n7618), .B(new_n7625), .C(new_n7623), .D(new_n7619), .Y(new_n7626));
  AOI22xp33_ASAP7_75t_L     g07370(.A1(new_n7623), .A2(new_n7625), .B1(new_n7619), .B2(new_n7618), .Y(new_n7627));
  OAI21xp33_ASAP7_75t_L     g07371(.A1(new_n7626), .A2(new_n7627), .B(new_n7607), .Y(new_n7628));
  AOI21xp33_ASAP7_75t_L     g07372(.A1(new_n7303), .A2(new_n7330), .B(new_n7345), .Y(new_n7629));
  NOR2xp33_ASAP7_75t_L      g07373(.A(new_n7627), .B(new_n7626), .Y(new_n7630));
  NAND2xp33_ASAP7_75t_L     g07374(.A(new_n7630), .B(new_n7629), .Y(new_n7631));
  NAND2xp33_ASAP7_75t_L     g07375(.A(new_n7628), .B(new_n7631), .Y(new_n7632));
  O2A1O1Ixp33_ASAP7_75t_L   g07376(.A1(new_n5626), .A2(new_n7602), .B(new_n7606), .C(new_n7632), .Y(new_n7633));
  NAND3xp33_ASAP7_75t_L     g07377(.A(new_n7631), .B(new_n7605), .C(new_n7628), .Y(new_n7634));
  O2A1O1Ixp33_ASAP7_75t_L   g07378(.A1(new_n7605), .A2(new_n7633), .B(new_n7634), .C(new_n7599), .Y(new_n7635));
  OAI21xp33_ASAP7_75t_L     g07379(.A1(new_n5626), .A2(new_n7602), .B(new_n7606), .Y(new_n7636));
  NOR2xp33_ASAP7_75t_L      g07380(.A(new_n7630), .B(new_n7629), .Y(new_n7637));
  NOR3xp33_ASAP7_75t_L      g07381(.A(new_n7607), .B(new_n7626), .C(new_n7627), .Y(new_n7638));
  NOR2xp33_ASAP7_75t_L      g07382(.A(new_n7638), .B(new_n7637), .Y(new_n7639));
  A2O1A1Ixp33_ASAP7_75t_L   g07383(.A1(new_n7603), .A2(\a[41] ), .B(new_n7604), .C(new_n7639), .Y(new_n7640));
  INVx1_ASAP7_75t_L         g07384(.A(new_n7634), .Y(new_n7641));
  A2O1A1Ixp33_ASAP7_75t_L   g07385(.A1(new_n7640), .A2(new_n7636), .B(new_n7641), .C(new_n7599), .Y(new_n7642));
  NOR2xp33_ASAP7_75t_L      g07386(.A(new_n748), .B(new_n4908), .Y(new_n7643));
  AOI221xp5_ASAP7_75t_L     g07387(.A1(\b[9] ), .A2(new_n5139), .B1(\b[10] ), .B2(new_n4916), .C(new_n7643), .Y(new_n7644));
  O2A1O1Ixp33_ASAP7_75t_L   g07388(.A1(new_n4911), .A2(new_n754), .B(new_n7644), .C(new_n4906), .Y(new_n7645));
  OAI21xp33_ASAP7_75t_L     g07389(.A1(new_n4911), .A2(new_n754), .B(new_n7644), .Y(new_n7646));
  NAND2xp33_ASAP7_75t_L     g07390(.A(new_n4906), .B(new_n7646), .Y(new_n7647));
  OAI21xp33_ASAP7_75t_L     g07391(.A1(new_n4906), .A2(new_n7645), .B(new_n7647), .Y(new_n7648));
  INVx1_ASAP7_75t_L         g07392(.A(new_n7648), .Y(new_n7649));
  OAI211xp5_ASAP7_75t_L     g07393(.A1(new_n7599), .A2(new_n7635), .B(new_n7642), .C(new_n7649), .Y(new_n7650));
  OAI21xp33_ASAP7_75t_L     g07394(.A1(new_n7638), .A2(new_n7637), .B(new_n7636), .Y(new_n7651));
  NAND2xp33_ASAP7_75t_L     g07395(.A(new_n7634), .B(new_n7651), .Y(new_n7652));
  A2O1A1Ixp33_ASAP7_75t_L   g07396(.A1(new_n7357), .A2(new_n7359), .B(new_n7598), .C(new_n7652), .Y(new_n7653));
  NOR2xp33_ASAP7_75t_L      g07397(.A(new_n7652), .B(new_n7599), .Y(new_n7654));
  A2O1A1Ixp33_ASAP7_75t_L   g07398(.A1(new_n7653), .A2(new_n7652), .B(new_n7654), .C(new_n7648), .Y(new_n7655));
  NAND3xp33_ASAP7_75t_L     g07399(.A(new_n7593), .B(new_n7650), .C(new_n7655), .Y(new_n7656));
  AO21x2_ASAP7_75t_L        g07400(.A1(new_n7357), .A2(new_n7359), .B(new_n7598), .Y(new_n7657));
  O2A1O1Ixp33_ASAP7_75t_L   g07401(.A1(new_n7605), .A2(new_n7633), .B(new_n7634), .C(new_n7657), .Y(new_n7658));
  NOR3xp33_ASAP7_75t_L      g07402(.A(new_n7658), .B(new_n7648), .C(new_n7654), .Y(new_n7659));
  O2A1O1Ixp33_ASAP7_75t_L   g07403(.A1(new_n7599), .A2(new_n7635), .B(new_n7642), .C(new_n7649), .Y(new_n7660));
  OAI21xp33_ASAP7_75t_L     g07404(.A1(new_n7659), .A2(new_n7660), .B(new_n7377), .Y(new_n7661));
  NAND2xp33_ASAP7_75t_L     g07405(.A(new_n7661), .B(new_n7656), .Y(new_n7662));
  NOR2xp33_ASAP7_75t_L      g07406(.A(new_n960), .B(new_n4147), .Y(new_n7663));
  AOI221xp5_ASAP7_75t_L     g07407(.A1(\b[12] ), .A2(new_n4402), .B1(\b[13] ), .B2(new_n4155), .C(new_n7663), .Y(new_n7664));
  O2A1O1Ixp33_ASAP7_75t_L   g07408(.A1(new_n4150), .A2(new_n1268), .B(new_n7664), .C(new_n4145), .Y(new_n7665));
  O2A1O1Ixp33_ASAP7_75t_L   g07409(.A1(new_n4150), .A2(new_n1268), .B(new_n7664), .C(\a[35] ), .Y(new_n7666));
  INVx1_ASAP7_75t_L         g07410(.A(new_n7666), .Y(new_n7667));
  OAI21xp33_ASAP7_75t_L     g07411(.A1(new_n4145), .A2(new_n7665), .B(new_n7667), .Y(new_n7668));
  NAND3xp33_ASAP7_75t_L     g07412(.A(new_n7656), .B(new_n7668), .C(new_n7661), .Y(new_n7669));
  INVx1_ASAP7_75t_L         g07413(.A(new_n7669), .Y(new_n7670));
  NOR3xp33_ASAP7_75t_L      g07414(.A(new_n7377), .B(new_n7660), .C(new_n7659), .Y(new_n7671));
  AOI21xp33_ASAP7_75t_L     g07415(.A1(new_n7655), .A2(new_n7650), .B(new_n7593), .Y(new_n7672));
  OAI21xp33_ASAP7_75t_L     g07416(.A1(new_n7671), .A2(new_n7672), .B(new_n7668), .Y(new_n7673));
  O2A1O1Ixp33_ASAP7_75t_L   g07417(.A1(new_n7662), .A2(new_n7670), .B(new_n7673), .C(new_n7595), .Y(new_n7674));
  NAND2xp33_ASAP7_75t_L     g07418(.A(new_n6990), .B(new_n7383), .Y(new_n7675));
  AOI211xp5_ASAP7_75t_L     g07419(.A1(new_n7377), .A2(new_n7366), .B(new_n7375), .C(new_n7380), .Y(new_n7676));
  A2O1A1Ixp33_ASAP7_75t_L   g07420(.A1(new_n7069), .A2(new_n7675), .B(new_n7676), .C(new_n7381), .Y(new_n7677));
  OAI211xp5_ASAP7_75t_L     g07421(.A1(new_n4150), .A2(new_n1268), .B(\a[35] ), .C(new_n7664), .Y(new_n7678));
  NAND4xp25_ASAP7_75t_L     g07422(.A(new_n7656), .B(new_n7667), .C(new_n7661), .D(new_n7678), .Y(new_n7679));
  NAND2xp33_ASAP7_75t_L     g07423(.A(new_n7679), .B(new_n7673), .Y(new_n7680));
  NOR2xp33_ASAP7_75t_L      g07424(.A(new_n7677), .B(new_n7680), .Y(new_n7681));
  OAI21xp33_ASAP7_75t_L     g07425(.A1(new_n7681), .A2(new_n7674), .B(new_n7590), .Y(new_n7682));
  XNOR2x2_ASAP7_75t_L       g07426(.A(new_n3493), .B(new_n7589), .Y(new_n7683));
  A2O1A1Ixp33_ASAP7_75t_L   g07427(.A1(new_n7374), .A2(new_n7300), .B(new_n7594), .C(new_n7680), .Y(new_n7684));
  NAND3xp33_ASAP7_75t_L     g07428(.A(new_n7595), .B(new_n7679), .C(new_n7673), .Y(new_n7685));
  NAND3xp33_ASAP7_75t_L     g07429(.A(new_n7684), .B(new_n7683), .C(new_n7685), .Y(new_n7686));
  AOI21xp33_ASAP7_75t_L     g07430(.A1(new_n7686), .A2(new_n7682), .B(new_n7587), .Y(new_n7687));
  NAND3xp33_ASAP7_75t_L     g07431(.A(new_n7684), .B(new_n7590), .C(new_n7685), .Y(new_n7688));
  NOR3xp33_ASAP7_75t_L      g07432(.A(new_n7674), .B(new_n7681), .C(new_n7590), .Y(new_n7689));
  A2O1A1Ixp33_ASAP7_75t_L   g07433(.A1(new_n7590), .A2(new_n7688), .B(new_n7689), .C(new_n7587), .Y(new_n7690));
  NOR2xp33_ASAP7_75t_L      g07434(.A(new_n1745), .B(new_n2930), .Y(new_n7691));
  AOI221xp5_ASAP7_75t_L     g07435(.A1(\b[18] ), .A2(new_n3129), .B1(\b[19] ), .B2(new_n2936), .C(new_n7691), .Y(new_n7692));
  O2A1O1Ixp33_ASAP7_75t_L   g07436(.A1(new_n2940), .A2(new_n1754), .B(new_n7692), .C(new_n2928), .Y(new_n7693));
  OAI21xp33_ASAP7_75t_L     g07437(.A1(new_n2940), .A2(new_n1754), .B(new_n7692), .Y(new_n7694));
  NAND2xp33_ASAP7_75t_L     g07438(.A(new_n2928), .B(new_n7694), .Y(new_n7695));
  OAI21xp33_ASAP7_75t_L     g07439(.A1(new_n2928), .A2(new_n7693), .B(new_n7695), .Y(new_n7696));
  O2A1O1Ixp33_ASAP7_75t_L   g07440(.A1(new_n7587), .A2(new_n7687), .B(new_n7690), .C(new_n7696), .Y(new_n7697));
  AOI21xp33_ASAP7_75t_L     g07441(.A1(new_n7684), .A2(new_n7685), .B(new_n7683), .Y(new_n7698));
  NOR3xp33_ASAP7_75t_L      g07442(.A(new_n7587), .B(new_n7698), .C(new_n7689), .Y(new_n7699));
  A2O1A1Ixp33_ASAP7_75t_L   g07443(.A1(new_n7396), .A2(new_n7395), .B(new_n7586), .C(new_n7392), .Y(new_n7700));
  AOI221xp5_ASAP7_75t_L     g07444(.A1(new_n7686), .A2(new_n7682), .B1(new_n7403), .B2(new_n7700), .C(new_n7586), .Y(new_n7701));
  OA21x2_ASAP7_75t_L        g07445(.A1(new_n2928), .A2(new_n7693), .B(new_n7695), .Y(new_n7702));
  NOR3xp33_ASAP7_75t_L      g07446(.A(new_n7702), .B(new_n7701), .C(new_n7699), .Y(new_n7703));
  NAND2xp33_ASAP7_75t_L     g07447(.A(new_n7404), .B(new_n7400), .Y(new_n7704));
  MAJIxp5_ASAP7_75t_L       g07448(.A(new_n7416), .B(new_n7410), .C(new_n7704), .Y(new_n7705));
  NOR3xp33_ASAP7_75t_L      g07449(.A(new_n7705), .B(new_n7703), .C(new_n7697), .Y(new_n7706));
  OAI21xp33_ASAP7_75t_L     g07450(.A1(new_n7697), .A2(new_n7703), .B(new_n7705), .Y(new_n7707));
  INVx1_ASAP7_75t_L         g07451(.A(new_n7707), .Y(new_n7708));
  NOR2xp33_ASAP7_75t_L      g07452(.A(new_n2188), .B(new_n2415), .Y(new_n7709));
  AOI221xp5_ASAP7_75t_L     g07453(.A1(\b[21] ), .A2(new_n2577), .B1(\b[22] ), .B2(new_n2421), .C(new_n7709), .Y(new_n7710));
  O2A1O1Ixp33_ASAP7_75t_L   g07454(.A1(new_n2425), .A2(new_n2194), .B(new_n7710), .C(new_n2413), .Y(new_n7711));
  OAI21xp33_ASAP7_75t_L     g07455(.A1(new_n2425), .A2(new_n2194), .B(new_n7710), .Y(new_n7712));
  NAND2xp33_ASAP7_75t_L     g07456(.A(new_n2413), .B(new_n7712), .Y(new_n7713));
  OAI21xp33_ASAP7_75t_L     g07457(.A1(new_n2413), .A2(new_n7711), .B(new_n7713), .Y(new_n7714));
  INVx1_ASAP7_75t_L         g07458(.A(new_n7714), .Y(new_n7715));
  OAI21xp33_ASAP7_75t_L     g07459(.A1(new_n7708), .A2(new_n7706), .B(new_n7715), .Y(new_n7716));
  INVx1_ASAP7_75t_L         g07460(.A(new_n7419), .Y(new_n7717));
  A2O1A1O1Ixp25_ASAP7_75t_L g07461(.A1(new_n7107), .A2(new_n7109), .B(new_n7112), .C(new_n7431), .D(new_n7717), .Y(new_n7718));
  O2A1O1Ixp33_ASAP7_75t_L   g07462(.A1(new_n7587), .A2(new_n7687), .B(new_n7690), .C(new_n7702), .Y(new_n7719));
  INVx1_ASAP7_75t_L         g07463(.A(new_n7697), .Y(new_n7720));
  NOR2xp33_ASAP7_75t_L      g07464(.A(new_n7412), .B(new_n7413), .Y(new_n7721));
  OAI21xp33_ASAP7_75t_L     g07465(.A1(new_n7088), .A2(new_n7091), .B(new_n7101), .Y(new_n7722));
  MAJIxp5_ASAP7_75t_L       g07466(.A(new_n7722), .B(new_n7721), .C(new_n7414), .Y(new_n7723));
  OAI211xp5_ASAP7_75t_L     g07467(.A1(new_n7702), .A2(new_n7719), .B(new_n7723), .C(new_n7720), .Y(new_n7724));
  NAND3xp33_ASAP7_75t_L     g07468(.A(new_n7724), .B(new_n7707), .C(new_n7714), .Y(new_n7725));
  AOI21xp33_ASAP7_75t_L     g07469(.A1(new_n7716), .A2(new_n7725), .B(new_n7718), .Y(new_n7726));
  OAI21xp33_ASAP7_75t_L     g07470(.A1(new_n7123), .A2(new_n7115), .B(new_n7441), .Y(new_n7727));
  NOR3xp33_ASAP7_75t_L      g07471(.A(new_n7715), .B(new_n7708), .C(new_n7706), .Y(new_n7728));
  A2O1A1O1Ixp25_ASAP7_75t_L g07472(.A1(new_n7431), .A2(new_n7727), .B(new_n7717), .C(new_n7716), .D(new_n7728), .Y(new_n7729));
  NAND2xp33_ASAP7_75t_L     g07473(.A(\b[26] ), .B(new_n1955), .Y(new_n7730));
  OAI221xp5_ASAP7_75t_L     g07474(.A1(new_n1962), .A2(new_n2377), .B1(new_n2205), .B2(new_n2089), .C(new_n7730), .Y(new_n7731));
  A2O1A1Ixp33_ASAP7_75t_L   g07475(.A1(new_n2709), .A2(new_n1964), .B(new_n7731), .C(\a[23] ), .Y(new_n7732));
  AOI211xp5_ASAP7_75t_L     g07476(.A1(new_n2709), .A2(new_n1964), .B(new_n7731), .C(new_n1952), .Y(new_n7733));
  A2O1A1O1Ixp25_ASAP7_75t_L g07477(.A1(new_n2709), .A2(new_n1964), .B(new_n7731), .C(new_n7732), .D(new_n7733), .Y(new_n7734));
  INVx1_ASAP7_75t_L         g07478(.A(new_n7734), .Y(new_n7735));
  AOI211xp5_ASAP7_75t_L     g07479(.A1(new_n7729), .A2(new_n7716), .B(new_n7726), .C(new_n7735), .Y(new_n7736));
  AOI21xp33_ASAP7_75t_L     g07480(.A1(new_n7724), .A2(new_n7707), .B(new_n7714), .Y(new_n7737));
  O2A1O1Ixp33_ASAP7_75t_L   g07481(.A1(new_n7423), .A2(new_n7424), .B(new_n7419), .C(new_n7737), .Y(new_n7738));
  NAND3xp33_ASAP7_75t_L     g07482(.A(new_n7718), .B(new_n7725), .C(new_n7716), .Y(new_n7739));
  A2O1A1O1Ixp25_ASAP7_75t_L g07483(.A1(new_n7725), .A2(new_n7738), .B(new_n7718), .C(new_n7739), .D(new_n7734), .Y(new_n7740));
  NOR3xp33_ASAP7_75t_L      g07484(.A(new_n7585), .B(new_n7736), .C(new_n7740), .Y(new_n7741));
  A2O1A1Ixp33_ASAP7_75t_L   g07485(.A1(new_n7437), .A2(new_n7438), .B(new_n7445), .C(new_n7454), .Y(new_n7742));
  A2O1A1Ixp33_ASAP7_75t_L   g07486(.A1(new_n7125), .A2(new_n7441), .B(new_n7423), .C(new_n7419), .Y(new_n7743));
  OAI21xp33_ASAP7_75t_L     g07487(.A1(new_n7728), .A2(new_n7737), .B(new_n7743), .Y(new_n7744));
  NAND3xp33_ASAP7_75t_L     g07488(.A(new_n7744), .B(new_n7739), .C(new_n7734), .Y(new_n7745));
  A2O1A1Ixp33_ASAP7_75t_L   g07489(.A1(new_n7729), .A2(new_n7716), .B(new_n7726), .C(new_n7735), .Y(new_n7746));
  AOI21xp33_ASAP7_75t_L     g07490(.A1(new_n7746), .A2(new_n7745), .B(new_n7742), .Y(new_n7747));
  OAI21xp33_ASAP7_75t_L     g07491(.A1(new_n7741), .A2(new_n7747), .B(new_n7584), .Y(new_n7748));
  AND2x2_ASAP7_75t_L        g07492(.A(\a[20] ), .B(new_n7583), .Y(new_n7749));
  NOR2xp33_ASAP7_75t_L      g07493(.A(\a[20] ), .B(new_n7583), .Y(new_n7750));
  NAND3xp33_ASAP7_75t_L     g07494(.A(new_n7742), .B(new_n7745), .C(new_n7746), .Y(new_n7751));
  OAI21xp33_ASAP7_75t_L     g07495(.A1(new_n7740), .A2(new_n7736), .B(new_n7585), .Y(new_n7752));
  OAI211xp5_ASAP7_75t_L     g07496(.A1(new_n7750), .A2(new_n7749), .B(new_n7751), .C(new_n7752), .Y(new_n7753));
  NAND2xp33_ASAP7_75t_L     g07497(.A(new_n7748), .B(new_n7753), .Y(new_n7754));
  NOR2xp33_ASAP7_75t_L      g07498(.A(new_n7754), .B(new_n7581), .Y(new_n7755));
  MAJIxp5_ASAP7_75t_L       g07499(.A(new_n7460), .B(new_n7291), .C(new_n7471), .Y(new_n7756));
  AOI21xp33_ASAP7_75t_L     g07500(.A1(new_n7753), .A2(new_n7748), .B(new_n7756), .Y(new_n7757));
  OAI21xp33_ASAP7_75t_L     g07501(.A1(new_n7757), .A2(new_n7755), .B(new_n7579), .Y(new_n7758));
  NAND3xp33_ASAP7_75t_L     g07502(.A(new_n7756), .B(new_n7748), .C(new_n7753), .Y(new_n7759));
  NAND2xp33_ASAP7_75t_L     g07503(.A(new_n7754), .B(new_n7581), .Y(new_n7760));
  NAND3xp33_ASAP7_75t_L     g07504(.A(new_n7760), .B(new_n7759), .C(new_n7578), .Y(new_n7761));
  NAND3xp33_ASAP7_75t_L     g07505(.A(new_n7572), .B(new_n7758), .C(new_n7761), .Y(new_n7762));
  INVx1_ASAP7_75t_L         g07506(.A(new_n6870), .Y(new_n7763));
  OAI21xp33_ASAP7_75t_L     g07507(.A1(new_n7763), .A2(new_n6877), .B(new_n6875), .Y(new_n7764));
  AOI21xp33_ASAP7_75t_L     g07508(.A1(new_n7458), .A2(new_n7462), .B(new_n7468), .Y(new_n7765));
  A2O1A1O1Ixp25_ASAP7_75t_L g07509(.A1(new_n7159), .A2(new_n7764), .B(new_n7154), .C(new_n7469), .D(new_n7765), .Y(new_n7766));
  AOI21xp33_ASAP7_75t_L     g07510(.A1(new_n7760), .A2(new_n7759), .B(new_n7578), .Y(new_n7767));
  NOR3xp33_ASAP7_75t_L      g07511(.A(new_n7755), .B(new_n7757), .C(new_n7579), .Y(new_n7768));
  OAI21xp33_ASAP7_75t_L     g07512(.A1(new_n7767), .A2(new_n7768), .B(new_n7766), .Y(new_n7769));
  NOR2xp33_ASAP7_75t_L      g07513(.A(new_n4344), .B(new_n864), .Y(new_n7770));
  AOI221xp5_ASAP7_75t_L     g07514(.A1(\b[33] ), .A2(new_n985), .B1(\b[35] ), .B2(new_n886), .C(new_n7770), .Y(new_n7771));
  OAI211xp5_ASAP7_75t_L     g07515(.A1(new_n872), .A2(new_n4589), .B(\a[14] ), .C(new_n7771), .Y(new_n7772));
  INVx1_ASAP7_75t_L         g07516(.A(new_n4589), .Y(new_n7773));
  INVx1_ASAP7_75t_L         g07517(.A(new_n7771), .Y(new_n7774));
  A2O1A1Ixp33_ASAP7_75t_L   g07518(.A1(new_n7773), .A2(new_n873), .B(new_n7774), .C(new_n867), .Y(new_n7775));
  NAND4xp25_ASAP7_75t_L     g07519(.A(new_n7762), .B(new_n7769), .C(new_n7775), .D(new_n7772), .Y(new_n7776));
  NOR3xp33_ASAP7_75t_L      g07520(.A(new_n7766), .B(new_n7767), .C(new_n7768), .Y(new_n7777));
  AOI21xp33_ASAP7_75t_L     g07521(.A1(new_n7761), .A2(new_n7758), .B(new_n7572), .Y(new_n7778));
  NAND2xp33_ASAP7_75t_L     g07522(.A(new_n7772), .B(new_n7775), .Y(new_n7779));
  OAI21xp33_ASAP7_75t_L     g07523(.A1(new_n7778), .A2(new_n7777), .B(new_n7779), .Y(new_n7780));
  NAND2xp33_ASAP7_75t_L     g07524(.A(new_n7776), .B(new_n7780), .Y(new_n7781));
  NAND2xp33_ASAP7_75t_L     g07525(.A(new_n7476), .B(new_n7479), .Y(new_n7782));
  MAJIxp5_ASAP7_75t_L       g07526(.A(new_n7489), .B(new_n7482), .C(new_n7782), .Y(new_n7783));
  NOR2xp33_ASAP7_75t_L      g07527(.A(new_n7783), .B(new_n7781), .Y(new_n7784));
  NOR2xp33_ASAP7_75t_L      g07528(.A(new_n7485), .B(new_n7484), .Y(new_n7785));
  MAJIxp5_ASAP7_75t_L       g07529(.A(new_n7494), .B(new_n7486), .C(new_n7785), .Y(new_n7786));
  AOI21xp33_ASAP7_75t_L     g07530(.A1(new_n7780), .A2(new_n7776), .B(new_n7786), .Y(new_n7787));
  OAI22xp33_ASAP7_75t_L     g07531(.A1(new_n1550), .A2(new_n5074), .B1(new_n4613), .B2(new_n712), .Y(new_n7788));
  AOI221xp5_ASAP7_75t_L     g07532(.A1(new_n640), .A2(\b[38] ), .B1(new_n718), .B2(new_n6083), .C(new_n7788), .Y(new_n7789));
  XNOR2x2_ASAP7_75t_L       g07533(.A(\a[11] ), .B(new_n7789), .Y(new_n7790));
  NOR3xp33_ASAP7_75t_L      g07534(.A(new_n7787), .B(new_n7784), .C(new_n7790), .Y(new_n7791));
  NAND3xp33_ASAP7_75t_L     g07535(.A(new_n7786), .B(new_n7780), .C(new_n7776), .Y(new_n7792));
  NAND2xp33_ASAP7_75t_L     g07536(.A(new_n7783), .B(new_n7781), .Y(new_n7793));
  XNOR2x2_ASAP7_75t_L       g07537(.A(new_n637), .B(new_n7789), .Y(new_n7794));
  AOI21xp33_ASAP7_75t_L     g07538(.A1(new_n7792), .A2(new_n7793), .B(new_n7794), .Y(new_n7795));
  NAND2xp33_ASAP7_75t_L     g07539(.A(new_n7490), .B(new_n7495), .Y(new_n7796));
  MAJIxp5_ASAP7_75t_L       g07540(.A(new_n7504), .B(new_n7796), .C(new_n7501), .Y(new_n7797));
  NOR3xp33_ASAP7_75t_L      g07541(.A(new_n7797), .B(new_n7795), .C(new_n7791), .Y(new_n7798));
  OA21x2_ASAP7_75t_L        g07542(.A1(new_n7791), .A2(new_n7795), .B(new_n7797), .Y(new_n7799));
  NOR2xp33_ASAP7_75t_L      g07543(.A(new_n5855), .B(new_n513), .Y(new_n7800));
  AOI221xp5_ASAP7_75t_L     g07544(.A1(\b[39] ), .A2(new_n560), .B1(\b[41] ), .B2(new_n475), .C(new_n7800), .Y(new_n7801));
  O2A1O1Ixp33_ASAP7_75t_L   g07545(.A1(new_n477), .A2(new_n6117), .B(new_n7801), .C(new_n466), .Y(new_n7802));
  INVx1_ASAP7_75t_L         g07546(.A(new_n7801), .Y(new_n7803));
  A2O1A1Ixp33_ASAP7_75t_L   g07547(.A1(new_n6118), .A2(new_n483), .B(new_n7803), .C(new_n466), .Y(new_n7804));
  OAI21xp33_ASAP7_75t_L     g07548(.A1(new_n466), .A2(new_n7802), .B(new_n7804), .Y(new_n7805));
  INVx1_ASAP7_75t_L         g07549(.A(new_n7805), .Y(new_n7806));
  NOR3xp33_ASAP7_75t_L      g07550(.A(new_n7799), .B(new_n7806), .C(new_n7798), .Y(new_n7807));
  INVx1_ASAP7_75t_L         g07551(.A(new_n7796), .Y(new_n7808));
  NAND2xp33_ASAP7_75t_L     g07552(.A(\a[11] ), .B(new_n7499), .Y(new_n7809));
  O2A1O1Ixp33_ASAP7_75t_L   g07553(.A1(new_n641), .A2(new_n5083), .B(new_n7497), .C(\a[11] ), .Y(new_n7810));
  A2O1A1Ixp33_ASAP7_75t_L   g07554(.A1(\a[11] ), .A2(new_n7809), .B(new_n7810), .C(new_n7808), .Y(new_n7811));
  NAND3xp33_ASAP7_75t_L     g07555(.A(new_n7792), .B(new_n7794), .C(new_n7793), .Y(new_n7812));
  OAI21xp33_ASAP7_75t_L     g07556(.A1(new_n7784), .A2(new_n7787), .B(new_n7790), .Y(new_n7813));
  NAND4xp25_ASAP7_75t_L     g07557(.A(new_n7533), .B(new_n7812), .C(new_n7813), .D(new_n7811), .Y(new_n7814));
  OAI21xp33_ASAP7_75t_L     g07558(.A1(new_n7791), .A2(new_n7795), .B(new_n7797), .Y(new_n7815));
  AOI21xp33_ASAP7_75t_L     g07559(.A1(new_n7814), .A2(new_n7815), .B(new_n7805), .Y(new_n7816));
  OAI22xp33_ASAP7_75t_L     g07560(.A1(new_n7566), .A2(new_n7517), .B1(new_n7816), .B2(new_n7807), .Y(new_n7817));
  NAND3xp33_ASAP7_75t_L     g07561(.A(new_n7814), .B(new_n7815), .C(new_n7805), .Y(new_n7818));
  OAI21xp33_ASAP7_75t_L     g07562(.A1(new_n7798), .A2(new_n7799), .B(new_n7806), .Y(new_n7819));
  NAND3xp33_ASAP7_75t_L     g07563(.A(new_n7520), .B(new_n7818), .C(new_n7819), .Y(new_n7820));
  NOR2xp33_ASAP7_75t_L      g07564(.A(new_n6378), .B(new_n375), .Y(new_n7821));
  AOI221xp5_ASAP7_75t_L     g07565(.A1(\b[44] ), .A2(new_n361), .B1(new_n349), .B2(\b[43] ), .C(new_n7821), .Y(new_n7822));
  O2A1O1Ixp33_ASAP7_75t_L   g07566(.A1(new_n356), .A2(new_n6951), .B(new_n7822), .C(new_n346), .Y(new_n7823));
  INVx1_ASAP7_75t_L         g07567(.A(new_n6951), .Y(new_n7824));
  INVx1_ASAP7_75t_L         g07568(.A(new_n7822), .Y(new_n7825));
  A2O1A1Ixp33_ASAP7_75t_L   g07569(.A1(new_n7824), .A2(new_n359), .B(new_n7825), .C(new_n346), .Y(new_n7826));
  OAI21xp33_ASAP7_75t_L     g07570(.A1(new_n346), .A2(new_n7823), .B(new_n7826), .Y(new_n7827));
  INVx1_ASAP7_75t_L         g07571(.A(new_n7827), .Y(new_n7828));
  NAND3xp33_ASAP7_75t_L     g07572(.A(new_n7817), .B(new_n7820), .C(new_n7828), .Y(new_n7829));
  A2O1A1Ixp33_ASAP7_75t_L   g07573(.A1(new_n7216), .A2(new_n7218), .B(new_n7515), .C(new_n7514), .Y(new_n7830));
  AOI22xp33_ASAP7_75t_L     g07574(.A1(new_n7818), .A2(new_n7819), .B1(new_n7518), .B2(new_n7830), .Y(new_n7831));
  AND4x1_ASAP7_75t_L        g07575(.A(new_n7830), .B(new_n7518), .C(new_n7819), .D(new_n7818), .Y(new_n7832));
  OAI21xp33_ASAP7_75t_L     g07576(.A1(new_n7831), .A2(new_n7832), .B(new_n7827), .Y(new_n7833));
  NAND2xp33_ASAP7_75t_L     g07577(.A(new_n7833), .B(new_n7829), .Y(new_n7834));
  O2A1O1Ixp33_ASAP7_75t_L   g07578(.A1(new_n7568), .A2(new_n7539), .B(new_n7565), .C(new_n7834), .Y(new_n7835));
  INVx1_ASAP7_75t_L         g07579(.A(new_n7565), .Y(new_n7836));
  A2O1A1Ixp33_ASAP7_75t_L   g07580(.A1(new_n7225), .A2(new_n7226), .B(new_n7241), .C(new_n7238), .Y(new_n7837));
  AOI221xp5_ASAP7_75t_L     g07581(.A1(new_n7833), .A2(new_n7829), .B1(new_n7538), .B2(new_n7837), .C(new_n7836), .Y(new_n7838));
  NOR3xp33_ASAP7_75t_L      g07582(.A(new_n7835), .B(new_n7564), .C(new_n7838), .Y(new_n7839));
  NOR3xp33_ASAP7_75t_L      g07583(.A(new_n7832), .B(new_n7827), .C(new_n7831), .Y(new_n7840));
  AOI21xp33_ASAP7_75t_L     g07584(.A1(new_n7817), .A2(new_n7820), .B(new_n7828), .Y(new_n7841));
  NOR2xp33_ASAP7_75t_L      g07585(.A(new_n7840), .B(new_n7841), .Y(new_n7842));
  A2O1A1Ixp33_ASAP7_75t_L   g07586(.A1(new_n7538), .A2(new_n7837), .B(new_n7836), .C(new_n7842), .Y(new_n7843));
  OAI221xp5_ASAP7_75t_L     g07587(.A1(new_n7840), .A2(new_n7841), .B1(new_n7539), .B2(new_n7568), .C(new_n7565), .Y(new_n7844));
  NAND3xp33_ASAP7_75t_L     g07588(.A(new_n7843), .B(new_n7844), .C(new_n7564), .Y(new_n7845));
  AOI21xp33_ASAP7_75t_L     g07589(.A1(new_n7281), .A2(\a[2] ), .B(new_n7282), .Y(new_n7846));
  MAJIxp5_ASAP7_75t_L       g07590(.A(new_n7546), .B(new_n7540), .C(new_n7846), .Y(new_n7847));
  INVx1_ASAP7_75t_L         g07591(.A(new_n7847), .Y(new_n7848));
  O2A1O1Ixp33_ASAP7_75t_L   g07592(.A1(new_n7564), .A2(new_n7839), .B(new_n7845), .C(new_n7848), .Y(new_n7849));
  INVx1_ASAP7_75t_L         g07593(.A(new_n7564), .Y(new_n7850));
  OAI21xp33_ASAP7_75t_L     g07594(.A1(new_n7838), .A2(new_n7835), .B(new_n7850), .Y(new_n7851));
  NAND2xp33_ASAP7_75t_L     g07595(.A(new_n7851), .B(new_n7845), .Y(new_n7852));
  NOR2xp33_ASAP7_75t_L      g07596(.A(new_n7852), .B(new_n7847), .Y(new_n7853));
  NOR2xp33_ASAP7_75t_L      g07597(.A(new_n7853), .B(new_n7849), .Y(\f[47] ));
  AO21x2_ASAP7_75t_L        g07598(.A1(new_n7852), .A2(new_n7847), .B(new_n7839), .Y(new_n7855));
  NOR2xp33_ASAP7_75t_L      g07599(.A(new_n7270), .B(new_n287), .Y(new_n7856));
  AOI221xp5_ASAP7_75t_L     g07600(.A1(\b[47] ), .A2(new_n264), .B1(\b[48] ), .B2(new_n283), .C(new_n7856), .Y(new_n7857));
  INVx1_ASAP7_75t_L         g07601(.A(new_n7553), .Y(new_n7858));
  NOR2xp33_ASAP7_75t_L      g07602(.A(\b[47] ), .B(\b[48] ), .Y(new_n7859));
  INVx1_ASAP7_75t_L         g07603(.A(\b[48] ), .Y(new_n7860));
  NOR2xp33_ASAP7_75t_L      g07604(.A(new_n7552), .B(new_n7860), .Y(new_n7861));
  NOR2xp33_ASAP7_75t_L      g07605(.A(new_n7859), .B(new_n7861), .Y(new_n7862));
  INVx1_ASAP7_75t_L         g07606(.A(new_n7862), .Y(new_n7863));
  O2A1O1Ixp33_ASAP7_75t_L   g07607(.A1(new_n7555), .A2(new_n7558), .B(new_n7858), .C(new_n7863), .Y(new_n7864));
  INVx1_ASAP7_75t_L         g07608(.A(new_n7864), .Y(new_n7865));
  A2O1A1O1Ixp25_ASAP7_75t_L g07609(.A1(new_n7272), .A2(new_n7276), .B(new_n7271), .C(new_n7554), .D(new_n7553), .Y(new_n7866));
  NAND2xp33_ASAP7_75t_L     g07610(.A(new_n7863), .B(new_n7866), .Y(new_n7867));
  NAND2xp33_ASAP7_75t_L     g07611(.A(new_n7865), .B(new_n7867), .Y(new_n7868));
  O2A1O1Ixp33_ASAP7_75t_L   g07612(.A1(new_n279), .A2(new_n7868), .B(new_n7857), .C(new_n257), .Y(new_n7869));
  OAI21xp33_ASAP7_75t_L     g07613(.A1(new_n279), .A2(new_n7868), .B(new_n7857), .Y(new_n7870));
  NAND2xp33_ASAP7_75t_L     g07614(.A(new_n257), .B(new_n7870), .Y(new_n7871));
  OAI21xp33_ASAP7_75t_L     g07615(.A1(new_n257), .A2(new_n7869), .B(new_n7871), .Y(new_n7872));
  A2O1A1Ixp33_ASAP7_75t_L   g07616(.A1(new_n7830), .A2(new_n7518), .B(new_n7816), .C(new_n7818), .Y(new_n7873));
  NAND2xp33_ASAP7_75t_L     g07617(.A(new_n7769), .B(new_n7762), .Y(new_n7874));
  O2A1O1Ixp33_ASAP7_75t_L   g07618(.A1(new_n872), .A2(new_n4589), .B(new_n7771), .C(new_n867), .Y(new_n7875));
  O2A1O1Ixp33_ASAP7_75t_L   g07619(.A1(new_n7875), .A2(new_n867), .B(new_n7775), .C(new_n7874), .Y(new_n7876));
  NOR3xp33_ASAP7_75t_L      g07620(.A(new_n7777), .B(new_n7778), .C(new_n7779), .Y(new_n7877));
  O2A1O1Ixp33_ASAP7_75t_L   g07621(.A1(new_n7877), .A2(new_n7779), .B(new_n7783), .C(new_n7876), .Y(new_n7878));
  A2O1A1O1Ixp25_ASAP7_75t_L g07622(.A1(new_n7469), .A2(new_n7283), .B(new_n7765), .C(new_n7758), .D(new_n7768), .Y(new_n7879));
  INVx1_ASAP7_75t_L         g07623(.A(new_n7719), .Y(new_n7880));
  INVx1_ASAP7_75t_L         g07624(.A(new_n7586), .Y(new_n7881));
  AO22x1_ASAP7_75t_L        g07625(.A1(new_n7686), .A2(new_n7682), .B1(new_n7881), .B2(new_n7404), .Y(new_n7882));
  A2O1A1Ixp33_ASAP7_75t_L   g07626(.A1(new_n7673), .A2(new_n7662), .B(new_n7595), .C(new_n7669), .Y(new_n7883));
  NOR2xp33_ASAP7_75t_L      g07627(.A(new_n960), .B(new_n4142), .Y(new_n7884));
  AOI221xp5_ASAP7_75t_L     g07628(.A1(\b[13] ), .A2(new_n4402), .B1(\b[15] ), .B2(new_n4156), .C(new_n7884), .Y(new_n7885));
  INVx1_ASAP7_75t_L         g07629(.A(new_n7885), .Y(new_n7886));
  A2O1A1Ixp33_ASAP7_75t_L   g07630(.A1(new_n1052), .A2(new_n4151), .B(new_n7886), .C(\a[35] ), .Y(new_n7887));
  O2A1O1Ixp33_ASAP7_75t_L   g07631(.A1(new_n4150), .A2(new_n1774), .B(new_n7885), .C(\a[35] ), .Y(new_n7888));
  AOI21xp33_ASAP7_75t_L     g07632(.A1(new_n7887), .A2(\a[35] ), .B(new_n7888), .Y(new_n7889));
  A2O1A1Ixp33_ASAP7_75t_L   g07633(.A1(new_n7049), .A2(new_n7052), .B(new_n7051), .C(new_n7366), .Y(new_n7890));
  A2O1A1Ixp33_ASAP7_75t_L   g07634(.A1(new_n7890), .A2(new_n7365), .B(new_n7659), .C(new_n7655), .Y(new_n7891));
  NOR2xp33_ASAP7_75t_L      g07635(.A(new_n748), .B(new_n4903), .Y(new_n7892));
  AOI221xp5_ASAP7_75t_L     g07636(.A1(\b[10] ), .A2(new_n5139), .B1(\b[12] ), .B2(new_n4917), .C(new_n7892), .Y(new_n7893));
  O2A1O1Ixp33_ASAP7_75t_L   g07637(.A1(new_n4911), .A2(new_n841), .B(new_n7893), .C(new_n4906), .Y(new_n7894));
  O2A1O1Ixp33_ASAP7_75t_L   g07638(.A1(new_n4911), .A2(new_n841), .B(new_n7893), .C(\a[38] ), .Y(new_n7895));
  INVx1_ASAP7_75t_L         g07639(.A(new_n7895), .Y(new_n7896));
  OAI21xp33_ASAP7_75t_L     g07640(.A1(new_n4906), .A2(new_n7894), .B(new_n7896), .Y(new_n7897));
  INVx1_ASAP7_75t_L         g07641(.A(new_n7652), .Y(new_n7898));
  NAND2xp33_ASAP7_75t_L     g07642(.A(new_n7619), .B(new_n7618), .Y(new_n7899));
  O2A1O1Ixp33_ASAP7_75t_L   g07643(.A1(new_n728), .A2(new_n6443), .B(new_n7621), .C(new_n6439), .Y(new_n7900));
  O2A1O1Ixp33_ASAP7_75t_L   g07644(.A1(new_n7900), .A2(new_n6439), .B(new_n7625), .C(new_n7899), .Y(new_n7901));
  INVx1_ASAP7_75t_L         g07645(.A(new_n7901), .Y(new_n7902));
  INVx1_ASAP7_75t_L         g07646(.A(\a[48] ), .Y(new_n7903));
  NAND2xp33_ASAP7_75t_L     g07647(.A(\a[47] ), .B(new_n7903), .Y(new_n7904));
  NAND2xp33_ASAP7_75t_L     g07648(.A(\a[48] ), .B(new_n7316), .Y(new_n7905));
  AND2x2_ASAP7_75t_L        g07649(.A(new_n7904), .B(new_n7905), .Y(new_n7906));
  NOR2xp33_ASAP7_75t_L      g07650(.A(new_n284), .B(new_n7906), .Y(new_n7907));
  A2O1A1Ixp33_ASAP7_75t_L   g07651(.A1(new_n7617), .A2(new_n7613), .B(new_n7324), .C(new_n7907), .Y(new_n7908));
  OAI21xp33_ASAP7_75t_L     g07652(.A1(new_n7321), .A2(new_n274), .B(new_n7335), .Y(new_n7909));
  NOR5xp2_ASAP7_75t_L       g07653(.A(new_n7909), .B(new_n7616), .C(new_n7611), .D(new_n7001), .E(new_n7316), .Y(new_n7910));
  A2O1A1Ixp33_ASAP7_75t_L   g07654(.A1(new_n7904), .A2(new_n7905), .B(new_n284), .C(new_n7910), .Y(new_n7911));
  NAND2xp33_ASAP7_75t_L     g07655(.A(\b[3] ), .B(new_n7334), .Y(new_n7912));
  NAND2xp33_ASAP7_75t_L     g07656(.A(\b[1] ), .B(new_n7609), .Y(new_n7913));
  NAND2xp33_ASAP7_75t_L     g07657(.A(\b[2] ), .B(new_n7333), .Y(new_n7914));
  NAND2xp33_ASAP7_75t_L     g07658(.A(new_n7322), .B(new_n312), .Y(new_n7915));
  NAND5xp2_ASAP7_75t_L      g07659(.A(new_n7915), .B(new_n7914), .C(new_n7913), .D(new_n7912), .E(\a[47] ), .Y(new_n7916));
  NAND3xp33_ASAP7_75t_L     g07660(.A(new_n7913), .B(new_n7912), .C(new_n7914), .Y(new_n7917));
  A2O1A1Ixp33_ASAP7_75t_L   g07661(.A1(new_n312), .A2(new_n7322), .B(new_n7917), .C(new_n7316), .Y(new_n7918));
  AND2x2_ASAP7_75t_L        g07662(.A(new_n7916), .B(new_n7918), .Y(new_n7919));
  AO21x2_ASAP7_75t_L        g07663(.A1(new_n7908), .A2(new_n7911), .B(new_n7919), .Y(new_n7920));
  NAND3xp33_ASAP7_75t_L     g07664(.A(new_n7911), .B(new_n7908), .C(new_n7919), .Y(new_n7921));
  NAND2xp33_ASAP7_75t_L     g07665(.A(\b[6] ), .B(new_n6442), .Y(new_n7922));
  OAI221xp5_ASAP7_75t_L     g07666(.A1(new_n7304), .A2(new_n384), .B1(new_n332), .B2(new_n6741), .C(new_n7922), .Y(new_n7923));
  A2O1A1Ixp33_ASAP7_75t_L   g07667(.A1(new_n5363), .A2(new_n6450), .B(new_n7923), .C(\a[44] ), .Y(new_n7924));
  AOI211xp5_ASAP7_75t_L     g07668(.A1(new_n5363), .A2(new_n6450), .B(new_n7923), .C(new_n6439), .Y(new_n7925));
  A2O1A1O1Ixp25_ASAP7_75t_L g07669(.A1(new_n6450), .A2(new_n5363), .B(new_n7923), .C(new_n7924), .D(new_n7925), .Y(new_n7926));
  NAND3xp33_ASAP7_75t_L     g07670(.A(new_n7920), .B(new_n7921), .C(new_n7926), .Y(new_n7927));
  AOI21xp33_ASAP7_75t_L     g07671(.A1(new_n7911), .A2(new_n7908), .B(new_n7919), .Y(new_n7928));
  AND3x1_ASAP7_75t_L        g07672(.A(new_n7911), .B(new_n7919), .C(new_n7908), .Y(new_n7929));
  INVx1_ASAP7_75t_L         g07673(.A(new_n7926), .Y(new_n7930));
  OAI21xp33_ASAP7_75t_L     g07674(.A1(new_n7928), .A2(new_n7929), .B(new_n7930), .Y(new_n7931));
  AND4x1_ASAP7_75t_L        g07675(.A(new_n7628), .B(new_n7902), .C(new_n7931), .D(new_n7927), .Y(new_n7932));
  A2O1A1Ixp33_ASAP7_75t_L   g07676(.A1(new_n7622), .A2(new_n7621), .B(new_n7900), .C(new_n7623), .Y(new_n7933));
  O2A1O1Ixp33_ASAP7_75t_L   g07677(.A1(new_n7626), .A2(new_n7933), .B(new_n7607), .C(new_n7901), .Y(new_n7934));
  AOI21xp33_ASAP7_75t_L     g07678(.A1(new_n7931), .A2(new_n7927), .B(new_n7934), .Y(new_n7935));
  NOR2xp33_ASAP7_75t_L      g07679(.A(new_n534), .B(new_n5640), .Y(new_n7936));
  AOI221xp5_ASAP7_75t_L     g07680(.A1(\b[7] ), .A2(new_n5920), .B1(\b[9] ), .B2(new_n5629), .C(new_n7936), .Y(new_n7937));
  INVx1_ASAP7_75t_L         g07681(.A(new_n7937), .Y(new_n7938));
  A2O1A1Ixp33_ASAP7_75t_L   g07682(.A1(new_n602), .A2(new_n5637), .B(new_n7938), .C(\a[41] ), .Y(new_n7939));
  O2A1O1Ixp33_ASAP7_75t_L   g07683(.A1(new_n5630), .A2(new_n1066), .B(new_n7937), .C(\a[41] ), .Y(new_n7940));
  AOI21xp33_ASAP7_75t_L     g07684(.A1(new_n7939), .A2(\a[41] ), .B(new_n7940), .Y(new_n7941));
  OAI21xp33_ASAP7_75t_L     g07685(.A1(new_n7935), .A2(new_n7932), .B(new_n7941), .Y(new_n7942));
  NAND3xp33_ASAP7_75t_L     g07686(.A(new_n7934), .B(new_n7931), .C(new_n7927), .Y(new_n7943));
  AO22x1_ASAP7_75t_L        g07687(.A1(new_n7927), .A2(new_n7931), .B1(new_n7902), .B2(new_n7628), .Y(new_n7944));
  AO21x2_ASAP7_75t_L        g07688(.A1(\a[41] ), .A2(new_n7939), .B(new_n7940), .Y(new_n7945));
  NAND3xp33_ASAP7_75t_L     g07689(.A(new_n7944), .B(new_n7943), .C(new_n7945), .Y(new_n7946));
  NAND2xp33_ASAP7_75t_L     g07690(.A(new_n7942), .B(new_n7946), .Y(new_n7947));
  O2A1O1Ixp33_ASAP7_75t_L   g07691(.A1(new_n7599), .A2(new_n7898), .B(new_n7640), .C(new_n7947), .Y(new_n7948));
  AOI221xp5_ASAP7_75t_L     g07692(.A1(new_n7942), .A2(new_n7946), .B1(new_n7652), .B2(new_n7657), .C(new_n7633), .Y(new_n7949));
  OAI21xp33_ASAP7_75t_L     g07693(.A1(new_n7949), .A2(new_n7948), .B(new_n7897), .Y(new_n7950));
  INVx1_ASAP7_75t_L         g07694(.A(new_n7894), .Y(new_n7951));
  AOI21xp33_ASAP7_75t_L     g07695(.A1(new_n7951), .A2(\a[38] ), .B(new_n7895), .Y(new_n7952));
  AOI21xp33_ASAP7_75t_L     g07696(.A1(new_n7944), .A2(new_n7943), .B(new_n7945), .Y(new_n7953));
  NOR3xp33_ASAP7_75t_L      g07697(.A(new_n7932), .B(new_n7935), .C(new_n7941), .Y(new_n7954));
  NOR2xp33_ASAP7_75t_L      g07698(.A(new_n7954), .B(new_n7953), .Y(new_n7955));
  A2O1A1Ixp33_ASAP7_75t_L   g07699(.A1(new_n7652), .A2(new_n7657), .B(new_n7633), .C(new_n7955), .Y(new_n7956));
  A2O1A1O1Ixp25_ASAP7_75t_L g07700(.A1(new_n7357), .A2(new_n7359), .B(new_n7598), .C(new_n7652), .D(new_n7633), .Y(new_n7957));
  NAND2xp33_ASAP7_75t_L     g07701(.A(new_n7947), .B(new_n7957), .Y(new_n7958));
  NAND3xp33_ASAP7_75t_L     g07702(.A(new_n7958), .B(new_n7956), .C(new_n7952), .Y(new_n7959));
  NAND2xp33_ASAP7_75t_L     g07703(.A(new_n7950), .B(new_n7959), .Y(new_n7960));
  NOR3xp33_ASAP7_75t_L      g07704(.A(new_n7948), .B(new_n7949), .C(new_n7897), .Y(new_n7961));
  AOI211xp5_ASAP7_75t_L     g07705(.A1(new_n7593), .A2(new_n7650), .B(new_n7660), .C(new_n7961), .Y(new_n7962));
  AOI221xp5_ASAP7_75t_L     g07706(.A1(new_n7891), .A2(new_n7960), .B1(new_n7950), .B2(new_n7962), .C(new_n7889), .Y(new_n7963));
  O2A1O1Ixp33_ASAP7_75t_L   g07707(.A1(new_n4150), .A2(new_n1774), .B(new_n7885), .C(new_n4145), .Y(new_n7964));
  A2O1A1Ixp33_ASAP7_75t_L   g07708(.A1(new_n1052), .A2(new_n4151), .B(new_n7886), .C(new_n4145), .Y(new_n7965));
  OAI21xp33_ASAP7_75t_L     g07709(.A1(new_n4145), .A2(new_n7964), .B(new_n7965), .Y(new_n7966));
  AOI21xp33_ASAP7_75t_L     g07710(.A1(new_n7958), .A2(new_n7956), .B(new_n7952), .Y(new_n7967));
  OAI21xp33_ASAP7_75t_L     g07711(.A1(new_n7967), .A2(new_n7961), .B(new_n7891), .Y(new_n7968));
  OAI211xp5_ASAP7_75t_L     g07712(.A1(new_n7377), .A2(new_n7659), .B(new_n7959), .C(new_n7655), .Y(new_n7969));
  O2A1O1Ixp33_ASAP7_75t_L   g07713(.A1(new_n7967), .A2(new_n7969), .B(new_n7968), .C(new_n7966), .Y(new_n7970));
  NOR2xp33_ASAP7_75t_L      g07714(.A(new_n7970), .B(new_n7963), .Y(new_n7971));
  XOR2x2_ASAP7_75t_L        g07715(.A(new_n7883), .B(new_n7971), .Y(new_n7972));
  NAND2xp33_ASAP7_75t_L     g07716(.A(new_n7883), .B(new_n7971), .Y(new_n7973));
  AND2x2_ASAP7_75t_L        g07717(.A(new_n7679), .B(new_n7673), .Y(new_n7974));
  OAI221xp5_ASAP7_75t_L     g07718(.A1(new_n7963), .A2(new_n7970), .B1(new_n7595), .B2(new_n7974), .C(new_n7669), .Y(new_n7975));
  NOR2xp33_ASAP7_75t_L      g07719(.A(new_n1349), .B(new_n3509), .Y(new_n7976));
  AOI221xp5_ASAP7_75t_L     g07720(.A1(\b[16] ), .A2(new_n3708), .B1(\b[18] ), .B2(new_n3503), .C(new_n7976), .Y(new_n7977));
  O2A1O1Ixp33_ASAP7_75t_L   g07721(.A1(new_n3513), .A2(new_n1464), .B(new_n7977), .C(new_n3493), .Y(new_n7978));
  INVx1_ASAP7_75t_L         g07722(.A(new_n7977), .Y(new_n7979));
  A2O1A1Ixp33_ASAP7_75t_L   g07723(.A1(new_n2329), .A2(new_n3505), .B(new_n7979), .C(new_n3493), .Y(new_n7980));
  OAI21xp33_ASAP7_75t_L     g07724(.A1(new_n3493), .A2(new_n7978), .B(new_n7980), .Y(new_n7981));
  NAND3xp33_ASAP7_75t_L     g07725(.A(new_n7973), .B(new_n7975), .C(new_n7981), .Y(new_n7982));
  INVx1_ASAP7_75t_L         g07726(.A(new_n7981), .Y(new_n7983));
  AOI21xp33_ASAP7_75t_L     g07727(.A1(new_n7973), .A2(new_n7975), .B(new_n7983), .Y(new_n7984));
  AOI21xp33_ASAP7_75t_L     g07728(.A1(new_n7982), .A2(new_n7972), .B(new_n7984), .Y(new_n7985));
  NAND3xp33_ASAP7_75t_L     g07729(.A(new_n7985), .B(new_n7882), .C(new_n7688), .Y(new_n7986));
  AND3x1_ASAP7_75t_L        g07730(.A(new_n7983), .B(new_n7973), .C(new_n7975), .Y(new_n7987));
  A2O1A1Ixp33_ASAP7_75t_L   g07731(.A1(new_n7686), .A2(new_n7683), .B(new_n7587), .C(new_n7688), .Y(new_n7988));
  OAI21xp33_ASAP7_75t_L     g07732(.A1(new_n7987), .A2(new_n7984), .B(new_n7988), .Y(new_n7989));
  NAND2xp33_ASAP7_75t_L     g07733(.A(\b[20] ), .B(new_n2936), .Y(new_n7990));
  OAI221xp5_ASAP7_75t_L     g07734(.A1(new_n2930), .A2(new_n1895), .B1(new_n1599), .B2(new_n3133), .C(new_n7990), .Y(new_n7991));
  A2O1A1Ixp33_ASAP7_75t_L   g07735(.A1(new_n2836), .A2(new_n2932), .B(new_n7991), .C(\a[29] ), .Y(new_n7992));
  AOI211xp5_ASAP7_75t_L     g07736(.A1(new_n2836), .A2(new_n2932), .B(new_n7991), .C(new_n2928), .Y(new_n7993));
  A2O1A1O1Ixp25_ASAP7_75t_L g07737(.A1(new_n2932), .A2(new_n2836), .B(new_n7991), .C(new_n7992), .D(new_n7993), .Y(new_n7994));
  NAND3xp33_ASAP7_75t_L     g07738(.A(new_n7986), .B(new_n7989), .C(new_n7994), .Y(new_n7995));
  NOR3xp33_ASAP7_75t_L      g07739(.A(new_n7988), .B(new_n7984), .C(new_n7987), .Y(new_n7996));
  NOR2xp33_ASAP7_75t_L      g07740(.A(new_n7698), .B(new_n7689), .Y(new_n7997));
  O2A1O1Ixp33_ASAP7_75t_L   g07741(.A1(new_n7587), .A2(new_n7997), .B(new_n7688), .C(new_n7985), .Y(new_n7998));
  INVx1_ASAP7_75t_L         g07742(.A(new_n7994), .Y(new_n7999));
  OAI21xp33_ASAP7_75t_L     g07743(.A1(new_n7996), .A2(new_n7998), .B(new_n7999), .Y(new_n8000));
  AND4x1_ASAP7_75t_L        g07744(.A(new_n7707), .B(new_n7880), .C(new_n8000), .D(new_n7995), .Y(new_n8001));
  O2A1O1Ixp33_ASAP7_75t_L   g07745(.A1(new_n7697), .A2(new_n7696), .B(new_n7705), .C(new_n7719), .Y(new_n8002));
  AOI21xp33_ASAP7_75t_L     g07746(.A1(new_n8000), .A2(new_n7995), .B(new_n8002), .Y(new_n8003));
  NOR2xp33_ASAP7_75t_L      g07747(.A(new_n2205), .B(new_n2415), .Y(new_n8004));
  AOI221xp5_ASAP7_75t_L     g07748(.A1(\b[22] ), .A2(new_n2577), .B1(\b[23] ), .B2(new_n2421), .C(new_n8004), .Y(new_n8005));
  OA21x2_ASAP7_75t_L        g07749(.A1(new_n2425), .A2(new_n2853), .B(new_n8005), .Y(new_n8006));
  O2A1O1Ixp33_ASAP7_75t_L   g07750(.A1(new_n2425), .A2(new_n2853), .B(new_n8005), .C(new_n2413), .Y(new_n8007));
  NAND2xp33_ASAP7_75t_L     g07751(.A(\a[26] ), .B(new_n8006), .Y(new_n8008));
  OA21x2_ASAP7_75t_L        g07752(.A1(new_n8006), .A2(new_n8007), .B(new_n8008), .Y(new_n8009));
  OAI21xp33_ASAP7_75t_L     g07753(.A1(new_n8003), .A2(new_n8001), .B(new_n8009), .Y(new_n8010));
  NAND3xp33_ASAP7_75t_L     g07754(.A(new_n8002), .B(new_n8000), .C(new_n7995), .Y(new_n8011));
  NOR3xp33_ASAP7_75t_L      g07755(.A(new_n7999), .B(new_n7998), .C(new_n7996), .Y(new_n8012));
  AOI21xp33_ASAP7_75t_L     g07756(.A1(new_n7986), .A2(new_n7989), .B(new_n7994), .Y(new_n8013));
  NOR2xp33_ASAP7_75t_L      g07757(.A(new_n7699), .B(new_n7701), .Y(new_n8014));
  MAJIxp5_ASAP7_75t_L       g07758(.A(new_n7723), .B(new_n8014), .C(new_n7702), .Y(new_n8015));
  OAI21xp33_ASAP7_75t_L     g07759(.A1(new_n8012), .A2(new_n8013), .B(new_n8015), .Y(new_n8016));
  NAND2xp33_ASAP7_75t_L     g07760(.A(new_n2417), .B(new_n2216), .Y(new_n8017));
  A2O1A1Ixp33_ASAP7_75t_L   g07761(.A1(new_n8017), .A2(new_n8005), .B(new_n8007), .C(new_n8008), .Y(new_n8018));
  NAND3xp33_ASAP7_75t_L     g07762(.A(new_n8016), .B(new_n8011), .C(new_n8018), .Y(new_n8019));
  OAI211xp5_ASAP7_75t_L     g07763(.A1(new_n7728), .A2(new_n7738), .B(new_n8010), .C(new_n8019), .Y(new_n8020));
  NAND2xp33_ASAP7_75t_L     g07764(.A(new_n8019), .B(new_n8010), .Y(new_n8021));
  NAND2xp33_ASAP7_75t_L     g07765(.A(new_n7729), .B(new_n8021), .Y(new_n8022));
  NOR2xp33_ASAP7_75t_L      g07766(.A(new_n2703), .B(new_n1962), .Y(new_n8023));
  AOI221xp5_ASAP7_75t_L     g07767(.A1(new_n1955), .A2(\b[27] ), .B1(new_n2093), .B2(\b[25] ), .C(new_n8023), .Y(new_n8024));
  INVx1_ASAP7_75t_L         g07768(.A(new_n8024), .Y(new_n8025));
  A2O1A1Ixp33_ASAP7_75t_L   g07769(.A1(new_n2887), .A2(new_n1964), .B(new_n8025), .C(\a[23] ), .Y(new_n8026));
  O2A1O1Ixp33_ASAP7_75t_L   g07770(.A1(new_n1956), .A2(new_n2889), .B(new_n8024), .C(\a[23] ), .Y(new_n8027));
  AOI21xp33_ASAP7_75t_L     g07771(.A1(new_n8026), .A2(\a[23] ), .B(new_n8027), .Y(new_n8028));
  NAND3xp33_ASAP7_75t_L     g07772(.A(new_n8022), .B(new_n8020), .C(new_n8028), .Y(new_n8029));
  NOR2xp33_ASAP7_75t_L      g07773(.A(new_n7729), .B(new_n8021), .Y(new_n8030));
  AOI211xp5_ASAP7_75t_L     g07774(.A1(new_n8019), .A2(new_n8010), .B(new_n7728), .C(new_n7738), .Y(new_n8031));
  O2A1O1Ixp33_ASAP7_75t_L   g07775(.A1(new_n1956), .A2(new_n2889), .B(new_n8024), .C(new_n1952), .Y(new_n8032));
  INVx1_ASAP7_75t_L         g07776(.A(new_n8027), .Y(new_n8033));
  OAI21xp33_ASAP7_75t_L     g07777(.A1(new_n1952), .A2(new_n8032), .B(new_n8033), .Y(new_n8034));
  OAI21xp33_ASAP7_75t_L     g07778(.A1(new_n8031), .A2(new_n8030), .B(new_n8034), .Y(new_n8035));
  NAND2xp33_ASAP7_75t_L     g07779(.A(new_n8029), .B(new_n8035), .Y(new_n8036));
  O2A1O1Ixp33_ASAP7_75t_L   g07780(.A1(new_n7585), .A2(new_n7736), .B(new_n7746), .C(new_n8036), .Y(new_n8037));
  OAI21xp33_ASAP7_75t_L     g07781(.A1(new_n7736), .A2(new_n7585), .B(new_n7746), .Y(new_n8038));
  NAND3xp33_ASAP7_75t_L     g07782(.A(new_n8022), .B(new_n8020), .C(new_n8034), .Y(new_n8039));
  INVx1_ASAP7_75t_L         g07783(.A(new_n8039), .Y(new_n8040));
  O2A1O1Ixp33_ASAP7_75t_L   g07784(.A1(new_n8028), .A2(new_n8040), .B(new_n8029), .C(new_n8038), .Y(new_n8041));
  NOR2xp33_ASAP7_75t_L      g07785(.A(new_n3456), .B(new_n1518), .Y(new_n8042));
  AOI221xp5_ASAP7_75t_L     g07786(.A1(\b[28] ), .A2(new_n1659), .B1(\b[29] ), .B2(new_n1507), .C(new_n8042), .Y(new_n8043));
  NAND2xp33_ASAP7_75t_L     g07787(.A(new_n1513), .B(new_n4813), .Y(new_n8044));
  O2A1O1Ixp33_ASAP7_75t_L   g07788(.A1(new_n1521), .A2(new_n3464), .B(new_n8043), .C(new_n1501), .Y(new_n8045));
  OA21x2_ASAP7_75t_L        g07789(.A1(new_n1521), .A2(new_n3464), .B(new_n8043), .Y(new_n8046));
  NAND2xp33_ASAP7_75t_L     g07790(.A(\a[20] ), .B(new_n8046), .Y(new_n8047));
  A2O1A1Ixp33_ASAP7_75t_L   g07791(.A1(new_n8044), .A2(new_n8043), .B(new_n8045), .C(new_n8047), .Y(new_n8048));
  OAI21xp33_ASAP7_75t_L     g07792(.A1(new_n8041), .A2(new_n8037), .B(new_n8048), .Y(new_n8049));
  NAND3xp33_ASAP7_75t_L     g07793(.A(new_n8038), .B(new_n8029), .C(new_n8035), .Y(new_n8050));
  INVx1_ASAP7_75t_L         g07794(.A(new_n7454), .Y(new_n8051));
  NAND2xp33_ASAP7_75t_L     g07795(.A(new_n7438), .B(new_n7444), .Y(new_n8052));
  A2O1A1O1Ixp25_ASAP7_75t_L g07796(.A1(new_n7450), .A2(new_n8052), .B(new_n8051), .C(new_n7745), .D(new_n7740), .Y(new_n8053));
  NAND2xp33_ASAP7_75t_L     g07797(.A(new_n8053), .B(new_n8036), .Y(new_n8054));
  OA21x2_ASAP7_75t_L        g07798(.A1(new_n8046), .A2(new_n8045), .B(new_n8047), .Y(new_n8055));
  NAND3xp33_ASAP7_75t_L     g07799(.A(new_n8055), .B(new_n8050), .C(new_n8054), .Y(new_n8056));
  NAND2xp33_ASAP7_75t_L     g07800(.A(new_n8056), .B(new_n8049), .Y(new_n8057));
  O2A1O1Ixp33_ASAP7_75t_L   g07801(.A1(new_n7581), .A2(new_n7754), .B(new_n7753), .C(new_n8057), .Y(new_n8058));
  NOR3xp33_ASAP7_75t_L      g07802(.A(new_n7747), .B(new_n7584), .C(new_n7741), .Y(new_n8059));
  AOI221xp5_ASAP7_75t_L     g07803(.A1(new_n7756), .A2(new_n7748), .B1(new_n8049), .B2(new_n8056), .C(new_n8059), .Y(new_n8060));
  NOR2xp33_ASAP7_75t_L      g07804(.A(new_n4101), .B(new_n1284), .Y(new_n8061));
  AOI221xp5_ASAP7_75t_L     g07805(.A1(\b[31] ), .A2(new_n1290), .B1(\b[32] ), .B2(new_n1204), .C(new_n8061), .Y(new_n8062));
  NAND2xp33_ASAP7_75t_L     g07806(.A(new_n1216), .B(new_n4831), .Y(new_n8063));
  O2A1O1Ixp33_ASAP7_75t_L   g07807(.A1(new_n1210), .A2(new_n4108), .B(new_n8062), .C(new_n1206), .Y(new_n8064));
  OA21x2_ASAP7_75t_L        g07808(.A1(new_n1210), .A2(new_n4108), .B(new_n8062), .Y(new_n8065));
  NAND2xp33_ASAP7_75t_L     g07809(.A(\a[17] ), .B(new_n8065), .Y(new_n8066));
  A2O1A1Ixp33_ASAP7_75t_L   g07810(.A1(new_n8063), .A2(new_n8062), .B(new_n8064), .C(new_n8066), .Y(new_n8067));
  NOR3xp33_ASAP7_75t_L      g07811(.A(new_n8058), .B(new_n8060), .C(new_n8067), .Y(new_n8068));
  A2O1A1O1Ixp25_ASAP7_75t_L g07812(.A1(new_n7461), .A2(new_n7285), .B(new_n7472), .C(new_n7748), .D(new_n8059), .Y(new_n8069));
  AOI21xp33_ASAP7_75t_L     g07813(.A1(new_n8050), .A2(new_n8054), .B(new_n8055), .Y(new_n8070));
  NOR3xp33_ASAP7_75t_L      g07814(.A(new_n8037), .B(new_n8041), .C(new_n8048), .Y(new_n8071));
  OR3x1_ASAP7_75t_L         g07815(.A(new_n8069), .B(new_n8070), .C(new_n8071), .Y(new_n8072));
  NAND2xp33_ASAP7_75t_L     g07816(.A(new_n8069), .B(new_n8057), .Y(new_n8073));
  OA21x2_ASAP7_75t_L        g07817(.A1(new_n8065), .A2(new_n8064), .B(new_n8066), .Y(new_n8074));
  AOI21xp33_ASAP7_75t_L     g07818(.A1(new_n8072), .A2(new_n8073), .B(new_n8074), .Y(new_n8075));
  NOR3xp33_ASAP7_75t_L      g07819(.A(new_n7879), .B(new_n8075), .C(new_n8068), .Y(new_n8076));
  NAND3xp33_ASAP7_75t_L     g07820(.A(new_n8072), .B(new_n8073), .C(new_n8074), .Y(new_n8077));
  OAI21xp33_ASAP7_75t_L     g07821(.A1(new_n8060), .A2(new_n8058), .B(new_n8067), .Y(new_n8078));
  AOI221xp5_ASAP7_75t_L     g07822(.A1(new_n7572), .A2(new_n7758), .B1(new_n8077), .B2(new_n8078), .C(new_n7768), .Y(new_n8079));
  OAI22xp33_ASAP7_75t_L     g07823(.A1(new_n980), .A2(new_n4344), .B1(new_n4581), .B2(new_n864), .Y(new_n8080));
  AOI221xp5_ASAP7_75t_L     g07824(.A1(new_n886), .A2(\b[36] ), .B1(new_n873), .B2(new_n4621), .C(new_n8080), .Y(new_n8081));
  XNOR2x2_ASAP7_75t_L       g07825(.A(\a[14] ), .B(new_n8081), .Y(new_n8082));
  OAI21xp33_ASAP7_75t_L     g07826(.A1(new_n8076), .A2(new_n8079), .B(new_n8082), .Y(new_n8083));
  OAI21xp33_ASAP7_75t_L     g07827(.A1(new_n7767), .A2(new_n7766), .B(new_n7761), .Y(new_n8084));
  NAND3xp33_ASAP7_75t_L     g07828(.A(new_n8084), .B(new_n8077), .C(new_n8078), .Y(new_n8085));
  OAI21xp33_ASAP7_75t_L     g07829(.A1(new_n8068), .A2(new_n8075), .B(new_n7879), .Y(new_n8086));
  XNOR2x2_ASAP7_75t_L       g07830(.A(new_n867), .B(new_n8081), .Y(new_n8087));
  NAND3xp33_ASAP7_75t_L     g07831(.A(new_n8085), .B(new_n8086), .C(new_n8087), .Y(new_n8088));
  NAND2xp33_ASAP7_75t_L     g07832(.A(new_n8083), .B(new_n8088), .Y(new_n8089));
  NAND2xp33_ASAP7_75t_L     g07833(.A(new_n8089), .B(new_n7878), .Y(new_n8090));
  AOI21xp33_ASAP7_75t_L     g07834(.A1(new_n8085), .A2(new_n8086), .B(new_n8087), .Y(new_n8091));
  NOR3xp33_ASAP7_75t_L      g07835(.A(new_n8079), .B(new_n8076), .C(new_n8082), .Y(new_n8092));
  NOR2xp33_ASAP7_75t_L      g07836(.A(new_n8091), .B(new_n8092), .Y(new_n8093));
  OAI21xp33_ASAP7_75t_L     g07837(.A1(new_n7876), .A2(new_n7787), .B(new_n8093), .Y(new_n8094));
  NOR2xp33_ASAP7_75t_L      g07838(.A(new_n5311), .B(new_n1550), .Y(new_n8095));
  AOI221xp5_ASAP7_75t_L     g07839(.A1(\b[37] ), .A2(new_n713), .B1(\b[39] ), .B2(new_n640), .C(new_n8095), .Y(new_n8096));
  O2A1O1Ixp33_ASAP7_75t_L   g07840(.A1(new_n641), .A2(new_n5578), .B(new_n8096), .C(new_n637), .Y(new_n8097));
  INVx1_ASAP7_75t_L         g07841(.A(new_n8097), .Y(new_n8098));
  O2A1O1Ixp33_ASAP7_75t_L   g07842(.A1(new_n641), .A2(new_n5578), .B(new_n8096), .C(\a[11] ), .Y(new_n8099));
  AOI21xp33_ASAP7_75t_L     g07843(.A1(new_n8098), .A2(\a[11] ), .B(new_n8099), .Y(new_n8100));
  NAND3xp33_ASAP7_75t_L     g07844(.A(new_n8094), .B(new_n8090), .C(new_n8100), .Y(new_n8101));
  AOI221xp5_ASAP7_75t_L     g07845(.A1(new_n7781), .A2(new_n7783), .B1(new_n8088), .B2(new_n8083), .C(new_n7876), .Y(new_n8102));
  NOR2xp33_ASAP7_75t_L      g07846(.A(new_n8089), .B(new_n7878), .Y(new_n8103));
  AO21x2_ASAP7_75t_L        g07847(.A1(\a[11] ), .A2(new_n8098), .B(new_n8099), .Y(new_n8104));
  OAI21xp33_ASAP7_75t_L     g07848(.A1(new_n8102), .A2(new_n8103), .B(new_n8104), .Y(new_n8105));
  NOR2xp33_ASAP7_75t_L      g07849(.A(new_n7784), .B(new_n7787), .Y(new_n8106));
  MAJIxp5_ASAP7_75t_L       g07850(.A(new_n7797), .B(new_n7790), .C(new_n8106), .Y(new_n8107));
  NAND3xp33_ASAP7_75t_L     g07851(.A(new_n8107), .B(new_n8105), .C(new_n8101), .Y(new_n8108));
  NOR3xp33_ASAP7_75t_L      g07852(.A(new_n7787), .B(new_n7784), .C(new_n7794), .Y(new_n8109));
  NAND2xp33_ASAP7_75t_L     g07853(.A(new_n8105), .B(new_n8101), .Y(new_n8110));
  OAI21xp33_ASAP7_75t_L     g07854(.A1(new_n8109), .A2(new_n7799), .B(new_n8110), .Y(new_n8111));
  NOR2xp33_ASAP7_75t_L      g07855(.A(new_n5855), .B(new_n506), .Y(new_n8112));
  AOI221xp5_ASAP7_75t_L     g07856(.A1(\b[42] ), .A2(new_n475), .B1(new_n470), .B2(\b[41] ), .C(new_n8112), .Y(new_n8113));
  OA21x2_ASAP7_75t_L        g07857(.A1(new_n477), .A2(new_n6386), .B(new_n8113), .Y(new_n8114));
  O2A1O1Ixp33_ASAP7_75t_L   g07858(.A1(new_n477), .A2(new_n6386), .B(new_n8113), .C(new_n466), .Y(new_n8115));
  NAND2xp33_ASAP7_75t_L     g07859(.A(\a[8] ), .B(new_n8114), .Y(new_n8116));
  OA21x2_ASAP7_75t_L        g07860(.A1(new_n8114), .A2(new_n8115), .B(new_n8116), .Y(new_n8117));
  NAND3xp33_ASAP7_75t_L     g07861(.A(new_n8111), .B(new_n8117), .C(new_n8108), .Y(new_n8118));
  AO21x2_ASAP7_75t_L        g07862(.A1(new_n8108), .A2(new_n8111), .B(new_n8117), .Y(new_n8119));
  NAND3xp33_ASAP7_75t_L     g07863(.A(new_n7873), .B(new_n8119), .C(new_n8118), .Y(new_n8120));
  A2O1A1O1Ixp25_ASAP7_75t_L g07864(.A1(new_n7514), .A2(new_n7531), .B(new_n7517), .C(new_n7819), .D(new_n7807), .Y(new_n8121));
  AND3x1_ASAP7_75t_L        g07865(.A(new_n8111), .B(new_n8117), .C(new_n8108), .Y(new_n8122));
  AOI21xp33_ASAP7_75t_L     g07866(.A1(new_n8111), .A2(new_n8108), .B(new_n8117), .Y(new_n8123));
  OAI21xp33_ASAP7_75t_L     g07867(.A1(new_n8122), .A2(new_n8123), .B(new_n8121), .Y(new_n8124));
  NOR2xp33_ASAP7_75t_L      g07868(.A(new_n6671), .B(new_n375), .Y(new_n8125));
  AOI221xp5_ASAP7_75t_L     g07869(.A1(\b[45] ), .A2(new_n361), .B1(new_n349), .B2(\b[44] ), .C(new_n8125), .Y(new_n8126));
  O2A1O1Ixp33_ASAP7_75t_L   g07870(.A1(new_n356), .A2(new_n7255), .B(new_n8126), .C(new_n346), .Y(new_n8127));
  NOR2xp33_ASAP7_75t_L      g07871(.A(new_n346), .B(new_n8127), .Y(new_n8128));
  O2A1O1Ixp33_ASAP7_75t_L   g07872(.A1(new_n356), .A2(new_n7255), .B(new_n8126), .C(\a[5] ), .Y(new_n8129));
  NOR2xp33_ASAP7_75t_L      g07873(.A(new_n8129), .B(new_n8128), .Y(new_n8130));
  AOI21xp33_ASAP7_75t_L     g07874(.A1(new_n8124), .A2(new_n8120), .B(new_n8130), .Y(new_n8131));
  AND3x1_ASAP7_75t_L        g07875(.A(new_n8124), .B(new_n8130), .C(new_n8120), .Y(new_n8132));
  NOR2xp33_ASAP7_75t_L      g07876(.A(new_n8131), .B(new_n8132), .Y(new_n8133));
  OAI21xp33_ASAP7_75t_L     g07877(.A1(new_n7841), .A2(new_n7835), .B(new_n8133), .Y(new_n8134));
  A2O1A1O1Ixp25_ASAP7_75t_L g07878(.A1(new_n7538), .A2(new_n7837), .B(new_n7836), .C(new_n7829), .D(new_n7841), .Y(new_n8135));
  OAI21xp33_ASAP7_75t_L     g07879(.A1(new_n8131), .A2(new_n8132), .B(new_n8135), .Y(new_n8136));
  AOI21xp33_ASAP7_75t_L     g07880(.A1(new_n8134), .A2(new_n8136), .B(new_n7872), .Y(new_n8137));
  INVx1_ASAP7_75t_L         g07881(.A(new_n7872), .Y(new_n8138));
  NOR3xp33_ASAP7_75t_L      g07882(.A(new_n8135), .B(new_n8131), .C(new_n8132), .Y(new_n8139));
  A2O1A1O1Ixp25_ASAP7_75t_L g07883(.A1(new_n7533), .A2(new_n7532), .B(new_n7512), .C(new_n7520), .D(new_n7519), .Y(new_n8140));
  MAJIxp5_ASAP7_75t_L       g07884(.A(new_n7539), .B(new_n8140), .C(new_n7527), .Y(new_n8141));
  AO21x2_ASAP7_75t_L        g07885(.A1(new_n8120), .A2(new_n8124), .B(new_n8130), .Y(new_n8142));
  NAND3xp33_ASAP7_75t_L     g07886(.A(new_n8124), .B(new_n8120), .C(new_n8130), .Y(new_n8143));
  AOI221xp5_ASAP7_75t_L     g07887(.A1(new_n8142), .A2(new_n8143), .B1(new_n7842), .B2(new_n8141), .C(new_n7841), .Y(new_n8144));
  NOR3xp33_ASAP7_75t_L      g07888(.A(new_n8139), .B(new_n8144), .C(new_n8138), .Y(new_n8145));
  NOR2xp33_ASAP7_75t_L      g07889(.A(new_n8145), .B(new_n8137), .Y(new_n8146));
  XOR2x2_ASAP7_75t_L        g07890(.A(new_n8146), .B(new_n7855), .Y(\f[48] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g07891(.A1(new_n7852), .A2(new_n7847), .B(new_n7839), .C(new_n8146), .D(new_n8145), .Y(new_n8148));
  NAND2xp33_ASAP7_75t_L     g07892(.A(new_n8090), .B(new_n8094), .Y(new_n8149));
  INVx1_ASAP7_75t_L         g07893(.A(new_n8149), .Y(new_n8150));
  A2O1A1Ixp33_ASAP7_75t_L   g07894(.A1(\a[11] ), .A2(new_n8098), .B(new_n8099), .C(new_n8150), .Y(new_n8151));
  NAND2xp33_ASAP7_75t_L     g07895(.A(new_n8020), .B(new_n8022), .Y(new_n8152));
  A2O1A1Ixp33_ASAP7_75t_L   g07896(.A1(new_n8035), .A2(new_n8152), .B(new_n8053), .C(new_n8039), .Y(new_n8153));
  OAI22xp33_ASAP7_75t_L     g07897(.A1(new_n2089), .A2(new_n2703), .B1(new_n2879), .B2(new_n1962), .Y(new_n8154));
  AOI221xp5_ASAP7_75t_L     g07898(.A1(new_n1955), .A2(\b[28] ), .B1(new_n1964), .B2(new_n3085), .C(new_n8154), .Y(new_n8155));
  XNOR2x2_ASAP7_75t_L       g07899(.A(new_n1952), .B(new_n8155), .Y(new_n8156));
  NAND2xp33_ASAP7_75t_L     g07900(.A(new_n7956), .B(new_n7958), .Y(new_n8157));
  O2A1O1Ixp33_ASAP7_75t_L   g07901(.A1(new_n4906), .A2(new_n7894), .B(new_n7896), .C(new_n8157), .Y(new_n8158));
  NAND3xp33_ASAP7_75t_L     g07902(.A(new_n7920), .B(new_n7921), .C(new_n7930), .Y(new_n8159));
  INVx1_ASAP7_75t_L         g07903(.A(new_n7907), .Y(new_n8160));
  MAJIxp5_ASAP7_75t_L       g07904(.A(new_n7919), .B(new_n7619), .C(new_n8160), .Y(new_n8161));
  NAND2xp33_ASAP7_75t_L     g07905(.A(\b[3] ), .B(new_n7333), .Y(new_n8162));
  OAI221xp5_ASAP7_75t_L     g07906(.A1(new_n7318), .A2(new_n332), .B1(new_n289), .B2(new_n7614), .C(new_n8162), .Y(new_n8163));
  A2O1A1Ixp33_ASAP7_75t_L   g07907(.A1(new_n342), .A2(new_n7322), .B(new_n8163), .C(\a[47] ), .Y(new_n8164));
  AOI211xp5_ASAP7_75t_L     g07908(.A1(new_n342), .A2(new_n7322), .B(new_n7316), .C(new_n8163), .Y(new_n8165));
  A2O1A1O1Ixp25_ASAP7_75t_L g07909(.A1(new_n7322), .A2(new_n342), .B(new_n8163), .C(new_n8164), .D(new_n8165), .Y(new_n8166));
  NAND2xp33_ASAP7_75t_L     g07910(.A(new_n7905), .B(new_n7904), .Y(new_n8167));
  XNOR2x2_ASAP7_75t_L       g07911(.A(\a[49] ), .B(\a[48] ), .Y(new_n8168));
  NOR2xp33_ASAP7_75t_L      g07912(.A(new_n8168), .B(new_n8167), .Y(new_n8169));
  INVx1_ASAP7_75t_L         g07913(.A(\a[49] ), .Y(new_n8170));
  NAND2xp33_ASAP7_75t_L     g07914(.A(\a[50] ), .B(new_n8170), .Y(new_n8171));
  INVx1_ASAP7_75t_L         g07915(.A(\a[50] ), .Y(new_n8172));
  NAND2xp33_ASAP7_75t_L     g07916(.A(\a[49] ), .B(new_n8172), .Y(new_n8173));
  NAND2xp33_ASAP7_75t_L     g07917(.A(new_n8173), .B(new_n8171), .Y(new_n8174));
  NOR2xp33_ASAP7_75t_L      g07918(.A(new_n8174), .B(new_n7906), .Y(new_n8175));
  NAND2xp33_ASAP7_75t_L     g07919(.A(new_n8174), .B(new_n8167), .Y(new_n8176));
  NOR2xp33_ASAP7_75t_L      g07920(.A(new_n274), .B(new_n8176), .Y(new_n8177));
  AOI221xp5_ASAP7_75t_L     g07921(.A1(\b[1] ), .A2(new_n8175), .B1(new_n8169), .B2(\b[0] ), .C(new_n8177), .Y(new_n8178));
  NAND3xp33_ASAP7_75t_L     g07922(.A(new_n8178), .B(new_n8160), .C(\a[50] ), .Y(new_n8179));
  INVx1_ASAP7_75t_L         g07923(.A(new_n8179), .Y(new_n8180));
  AOI22xp33_ASAP7_75t_L     g07924(.A1(new_n8169), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n8175), .Y(new_n8181));
  OAI21xp33_ASAP7_75t_L     g07925(.A1(new_n8176), .A2(new_n274), .B(new_n8181), .Y(new_n8182));
  NAND2xp33_ASAP7_75t_L     g07926(.A(\a[50] ), .B(new_n8182), .Y(new_n8183));
  O2A1O1Ixp33_ASAP7_75t_L   g07927(.A1(new_n8176), .A2(new_n274), .B(new_n8181), .C(\a[50] ), .Y(new_n8184));
  O2A1O1Ixp33_ASAP7_75t_L   g07928(.A1(new_n8160), .A2(new_n8183), .B(\a[50] ), .C(new_n8184), .Y(new_n8185));
  OAI21xp33_ASAP7_75t_L     g07929(.A1(new_n8180), .A2(new_n8185), .B(new_n8166), .Y(new_n8186));
  A2O1A1Ixp33_ASAP7_75t_L   g07930(.A1(new_n342), .A2(new_n7322), .B(new_n8163), .C(new_n7316), .Y(new_n8187));
  INVx1_ASAP7_75t_L         g07931(.A(new_n8187), .Y(new_n8188));
  A2O1A1Ixp33_ASAP7_75t_L   g07932(.A1(new_n7904), .A2(new_n7905), .B(new_n284), .C(\a[50] ), .Y(new_n8189));
  O2A1O1Ixp33_ASAP7_75t_L   g07933(.A1(new_n8176), .A2(new_n274), .B(new_n8181), .C(new_n8172), .Y(new_n8190));
  NAND2xp33_ASAP7_75t_L     g07934(.A(\a[50] ), .B(new_n8178), .Y(new_n8191));
  OAI211xp5_ASAP7_75t_L     g07935(.A1(new_n8178), .A2(new_n8190), .B(new_n8191), .C(new_n8189), .Y(new_n8192));
  OAI211xp5_ASAP7_75t_L     g07936(.A1(new_n8165), .A2(new_n8188), .B(new_n8179), .C(new_n8192), .Y(new_n8193));
  NAND3xp33_ASAP7_75t_L     g07937(.A(new_n8161), .B(new_n8186), .C(new_n8193), .Y(new_n8194));
  NAND2xp33_ASAP7_75t_L     g07938(.A(new_n7916), .B(new_n7918), .Y(new_n8195));
  MAJIxp5_ASAP7_75t_L       g07939(.A(new_n8195), .B(new_n7907), .C(new_n7910), .Y(new_n8196));
  AOI211xp5_ASAP7_75t_L     g07940(.A1(new_n8192), .A2(new_n8179), .B(new_n8165), .C(new_n8188), .Y(new_n8197));
  INVx1_ASAP7_75t_L         g07941(.A(new_n8165), .Y(new_n8198));
  AOI211xp5_ASAP7_75t_L     g07942(.A1(new_n8198), .A2(new_n8187), .B(new_n8180), .C(new_n8185), .Y(new_n8199));
  OAI21xp33_ASAP7_75t_L     g07943(.A1(new_n8197), .A2(new_n8199), .B(new_n8196), .Y(new_n8200));
  NOR2xp33_ASAP7_75t_L      g07944(.A(new_n384), .B(new_n6741), .Y(new_n8201));
  AOI221xp5_ASAP7_75t_L     g07945(.A1(\b[7] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[6] ), .C(new_n8201), .Y(new_n8202));
  O2A1O1Ixp33_ASAP7_75t_L   g07946(.A1(new_n6443), .A2(new_n456), .B(new_n8202), .C(new_n6439), .Y(new_n8203));
  OAI21xp33_ASAP7_75t_L     g07947(.A1(new_n6443), .A2(new_n456), .B(new_n8202), .Y(new_n8204));
  NAND2xp33_ASAP7_75t_L     g07948(.A(new_n6439), .B(new_n8204), .Y(new_n8205));
  OA21x2_ASAP7_75t_L        g07949(.A1(new_n6439), .A2(new_n8203), .B(new_n8205), .Y(new_n8206));
  NAND3xp33_ASAP7_75t_L     g07950(.A(new_n8200), .B(new_n8194), .C(new_n8206), .Y(new_n8207));
  NOR3xp33_ASAP7_75t_L      g07951(.A(new_n8199), .B(new_n8197), .C(new_n8196), .Y(new_n8208));
  AOI21xp33_ASAP7_75t_L     g07952(.A1(new_n8186), .A2(new_n8193), .B(new_n8161), .Y(new_n8209));
  OAI21xp33_ASAP7_75t_L     g07953(.A1(new_n6439), .A2(new_n8203), .B(new_n8205), .Y(new_n8210));
  OAI21xp33_ASAP7_75t_L     g07954(.A1(new_n8209), .A2(new_n8208), .B(new_n8210), .Y(new_n8211));
  NAND4xp25_ASAP7_75t_L     g07955(.A(new_n7944), .B(new_n8207), .C(new_n8211), .D(new_n8159), .Y(new_n8212));
  NAND2xp33_ASAP7_75t_L     g07956(.A(new_n8207), .B(new_n8211), .Y(new_n8213));
  A2O1A1Ixp33_ASAP7_75t_L   g07957(.A1(new_n7926), .A2(new_n7927), .B(new_n7934), .C(new_n8159), .Y(new_n8214));
  NAND2xp33_ASAP7_75t_L     g07958(.A(new_n8214), .B(new_n8213), .Y(new_n8215));
  OAI22xp33_ASAP7_75t_L     g07959(.A1(new_n5640), .A2(new_n590), .B1(new_n534), .B2(new_n5925), .Y(new_n8216));
  AOI221xp5_ASAP7_75t_L     g07960(.A1(new_n5629), .A2(\b[10] ), .B1(new_n5637), .B2(new_n690), .C(new_n8216), .Y(new_n8217));
  XNOR2x2_ASAP7_75t_L       g07961(.A(\a[41] ), .B(new_n8217), .Y(new_n8218));
  NAND3xp33_ASAP7_75t_L     g07962(.A(new_n8212), .B(new_n8215), .C(new_n8218), .Y(new_n8219));
  AO21x2_ASAP7_75t_L        g07963(.A1(new_n8215), .A2(new_n8212), .B(new_n8218), .Y(new_n8220));
  A2O1A1Ixp33_ASAP7_75t_L   g07964(.A1(new_n7634), .A2(new_n7605), .B(new_n7599), .C(new_n7640), .Y(new_n8221));
  A2O1A1Ixp33_ASAP7_75t_L   g07965(.A1(new_n8221), .A2(new_n7955), .B(new_n7954), .C(new_n8220), .Y(new_n8222));
  A2O1A1O1Ixp25_ASAP7_75t_L g07966(.A1(new_n7652), .A2(new_n7657), .B(new_n7633), .C(new_n7942), .D(new_n7954), .Y(new_n8223));
  AOI21xp33_ASAP7_75t_L     g07967(.A1(new_n8219), .A2(new_n8220), .B(new_n8223), .Y(new_n8224));
  NAND2xp33_ASAP7_75t_L     g07968(.A(\b[12] ), .B(new_n4916), .Y(new_n8225));
  OAI221xp5_ASAP7_75t_L     g07969(.A1(new_n4908), .A2(new_n936), .B1(new_n748), .B2(new_n5144), .C(new_n8225), .Y(new_n8226));
  AOI211xp5_ASAP7_75t_L     g07970(.A1(new_n1166), .A2(new_n4912), .B(new_n8226), .C(new_n4906), .Y(new_n8227));
  INVx1_ASAP7_75t_L         g07971(.A(new_n8227), .Y(new_n8228));
  A2O1A1Ixp33_ASAP7_75t_L   g07972(.A1(new_n1166), .A2(new_n4912), .B(new_n8226), .C(new_n4906), .Y(new_n8229));
  NAND2xp33_ASAP7_75t_L     g07973(.A(new_n8229), .B(new_n8228), .Y(new_n8230));
  AOI311xp33_ASAP7_75t_L    g07974(.A1(new_n8219), .A2(new_n8222), .A3(new_n8220), .B(new_n8230), .C(new_n8224), .Y(new_n8231));
  AOI21xp33_ASAP7_75t_L     g07975(.A1(new_n8212), .A2(new_n8215), .B(new_n8218), .Y(new_n8232));
  O2A1O1Ixp33_ASAP7_75t_L   g07976(.A1(new_n7953), .A2(new_n7957), .B(new_n7946), .C(new_n8232), .Y(new_n8233));
  NAND3xp33_ASAP7_75t_L     g07977(.A(new_n8223), .B(new_n8219), .C(new_n8220), .Y(new_n8234));
  A2O1A1Ixp33_ASAP7_75t_L   g07978(.A1(new_n1166), .A2(new_n4912), .B(new_n8226), .C(\a[38] ), .Y(new_n8235));
  A2O1A1O1Ixp25_ASAP7_75t_L g07979(.A1(new_n4912), .A2(new_n1166), .B(new_n8226), .C(new_n8235), .D(new_n8227), .Y(new_n8236));
  A2O1A1O1Ixp25_ASAP7_75t_L g07980(.A1(new_n8219), .A2(new_n8233), .B(new_n8223), .C(new_n8234), .D(new_n8236), .Y(new_n8237));
  NOR2xp33_ASAP7_75t_L      g07981(.A(new_n8231), .B(new_n8237), .Y(new_n8238));
  A2O1A1Ixp33_ASAP7_75t_L   g07982(.A1(new_n7960), .A2(new_n7891), .B(new_n8158), .C(new_n8238), .Y(new_n8239));
  NOR2xp33_ASAP7_75t_L      g07983(.A(new_n7949), .B(new_n7948), .Y(new_n8240));
  O2A1O1Ixp33_ASAP7_75t_L   g07984(.A1(new_n7967), .A2(new_n8240), .B(new_n7891), .C(new_n8158), .Y(new_n8241));
  A2O1A1Ixp33_ASAP7_75t_L   g07985(.A1(new_n7653), .A2(new_n7640), .B(new_n7947), .C(new_n7946), .Y(new_n8242));
  INVx1_ASAP7_75t_L         g07986(.A(new_n8219), .Y(new_n8243));
  OAI21xp33_ASAP7_75t_L     g07987(.A1(new_n8243), .A2(new_n8232), .B(new_n8242), .Y(new_n8244));
  NAND3xp33_ASAP7_75t_L     g07988(.A(new_n8244), .B(new_n8234), .C(new_n8236), .Y(new_n8245));
  A2O1A1O1Ixp25_ASAP7_75t_L g07989(.A1(new_n7942), .A2(new_n8221), .B(new_n7954), .C(new_n8220), .D(new_n8243), .Y(new_n8246));
  A2O1A1Ixp33_ASAP7_75t_L   g07990(.A1(new_n8246), .A2(new_n8220), .B(new_n8224), .C(new_n8230), .Y(new_n8247));
  NAND2xp33_ASAP7_75t_L     g07991(.A(new_n8245), .B(new_n8247), .Y(new_n8248));
  NAND2xp33_ASAP7_75t_L     g07992(.A(new_n8248), .B(new_n8241), .Y(new_n8249));
  OAI22xp33_ASAP7_75t_L     g07993(.A1(new_n4397), .A2(new_n960), .B1(new_n1043), .B2(new_n4142), .Y(new_n8250));
  AOI221xp5_ASAP7_75t_L     g07994(.A1(new_n4156), .A2(\b[16] ), .B1(new_n4151), .B2(new_n1156), .C(new_n8250), .Y(new_n8251));
  XNOR2x2_ASAP7_75t_L       g07995(.A(new_n4145), .B(new_n8251), .Y(new_n8252));
  NAND3xp33_ASAP7_75t_L     g07996(.A(new_n8249), .B(new_n8239), .C(new_n8252), .Y(new_n8253));
  O2A1O1Ixp33_ASAP7_75t_L   g07997(.A1(new_n7952), .A2(new_n8157), .B(new_n7968), .C(new_n8248), .Y(new_n8254));
  O2A1O1Ixp33_ASAP7_75t_L   g07998(.A1(new_n7360), .A2(new_n7361), .B(new_n7364), .C(new_n7301), .Y(new_n8255));
  O2A1O1Ixp33_ASAP7_75t_L   g07999(.A1(new_n7376), .A2(new_n8255), .B(new_n7650), .C(new_n7660), .Y(new_n8256));
  A2O1A1Ixp33_ASAP7_75t_L   g08000(.A1(new_n7951), .A2(\a[38] ), .B(new_n7895), .C(new_n8240), .Y(new_n8257));
  A2O1A1Ixp33_ASAP7_75t_L   g08001(.A1(new_n7950), .A2(new_n8157), .B(new_n8256), .C(new_n8257), .Y(new_n8258));
  NOR2xp33_ASAP7_75t_L      g08002(.A(new_n8238), .B(new_n8258), .Y(new_n8259));
  XNOR2x2_ASAP7_75t_L       g08003(.A(\a[35] ), .B(new_n8251), .Y(new_n8260));
  OAI21xp33_ASAP7_75t_L     g08004(.A1(new_n8259), .A2(new_n8254), .B(new_n8260), .Y(new_n8261));
  NOR3xp33_ASAP7_75t_L      g08005(.A(new_n7891), .B(new_n7967), .C(new_n7961), .Y(new_n8262));
  A2O1A1Ixp33_ASAP7_75t_L   g08006(.A1(new_n7891), .A2(new_n7960), .B(new_n8262), .C(new_n7889), .Y(new_n8263));
  A2O1A1O1Ixp25_ASAP7_75t_L g08007(.A1(new_n7677), .A2(new_n7680), .B(new_n7670), .C(new_n8263), .D(new_n7963), .Y(new_n8264));
  NAND3xp33_ASAP7_75t_L     g08008(.A(new_n8264), .B(new_n8261), .C(new_n8253), .Y(new_n8265));
  AO21x2_ASAP7_75t_L        g08009(.A1(new_n8253), .A2(new_n8261), .B(new_n8264), .Y(new_n8266));
  NOR2xp33_ASAP7_75t_L      g08010(.A(new_n1458), .B(new_n3509), .Y(new_n8267));
  AOI221xp5_ASAP7_75t_L     g08011(.A1(\b[17] ), .A2(new_n3708), .B1(\b[19] ), .B2(new_n3503), .C(new_n8267), .Y(new_n8268));
  INVx1_ASAP7_75t_L         g08012(.A(new_n8268), .Y(new_n8269));
  A2O1A1Ixp33_ASAP7_75t_L   g08013(.A1(new_n1607), .A2(new_n3505), .B(new_n8269), .C(\a[32] ), .Y(new_n8270));
  O2A1O1Ixp33_ASAP7_75t_L   g08014(.A1(new_n3513), .A2(new_n1628), .B(new_n8268), .C(\a[32] ), .Y(new_n8271));
  AOI21xp33_ASAP7_75t_L     g08015(.A1(new_n8270), .A2(\a[32] ), .B(new_n8271), .Y(new_n8272));
  NAND3xp33_ASAP7_75t_L     g08016(.A(new_n8266), .B(new_n8265), .C(new_n8272), .Y(new_n8273));
  AND3x1_ASAP7_75t_L        g08017(.A(new_n8264), .B(new_n8261), .C(new_n8253), .Y(new_n8274));
  AOI21xp33_ASAP7_75t_L     g08018(.A1(new_n8261), .A2(new_n8253), .B(new_n8264), .Y(new_n8275));
  INVx1_ASAP7_75t_L         g08019(.A(new_n8272), .Y(new_n8276));
  OAI21xp33_ASAP7_75t_L     g08020(.A1(new_n8275), .A2(new_n8274), .B(new_n8276), .Y(new_n8277));
  AND4x1_ASAP7_75t_L        g08021(.A(new_n7989), .B(new_n7982), .C(new_n8277), .D(new_n8273), .Y(new_n8278));
  MAJIxp5_ASAP7_75t_L       g08022(.A(new_n7988), .B(new_n7972), .C(new_n7981), .Y(new_n8279));
  AOI21xp33_ASAP7_75t_L     g08023(.A1(new_n8277), .A2(new_n8273), .B(new_n8279), .Y(new_n8280));
  NAND2xp33_ASAP7_75t_L     g08024(.A(\b[21] ), .B(new_n2936), .Y(new_n8281));
  OAI221xp5_ASAP7_75t_L     g08025(.A1(new_n2930), .A2(new_n2045), .B1(new_n1745), .B2(new_n3133), .C(new_n8281), .Y(new_n8282));
  A2O1A1Ixp33_ASAP7_75t_L   g08026(.A1(new_n2056), .A2(new_n2932), .B(new_n8282), .C(\a[29] ), .Y(new_n8283));
  AOI211xp5_ASAP7_75t_L     g08027(.A1(new_n2056), .A2(new_n2932), .B(new_n8282), .C(new_n2928), .Y(new_n8284));
  A2O1A1O1Ixp25_ASAP7_75t_L g08028(.A1(new_n2932), .A2(new_n2056), .B(new_n8282), .C(new_n8283), .D(new_n8284), .Y(new_n8285));
  INVx1_ASAP7_75t_L         g08029(.A(new_n8285), .Y(new_n8286));
  NOR3xp33_ASAP7_75t_L      g08030(.A(new_n8286), .B(new_n8280), .C(new_n8278), .Y(new_n8287));
  NAND3xp33_ASAP7_75t_L     g08031(.A(new_n8279), .B(new_n8277), .C(new_n8273), .Y(new_n8288));
  NAND2xp33_ASAP7_75t_L     g08032(.A(new_n8273), .B(new_n8277), .Y(new_n8289));
  A2O1A1Ixp33_ASAP7_75t_L   g08033(.A1(new_n7688), .A2(new_n7882), .B(new_n7985), .C(new_n7982), .Y(new_n8290));
  NAND2xp33_ASAP7_75t_L     g08034(.A(new_n8289), .B(new_n8290), .Y(new_n8291));
  AOI21xp33_ASAP7_75t_L     g08035(.A1(new_n8291), .A2(new_n8288), .B(new_n8285), .Y(new_n8292));
  NAND2xp33_ASAP7_75t_L     g08036(.A(new_n7989), .B(new_n7986), .Y(new_n8293));
  MAJIxp5_ASAP7_75t_L       g08037(.A(new_n8002), .B(new_n7994), .C(new_n8293), .Y(new_n8294));
  NOR3xp33_ASAP7_75t_L      g08038(.A(new_n8294), .B(new_n8292), .C(new_n8287), .Y(new_n8295));
  NOR2xp33_ASAP7_75t_L      g08039(.A(new_n7996), .B(new_n7998), .Y(new_n8296));
  NAND2xp33_ASAP7_75t_L     g08040(.A(new_n7999), .B(new_n8296), .Y(new_n8297));
  NAND3xp33_ASAP7_75t_L     g08041(.A(new_n8291), .B(new_n8288), .C(new_n8285), .Y(new_n8298));
  OAI21xp33_ASAP7_75t_L     g08042(.A1(new_n8280), .A2(new_n8278), .B(new_n8286), .Y(new_n8299));
  AOI22xp33_ASAP7_75t_L     g08043(.A1(new_n8298), .A2(new_n8299), .B1(new_n8297), .B2(new_n8016), .Y(new_n8300));
  NAND2xp33_ASAP7_75t_L     g08044(.A(\b[24] ), .B(new_n2421), .Y(new_n8301));
  OAI221xp5_ASAP7_75t_L     g08045(.A1(new_n2415), .A2(new_n2377), .B1(new_n2188), .B2(new_n2572), .C(new_n8301), .Y(new_n8302));
  A2O1A1Ixp33_ASAP7_75t_L   g08046(.A1(new_n5001), .A2(new_n2417), .B(new_n8302), .C(\a[26] ), .Y(new_n8303));
  AOI211xp5_ASAP7_75t_L     g08047(.A1(new_n5001), .A2(new_n2417), .B(new_n8302), .C(new_n2413), .Y(new_n8304));
  A2O1A1O1Ixp25_ASAP7_75t_L g08048(.A1(new_n2417), .A2(new_n5001), .B(new_n8302), .C(new_n8303), .D(new_n8304), .Y(new_n8305));
  INVx1_ASAP7_75t_L         g08049(.A(new_n8305), .Y(new_n8306));
  NOR3xp33_ASAP7_75t_L      g08050(.A(new_n8300), .B(new_n8295), .C(new_n8306), .Y(new_n8307));
  NAND4xp25_ASAP7_75t_L     g08051(.A(new_n8016), .B(new_n8298), .C(new_n8299), .D(new_n8297), .Y(new_n8308));
  OAI21xp33_ASAP7_75t_L     g08052(.A1(new_n8287), .A2(new_n8292), .B(new_n8294), .Y(new_n8309));
  AOI21xp33_ASAP7_75t_L     g08053(.A1(new_n8308), .A2(new_n8309), .B(new_n8305), .Y(new_n8310));
  A2O1A1Ixp33_ASAP7_75t_L   g08054(.A1(new_n7727), .A2(new_n7431), .B(new_n7717), .C(new_n7716), .Y(new_n8311));
  AOI21xp33_ASAP7_75t_L     g08055(.A1(new_n8016), .A2(new_n8011), .B(new_n8018), .Y(new_n8312));
  A2O1A1Ixp33_ASAP7_75t_L   g08056(.A1(new_n8311), .A2(new_n7725), .B(new_n8312), .C(new_n8019), .Y(new_n8313));
  OAI21xp33_ASAP7_75t_L     g08057(.A1(new_n8307), .A2(new_n8310), .B(new_n8313), .Y(new_n8314));
  NAND3xp33_ASAP7_75t_L     g08058(.A(new_n8308), .B(new_n8305), .C(new_n8309), .Y(new_n8315));
  OAI21xp33_ASAP7_75t_L     g08059(.A1(new_n8295), .A2(new_n8300), .B(new_n8306), .Y(new_n8316));
  NOR3xp33_ASAP7_75t_L      g08060(.A(new_n8001), .B(new_n8009), .C(new_n8003), .Y(new_n8317));
  A2O1A1O1Ixp25_ASAP7_75t_L g08061(.A1(new_n7716), .A2(new_n7743), .B(new_n7728), .C(new_n8010), .D(new_n8317), .Y(new_n8318));
  NAND3xp33_ASAP7_75t_L     g08062(.A(new_n8318), .B(new_n8316), .C(new_n8315), .Y(new_n8319));
  AOI21xp33_ASAP7_75t_L     g08063(.A1(new_n8319), .A2(new_n8314), .B(new_n8156), .Y(new_n8320));
  XNOR2x2_ASAP7_75t_L       g08064(.A(\a[23] ), .B(new_n8155), .Y(new_n8321));
  AOI21xp33_ASAP7_75t_L     g08065(.A1(new_n8316), .A2(new_n8315), .B(new_n8318), .Y(new_n8322));
  NOR3xp33_ASAP7_75t_L      g08066(.A(new_n8313), .B(new_n8310), .C(new_n8307), .Y(new_n8323));
  NOR3xp33_ASAP7_75t_L      g08067(.A(new_n8323), .B(new_n8322), .C(new_n8321), .Y(new_n8324));
  NOR2xp33_ASAP7_75t_L      g08068(.A(new_n8320), .B(new_n8324), .Y(new_n8325));
  NAND2xp33_ASAP7_75t_L     g08069(.A(new_n8153), .B(new_n8325), .Y(new_n8326));
  OAI21xp33_ASAP7_75t_L     g08070(.A1(new_n8322), .A2(new_n8323), .B(new_n8321), .Y(new_n8327));
  NAND3xp33_ASAP7_75t_L     g08071(.A(new_n8319), .B(new_n8314), .C(new_n8156), .Y(new_n8328));
  AO221x2_ASAP7_75t_L       g08072(.A1(new_n8036), .A2(new_n8038), .B1(new_n8327), .B2(new_n8328), .C(new_n8040), .Y(new_n8329));
  NOR2xp33_ASAP7_75t_L      g08073(.A(new_n3456), .B(new_n1517), .Y(new_n8330));
  AOI221xp5_ASAP7_75t_L     g08074(.A1(\b[29] ), .A2(new_n1659), .B1(\b[31] ), .B2(new_n1511), .C(new_n8330), .Y(new_n8331));
  O2A1O1Ixp33_ASAP7_75t_L   g08075(.A1(new_n1521), .A2(new_n3681), .B(new_n8331), .C(new_n1501), .Y(new_n8332));
  INVx1_ASAP7_75t_L         g08076(.A(new_n8332), .Y(new_n8333));
  O2A1O1Ixp33_ASAP7_75t_L   g08077(.A1(new_n1521), .A2(new_n3681), .B(new_n8331), .C(\a[20] ), .Y(new_n8334));
  AO21x2_ASAP7_75t_L        g08078(.A1(\a[20] ), .A2(new_n8333), .B(new_n8334), .Y(new_n8335));
  AOI21xp33_ASAP7_75t_L     g08079(.A1(new_n8326), .A2(new_n8329), .B(new_n8335), .Y(new_n8336));
  A2O1A1Ixp33_ASAP7_75t_L   g08080(.A1(new_n7745), .A2(new_n7742), .B(new_n7740), .C(new_n8036), .Y(new_n8337));
  NAND2xp33_ASAP7_75t_L     g08081(.A(new_n8328), .B(new_n8327), .Y(new_n8338));
  O2A1O1Ixp33_ASAP7_75t_L   g08082(.A1(new_n8152), .A2(new_n8028), .B(new_n8337), .C(new_n8338), .Y(new_n8339));
  AOI21xp33_ASAP7_75t_L     g08083(.A1(new_n8328), .A2(new_n8327), .B(new_n8153), .Y(new_n8340));
  AOI21xp33_ASAP7_75t_L     g08084(.A1(new_n8333), .A2(\a[20] ), .B(new_n8334), .Y(new_n8341));
  NOR3xp33_ASAP7_75t_L      g08085(.A(new_n8339), .B(new_n8340), .C(new_n8341), .Y(new_n8342));
  OAI21xp33_ASAP7_75t_L     g08086(.A1(new_n8071), .A2(new_n8069), .B(new_n8049), .Y(new_n8343));
  NOR3xp33_ASAP7_75t_L      g08087(.A(new_n8343), .B(new_n8342), .C(new_n8336), .Y(new_n8344));
  OAI21xp33_ASAP7_75t_L     g08088(.A1(new_n8320), .A2(new_n8324), .B(new_n8153), .Y(new_n8345));
  A2O1A1Ixp33_ASAP7_75t_L   g08089(.A1(new_n8345), .A2(new_n8153), .B(new_n8340), .C(new_n8341), .Y(new_n8346));
  NAND3xp33_ASAP7_75t_L     g08090(.A(new_n8326), .B(new_n8329), .C(new_n8335), .Y(new_n8347));
  A2O1A1O1Ixp25_ASAP7_75t_L g08091(.A1(new_n7748), .A2(new_n7756), .B(new_n8059), .C(new_n8056), .D(new_n8070), .Y(new_n8348));
  AOI21xp33_ASAP7_75t_L     g08092(.A1(new_n8347), .A2(new_n8346), .B(new_n8348), .Y(new_n8349));
  NOR2xp33_ASAP7_75t_L      g08093(.A(new_n4101), .B(new_n2118), .Y(new_n8350));
  AOI221xp5_ASAP7_75t_L     g08094(.A1(\b[32] ), .A2(new_n1290), .B1(\b[34] ), .B2(new_n1209), .C(new_n8350), .Y(new_n8351));
  O2A1O1Ixp33_ASAP7_75t_L   g08095(.A1(new_n1210), .A2(new_n4352), .B(new_n8351), .C(new_n1206), .Y(new_n8352));
  O2A1O1Ixp33_ASAP7_75t_L   g08096(.A1(new_n1210), .A2(new_n4352), .B(new_n8351), .C(\a[17] ), .Y(new_n8353));
  INVx1_ASAP7_75t_L         g08097(.A(new_n8353), .Y(new_n8354));
  OAI21xp33_ASAP7_75t_L     g08098(.A1(new_n1206), .A2(new_n8352), .B(new_n8354), .Y(new_n8355));
  NOR3xp33_ASAP7_75t_L      g08099(.A(new_n8344), .B(new_n8349), .C(new_n8355), .Y(new_n8356));
  NAND3xp33_ASAP7_75t_L     g08100(.A(new_n8348), .B(new_n8347), .C(new_n8346), .Y(new_n8357));
  OAI21xp33_ASAP7_75t_L     g08101(.A1(new_n8336), .A2(new_n8342), .B(new_n8343), .Y(new_n8358));
  OA21x2_ASAP7_75t_L        g08102(.A1(new_n1206), .A2(new_n8352), .B(new_n8354), .Y(new_n8359));
  AOI21xp33_ASAP7_75t_L     g08103(.A1(new_n8357), .A2(new_n8358), .B(new_n8359), .Y(new_n8360));
  NOR2xp33_ASAP7_75t_L      g08104(.A(new_n8360), .B(new_n8356), .Y(new_n8361));
  NOR2xp33_ASAP7_75t_L      g08105(.A(new_n8060), .B(new_n8058), .Y(new_n8362));
  MAJIxp5_ASAP7_75t_L       g08106(.A(new_n8084), .B(new_n8067), .C(new_n8362), .Y(new_n8363));
  NAND2xp33_ASAP7_75t_L     g08107(.A(new_n8361), .B(new_n8363), .Y(new_n8364));
  NAND3xp33_ASAP7_75t_L     g08108(.A(new_n8357), .B(new_n8358), .C(new_n8355), .Y(new_n8365));
  NAND2xp33_ASAP7_75t_L     g08109(.A(new_n8073), .B(new_n8072), .Y(new_n8366));
  MAJIxp5_ASAP7_75t_L       g08110(.A(new_n7879), .B(new_n8074), .C(new_n8366), .Y(new_n8367));
  A2O1A1Ixp33_ASAP7_75t_L   g08111(.A1(new_n8365), .A2(new_n8355), .B(new_n8356), .C(new_n8367), .Y(new_n8368));
  NOR2xp33_ASAP7_75t_L      g08112(.A(new_n5074), .B(new_n869), .Y(new_n8369));
  AOI221xp5_ASAP7_75t_L     g08113(.A1(\b[35] ), .A2(new_n985), .B1(\b[36] ), .B2(new_n885), .C(new_n8369), .Y(new_n8370));
  O2A1O1Ixp33_ASAP7_75t_L   g08114(.A1(new_n872), .A2(new_n5083), .B(new_n8370), .C(new_n867), .Y(new_n8371));
  NOR2xp33_ASAP7_75t_L      g08115(.A(new_n867), .B(new_n8371), .Y(new_n8372));
  O2A1O1Ixp33_ASAP7_75t_L   g08116(.A1(new_n872), .A2(new_n5083), .B(new_n8370), .C(\a[14] ), .Y(new_n8373));
  NOR2xp33_ASAP7_75t_L      g08117(.A(new_n8373), .B(new_n8372), .Y(new_n8374));
  NAND3xp33_ASAP7_75t_L     g08118(.A(new_n8364), .B(new_n8368), .C(new_n8374), .Y(new_n8375));
  AO21x2_ASAP7_75t_L        g08119(.A1(new_n8368), .A2(new_n8364), .B(new_n8374), .Y(new_n8376));
  A2O1A1O1Ixp25_ASAP7_75t_L g08120(.A1(new_n7783), .A2(new_n7781), .B(new_n7876), .C(new_n8088), .D(new_n8091), .Y(new_n8377));
  AND3x1_ASAP7_75t_L        g08121(.A(new_n8377), .B(new_n8376), .C(new_n8375), .Y(new_n8378));
  AOI21xp33_ASAP7_75t_L     g08122(.A1(new_n8376), .A2(new_n8375), .B(new_n8377), .Y(new_n8379));
  NOR2xp33_ASAP7_75t_L      g08123(.A(new_n5570), .B(new_n1550), .Y(new_n8380));
  AOI221xp5_ASAP7_75t_L     g08124(.A1(\b[38] ), .A2(new_n713), .B1(\b[40] ), .B2(new_n640), .C(new_n8380), .Y(new_n8381));
  O2A1O1Ixp33_ASAP7_75t_L   g08125(.A1(new_n641), .A2(new_n5862), .B(new_n8381), .C(new_n637), .Y(new_n8382));
  INVx1_ASAP7_75t_L         g08126(.A(new_n8382), .Y(new_n8383));
  O2A1O1Ixp33_ASAP7_75t_L   g08127(.A1(new_n641), .A2(new_n5862), .B(new_n8381), .C(\a[11] ), .Y(new_n8384));
  AOI21xp33_ASAP7_75t_L     g08128(.A1(new_n8383), .A2(\a[11] ), .B(new_n8384), .Y(new_n8385));
  INVx1_ASAP7_75t_L         g08129(.A(new_n8385), .Y(new_n8386));
  NOR3xp33_ASAP7_75t_L      g08130(.A(new_n8378), .B(new_n8386), .C(new_n8379), .Y(new_n8387));
  NAND3xp33_ASAP7_75t_L     g08131(.A(new_n8377), .B(new_n8376), .C(new_n8375), .Y(new_n8388));
  AO21x2_ASAP7_75t_L        g08132(.A1(new_n8375), .A2(new_n8376), .B(new_n8377), .Y(new_n8389));
  AOI21xp33_ASAP7_75t_L     g08133(.A1(new_n8389), .A2(new_n8388), .B(new_n8385), .Y(new_n8390));
  NOR2xp33_ASAP7_75t_L      g08134(.A(new_n8390), .B(new_n8387), .Y(new_n8391));
  NAND3xp33_ASAP7_75t_L     g08135(.A(new_n8391), .B(new_n8111), .C(new_n8151), .Y(new_n8392));
  NAND3xp33_ASAP7_75t_L     g08136(.A(new_n8389), .B(new_n8388), .C(new_n8385), .Y(new_n8393));
  OAI21xp33_ASAP7_75t_L     g08137(.A1(new_n8379), .A2(new_n8378), .B(new_n8386), .Y(new_n8394));
  NAND2xp33_ASAP7_75t_L     g08138(.A(new_n8393), .B(new_n8394), .Y(new_n8395));
  MAJIxp5_ASAP7_75t_L       g08139(.A(new_n8107), .B(new_n8100), .C(new_n8149), .Y(new_n8396));
  NAND2xp33_ASAP7_75t_L     g08140(.A(new_n8396), .B(new_n8395), .Y(new_n8397));
  NOR2xp33_ASAP7_75t_L      g08141(.A(new_n6378), .B(new_n513), .Y(new_n8398));
  AOI221xp5_ASAP7_75t_L     g08142(.A1(\b[41] ), .A2(new_n560), .B1(\b[43] ), .B2(new_n475), .C(new_n8398), .Y(new_n8399));
  O2A1O1Ixp33_ASAP7_75t_L   g08143(.A1(new_n477), .A2(new_n6679), .B(new_n8399), .C(new_n466), .Y(new_n8400));
  INVx1_ASAP7_75t_L         g08144(.A(new_n8400), .Y(new_n8401));
  O2A1O1Ixp33_ASAP7_75t_L   g08145(.A1(new_n477), .A2(new_n6679), .B(new_n8399), .C(\a[8] ), .Y(new_n8402));
  AOI21xp33_ASAP7_75t_L     g08146(.A1(new_n8401), .A2(\a[8] ), .B(new_n8402), .Y(new_n8403));
  NAND3xp33_ASAP7_75t_L     g08147(.A(new_n8392), .B(new_n8397), .C(new_n8403), .Y(new_n8404));
  NOR2xp33_ASAP7_75t_L      g08148(.A(new_n8396), .B(new_n8395), .Y(new_n8405));
  AOI21xp33_ASAP7_75t_L     g08149(.A1(new_n8111), .A2(new_n8151), .B(new_n8391), .Y(new_n8406));
  INVx1_ASAP7_75t_L         g08150(.A(new_n8403), .Y(new_n8407));
  OAI21xp33_ASAP7_75t_L     g08151(.A1(new_n8405), .A2(new_n8406), .B(new_n8407), .Y(new_n8408));
  XNOR2x2_ASAP7_75t_L       g08152(.A(new_n8107), .B(new_n8110), .Y(new_n8409));
  INVx1_ASAP7_75t_L         g08153(.A(new_n8117), .Y(new_n8410));
  MAJIxp5_ASAP7_75t_L       g08154(.A(new_n7873), .B(new_n8410), .C(new_n8409), .Y(new_n8411));
  NAND3xp33_ASAP7_75t_L     g08155(.A(new_n8411), .B(new_n8408), .C(new_n8404), .Y(new_n8412));
  NOR3xp33_ASAP7_75t_L      g08156(.A(new_n8406), .B(new_n8407), .C(new_n8405), .Y(new_n8413));
  AOI21xp33_ASAP7_75t_L     g08157(.A1(new_n8392), .A2(new_n8397), .B(new_n8403), .Y(new_n8414));
  NAND2xp33_ASAP7_75t_L     g08158(.A(new_n8108), .B(new_n8111), .Y(new_n8415));
  MAJIxp5_ASAP7_75t_L       g08159(.A(new_n8121), .B(new_n8415), .C(new_n8117), .Y(new_n8416));
  OAI21xp33_ASAP7_75t_L     g08160(.A1(new_n8413), .A2(new_n8414), .B(new_n8416), .Y(new_n8417));
  OAI22xp33_ASAP7_75t_L     g08161(.A1(new_n350), .A2(new_n7249), .B1(new_n6944), .B2(new_n375), .Y(new_n8418));
  AOI221xp5_ASAP7_75t_L     g08162(.A1(new_n361), .A2(\b[46] ), .B1(new_n359), .B2(new_n7278), .C(new_n8418), .Y(new_n8419));
  XNOR2x2_ASAP7_75t_L       g08163(.A(new_n346), .B(new_n8419), .Y(new_n8420));
  AND3x1_ASAP7_75t_L        g08164(.A(new_n8417), .B(new_n8412), .C(new_n8420), .Y(new_n8421));
  AOI21xp33_ASAP7_75t_L     g08165(.A1(new_n8417), .A2(new_n8412), .B(new_n8420), .Y(new_n8422));
  OAI21xp33_ASAP7_75t_L     g08166(.A1(new_n8132), .A2(new_n8135), .B(new_n8142), .Y(new_n8423));
  NOR3xp33_ASAP7_75t_L      g08167(.A(new_n8423), .B(new_n8421), .C(new_n8422), .Y(new_n8424));
  NOR2xp33_ASAP7_75t_L      g08168(.A(new_n8422), .B(new_n8421), .Y(new_n8425));
  O2A1O1Ixp33_ASAP7_75t_L   g08169(.A1(new_n8135), .A2(new_n8132), .B(new_n8142), .C(new_n8425), .Y(new_n8426));
  INVx1_ASAP7_75t_L         g08170(.A(\b[49] ), .Y(new_n8427));
  NAND2xp33_ASAP7_75t_L     g08171(.A(\b[47] ), .B(new_n286), .Y(new_n8428));
  OAI221xp5_ASAP7_75t_L     g08172(.A1(new_n285), .A2(new_n7860), .B1(new_n8427), .B2(new_n269), .C(new_n8428), .Y(new_n8429));
  NOR2xp33_ASAP7_75t_L      g08173(.A(\b[48] ), .B(\b[49] ), .Y(new_n8430));
  NOR2xp33_ASAP7_75t_L      g08174(.A(new_n7860), .B(new_n8427), .Y(new_n8431));
  NOR2xp33_ASAP7_75t_L      g08175(.A(new_n8430), .B(new_n8431), .Y(new_n8432));
  A2O1A1Ixp33_ASAP7_75t_L   g08176(.A1(\b[48] ), .A2(\b[47] ), .B(new_n7864), .C(new_n8432), .Y(new_n8433));
  INVx1_ASAP7_75t_L         g08177(.A(new_n8433), .Y(new_n8434));
  O2A1O1Ixp33_ASAP7_75t_L   g08178(.A1(new_n7553), .A2(new_n7556), .B(new_n7862), .C(new_n7861), .Y(new_n8435));
  INVx1_ASAP7_75t_L         g08179(.A(new_n8435), .Y(new_n8436));
  NOR2xp33_ASAP7_75t_L      g08180(.A(new_n8432), .B(new_n8436), .Y(new_n8437));
  NOR2xp33_ASAP7_75t_L      g08181(.A(new_n8434), .B(new_n8437), .Y(new_n8438));
  A2O1A1Ixp33_ASAP7_75t_L   g08182(.A1(new_n8438), .A2(new_n273), .B(new_n8429), .C(\a[2] ), .Y(new_n8439));
  AOI211xp5_ASAP7_75t_L     g08183(.A1(new_n8438), .A2(new_n273), .B(new_n8429), .C(new_n257), .Y(new_n8440));
  A2O1A1O1Ixp25_ASAP7_75t_L g08184(.A1(new_n273), .A2(new_n8438), .B(new_n8429), .C(new_n8439), .D(new_n8440), .Y(new_n8441));
  OAI21xp33_ASAP7_75t_L     g08185(.A1(new_n8424), .A2(new_n8426), .B(new_n8441), .Y(new_n8442));
  NOR3xp33_ASAP7_75t_L      g08186(.A(new_n8426), .B(new_n8441), .C(new_n8424), .Y(new_n8443));
  INVx1_ASAP7_75t_L         g08187(.A(new_n8443), .Y(new_n8444));
  NAND2xp33_ASAP7_75t_L     g08188(.A(new_n8442), .B(new_n8444), .Y(new_n8445));
  XOR2x2_ASAP7_75t_L        g08189(.A(new_n8148), .B(new_n8445), .Y(\f[49] ));
  OAI211xp5_ASAP7_75t_L     g08190(.A1(new_n8372), .A2(new_n8373), .B(new_n8364), .C(new_n8368), .Y(new_n8447));
  A2O1A1Ixp33_ASAP7_75t_L   g08191(.A1(new_n8345), .A2(new_n8153), .B(new_n8340), .C(new_n8335), .Y(new_n8448));
  A2O1A1Ixp33_ASAP7_75t_L   g08192(.A1(new_n8341), .A2(new_n8346), .B(new_n8348), .C(new_n8448), .Y(new_n8449));
  NOR2xp33_ASAP7_75t_L      g08193(.A(new_n3674), .B(new_n1517), .Y(new_n8450));
  AOI221xp5_ASAP7_75t_L     g08194(.A1(\b[30] ), .A2(new_n1659), .B1(\b[32] ), .B2(new_n1511), .C(new_n8450), .Y(new_n8451));
  O2A1O1Ixp33_ASAP7_75t_L   g08195(.A1(new_n1521), .A2(new_n3897), .B(new_n8451), .C(new_n1501), .Y(new_n8452));
  INVx1_ASAP7_75t_L         g08196(.A(new_n8452), .Y(new_n8453));
  O2A1O1Ixp33_ASAP7_75t_L   g08197(.A1(new_n1521), .A2(new_n3897), .B(new_n8451), .C(\a[20] ), .Y(new_n8454));
  AOI21xp33_ASAP7_75t_L     g08198(.A1(new_n8453), .A2(\a[20] ), .B(new_n8454), .Y(new_n8455));
  NOR3xp33_ASAP7_75t_L      g08199(.A(new_n8323), .B(new_n8322), .C(new_n8156), .Y(new_n8456));
  O2A1O1Ixp33_ASAP7_75t_L   g08200(.A1(new_n8320), .A2(new_n8324), .B(new_n8153), .C(new_n8456), .Y(new_n8457));
  OAI22xp33_ASAP7_75t_L     g08201(.A1(new_n2089), .A2(new_n2879), .B1(new_n3079), .B2(new_n1962), .Y(new_n8458));
  AOI221xp5_ASAP7_75t_L     g08202(.A1(new_n1955), .A2(\b[29] ), .B1(new_n1964), .B2(new_n3873), .C(new_n8458), .Y(new_n8459));
  XNOR2x2_ASAP7_75t_L       g08203(.A(new_n1952), .B(new_n8459), .Y(new_n8460));
  NAND2xp33_ASAP7_75t_L     g08204(.A(new_n8309), .B(new_n8308), .Y(new_n8461));
  NOR2xp33_ASAP7_75t_L      g08205(.A(new_n8305), .B(new_n8461), .Y(new_n8462));
  O2A1O1Ixp33_ASAP7_75t_L   g08206(.A1(new_n8307), .A2(new_n8306), .B(new_n8313), .C(new_n8462), .Y(new_n8463));
  NAND3xp33_ASAP7_75t_L     g08207(.A(new_n8249), .B(new_n8239), .C(new_n8260), .Y(new_n8464));
  A2O1A1Ixp33_ASAP7_75t_L   g08208(.A1(new_n8252), .A2(new_n8253), .B(new_n8264), .C(new_n8464), .Y(new_n8465));
  NAND2xp33_ASAP7_75t_L     g08209(.A(\b[16] ), .B(new_n4155), .Y(new_n8466));
  OAI221xp5_ASAP7_75t_L     g08210(.A1(new_n4147), .A2(new_n1349), .B1(new_n1043), .B2(new_n4397), .C(new_n8466), .Y(new_n8467));
  A2O1A1Ixp33_ASAP7_75t_L   g08211(.A1(new_n1633), .A2(new_n4151), .B(new_n8467), .C(\a[35] ), .Y(new_n8468));
  AOI211xp5_ASAP7_75t_L     g08212(.A1(new_n1633), .A2(new_n4151), .B(new_n8467), .C(new_n4145), .Y(new_n8469));
  A2O1A1O1Ixp25_ASAP7_75t_L g08213(.A1(new_n4151), .A2(new_n1633), .B(new_n8467), .C(new_n8468), .D(new_n8469), .Y(new_n8470));
  A2O1A1Ixp33_ASAP7_75t_L   g08214(.A1(new_n7968), .A2(new_n8257), .B(new_n8231), .C(new_n8247), .Y(new_n8471));
  OAI21xp33_ASAP7_75t_L     g08215(.A1(new_n8232), .A2(new_n8223), .B(new_n8219), .Y(new_n8472));
  NAND2xp33_ASAP7_75t_L     g08216(.A(new_n8194), .B(new_n8200), .Y(new_n8473));
  O2A1O1Ixp33_ASAP7_75t_L   g08217(.A1(new_n8203), .A2(new_n6439), .B(new_n8205), .C(new_n8473), .Y(new_n8474));
  NOR2xp33_ASAP7_75t_L      g08218(.A(new_n448), .B(new_n7304), .Y(new_n8475));
  AOI221xp5_ASAP7_75t_L     g08219(.A1(\b[6] ), .A2(new_n6742), .B1(\b[8] ), .B2(new_n6442), .C(new_n8475), .Y(new_n8476));
  O2A1O1Ixp33_ASAP7_75t_L   g08220(.A1(new_n6443), .A2(new_n540), .B(new_n8476), .C(new_n6439), .Y(new_n8477));
  INVx1_ASAP7_75t_L         g08221(.A(new_n8477), .Y(new_n8478));
  O2A1O1Ixp33_ASAP7_75t_L   g08222(.A1(new_n6443), .A2(new_n540), .B(new_n8476), .C(\a[44] ), .Y(new_n8479));
  AOI21xp33_ASAP7_75t_L     g08223(.A1(new_n8478), .A2(\a[44] ), .B(new_n8479), .Y(new_n8480));
  OAI21xp33_ASAP7_75t_L     g08224(.A1(new_n8196), .A2(new_n8197), .B(new_n8193), .Y(new_n8481));
  NAND2xp33_ASAP7_75t_L     g08225(.A(\b[2] ), .B(new_n8175), .Y(new_n8482));
  NAND3xp33_ASAP7_75t_L     g08226(.A(new_n7906), .B(new_n8168), .C(new_n8174), .Y(new_n8483));
  INVx1_ASAP7_75t_L         g08227(.A(new_n8483), .Y(new_n8484));
  NAND2xp33_ASAP7_75t_L     g08228(.A(\b[0] ), .B(new_n8484), .Y(new_n8485));
  NAND2xp33_ASAP7_75t_L     g08229(.A(\b[1] ), .B(new_n8169), .Y(new_n8486));
  NOR2xp33_ASAP7_75t_L      g08230(.A(new_n8176), .B(new_n509), .Y(new_n8487));
  INVx1_ASAP7_75t_L         g08231(.A(new_n8487), .Y(new_n8488));
  NAND5xp2_ASAP7_75t_L      g08232(.A(\a[50] ), .B(new_n8485), .C(new_n8488), .D(new_n8486), .E(new_n8482), .Y(new_n8489));
  INVx1_ASAP7_75t_L         g08233(.A(new_n8176), .Y(new_n8490));
  OAI211xp5_ASAP7_75t_L     g08234(.A1(new_n284), .A2(new_n8483), .B(new_n8482), .C(new_n8486), .Y(new_n8491));
  A2O1A1Ixp33_ASAP7_75t_L   g08235(.A1(new_n294), .A2(new_n8490), .B(new_n8491), .C(new_n8172), .Y(new_n8492));
  NAND3xp33_ASAP7_75t_L     g08236(.A(new_n8492), .B(new_n8489), .C(new_n8179), .Y(new_n8493));
  NOR2xp33_ASAP7_75t_L      g08237(.A(new_n8487), .B(new_n8491), .Y(new_n8494));
  NAND4xp25_ASAP7_75t_L     g08238(.A(new_n8494), .B(\a[50] ), .C(new_n8160), .D(new_n8178), .Y(new_n8495));
  NOR2xp33_ASAP7_75t_L      g08239(.A(new_n384), .B(new_n7318), .Y(new_n8496));
  AOI221xp5_ASAP7_75t_L     g08240(.A1(new_n7333), .A2(\b[4] ), .B1(new_n7609), .B2(\b[3] ), .C(new_n8496), .Y(new_n8497));
  OAI211xp5_ASAP7_75t_L     g08241(.A1(new_n7321), .A2(new_n728), .B(\a[47] ), .C(new_n8497), .Y(new_n8498));
  OAI21xp33_ASAP7_75t_L     g08242(.A1(new_n7321), .A2(new_n728), .B(new_n8497), .Y(new_n8499));
  NAND2xp33_ASAP7_75t_L     g08243(.A(new_n7316), .B(new_n8499), .Y(new_n8500));
  AND4x1_ASAP7_75t_L        g08244(.A(new_n8493), .B(new_n8500), .C(new_n8495), .D(new_n8498), .Y(new_n8501));
  AOI22xp33_ASAP7_75t_L     g08245(.A1(new_n8498), .A2(new_n8500), .B1(new_n8495), .B2(new_n8493), .Y(new_n8502));
  OAI21xp33_ASAP7_75t_L     g08246(.A1(new_n8501), .A2(new_n8502), .B(new_n8481), .Y(new_n8503));
  NOR2xp33_ASAP7_75t_L      g08247(.A(new_n8502), .B(new_n8501), .Y(new_n8504));
  NAND3xp33_ASAP7_75t_L     g08248(.A(new_n8194), .B(new_n8504), .C(new_n8193), .Y(new_n8505));
  AOI21xp33_ASAP7_75t_L     g08249(.A1(new_n8505), .A2(new_n8503), .B(new_n8480), .Y(new_n8506));
  INVx1_ASAP7_75t_L         g08250(.A(new_n8479), .Y(new_n8507));
  OAI21xp33_ASAP7_75t_L     g08251(.A1(new_n6439), .A2(new_n8477), .B(new_n8507), .Y(new_n8508));
  O2A1O1Ixp33_ASAP7_75t_L   g08252(.A1(new_n8196), .A2(new_n8197), .B(new_n8193), .C(new_n8504), .Y(new_n8509));
  NOR3xp33_ASAP7_75t_L      g08253(.A(new_n8481), .B(new_n8501), .C(new_n8502), .Y(new_n8510));
  NOR3xp33_ASAP7_75t_L      g08254(.A(new_n8509), .B(new_n8510), .C(new_n8508), .Y(new_n8511));
  NOR2xp33_ASAP7_75t_L      g08255(.A(new_n8506), .B(new_n8511), .Y(new_n8512));
  A2O1A1Ixp33_ASAP7_75t_L   g08256(.A1(new_n8213), .A2(new_n8214), .B(new_n8474), .C(new_n8512), .Y(new_n8513));
  NOR2xp33_ASAP7_75t_L      g08257(.A(new_n8210), .B(new_n8473), .Y(new_n8514));
  O2A1O1Ixp33_ASAP7_75t_L   g08258(.A1(new_n8210), .A2(new_n8514), .B(new_n8214), .C(new_n8474), .Y(new_n8515));
  NOR2xp33_ASAP7_75t_L      g08259(.A(new_n8510), .B(new_n8509), .Y(new_n8516));
  A2O1A1Ixp33_ASAP7_75t_L   g08260(.A1(new_n8478), .A2(\a[44] ), .B(new_n8479), .C(new_n8516), .Y(new_n8517));
  A2O1A1Ixp33_ASAP7_75t_L   g08261(.A1(new_n8517), .A2(new_n8508), .B(new_n8511), .C(new_n8515), .Y(new_n8518));
  NOR2xp33_ASAP7_75t_L      g08262(.A(new_n748), .B(new_n5641), .Y(new_n8519));
  AOI221xp5_ASAP7_75t_L     g08263(.A1(\b[9] ), .A2(new_n5920), .B1(\b[10] ), .B2(new_n5623), .C(new_n8519), .Y(new_n8520));
  O2A1O1Ixp33_ASAP7_75t_L   g08264(.A1(new_n5630), .A2(new_n754), .B(new_n8520), .C(new_n5626), .Y(new_n8521));
  OAI21xp33_ASAP7_75t_L     g08265(.A1(new_n5630), .A2(new_n754), .B(new_n8520), .Y(new_n8522));
  NAND2xp33_ASAP7_75t_L     g08266(.A(new_n5626), .B(new_n8522), .Y(new_n8523));
  OAI21xp33_ASAP7_75t_L     g08267(.A1(new_n5626), .A2(new_n8521), .B(new_n8523), .Y(new_n8524));
  INVx1_ASAP7_75t_L         g08268(.A(new_n8524), .Y(new_n8525));
  NAND3xp33_ASAP7_75t_L     g08269(.A(new_n8518), .B(new_n8513), .C(new_n8525), .Y(new_n8526));
  OAI21xp33_ASAP7_75t_L     g08270(.A1(new_n8510), .A2(new_n8509), .B(new_n8508), .Y(new_n8527));
  NAND3xp33_ASAP7_75t_L     g08271(.A(new_n8505), .B(new_n8503), .C(new_n8480), .Y(new_n8528));
  NAND2xp33_ASAP7_75t_L     g08272(.A(new_n8528), .B(new_n8527), .Y(new_n8529));
  A2O1A1Ixp33_ASAP7_75t_L   g08273(.A1(new_n8213), .A2(new_n8214), .B(new_n8474), .C(new_n8529), .Y(new_n8530));
  O2A1O1Ixp33_ASAP7_75t_L   g08274(.A1(new_n8473), .A2(new_n8206), .B(new_n8215), .C(new_n8529), .Y(new_n8531));
  A2O1A1Ixp33_ASAP7_75t_L   g08275(.A1(new_n8530), .A2(new_n8529), .B(new_n8531), .C(new_n8524), .Y(new_n8532));
  NAND3xp33_ASAP7_75t_L     g08276(.A(new_n8472), .B(new_n8526), .C(new_n8532), .Y(new_n8533));
  AO21x2_ASAP7_75t_L        g08277(.A1(new_n8214), .A2(new_n8213), .B(new_n8474), .Y(new_n8534));
  NAND2xp33_ASAP7_75t_L     g08278(.A(new_n8503), .B(new_n8505), .Y(new_n8535));
  O2A1O1Ixp33_ASAP7_75t_L   g08279(.A1(new_n6439), .A2(new_n8477), .B(new_n8507), .C(new_n8535), .Y(new_n8536));
  O2A1O1Ixp33_ASAP7_75t_L   g08280(.A1(new_n8480), .A2(new_n8536), .B(new_n8528), .C(new_n8534), .Y(new_n8537));
  NOR3xp33_ASAP7_75t_L      g08281(.A(new_n8537), .B(new_n8524), .C(new_n8531), .Y(new_n8538));
  O2A1O1Ixp33_ASAP7_75t_L   g08282(.A1(new_n8473), .A2(new_n8206), .B(new_n8215), .C(new_n8512), .Y(new_n8539));
  O2A1O1Ixp33_ASAP7_75t_L   g08283(.A1(new_n8515), .A2(new_n8539), .B(new_n8518), .C(new_n8525), .Y(new_n8540));
  OAI211xp5_ASAP7_75t_L     g08284(.A1(new_n8540), .A2(new_n8538), .B(new_n8222), .C(new_n8219), .Y(new_n8541));
  NOR2xp33_ASAP7_75t_L      g08285(.A(new_n936), .B(new_n4903), .Y(new_n8542));
  AOI221xp5_ASAP7_75t_L     g08286(.A1(\b[12] ), .A2(new_n5139), .B1(\b[14] ), .B2(new_n4917), .C(new_n8542), .Y(new_n8543));
  INVx1_ASAP7_75t_L         g08287(.A(new_n8543), .Y(new_n8544));
  A2O1A1Ixp33_ASAP7_75t_L   g08288(.A1(new_n971), .A2(new_n4912), .B(new_n8544), .C(\a[38] ), .Y(new_n8545));
  O2A1O1Ixp33_ASAP7_75t_L   g08289(.A1(new_n4911), .A2(new_n1268), .B(new_n8543), .C(\a[38] ), .Y(new_n8546));
  AOI21xp33_ASAP7_75t_L     g08290(.A1(new_n8545), .A2(\a[38] ), .B(new_n8546), .Y(new_n8547));
  NAND3xp33_ASAP7_75t_L     g08291(.A(new_n8533), .B(new_n8547), .C(new_n8541), .Y(new_n8548));
  AOI211xp5_ASAP7_75t_L     g08292(.A1(new_n8222), .A2(new_n8219), .B(new_n8538), .C(new_n8540), .Y(new_n8549));
  AOI211xp5_ASAP7_75t_L     g08293(.A1(new_n8532), .A2(new_n8526), .B(new_n8243), .C(new_n8233), .Y(new_n8550));
  INVx1_ASAP7_75t_L         g08294(.A(new_n8547), .Y(new_n8551));
  OAI21xp33_ASAP7_75t_L     g08295(.A1(new_n8550), .A2(new_n8549), .B(new_n8551), .Y(new_n8552));
  NAND2xp33_ASAP7_75t_L     g08296(.A(new_n8552), .B(new_n8548), .Y(new_n8553));
  NAND2xp33_ASAP7_75t_L     g08297(.A(new_n8471), .B(new_n8553), .Y(new_n8554));
  A2O1A1O1Ixp25_ASAP7_75t_L g08298(.A1(new_n7891), .A2(new_n7960), .B(new_n8158), .C(new_n8245), .D(new_n8237), .Y(new_n8555));
  NAND3xp33_ASAP7_75t_L     g08299(.A(new_n8555), .B(new_n8548), .C(new_n8552), .Y(new_n8556));
  AOI21xp33_ASAP7_75t_L     g08300(.A1(new_n8554), .A2(new_n8556), .B(new_n8470), .Y(new_n8557));
  INVx1_ASAP7_75t_L         g08301(.A(new_n8469), .Y(new_n8558));
  A2O1A1Ixp33_ASAP7_75t_L   g08302(.A1(new_n1633), .A2(new_n4151), .B(new_n8467), .C(new_n4145), .Y(new_n8559));
  NAND2xp33_ASAP7_75t_L     g08303(.A(new_n8559), .B(new_n8558), .Y(new_n8560));
  AOI21xp33_ASAP7_75t_L     g08304(.A1(new_n8552), .A2(new_n8548), .B(new_n8555), .Y(new_n8561));
  NOR2xp33_ASAP7_75t_L      g08305(.A(new_n8471), .B(new_n8553), .Y(new_n8562));
  NOR3xp33_ASAP7_75t_L      g08306(.A(new_n8562), .B(new_n8561), .C(new_n8560), .Y(new_n8563));
  OAI21xp33_ASAP7_75t_L     g08307(.A1(new_n8557), .A2(new_n8563), .B(new_n8465), .Y(new_n8564));
  NOR3xp33_ASAP7_75t_L      g08308(.A(new_n8562), .B(new_n8561), .C(new_n8470), .Y(new_n8565));
  NAND3xp33_ASAP7_75t_L     g08309(.A(new_n8554), .B(new_n8470), .C(new_n8556), .Y(new_n8566));
  O2A1O1Ixp33_ASAP7_75t_L   g08310(.A1(new_n8470), .A2(new_n8565), .B(new_n8566), .C(new_n8465), .Y(new_n8567));
  NOR2xp33_ASAP7_75t_L      g08311(.A(new_n1745), .B(new_n3510), .Y(new_n8568));
  AOI221xp5_ASAP7_75t_L     g08312(.A1(\b[18] ), .A2(new_n3708), .B1(\b[19] ), .B2(new_n3499), .C(new_n8568), .Y(new_n8569));
  OAI21xp33_ASAP7_75t_L     g08313(.A1(new_n3513), .A2(new_n1754), .B(new_n8569), .Y(new_n8570));
  NOR2xp33_ASAP7_75t_L      g08314(.A(new_n3493), .B(new_n8570), .Y(new_n8571));
  O2A1O1Ixp33_ASAP7_75t_L   g08315(.A1(new_n3513), .A2(new_n1754), .B(new_n8569), .C(\a[32] ), .Y(new_n8572));
  NOR2xp33_ASAP7_75t_L      g08316(.A(new_n8572), .B(new_n8571), .Y(new_n8573));
  A2O1A1Ixp33_ASAP7_75t_L   g08317(.A1(new_n8564), .A2(new_n8465), .B(new_n8567), .C(new_n8573), .Y(new_n8574));
  NOR2xp33_ASAP7_75t_L      g08318(.A(new_n8557), .B(new_n8563), .Y(new_n8575));
  NAND2xp33_ASAP7_75t_L     g08319(.A(new_n8465), .B(new_n8575), .Y(new_n8576));
  NOR3xp33_ASAP7_75t_L      g08320(.A(new_n8254), .B(new_n8259), .C(new_n8260), .Y(new_n8577));
  AOI21xp33_ASAP7_75t_L     g08321(.A1(new_n8464), .A2(new_n8260), .B(new_n8577), .Y(new_n8578));
  OAI221xp5_ASAP7_75t_L     g08322(.A1(new_n8557), .A2(new_n8563), .B1(new_n8264), .B2(new_n8578), .C(new_n8464), .Y(new_n8579));
  O2A1O1Ixp33_ASAP7_75t_L   g08323(.A1(new_n3513), .A2(new_n1754), .B(new_n8569), .C(new_n3493), .Y(new_n8580));
  INVx1_ASAP7_75t_L         g08324(.A(new_n8572), .Y(new_n8581));
  OAI21xp33_ASAP7_75t_L     g08325(.A1(new_n3493), .A2(new_n8580), .B(new_n8581), .Y(new_n8582));
  NAND3xp33_ASAP7_75t_L     g08326(.A(new_n8576), .B(new_n8579), .C(new_n8582), .Y(new_n8583));
  NAND2xp33_ASAP7_75t_L     g08327(.A(new_n8574), .B(new_n8583), .Y(new_n8584));
  NAND2xp33_ASAP7_75t_L     g08328(.A(new_n8265), .B(new_n8266), .Y(new_n8585));
  MAJIxp5_ASAP7_75t_L       g08329(.A(new_n8279), .B(new_n8272), .C(new_n8585), .Y(new_n8586));
  NOR2xp33_ASAP7_75t_L      g08330(.A(new_n8584), .B(new_n8586), .Y(new_n8587));
  INVx1_ASAP7_75t_L         g08331(.A(new_n8585), .Y(new_n8588));
  A2O1A1Ixp33_ASAP7_75t_L   g08332(.A1(\a[32] ), .A2(new_n8270), .B(new_n8271), .C(new_n8588), .Y(new_n8589));
  AOI22xp33_ASAP7_75t_L     g08333(.A1(new_n8574), .A2(new_n8583), .B1(new_n8589), .B2(new_n8291), .Y(new_n8590));
  NAND2xp33_ASAP7_75t_L     g08334(.A(\b[22] ), .B(new_n2936), .Y(new_n8591));
  OAI221xp5_ASAP7_75t_L     g08335(.A1(new_n2930), .A2(new_n2188), .B1(new_n1895), .B2(new_n3133), .C(new_n8591), .Y(new_n8592));
  A2O1A1Ixp33_ASAP7_75t_L   g08336(.A1(new_n2679), .A2(new_n2932), .B(new_n8592), .C(\a[29] ), .Y(new_n8593));
  AOI211xp5_ASAP7_75t_L     g08337(.A1(new_n2679), .A2(new_n2932), .B(new_n8592), .C(new_n2928), .Y(new_n8594));
  A2O1A1O1Ixp25_ASAP7_75t_L g08338(.A1(new_n2932), .A2(new_n2679), .B(new_n8592), .C(new_n8593), .D(new_n8594), .Y(new_n8595));
  OAI21xp33_ASAP7_75t_L     g08339(.A1(new_n8587), .A2(new_n8590), .B(new_n8595), .Y(new_n8596));
  NOR3xp33_ASAP7_75t_L      g08340(.A(new_n8278), .B(new_n8280), .C(new_n8285), .Y(new_n8597));
  O2A1O1Ixp33_ASAP7_75t_L   g08341(.A1(new_n8287), .A2(new_n8286), .B(new_n8294), .C(new_n8597), .Y(new_n8598));
  NAND4xp25_ASAP7_75t_L     g08342(.A(new_n8291), .B(new_n8574), .C(new_n8583), .D(new_n8589), .Y(new_n8599));
  A2O1A1Ixp33_ASAP7_75t_L   g08343(.A1(new_n8276), .A2(new_n8588), .B(new_n8280), .C(new_n8584), .Y(new_n8600));
  INVx1_ASAP7_75t_L         g08344(.A(new_n8594), .Y(new_n8601));
  A2O1A1Ixp33_ASAP7_75t_L   g08345(.A1(new_n2679), .A2(new_n2932), .B(new_n8592), .C(new_n2928), .Y(new_n8602));
  NAND2xp33_ASAP7_75t_L     g08346(.A(new_n8602), .B(new_n8601), .Y(new_n8603));
  NAND3xp33_ASAP7_75t_L     g08347(.A(new_n8599), .B(new_n8600), .C(new_n8603), .Y(new_n8604));
  AOI21xp33_ASAP7_75t_L     g08348(.A1(new_n8596), .A2(new_n8604), .B(new_n8598), .Y(new_n8605));
  NAND2xp33_ASAP7_75t_L     g08349(.A(new_n8298), .B(new_n8299), .Y(new_n8606));
  NOR3xp33_ASAP7_75t_L      g08350(.A(new_n8590), .B(new_n8595), .C(new_n8587), .Y(new_n8607));
  A2O1A1O1Ixp25_ASAP7_75t_L g08351(.A1(new_n8294), .A2(new_n8606), .B(new_n8597), .C(new_n8596), .D(new_n8607), .Y(new_n8608));
  NAND2xp33_ASAP7_75t_L     g08352(.A(\b[25] ), .B(new_n2421), .Y(new_n8609));
  OAI221xp5_ASAP7_75t_L     g08353(.A1(new_n2415), .A2(new_n2703), .B1(new_n2205), .B2(new_n2572), .C(new_n8609), .Y(new_n8610));
  A2O1A1Ixp33_ASAP7_75t_L   g08354(.A1(new_n2709), .A2(new_n2417), .B(new_n8610), .C(\a[26] ), .Y(new_n8611));
  AOI211xp5_ASAP7_75t_L     g08355(.A1(new_n2709), .A2(new_n2417), .B(new_n8610), .C(new_n2413), .Y(new_n8612));
  A2O1A1O1Ixp25_ASAP7_75t_L g08356(.A1(new_n2709), .A2(new_n2417), .B(new_n8610), .C(new_n8611), .D(new_n8612), .Y(new_n8613));
  INVx1_ASAP7_75t_L         g08357(.A(new_n8613), .Y(new_n8614));
  AOI211xp5_ASAP7_75t_L     g08358(.A1(new_n8608), .A2(new_n8596), .B(new_n8605), .C(new_n8614), .Y(new_n8615));
  INVx1_ASAP7_75t_L         g08359(.A(new_n8597), .Y(new_n8616));
  MAJIxp5_ASAP7_75t_L       g08360(.A(new_n8015), .B(new_n8296), .C(new_n7999), .Y(new_n8617));
  AOI21xp33_ASAP7_75t_L     g08361(.A1(new_n8599), .A2(new_n8600), .B(new_n8603), .Y(new_n8618));
  A2O1A1O1Ixp25_ASAP7_75t_L g08362(.A1(new_n8298), .A2(new_n8285), .B(new_n8617), .C(new_n8616), .D(new_n8618), .Y(new_n8619));
  NAND3xp33_ASAP7_75t_L     g08363(.A(new_n8598), .B(new_n8604), .C(new_n8596), .Y(new_n8620));
  A2O1A1O1Ixp25_ASAP7_75t_L g08364(.A1(new_n8604), .A2(new_n8619), .B(new_n8598), .C(new_n8620), .D(new_n8613), .Y(new_n8621));
  NOR3xp33_ASAP7_75t_L      g08365(.A(new_n8463), .B(new_n8615), .C(new_n8621), .Y(new_n8622));
  MAJIxp5_ASAP7_75t_L       g08366(.A(new_n8318), .B(new_n8305), .C(new_n8461), .Y(new_n8623));
  A2O1A1Ixp33_ASAP7_75t_L   g08367(.A1(new_n8285), .A2(new_n8298), .B(new_n8617), .C(new_n8616), .Y(new_n8624));
  OAI21xp33_ASAP7_75t_L     g08368(.A1(new_n8607), .A2(new_n8618), .B(new_n8624), .Y(new_n8625));
  NAND3xp33_ASAP7_75t_L     g08369(.A(new_n8625), .B(new_n8620), .C(new_n8613), .Y(new_n8626));
  A2O1A1Ixp33_ASAP7_75t_L   g08370(.A1(new_n8608), .A2(new_n8596), .B(new_n8605), .C(new_n8614), .Y(new_n8627));
  AOI21xp33_ASAP7_75t_L     g08371(.A1(new_n8627), .A2(new_n8626), .B(new_n8623), .Y(new_n8628));
  OAI21xp33_ASAP7_75t_L     g08372(.A1(new_n8628), .A2(new_n8622), .B(new_n8460), .Y(new_n8629));
  AND2x2_ASAP7_75t_L        g08373(.A(\a[23] ), .B(new_n8459), .Y(new_n8630));
  NOR2xp33_ASAP7_75t_L      g08374(.A(\a[23] ), .B(new_n8459), .Y(new_n8631));
  NAND3xp33_ASAP7_75t_L     g08375(.A(new_n8623), .B(new_n8626), .C(new_n8627), .Y(new_n8632));
  OAI21xp33_ASAP7_75t_L     g08376(.A1(new_n8615), .A2(new_n8621), .B(new_n8463), .Y(new_n8633));
  OAI211xp5_ASAP7_75t_L     g08377(.A1(new_n8631), .A2(new_n8630), .B(new_n8632), .C(new_n8633), .Y(new_n8634));
  NAND2xp33_ASAP7_75t_L     g08378(.A(new_n8634), .B(new_n8629), .Y(new_n8635));
  NOR2xp33_ASAP7_75t_L      g08379(.A(new_n8457), .B(new_n8635), .Y(new_n8636));
  AOI221xp5_ASAP7_75t_L     g08380(.A1(new_n8338), .A2(new_n8153), .B1(new_n8634), .B2(new_n8629), .C(new_n8456), .Y(new_n8637));
  OAI21xp33_ASAP7_75t_L     g08381(.A1(new_n8637), .A2(new_n8636), .B(new_n8455), .Y(new_n8638));
  INVx1_ASAP7_75t_L         g08382(.A(new_n8455), .Y(new_n8639));
  AOI21xp33_ASAP7_75t_L     g08383(.A1(new_n8036), .A2(new_n8038), .B(new_n8040), .Y(new_n8640));
  INVx1_ASAP7_75t_L         g08384(.A(new_n8456), .Y(new_n8641));
  OAI21xp33_ASAP7_75t_L     g08385(.A1(new_n8640), .A2(new_n8325), .B(new_n8641), .Y(new_n8642));
  NAND3xp33_ASAP7_75t_L     g08386(.A(new_n8642), .B(new_n8629), .C(new_n8634), .Y(new_n8643));
  INVx1_ASAP7_75t_L         g08387(.A(new_n8637), .Y(new_n8644));
  NAND3xp33_ASAP7_75t_L     g08388(.A(new_n8644), .B(new_n8643), .C(new_n8639), .Y(new_n8645));
  NAND3xp33_ASAP7_75t_L     g08389(.A(new_n8449), .B(new_n8638), .C(new_n8645), .Y(new_n8646));
  O2A1O1Ixp33_ASAP7_75t_L   g08390(.A1(new_n8156), .A2(new_n8456), .B(new_n8328), .C(new_n8640), .Y(new_n8647));
  O2A1O1Ixp33_ASAP7_75t_L   g08391(.A1(new_n8640), .A2(new_n8647), .B(new_n8329), .C(new_n8341), .Y(new_n8648));
  O2A1O1Ixp33_ASAP7_75t_L   g08392(.A1(new_n8336), .A2(new_n8335), .B(new_n8343), .C(new_n8648), .Y(new_n8649));
  AOI21xp33_ASAP7_75t_L     g08393(.A1(new_n8644), .A2(new_n8643), .B(new_n8639), .Y(new_n8650));
  NOR3xp33_ASAP7_75t_L      g08394(.A(new_n8636), .B(new_n8637), .C(new_n8455), .Y(new_n8651));
  OAI21xp33_ASAP7_75t_L     g08395(.A1(new_n8650), .A2(new_n8651), .B(new_n8649), .Y(new_n8652));
  NOR2xp33_ASAP7_75t_L      g08396(.A(new_n4344), .B(new_n2118), .Y(new_n8653));
  AOI221xp5_ASAP7_75t_L     g08397(.A1(\b[33] ), .A2(new_n1290), .B1(\b[35] ), .B2(new_n1209), .C(new_n8653), .Y(new_n8654));
  O2A1O1Ixp33_ASAP7_75t_L   g08398(.A1(new_n1210), .A2(new_n4589), .B(new_n8654), .C(new_n1206), .Y(new_n8655));
  INVx1_ASAP7_75t_L         g08399(.A(new_n8655), .Y(new_n8656));
  O2A1O1Ixp33_ASAP7_75t_L   g08400(.A1(new_n1210), .A2(new_n4589), .B(new_n8654), .C(\a[17] ), .Y(new_n8657));
  AOI21xp33_ASAP7_75t_L     g08401(.A1(new_n8656), .A2(\a[17] ), .B(new_n8657), .Y(new_n8658));
  NAND3xp33_ASAP7_75t_L     g08402(.A(new_n8646), .B(new_n8652), .C(new_n8658), .Y(new_n8659));
  NOR3xp33_ASAP7_75t_L      g08403(.A(new_n8649), .B(new_n8650), .C(new_n8651), .Y(new_n8660));
  AOI21xp33_ASAP7_75t_L     g08404(.A1(new_n8645), .A2(new_n8638), .B(new_n8449), .Y(new_n8661));
  INVx1_ASAP7_75t_L         g08405(.A(new_n8658), .Y(new_n8662));
  OAI21xp33_ASAP7_75t_L     g08406(.A1(new_n8661), .A2(new_n8660), .B(new_n8662), .Y(new_n8663));
  AND2x2_ASAP7_75t_L        g08407(.A(new_n8659), .B(new_n8663), .Y(new_n8664));
  INVx1_ASAP7_75t_L         g08408(.A(new_n8365), .Y(new_n8665));
  O2A1O1Ixp33_ASAP7_75t_L   g08409(.A1(new_n8356), .A2(new_n8360), .B(new_n8367), .C(new_n8665), .Y(new_n8666));
  NAND2xp33_ASAP7_75t_L     g08410(.A(new_n8666), .B(new_n8664), .Y(new_n8667));
  NAND2xp33_ASAP7_75t_L     g08411(.A(new_n8659), .B(new_n8663), .Y(new_n8668));
  OAI21xp33_ASAP7_75t_L     g08412(.A1(new_n8361), .A2(new_n8363), .B(new_n8365), .Y(new_n8669));
  NAND2xp33_ASAP7_75t_L     g08413(.A(new_n8668), .B(new_n8669), .Y(new_n8670));
  OAI22xp33_ASAP7_75t_L     g08414(.A1(new_n980), .A2(new_n4613), .B1(new_n5074), .B2(new_n864), .Y(new_n8671));
  AOI221xp5_ASAP7_75t_L     g08415(.A1(new_n886), .A2(\b[38] ), .B1(new_n873), .B2(new_n6083), .C(new_n8671), .Y(new_n8672));
  XNOR2x2_ASAP7_75t_L       g08416(.A(\a[14] ), .B(new_n8672), .Y(new_n8673));
  INVx1_ASAP7_75t_L         g08417(.A(new_n8673), .Y(new_n8674));
  NAND3xp33_ASAP7_75t_L     g08418(.A(new_n8674), .B(new_n8670), .C(new_n8667), .Y(new_n8675));
  NOR2xp33_ASAP7_75t_L      g08419(.A(new_n8668), .B(new_n8669), .Y(new_n8676));
  NOR3xp33_ASAP7_75t_L      g08420(.A(new_n8660), .B(new_n8661), .C(new_n8658), .Y(new_n8677));
  O2A1O1Ixp33_ASAP7_75t_L   g08421(.A1(new_n8658), .A2(new_n8677), .B(new_n8659), .C(new_n8666), .Y(new_n8678));
  OAI21xp33_ASAP7_75t_L     g08422(.A1(new_n8676), .A2(new_n8678), .B(new_n8673), .Y(new_n8679));
  NAND4xp25_ASAP7_75t_L     g08423(.A(new_n8389), .B(new_n8675), .C(new_n8679), .D(new_n8447), .Y(new_n8680));
  NOR3xp33_ASAP7_75t_L      g08424(.A(new_n8678), .B(new_n8676), .C(new_n8673), .Y(new_n8681));
  AOI21xp33_ASAP7_75t_L     g08425(.A1(new_n8667), .A2(new_n8670), .B(new_n8674), .Y(new_n8682));
  A2O1A1Ixp33_ASAP7_75t_L   g08426(.A1(new_n8375), .A2(new_n8376), .B(new_n8377), .C(new_n8447), .Y(new_n8683));
  OAI21xp33_ASAP7_75t_L     g08427(.A1(new_n8681), .A2(new_n8682), .B(new_n8683), .Y(new_n8684));
  NOR2xp33_ASAP7_75t_L      g08428(.A(new_n5570), .B(new_n712), .Y(new_n8685));
  AOI221xp5_ASAP7_75t_L     g08429(.A1(\b[41] ), .A2(new_n640), .B1(new_n635), .B2(\b[40] ), .C(new_n8685), .Y(new_n8686));
  OA21x2_ASAP7_75t_L        g08430(.A1(new_n641), .A2(new_n6117), .B(new_n8686), .Y(new_n8687));
  O2A1O1Ixp33_ASAP7_75t_L   g08431(.A1(new_n641), .A2(new_n6117), .B(new_n8686), .C(new_n637), .Y(new_n8688));
  NAND2xp33_ASAP7_75t_L     g08432(.A(\a[11] ), .B(new_n8687), .Y(new_n8689));
  OA21x2_ASAP7_75t_L        g08433(.A1(new_n8687), .A2(new_n8688), .B(new_n8689), .Y(new_n8690));
  NAND3xp33_ASAP7_75t_L     g08434(.A(new_n8680), .B(new_n8684), .C(new_n8690), .Y(new_n8691));
  NOR3xp33_ASAP7_75t_L      g08435(.A(new_n8683), .B(new_n8682), .C(new_n8681), .Y(new_n8692));
  OA21x2_ASAP7_75t_L        g08436(.A1(new_n8681), .A2(new_n8682), .B(new_n8683), .Y(new_n8693));
  INVx1_ASAP7_75t_L         g08437(.A(new_n8690), .Y(new_n8694));
  OAI21xp33_ASAP7_75t_L     g08438(.A1(new_n8692), .A2(new_n8693), .B(new_n8694), .Y(new_n8695));
  NAND2xp33_ASAP7_75t_L     g08439(.A(new_n8691), .B(new_n8695), .Y(new_n8696));
  NOR2xp33_ASAP7_75t_L      g08440(.A(new_n8379), .B(new_n8378), .Y(new_n8697));
  A2O1A1Ixp33_ASAP7_75t_L   g08441(.A1(\a[11] ), .A2(new_n8383), .B(new_n8384), .C(new_n8697), .Y(new_n8698));
  A2O1A1Ixp33_ASAP7_75t_L   g08442(.A1(new_n8111), .A2(new_n8151), .B(new_n8391), .C(new_n8698), .Y(new_n8699));
  NOR2xp33_ASAP7_75t_L      g08443(.A(new_n8696), .B(new_n8699), .Y(new_n8700));
  MAJIxp5_ASAP7_75t_L       g08444(.A(new_n8396), .B(new_n8697), .C(new_n8386), .Y(new_n8701));
  AOI21xp33_ASAP7_75t_L     g08445(.A1(new_n8695), .A2(new_n8691), .B(new_n8701), .Y(new_n8702));
  NOR2xp33_ASAP7_75t_L      g08446(.A(new_n6378), .B(new_n506), .Y(new_n8703));
  AOI221xp5_ASAP7_75t_L     g08447(.A1(\b[44] ), .A2(new_n475), .B1(new_n470), .B2(\b[43] ), .C(new_n8703), .Y(new_n8704));
  O2A1O1Ixp33_ASAP7_75t_L   g08448(.A1(new_n477), .A2(new_n6951), .B(new_n8704), .C(new_n466), .Y(new_n8705));
  OAI21xp33_ASAP7_75t_L     g08449(.A1(new_n477), .A2(new_n6951), .B(new_n8704), .Y(new_n8706));
  NAND2xp33_ASAP7_75t_L     g08450(.A(new_n466), .B(new_n8706), .Y(new_n8707));
  OAI21xp33_ASAP7_75t_L     g08451(.A1(new_n466), .A2(new_n8705), .B(new_n8707), .Y(new_n8708));
  INVx1_ASAP7_75t_L         g08452(.A(new_n8708), .Y(new_n8709));
  OAI21xp33_ASAP7_75t_L     g08453(.A1(new_n8702), .A2(new_n8700), .B(new_n8709), .Y(new_n8710));
  NOR2xp33_ASAP7_75t_L      g08454(.A(new_n8405), .B(new_n8406), .Y(new_n8711));
  A2O1A1Ixp33_ASAP7_75t_L   g08455(.A1(\a[8] ), .A2(new_n8401), .B(new_n8402), .C(new_n8711), .Y(new_n8712));
  NAND3xp33_ASAP7_75t_L     g08456(.A(new_n8701), .B(new_n8695), .C(new_n8691), .Y(new_n8713));
  INVx1_ASAP7_75t_L         g08457(.A(new_n8698), .Y(new_n8714));
  A2O1A1Ixp33_ASAP7_75t_L   g08458(.A1(new_n8395), .A2(new_n8396), .B(new_n8714), .C(new_n8696), .Y(new_n8715));
  NAND3xp33_ASAP7_75t_L     g08459(.A(new_n8715), .B(new_n8713), .C(new_n8708), .Y(new_n8716));
  AOI22xp33_ASAP7_75t_L     g08460(.A1(new_n8716), .A2(new_n8710), .B1(new_n8712), .B2(new_n8417), .Y(new_n8717));
  NAND2xp33_ASAP7_75t_L     g08461(.A(new_n8397), .B(new_n8392), .Y(new_n8718));
  INVx1_ASAP7_75t_L         g08462(.A(new_n8402), .Y(new_n8719));
  O2A1O1Ixp33_ASAP7_75t_L   g08463(.A1(new_n8400), .A2(new_n466), .B(new_n8719), .C(new_n8718), .Y(new_n8720));
  NAND2xp33_ASAP7_75t_L     g08464(.A(new_n8404), .B(new_n8408), .Y(new_n8721));
  NOR3xp33_ASAP7_75t_L      g08465(.A(new_n8700), .B(new_n8702), .C(new_n8709), .Y(new_n8722));
  A2O1A1O1Ixp25_ASAP7_75t_L g08466(.A1(new_n8416), .A2(new_n8721), .B(new_n8720), .C(new_n8710), .D(new_n8722), .Y(new_n8723));
  NOR2xp33_ASAP7_75t_L      g08467(.A(new_n7249), .B(new_n375), .Y(new_n8724));
  AOI221xp5_ASAP7_75t_L     g08468(.A1(\b[47] ), .A2(new_n361), .B1(new_n349), .B2(\b[46] ), .C(new_n8724), .Y(new_n8725));
  INVx1_ASAP7_75t_L         g08469(.A(new_n7560), .Y(new_n8726));
  NAND2xp33_ASAP7_75t_L     g08470(.A(new_n359), .B(new_n8726), .Y(new_n8727));
  O2A1O1Ixp33_ASAP7_75t_L   g08471(.A1(new_n356), .A2(new_n7560), .B(new_n8725), .C(new_n346), .Y(new_n8728));
  OA21x2_ASAP7_75t_L        g08472(.A1(new_n356), .A2(new_n7560), .B(new_n8725), .Y(new_n8729));
  NAND2xp33_ASAP7_75t_L     g08473(.A(\a[5] ), .B(new_n8729), .Y(new_n8730));
  A2O1A1Ixp33_ASAP7_75t_L   g08474(.A1(new_n8727), .A2(new_n8725), .B(new_n8728), .C(new_n8730), .Y(new_n8731));
  INVx1_ASAP7_75t_L         g08475(.A(new_n8731), .Y(new_n8732));
  A2O1A1Ixp33_ASAP7_75t_L   g08476(.A1(new_n8723), .A2(new_n8710), .B(new_n8717), .C(new_n8732), .Y(new_n8733));
  MAJIxp5_ASAP7_75t_L       g08477(.A(new_n8411), .B(new_n8403), .C(new_n8718), .Y(new_n8734));
  AOI21xp33_ASAP7_75t_L     g08478(.A1(new_n8715), .A2(new_n8713), .B(new_n8708), .Y(new_n8735));
  OAI21xp33_ASAP7_75t_L     g08479(.A1(new_n8722), .A2(new_n8735), .B(new_n8734), .Y(new_n8736));
  NAND4xp25_ASAP7_75t_L     g08480(.A(new_n8417), .B(new_n8716), .C(new_n8710), .D(new_n8712), .Y(new_n8737));
  NAND3xp33_ASAP7_75t_L     g08481(.A(new_n8737), .B(new_n8736), .C(new_n8731), .Y(new_n8738));
  NAND2xp33_ASAP7_75t_L     g08482(.A(new_n8412), .B(new_n8417), .Y(new_n8739));
  NOR2xp33_ASAP7_75t_L      g08483(.A(new_n8420), .B(new_n8739), .Y(new_n8740));
  O2A1O1Ixp33_ASAP7_75t_L   g08484(.A1(new_n8421), .A2(new_n8422), .B(new_n8423), .C(new_n8740), .Y(new_n8741));
  NAND3xp33_ASAP7_75t_L     g08485(.A(new_n8741), .B(new_n8738), .C(new_n8733), .Y(new_n8742));
  INVx1_ASAP7_75t_L         g08486(.A(new_n8734), .Y(new_n8743));
  A2O1A1O1Ixp25_ASAP7_75t_L g08487(.A1(new_n8404), .A2(new_n8403), .B(new_n8411), .C(new_n8712), .D(new_n8735), .Y(new_n8744));
  A2O1A1O1Ixp25_ASAP7_75t_L g08488(.A1(new_n8716), .A2(new_n8744), .B(new_n8743), .C(new_n8737), .D(new_n8731), .Y(new_n8745));
  INVx1_ASAP7_75t_L         g08489(.A(new_n8738), .Y(new_n8746));
  A2O1A1O1Ixp25_ASAP7_75t_L g08490(.A1(new_n7842), .A2(new_n8141), .B(new_n7841), .C(new_n8143), .D(new_n8131), .Y(new_n8747));
  MAJIxp5_ASAP7_75t_L       g08491(.A(new_n8747), .B(new_n8739), .C(new_n8420), .Y(new_n8748));
  OAI21xp33_ASAP7_75t_L     g08492(.A1(new_n8745), .A2(new_n8746), .B(new_n8748), .Y(new_n8749));
  NAND2xp33_ASAP7_75t_L     g08493(.A(new_n8749), .B(new_n8742), .Y(new_n8750));
  NOR2xp33_ASAP7_75t_L      g08494(.A(new_n7860), .B(new_n287), .Y(new_n8751));
  AOI221xp5_ASAP7_75t_L     g08495(.A1(\b[49] ), .A2(new_n264), .B1(\b[50] ), .B2(new_n283), .C(new_n8751), .Y(new_n8752));
  INVx1_ASAP7_75t_L         g08496(.A(new_n8431), .Y(new_n8753));
  NOR2xp33_ASAP7_75t_L      g08497(.A(\b[49] ), .B(\b[50] ), .Y(new_n8754));
  INVx1_ASAP7_75t_L         g08498(.A(\b[50] ), .Y(new_n8755));
  NOR2xp33_ASAP7_75t_L      g08499(.A(new_n8427), .B(new_n8755), .Y(new_n8756));
  NOR2xp33_ASAP7_75t_L      g08500(.A(new_n8754), .B(new_n8756), .Y(new_n8757));
  INVx1_ASAP7_75t_L         g08501(.A(new_n8757), .Y(new_n8758));
  O2A1O1Ixp33_ASAP7_75t_L   g08502(.A1(new_n8430), .A2(new_n8435), .B(new_n8753), .C(new_n8758), .Y(new_n8759));
  INVx1_ASAP7_75t_L         g08503(.A(new_n7861), .Y(new_n8760));
  A2O1A1Ixp33_ASAP7_75t_L   g08504(.A1(new_n7865), .A2(new_n8760), .B(new_n8430), .C(new_n8753), .Y(new_n8761));
  NOR2xp33_ASAP7_75t_L      g08505(.A(new_n8757), .B(new_n8761), .Y(new_n8762));
  NOR2xp33_ASAP7_75t_L      g08506(.A(new_n8759), .B(new_n8762), .Y(new_n8763));
  INVx1_ASAP7_75t_L         g08507(.A(new_n8763), .Y(new_n8764));
  O2A1O1Ixp33_ASAP7_75t_L   g08508(.A1(new_n279), .A2(new_n8764), .B(new_n8752), .C(new_n257), .Y(new_n8765));
  O2A1O1Ixp33_ASAP7_75t_L   g08509(.A1(new_n279), .A2(new_n8764), .B(new_n8752), .C(\a[2] ), .Y(new_n8766));
  INVx1_ASAP7_75t_L         g08510(.A(new_n8766), .Y(new_n8767));
  O2A1O1Ixp33_ASAP7_75t_L   g08511(.A1(new_n8765), .A2(new_n257), .B(new_n8767), .C(new_n8750), .Y(new_n8768));
  INVx1_ASAP7_75t_L         g08512(.A(new_n8765), .Y(new_n8769));
  A2O1A1Ixp33_ASAP7_75t_L   g08513(.A1(\a[2] ), .A2(new_n8769), .B(new_n8766), .C(new_n8750), .Y(new_n8770));
  A2O1A1O1Ixp25_ASAP7_75t_L g08514(.A1(new_n8146), .A2(new_n7855), .B(new_n8145), .C(new_n8442), .D(new_n8443), .Y(new_n8771));
  O2A1O1Ixp33_ASAP7_75t_L   g08515(.A1(new_n8750), .A2(new_n8768), .B(new_n8770), .C(new_n8771), .Y(new_n8772));
  OAI21xp33_ASAP7_75t_L     g08516(.A1(new_n8750), .A2(new_n8768), .B(new_n8770), .Y(new_n8773));
  INVx1_ASAP7_75t_L         g08517(.A(new_n8771), .Y(new_n8774));
  NOR2xp33_ASAP7_75t_L      g08518(.A(new_n8774), .B(new_n8773), .Y(new_n8775));
  NOR2xp33_ASAP7_75t_L      g08519(.A(new_n8772), .B(new_n8775), .Y(\f[50] ));
  AOI21xp33_ASAP7_75t_L     g08520(.A1(new_n8769), .A2(\a[2] ), .B(new_n8766), .Y(new_n8777));
  MAJIxp5_ASAP7_75t_L       g08521(.A(new_n8771), .B(new_n8750), .C(new_n8777), .Y(new_n8778));
  INVx1_ASAP7_75t_L         g08522(.A(\b[51] ), .Y(new_n8779));
  NAND2xp33_ASAP7_75t_L     g08523(.A(\b[49] ), .B(new_n286), .Y(new_n8780));
  OAI221xp5_ASAP7_75t_L     g08524(.A1(new_n285), .A2(new_n8755), .B1(new_n8779), .B2(new_n269), .C(new_n8780), .Y(new_n8781));
  NOR2xp33_ASAP7_75t_L      g08525(.A(\b[50] ), .B(\b[51] ), .Y(new_n8782));
  NOR2xp33_ASAP7_75t_L      g08526(.A(new_n8755), .B(new_n8779), .Y(new_n8783));
  NOR2xp33_ASAP7_75t_L      g08527(.A(new_n8782), .B(new_n8783), .Y(new_n8784));
  A2O1A1Ixp33_ASAP7_75t_L   g08528(.A1(new_n8761), .A2(new_n8757), .B(new_n8756), .C(new_n8784), .Y(new_n8785));
  INVx1_ASAP7_75t_L         g08529(.A(new_n8756), .Y(new_n8786));
  INVx1_ASAP7_75t_L         g08530(.A(new_n8759), .Y(new_n8787));
  OAI211xp5_ASAP7_75t_L     g08531(.A1(new_n8782), .A2(new_n8783), .B(new_n8787), .C(new_n8786), .Y(new_n8788));
  NAND2xp33_ASAP7_75t_L     g08532(.A(new_n8785), .B(new_n8788), .Y(new_n8789));
  INVx1_ASAP7_75t_L         g08533(.A(new_n8789), .Y(new_n8790));
  A2O1A1Ixp33_ASAP7_75t_L   g08534(.A1(new_n8790), .A2(new_n273), .B(new_n8781), .C(\a[2] ), .Y(new_n8791));
  AOI211xp5_ASAP7_75t_L     g08535(.A1(new_n8790), .A2(new_n273), .B(new_n8781), .C(new_n257), .Y(new_n8792));
  A2O1A1O1Ixp25_ASAP7_75t_L g08536(.A1(new_n273), .A2(new_n8790), .B(new_n8781), .C(new_n8791), .D(new_n8792), .Y(new_n8793));
  A2O1A1O1Ixp25_ASAP7_75t_L g08537(.A1(new_n8716), .A2(new_n8744), .B(new_n8743), .C(new_n8737), .D(new_n8732), .Y(new_n8794));
  INVx1_ASAP7_75t_L         g08538(.A(new_n8794), .Y(new_n8795));
  A2O1A1Ixp33_ASAP7_75t_L   g08539(.A1(new_n8417), .A2(new_n8712), .B(new_n8735), .C(new_n8716), .Y(new_n8796));
  XNOR2x2_ASAP7_75t_L       g08540(.A(new_n8666), .B(new_n8668), .Y(new_n8797));
  NAND2xp33_ASAP7_75t_L     g08541(.A(new_n8673), .B(new_n8797), .Y(new_n8798));
  INVx1_ASAP7_75t_L         g08542(.A(new_n8677), .Y(new_n8799));
  A2O1A1Ixp33_ASAP7_75t_L   g08543(.A1(new_n8358), .A2(new_n8448), .B(new_n8650), .C(new_n8645), .Y(new_n8800));
  NOR3xp33_ASAP7_75t_L      g08544(.A(new_n8622), .B(new_n8628), .C(new_n8460), .Y(new_n8801));
  A2O1A1O1Ixp25_ASAP7_75t_L g08545(.A1(new_n8153), .A2(new_n8338), .B(new_n8456), .C(new_n8629), .D(new_n8801), .Y(new_n8802));
  NAND2xp33_ASAP7_75t_L     g08546(.A(new_n8315), .B(new_n8316), .Y(new_n8803));
  A2O1A1O1Ixp25_ASAP7_75t_L g08547(.A1(new_n8313), .A2(new_n8803), .B(new_n8462), .C(new_n8626), .D(new_n8621), .Y(new_n8804));
  OAI21xp33_ASAP7_75t_L     g08548(.A1(new_n8561), .A2(new_n8562), .B(new_n8560), .Y(new_n8805));
  NAND2xp33_ASAP7_75t_L     g08549(.A(new_n8566), .B(new_n8805), .Y(new_n8806));
  NOR2xp33_ASAP7_75t_L      g08550(.A(new_n1349), .B(new_n4142), .Y(new_n8807));
  AOI221xp5_ASAP7_75t_L     g08551(.A1(\b[16] ), .A2(new_n4402), .B1(\b[18] ), .B2(new_n4156), .C(new_n8807), .Y(new_n8808));
  O2A1O1Ixp33_ASAP7_75t_L   g08552(.A1(new_n4150), .A2(new_n1464), .B(new_n8808), .C(new_n4145), .Y(new_n8809));
  INVx1_ASAP7_75t_L         g08553(.A(new_n8808), .Y(new_n8810));
  A2O1A1Ixp33_ASAP7_75t_L   g08554(.A1(new_n2329), .A2(new_n4151), .B(new_n8810), .C(new_n4145), .Y(new_n8811));
  OAI21xp33_ASAP7_75t_L     g08555(.A1(new_n4145), .A2(new_n8809), .B(new_n8811), .Y(new_n8812));
  NAND2xp33_ASAP7_75t_L     g08556(.A(new_n8541), .B(new_n8533), .Y(new_n8813));
  NOR2xp33_ASAP7_75t_L      g08557(.A(new_n8547), .B(new_n8813), .Y(new_n8814));
  NOR2xp33_ASAP7_75t_L      g08558(.A(new_n960), .B(new_n4903), .Y(new_n8815));
  AOI221xp5_ASAP7_75t_L     g08559(.A1(\b[13] ), .A2(new_n5139), .B1(\b[15] ), .B2(new_n4917), .C(new_n8815), .Y(new_n8816));
  INVx1_ASAP7_75t_L         g08560(.A(new_n8816), .Y(new_n8817));
  A2O1A1Ixp33_ASAP7_75t_L   g08561(.A1(new_n1052), .A2(new_n4912), .B(new_n8817), .C(\a[38] ), .Y(new_n8818));
  O2A1O1Ixp33_ASAP7_75t_L   g08562(.A1(new_n4911), .A2(new_n1774), .B(new_n8816), .C(\a[38] ), .Y(new_n8819));
  AOI21xp33_ASAP7_75t_L     g08563(.A1(new_n8818), .A2(\a[38] ), .B(new_n8819), .Y(new_n8820));
  A2O1A1Ixp33_ASAP7_75t_L   g08564(.A1(new_n8222), .A2(new_n8219), .B(new_n8538), .C(new_n8532), .Y(new_n8821));
  NOR2xp33_ASAP7_75t_L      g08565(.A(new_n833), .B(new_n5641), .Y(new_n8822));
  AOI221xp5_ASAP7_75t_L     g08566(.A1(\b[10] ), .A2(new_n5920), .B1(\b[11] ), .B2(new_n5623), .C(new_n8822), .Y(new_n8823));
  O2A1O1Ixp33_ASAP7_75t_L   g08567(.A1(new_n5630), .A2(new_n841), .B(new_n8823), .C(new_n5626), .Y(new_n8824));
  OAI21xp33_ASAP7_75t_L     g08568(.A1(new_n5630), .A2(new_n841), .B(new_n8823), .Y(new_n8825));
  NAND2xp33_ASAP7_75t_L     g08569(.A(new_n5626), .B(new_n8825), .Y(new_n8826));
  OAI21xp33_ASAP7_75t_L     g08570(.A1(new_n5626), .A2(new_n8824), .B(new_n8826), .Y(new_n8827));
  A2O1A1O1Ixp25_ASAP7_75t_L g08571(.A1(new_n8213), .A2(new_n8214), .B(new_n8474), .C(new_n8529), .D(new_n8536), .Y(new_n8828));
  NAND2xp33_ASAP7_75t_L     g08572(.A(new_n8495), .B(new_n8493), .Y(new_n8829));
  O2A1O1Ixp33_ASAP7_75t_L   g08573(.A1(new_n7321), .A2(new_n728), .B(new_n8497), .C(new_n7316), .Y(new_n8830));
  O2A1O1Ixp33_ASAP7_75t_L   g08574(.A1(new_n8830), .A2(new_n7316), .B(new_n8500), .C(new_n8829), .Y(new_n8831));
  INVx1_ASAP7_75t_L         g08575(.A(new_n8831), .Y(new_n8832));
  NOR5xp2_ASAP7_75t_L       g08576(.A(new_n8182), .B(new_n8491), .C(new_n8487), .D(new_n7907), .E(new_n8172), .Y(new_n8833));
  INVx1_ASAP7_75t_L         g08577(.A(\a[51] ), .Y(new_n8834));
  NAND2xp33_ASAP7_75t_L     g08578(.A(\a[50] ), .B(new_n8834), .Y(new_n8835));
  NAND2xp33_ASAP7_75t_L     g08579(.A(\a[51] ), .B(new_n8172), .Y(new_n8836));
  AND2x2_ASAP7_75t_L        g08580(.A(new_n8835), .B(new_n8836), .Y(new_n8837));
  NOR2xp33_ASAP7_75t_L      g08581(.A(new_n284), .B(new_n8837), .Y(new_n8838));
  INVx1_ASAP7_75t_L         g08582(.A(new_n8838), .Y(new_n8839));
  NOR2xp33_ASAP7_75t_L      g08583(.A(new_n8839), .B(new_n8833), .Y(new_n8840));
  NOR2xp33_ASAP7_75t_L      g08584(.A(new_n8838), .B(new_n8495), .Y(new_n8841));
  INVx1_ASAP7_75t_L         g08585(.A(new_n8174), .Y(new_n8842));
  NAND2xp33_ASAP7_75t_L     g08586(.A(new_n8167), .B(new_n8842), .Y(new_n8843));
  NAND2xp33_ASAP7_75t_L     g08587(.A(\b[2] ), .B(new_n8169), .Y(new_n8844));
  OAI221xp5_ASAP7_75t_L     g08588(.A1(new_n8483), .A2(new_n262), .B1(new_n301), .B2(new_n8843), .C(new_n8844), .Y(new_n8845));
  NOR2xp33_ASAP7_75t_L      g08589(.A(new_n8176), .B(new_n319), .Y(new_n8846));
  OR3x1_ASAP7_75t_L         g08590(.A(new_n8845), .B(new_n8846), .C(new_n8172), .Y(new_n8847));
  A2O1A1Ixp33_ASAP7_75t_L   g08591(.A1(new_n312), .A2(new_n8490), .B(new_n8845), .C(new_n8172), .Y(new_n8848));
  NAND2xp33_ASAP7_75t_L     g08592(.A(new_n8848), .B(new_n8847), .Y(new_n8849));
  OAI21xp33_ASAP7_75t_L     g08593(.A1(new_n8840), .A2(new_n8841), .B(new_n8849), .Y(new_n8850));
  A2O1A1Ixp33_ASAP7_75t_L   g08594(.A1(new_n8492), .A2(new_n8489), .B(new_n8179), .C(new_n8838), .Y(new_n8851));
  A2O1A1Ixp33_ASAP7_75t_L   g08595(.A1(new_n8835), .A2(new_n8836), .B(new_n284), .C(new_n8833), .Y(new_n8852));
  A2O1A1Ixp33_ASAP7_75t_L   g08596(.A1(new_n312), .A2(new_n8490), .B(new_n8845), .C(\a[50] ), .Y(new_n8853));
  NOR3xp33_ASAP7_75t_L      g08597(.A(new_n8845), .B(new_n8846), .C(new_n8172), .Y(new_n8854));
  O2A1O1Ixp33_ASAP7_75t_L   g08598(.A1(new_n8845), .A2(new_n8846), .B(new_n8853), .C(new_n8854), .Y(new_n8855));
  NAND3xp33_ASAP7_75t_L     g08599(.A(new_n8852), .B(new_n8851), .C(new_n8855), .Y(new_n8856));
  NAND2xp33_ASAP7_75t_L     g08600(.A(\b[5] ), .B(new_n7333), .Y(new_n8857));
  OAI221xp5_ASAP7_75t_L     g08601(.A1(new_n7318), .A2(new_n427), .B1(new_n332), .B2(new_n7614), .C(new_n8857), .Y(new_n8858));
  A2O1A1Ixp33_ASAP7_75t_L   g08602(.A1(new_n5363), .A2(new_n7322), .B(new_n8858), .C(\a[47] ), .Y(new_n8859));
  NAND2xp33_ASAP7_75t_L     g08603(.A(\a[47] ), .B(new_n8859), .Y(new_n8860));
  A2O1A1Ixp33_ASAP7_75t_L   g08604(.A1(new_n5363), .A2(new_n7322), .B(new_n8858), .C(new_n7316), .Y(new_n8861));
  NAND2xp33_ASAP7_75t_L     g08605(.A(new_n8861), .B(new_n8860), .Y(new_n8862));
  INVx1_ASAP7_75t_L         g08606(.A(new_n8862), .Y(new_n8863));
  NAND3xp33_ASAP7_75t_L     g08607(.A(new_n8863), .B(new_n8850), .C(new_n8856), .Y(new_n8864));
  AOI21xp33_ASAP7_75t_L     g08608(.A1(new_n8852), .A2(new_n8851), .B(new_n8855), .Y(new_n8865));
  NOR3xp33_ASAP7_75t_L      g08609(.A(new_n8841), .B(new_n8849), .C(new_n8840), .Y(new_n8866));
  OAI21xp33_ASAP7_75t_L     g08610(.A1(new_n8865), .A2(new_n8866), .B(new_n8862), .Y(new_n8867));
  AND4x1_ASAP7_75t_L        g08611(.A(new_n8503), .B(new_n8832), .C(new_n8864), .D(new_n8867), .Y(new_n8868));
  O2A1O1Ixp33_ASAP7_75t_L   g08612(.A1(new_n8501), .A2(new_n8502), .B(new_n8481), .C(new_n8831), .Y(new_n8869));
  AOI21xp33_ASAP7_75t_L     g08613(.A1(new_n8867), .A2(new_n8864), .B(new_n8869), .Y(new_n8870));
  NAND2xp33_ASAP7_75t_L     g08614(.A(\b[9] ), .B(new_n6442), .Y(new_n8871));
  OAI221xp5_ASAP7_75t_L     g08615(.A1(new_n7304), .A2(new_n534), .B1(new_n448), .B2(new_n6741), .C(new_n8871), .Y(new_n8872));
  A2O1A1Ixp33_ASAP7_75t_L   g08616(.A1(new_n602), .A2(new_n6450), .B(new_n8872), .C(\a[44] ), .Y(new_n8873));
  AOI211xp5_ASAP7_75t_L     g08617(.A1(new_n602), .A2(new_n6450), .B(new_n8872), .C(new_n6439), .Y(new_n8874));
  A2O1A1O1Ixp25_ASAP7_75t_L g08618(.A1(new_n6450), .A2(new_n602), .B(new_n8872), .C(new_n8873), .D(new_n8874), .Y(new_n8875));
  OAI21xp33_ASAP7_75t_L     g08619(.A1(new_n8870), .A2(new_n8868), .B(new_n8875), .Y(new_n8876));
  NAND3xp33_ASAP7_75t_L     g08620(.A(new_n8869), .B(new_n8867), .C(new_n8864), .Y(new_n8877));
  AO21x2_ASAP7_75t_L        g08621(.A1(new_n8864), .A2(new_n8867), .B(new_n8869), .Y(new_n8878));
  INVx1_ASAP7_75t_L         g08622(.A(new_n8874), .Y(new_n8879));
  A2O1A1Ixp33_ASAP7_75t_L   g08623(.A1(new_n602), .A2(new_n6450), .B(new_n8872), .C(new_n6439), .Y(new_n8880));
  NAND2xp33_ASAP7_75t_L     g08624(.A(new_n8880), .B(new_n8879), .Y(new_n8881));
  NAND3xp33_ASAP7_75t_L     g08625(.A(new_n8878), .B(new_n8881), .C(new_n8877), .Y(new_n8882));
  NAND2xp33_ASAP7_75t_L     g08626(.A(new_n8876), .B(new_n8882), .Y(new_n8883));
  NOR2xp33_ASAP7_75t_L      g08627(.A(new_n8883), .B(new_n8828), .Y(new_n8884));
  AOI221xp5_ASAP7_75t_L     g08628(.A1(new_n8882), .A2(new_n8876), .B1(new_n8529), .B2(new_n8534), .C(new_n8536), .Y(new_n8885));
  OAI21xp33_ASAP7_75t_L     g08629(.A1(new_n8885), .A2(new_n8884), .B(new_n8827), .Y(new_n8886));
  INVx1_ASAP7_75t_L         g08630(.A(new_n8827), .Y(new_n8887));
  AOI21xp33_ASAP7_75t_L     g08631(.A1(new_n8878), .A2(new_n8877), .B(new_n8881), .Y(new_n8888));
  NOR3xp33_ASAP7_75t_L      g08632(.A(new_n8868), .B(new_n8870), .C(new_n8875), .Y(new_n8889));
  NOR2xp33_ASAP7_75t_L      g08633(.A(new_n8889), .B(new_n8888), .Y(new_n8890));
  A2O1A1Ixp33_ASAP7_75t_L   g08634(.A1(new_n8516), .A2(new_n8508), .B(new_n8539), .C(new_n8890), .Y(new_n8891));
  NAND2xp33_ASAP7_75t_L     g08635(.A(new_n8883), .B(new_n8828), .Y(new_n8892));
  NAND3xp33_ASAP7_75t_L     g08636(.A(new_n8891), .B(new_n8892), .C(new_n8887), .Y(new_n8893));
  NAND2xp33_ASAP7_75t_L     g08637(.A(new_n8886), .B(new_n8893), .Y(new_n8894));
  NOR3xp33_ASAP7_75t_L      g08638(.A(new_n8884), .B(new_n8885), .C(new_n8827), .Y(new_n8895));
  AOI211xp5_ASAP7_75t_L     g08639(.A1(new_n8472), .A2(new_n8526), .B(new_n8540), .C(new_n8895), .Y(new_n8896));
  AOI221xp5_ASAP7_75t_L     g08640(.A1(new_n8821), .A2(new_n8894), .B1(new_n8886), .B2(new_n8896), .C(new_n8820), .Y(new_n8897));
  O2A1O1Ixp33_ASAP7_75t_L   g08641(.A1(new_n4911), .A2(new_n1774), .B(new_n8816), .C(new_n4906), .Y(new_n8898));
  A2O1A1Ixp33_ASAP7_75t_L   g08642(.A1(new_n1052), .A2(new_n4912), .B(new_n8817), .C(new_n4906), .Y(new_n8899));
  OAI21xp33_ASAP7_75t_L     g08643(.A1(new_n4906), .A2(new_n8898), .B(new_n8899), .Y(new_n8900));
  AOI21xp33_ASAP7_75t_L     g08644(.A1(new_n8891), .A2(new_n8892), .B(new_n8887), .Y(new_n8901));
  OAI21xp33_ASAP7_75t_L     g08645(.A1(new_n8901), .A2(new_n8895), .B(new_n8821), .Y(new_n8902));
  OAI211xp5_ASAP7_75t_L     g08646(.A1(new_n8246), .A2(new_n8538), .B(new_n8893), .C(new_n8532), .Y(new_n8903));
  O2A1O1Ixp33_ASAP7_75t_L   g08647(.A1(new_n8901), .A2(new_n8903), .B(new_n8902), .C(new_n8900), .Y(new_n8904));
  NOR2xp33_ASAP7_75t_L      g08648(.A(new_n8904), .B(new_n8897), .Y(new_n8905));
  OAI21xp33_ASAP7_75t_L     g08649(.A1(new_n8814), .A2(new_n8561), .B(new_n8905), .Y(new_n8906));
  INVx1_ASAP7_75t_L         g08650(.A(new_n8814), .Y(new_n8907));
  AND2x2_ASAP7_75t_L        g08651(.A(new_n8552), .B(new_n8548), .Y(new_n8908));
  OAI221xp5_ASAP7_75t_L     g08652(.A1(new_n8897), .A2(new_n8904), .B1(new_n8555), .B2(new_n8908), .C(new_n8907), .Y(new_n8909));
  AND3x1_ASAP7_75t_L        g08653(.A(new_n8906), .B(new_n8909), .C(new_n8812), .Y(new_n8910));
  AOI21xp33_ASAP7_75t_L     g08654(.A1(new_n8906), .A2(new_n8909), .B(new_n8812), .Y(new_n8911));
  NOR2xp33_ASAP7_75t_L      g08655(.A(new_n8911), .B(new_n8910), .Y(new_n8912));
  A2O1A1Ixp33_ASAP7_75t_L   g08656(.A1(new_n8806), .A2(new_n8465), .B(new_n8565), .C(new_n8912), .Y(new_n8913));
  O2A1O1Ixp33_ASAP7_75t_L   g08657(.A1(new_n8557), .A2(new_n8563), .B(new_n8465), .C(new_n8565), .Y(new_n8914));
  NAND3xp33_ASAP7_75t_L     g08658(.A(new_n8906), .B(new_n8909), .C(new_n8812), .Y(new_n8915));
  AO21x2_ASAP7_75t_L        g08659(.A1(new_n8909), .A2(new_n8906), .B(new_n8812), .Y(new_n8916));
  NAND2xp33_ASAP7_75t_L     g08660(.A(new_n8915), .B(new_n8916), .Y(new_n8917));
  NAND2xp33_ASAP7_75t_L     g08661(.A(new_n8914), .B(new_n8917), .Y(new_n8918));
  OAI22xp33_ASAP7_75t_L     g08662(.A1(new_n3703), .A2(new_n1599), .B1(new_n1745), .B2(new_n3509), .Y(new_n8919));
  AOI221xp5_ASAP7_75t_L     g08663(.A1(new_n3503), .A2(\b[21] ), .B1(new_n3505), .B2(new_n2836), .C(new_n8919), .Y(new_n8920));
  XNOR2x2_ASAP7_75t_L       g08664(.A(new_n3493), .B(new_n8920), .Y(new_n8921));
  NAND3xp33_ASAP7_75t_L     g08665(.A(new_n8913), .B(new_n8918), .C(new_n8921), .Y(new_n8922));
  NOR2xp33_ASAP7_75t_L      g08666(.A(new_n8914), .B(new_n8917), .Y(new_n8923));
  AOI221xp5_ASAP7_75t_L     g08667(.A1(new_n8465), .A2(new_n8806), .B1(new_n8915), .B2(new_n8916), .C(new_n8565), .Y(new_n8924));
  XNOR2x2_ASAP7_75t_L       g08668(.A(\a[32] ), .B(new_n8920), .Y(new_n8925));
  OAI21xp33_ASAP7_75t_L     g08669(.A1(new_n8924), .A2(new_n8923), .B(new_n8925), .Y(new_n8926));
  NAND2xp33_ASAP7_75t_L     g08670(.A(new_n8926), .B(new_n8922), .Y(new_n8927));
  INVx1_ASAP7_75t_L         g08671(.A(new_n8564), .Y(new_n8928));
  O2A1O1Ixp33_ASAP7_75t_L   g08672(.A1(new_n8575), .A2(new_n8928), .B(new_n8576), .C(new_n8573), .Y(new_n8929));
  AO21x2_ASAP7_75t_L        g08673(.A1(new_n8584), .A2(new_n8586), .B(new_n8929), .Y(new_n8930));
  NOR2xp33_ASAP7_75t_L      g08674(.A(new_n8927), .B(new_n8930), .Y(new_n8931));
  O2A1O1Ixp33_ASAP7_75t_L   g08675(.A1(new_n8575), .A2(new_n8928), .B(new_n8576), .C(new_n8582), .Y(new_n8932));
  O2A1O1Ixp33_ASAP7_75t_L   g08676(.A1(new_n8932), .A2(new_n8582), .B(new_n8586), .C(new_n8929), .Y(new_n8933));
  AOI21xp33_ASAP7_75t_L     g08677(.A1(new_n8926), .A2(new_n8922), .B(new_n8933), .Y(new_n8934));
  OAI22xp33_ASAP7_75t_L     g08678(.A1(new_n3133), .A2(new_n2045), .B1(new_n2188), .B2(new_n2925), .Y(new_n8935));
  AOI221xp5_ASAP7_75t_L     g08679(.A1(new_n2938), .A2(\b[24] ), .B1(new_n2932), .B2(new_n2216), .C(new_n8935), .Y(new_n8936));
  XNOR2x2_ASAP7_75t_L       g08680(.A(new_n2928), .B(new_n8936), .Y(new_n8937));
  OAI21xp33_ASAP7_75t_L     g08681(.A1(new_n8934), .A2(new_n8931), .B(new_n8937), .Y(new_n8938));
  NOR3xp33_ASAP7_75t_L      g08682(.A(new_n8923), .B(new_n8925), .C(new_n8924), .Y(new_n8939));
  AOI21xp33_ASAP7_75t_L     g08683(.A1(new_n8913), .A2(new_n8918), .B(new_n8921), .Y(new_n8940));
  NOR2xp33_ASAP7_75t_L      g08684(.A(new_n8939), .B(new_n8940), .Y(new_n8941));
  NAND2xp33_ASAP7_75t_L     g08685(.A(new_n8933), .B(new_n8941), .Y(new_n8942));
  A2O1A1Ixp33_ASAP7_75t_L   g08686(.A1(new_n8584), .A2(new_n8586), .B(new_n8929), .C(new_n8927), .Y(new_n8943));
  XNOR2x2_ASAP7_75t_L       g08687(.A(\a[29] ), .B(new_n8936), .Y(new_n8944));
  NAND3xp33_ASAP7_75t_L     g08688(.A(new_n8943), .B(new_n8942), .C(new_n8944), .Y(new_n8945));
  OAI211xp5_ASAP7_75t_L     g08689(.A1(new_n8607), .A2(new_n8619), .B(new_n8938), .C(new_n8945), .Y(new_n8946));
  AOI21xp33_ASAP7_75t_L     g08690(.A1(new_n8943), .A2(new_n8942), .B(new_n8944), .Y(new_n8947));
  NOR3xp33_ASAP7_75t_L      g08691(.A(new_n8931), .B(new_n8934), .C(new_n8937), .Y(new_n8948));
  OAI21xp33_ASAP7_75t_L     g08692(.A1(new_n8947), .A2(new_n8948), .B(new_n8608), .Y(new_n8949));
  NOR2xp33_ASAP7_75t_L      g08693(.A(new_n2703), .B(new_n2410), .Y(new_n8950));
  AOI221xp5_ASAP7_75t_L     g08694(.A1(\b[25] ), .A2(new_n2577), .B1(\b[27] ), .B2(new_n2423), .C(new_n8950), .Y(new_n8951));
  O2A1O1Ixp33_ASAP7_75t_L   g08695(.A1(new_n2425), .A2(new_n2889), .B(new_n8951), .C(new_n2413), .Y(new_n8952));
  INVx1_ASAP7_75t_L         g08696(.A(new_n8952), .Y(new_n8953));
  O2A1O1Ixp33_ASAP7_75t_L   g08697(.A1(new_n2425), .A2(new_n2889), .B(new_n8951), .C(\a[26] ), .Y(new_n8954));
  AOI21xp33_ASAP7_75t_L     g08698(.A1(new_n8953), .A2(\a[26] ), .B(new_n8954), .Y(new_n8955));
  NAND3xp33_ASAP7_75t_L     g08699(.A(new_n8946), .B(new_n8949), .C(new_n8955), .Y(new_n8956));
  NOR3xp33_ASAP7_75t_L      g08700(.A(new_n8608), .B(new_n8947), .C(new_n8948), .Y(new_n8957));
  AOI211xp5_ASAP7_75t_L     g08701(.A1(new_n8938), .A2(new_n8945), .B(new_n8619), .C(new_n8607), .Y(new_n8958));
  INVx1_ASAP7_75t_L         g08702(.A(new_n8954), .Y(new_n8959));
  OAI21xp33_ASAP7_75t_L     g08703(.A1(new_n2413), .A2(new_n8952), .B(new_n8959), .Y(new_n8960));
  OAI21xp33_ASAP7_75t_L     g08704(.A1(new_n8957), .A2(new_n8958), .B(new_n8960), .Y(new_n8961));
  NAND2xp33_ASAP7_75t_L     g08705(.A(new_n8956), .B(new_n8961), .Y(new_n8962));
  NOR2xp33_ASAP7_75t_L      g08706(.A(new_n8804), .B(new_n8962), .Y(new_n8963));
  INVx1_ASAP7_75t_L         g08707(.A(new_n8462), .Y(new_n8964));
  A2O1A1Ixp33_ASAP7_75t_L   g08708(.A1(new_n8314), .A2(new_n8964), .B(new_n8615), .C(new_n8627), .Y(new_n8965));
  AOI21xp33_ASAP7_75t_L     g08709(.A1(new_n8961), .A2(new_n8956), .B(new_n8965), .Y(new_n8966));
  NAND2xp33_ASAP7_75t_L     g08710(.A(\b[30] ), .B(new_n1955), .Y(new_n8967));
  OAI221xp5_ASAP7_75t_L     g08711(.A1(new_n1962), .A2(new_n3098), .B1(new_n3079), .B2(new_n2089), .C(new_n8967), .Y(new_n8968));
  A2O1A1Ixp33_ASAP7_75t_L   g08712(.A1(new_n4813), .A2(new_n1964), .B(new_n8968), .C(\a[23] ), .Y(new_n8969));
  AOI211xp5_ASAP7_75t_L     g08713(.A1(new_n4813), .A2(new_n1964), .B(new_n8968), .C(new_n1952), .Y(new_n8970));
  A2O1A1O1Ixp25_ASAP7_75t_L g08714(.A1(new_n4813), .A2(new_n1964), .B(new_n8968), .C(new_n8969), .D(new_n8970), .Y(new_n8971));
  INVx1_ASAP7_75t_L         g08715(.A(new_n8971), .Y(new_n8972));
  OAI21xp33_ASAP7_75t_L     g08716(.A1(new_n8963), .A2(new_n8966), .B(new_n8972), .Y(new_n8973));
  NAND3xp33_ASAP7_75t_L     g08717(.A(new_n8965), .B(new_n8956), .C(new_n8961), .Y(new_n8974));
  NAND2xp33_ASAP7_75t_L     g08718(.A(new_n8804), .B(new_n8962), .Y(new_n8975));
  NAND3xp33_ASAP7_75t_L     g08719(.A(new_n8974), .B(new_n8975), .C(new_n8971), .Y(new_n8976));
  NAND2xp33_ASAP7_75t_L     g08720(.A(new_n8976), .B(new_n8973), .Y(new_n8977));
  NOR2xp33_ASAP7_75t_L      g08721(.A(new_n8802), .B(new_n8977), .Y(new_n8978));
  AOI221xp5_ASAP7_75t_L     g08722(.A1(new_n8642), .A2(new_n8629), .B1(new_n8973), .B2(new_n8976), .C(new_n8801), .Y(new_n8979));
  NOR2xp33_ASAP7_75t_L      g08723(.A(new_n4101), .B(new_n1518), .Y(new_n8980));
  AOI221xp5_ASAP7_75t_L     g08724(.A1(\b[31] ), .A2(new_n1659), .B1(\b[32] ), .B2(new_n1507), .C(new_n8980), .Y(new_n8981));
  O2A1O1Ixp33_ASAP7_75t_L   g08725(.A1(new_n1521), .A2(new_n4108), .B(new_n8981), .C(new_n1501), .Y(new_n8982));
  OAI21xp33_ASAP7_75t_L     g08726(.A1(new_n1521), .A2(new_n4108), .B(new_n8981), .Y(new_n8983));
  NAND2xp33_ASAP7_75t_L     g08727(.A(new_n1501), .B(new_n8983), .Y(new_n8984));
  OAI21xp33_ASAP7_75t_L     g08728(.A1(new_n1501), .A2(new_n8982), .B(new_n8984), .Y(new_n8985));
  NOR3xp33_ASAP7_75t_L      g08729(.A(new_n8978), .B(new_n8979), .C(new_n8985), .Y(new_n8986));
  INVx1_ASAP7_75t_L         g08730(.A(new_n8986), .Y(new_n8987));
  OAI21xp33_ASAP7_75t_L     g08731(.A1(new_n8979), .A2(new_n8978), .B(new_n8985), .Y(new_n8988));
  NAND3xp33_ASAP7_75t_L     g08732(.A(new_n8987), .B(new_n8800), .C(new_n8988), .Y(new_n8989));
  NAND2xp33_ASAP7_75t_L     g08733(.A(new_n8347), .B(new_n8346), .Y(new_n8990));
  A2O1A1O1Ixp25_ASAP7_75t_L g08734(.A1(new_n8343), .A2(new_n8990), .B(new_n8648), .C(new_n8638), .D(new_n8651), .Y(new_n8991));
  OA21x2_ASAP7_75t_L        g08735(.A1(new_n8979), .A2(new_n8978), .B(new_n8985), .Y(new_n8992));
  OAI21xp33_ASAP7_75t_L     g08736(.A1(new_n8986), .A2(new_n8992), .B(new_n8991), .Y(new_n8993));
  OAI22xp33_ASAP7_75t_L     g08737(.A1(new_n1285), .A2(new_n4344), .B1(new_n4581), .B2(new_n2118), .Y(new_n8994));
  AOI221xp5_ASAP7_75t_L     g08738(.A1(new_n1209), .A2(\b[36] ), .B1(new_n1216), .B2(new_n4621), .C(new_n8994), .Y(new_n8995));
  XNOR2x2_ASAP7_75t_L       g08739(.A(\a[17] ), .B(new_n8995), .Y(new_n8996));
  INVx1_ASAP7_75t_L         g08740(.A(new_n8996), .Y(new_n8997));
  AOI21xp33_ASAP7_75t_L     g08741(.A1(new_n8989), .A2(new_n8993), .B(new_n8997), .Y(new_n8998));
  NOR3xp33_ASAP7_75t_L      g08742(.A(new_n8991), .B(new_n8992), .C(new_n8986), .Y(new_n8999));
  AOI21xp33_ASAP7_75t_L     g08743(.A1(new_n8987), .A2(new_n8988), .B(new_n8800), .Y(new_n9000));
  NOR3xp33_ASAP7_75t_L      g08744(.A(new_n9000), .B(new_n8996), .C(new_n8999), .Y(new_n9001));
  OAI211xp5_ASAP7_75t_L     g08745(.A1(new_n8998), .A2(new_n9001), .B(new_n8670), .C(new_n8799), .Y(new_n9002));
  A2O1A1Ixp33_ASAP7_75t_L   g08746(.A1(new_n8659), .A2(new_n8663), .B(new_n8666), .C(new_n8799), .Y(new_n9003));
  NOR2xp33_ASAP7_75t_L      g08747(.A(new_n8998), .B(new_n9001), .Y(new_n9004));
  NAND2xp33_ASAP7_75t_L     g08748(.A(new_n9003), .B(new_n9004), .Y(new_n9005));
  NOR2xp33_ASAP7_75t_L      g08749(.A(new_n5311), .B(new_n864), .Y(new_n9006));
  AOI221xp5_ASAP7_75t_L     g08750(.A1(\b[37] ), .A2(new_n985), .B1(\b[39] ), .B2(new_n886), .C(new_n9006), .Y(new_n9007));
  O2A1O1Ixp33_ASAP7_75t_L   g08751(.A1(new_n872), .A2(new_n5578), .B(new_n9007), .C(new_n867), .Y(new_n9008));
  INVx1_ASAP7_75t_L         g08752(.A(new_n9008), .Y(new_n9009));
  O2A1O1Ixp33_ASAP7_75t_L   g08753(.A1(new_n872), .A2(new_n5578), .B(new_n9007), .C(\a[14] ), .Y(new_n9010));
  AOI21xp33_ASAP7_75t_L     g08754(.A1(new_n9009), .A2(\a[14] ), .B(new_n9010), .Y(new_n9011));
  NAND3xp33_ASAP7_75t_L     g08755(.A(new_n9002), .B(new_n9005), .C(new_n9011), .Y(new_n9012));
  AO21x2_ASAP7_75t_L        g08756(.A1(new_n9005), .A2(new_n9002), .B(new_n9011), .Y(new_n9013));
  AND4x1_ASAP7_75t_L        g08757(.A(new_n8684), .B(new_n8798), .C(new_n9013), .D(new_n9012), .Y(new_n9014));
  MAJIxp5_ASAP7_75t_L       g08758(.A(new_n8683), .B(new_n8797), .C(new_n8673), .Y(new_n9015));
  AOI21xp33_ASAP7_75t_L     g08759(.A1(new_n9013), .A2(new_n9012), .B(new_n9015), .Y(new_n9016));
  OAI22xp33_ASAP7_75t_L     g08760(.A1(new_n1550), .A2(new_n6110), .B1(new_n5855), .B2(new_n712), .Y(new_n9017));
  AOI221xp5_ASAP7_75t_L     g08761(.A1(new_n640), .A2(\b[42] ), .B1(new_n718), .B2(new_n6389), .C(new_n9017), .Y(new_n9018));
  XNOR2x2_ASAP7_75t_L       g08762(.A(new_n637), .B(new_n9018), .Y(new_n9019));
  OAI21xp33_ASAP7_75t_L     g08763(.A1(new_n9016), .A2(new_n9014), .B(new_n9019), .Y(new_n9020));
  NAND3xp33_ASAP7_75t_L     g08764(.A(new_n9015), .B(new_n9013), .C(new_n9012), .Y(new_n9021));
  AO22x1_ASAP7_75t_L        g08765(.A1(new_n9013), .A2(new_n9012), .B1(new_n8798), .B2(new_n8684), .Y(new_n9022));
  XNOR2x2_ASAP7_75t_L       g08766(.A(\a[11] ), .B(new_n9018), .Y(new_n9023));
  NAND3xp33_ASAP7_75t_L     g08767(.A(new_n9022), .B(new_n9021), .C(new_n9023), .Y(new_n9024));
  NAND3xp33_ASAP7_75t_L     g08768(.A(new_n8694), .B(new_n8684), .C(new_n8680), .Y(new_n9025));
  A2O1A1Ixp33_ASAP7_75t_L   g08769(.A1(new_n8690), .A2(new_n8691), .B(new_n8701), .C(new_n9025), .Y(new_n9026));
  NAND3xp33_ASAP7_75t_L     g08770(.A(new_n9026), .B(new_n9024), .C(new_n9020), .Y(new_n9027));
  NAND2xp33_ASAP7_75t_L     g08771(.A(new_n9020), .B(new_n9024), .Y(new_n9028));
  INVx1_ASAP7_75t_L         g08772(.A(new_n9025), .Y(new_n9029));
  A2O1A1O1Ixp25_ASAP7_75t_L g08773(.A1(new_n8395), .A2(new_n8396), .B(new_n8714), .C(new_n8696), .D(new_n9029), .Y(new_n9030));
  NAND2xp33_ASAP7_75t_L     g08774(.A(new_n9028), .B(new_n9030), .Y(new_n9031));
  NOR2xp33_ASAP7_75t_L      g08775(.A(new_n6671), .B(new_n506), .Y(new_n9032));
  AOI221xp5_ASAP7_75t_L     g08776(.A1(\b[45] ), .A2(new_n475), .B1(new_n470), .B2(\b[44] ), .C(new_n9032), .Y(new_n9033));
  O2A1O1Ixp33_ASAP7_75t_L   g08777(.A1(new_n477), .A2(new_n7255), .B(new_n9033), .C(new_n466), .Y(new_n9034));
  OAI21xp33_ASAP7_75t_L     g08778(.A1(new_n477), .A2(new_n7255), .B(new_n9033), .Y(new_n9035));
  NAND2xp33_ASAP7_75t_L     g08779(.A(new_n466), .B(new_n9035), .Y(new_n9036));
  OAI21xp33_ASAP7_75t_L     g08780(.A1(new_n466), .A2(new_n9034), .B(new_n9036), .Y(new_n9037));
  INVx1_ASAP7_75t_L         g08781(.A(new_n9037), .Y(new_n9038));
  NAND3xp33_ASAP7_75t_L     g08782(.A(new_n9031), .B(new_n9027), .C(new_n9038), .Y(new_n9039));
  NOR2xp33_ASAP7_75t_L      g08783(.A(new_n9028), .B(new_n9030), .Y(new_n9040));
  AOI21xp33_ASAP7_75t_L     g08784(.A1(new_n9024), .A2(new_n9020), .B(new_n9026), .Y(new_n9041));
  OAI21xp33_ASAP7_75t_L     g08785(.A1(new_n9041), .A2(new_n9040), .B(new_n9037), .Y(new_n9042));
  NAND3xp33_ASAP7_75t_L     g08786(.A(new_n8796), .B(new_n9039), .C(new_n9042), .Y(new_n9043));
  NAND3xp33_ASAP7_75t_L     g08787(.A(new_n9031), .B(new_n9027), .C(new_n9037), .Y(new_n9044));
  NOR3xp33_ASAP7_75t_L      g08788(.A(new_n9040), .B(new_n9041), .C(new_n9037), .Y(new_n9045));
  A2O1A1Ixp33_ASAP7_75t_L   g08789(.A1(new_n9037), .A2(new_n9044), .B(new_n9045), .C(new_n8723), .Y(new_n9046));
  NOR2xp33_ASAP7_75t_L      g08790(.A(new_n7270), .B(new_n375), .Y(new_n9047));
  AOI221xp5_ASAP7_75t_L     g08791(.A1(\b[48] ), .A2(new_n361), .B1(new_n349), .B2(\b[47] ), .C(new_n9047), .Y(new_n9048));
  O2A1O1Ixp33_ASAP7_75t_L   g08792(.A1(new_n356), .A2(new_n7868), .B(new_n9048), .C(new_n346), .Y(new_n9049));
  INVx1_ASAP7_75t_L         g08793(.A(new_n9049), .Y(new_n9050));
  O2A1O1Ixp33_ASAP7_75t_L   g08794(.A1(new_n356), .A2(new_n7868), .B(new_n9048), .C(\a[5] ), .Y(new_n9051));
  AOI21xp33_ASAP7_75t_L     g08795(.A1(new_n9050), .A2(\a[5] ), .B(new_n9051), .Y(new_n9052));
  NAND3xp33_ASAP7_75t_L     g08796(.A(new_n9043), .B(new_n9046), .C(new_n9052), .Y(new_n9053));
  AO21x2_ASAP7_75t_L        g08797(.A1(new_n9046), .A2(new_n9043), .B(new_n9052), .Y(new_n9054));
  NAND2xp33_ASAP7_75t_L     g08798(.A(new_n9053), .B(new_n9054), .Y(new_n9055));
  A2O1A1O1Ixp25_ASAP7_75t_L g08799(.A1(new_n8738), .A2(new_n8733), .B(new_n8741), .C(new_n8795), .D(new_n9055), .Y(new_n9056));
  A2O1A1Ixp33_ASAP7_75t_L   g08800(.A1(new_n8732), .A2(new_n8733), .B(new_n8741), .C(new_n8795), .Y(new_n9057));
  AOI21xp33_ASAP7_75t_L     g08801(.A1(new_n9054), .A2(new_n9053), .B(new_n9057), .Y(new_n9058));
  NOR3xp33_ASAP7_75t_L      g08802(.A(new_n9056), .B(new_n9058), .C(new_n8793), .Y(new_n9059));
  INVx1_ASAP7_75t_L         g08803(.A(new_n9059), .Y(new_n9060));
  OAI21xp33_ASAP7_75t_L     g08804(.A1(new_n9058), .A2(new_n9056), .B(new_n8793), .Y(new_n9061));
  NAND2xp33_ASAP7_75t_L     g08805(.A(new_n9061), .B(new_n9060), .Y(new_n9062));
  XNOR2x2_ASAP7_75t_L       g08806(.A(new_n8778), .B(new_n9062), .Y(\f[51] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g08807(.A1(new_n8774), .A2(new_n8773), .B(new_n8768), .C(new_n9061), .D(new_n9059), .Y(new_n9064));
  NAND2xp33_ASAP7_75t_L     g08808(.A(new_n8738), .B(new_n8733), .Y(new_n9065));
  AOI21xp33_ASAP7_75t_L     g08809(.A1(new_n9043), .A2(new_n9046), .B(new_n9052), .Y(new_n9066));
  A2O1A1O1Ixp25_ASAP7_75t_L g08810(.A1(new_n8748), .A2(new_n9065), .B(new_n8794), .C(new_n9053), .D(new_n9066), .Y(new_n9067));
  INVx1_ASAP7_75t_L         g08811(.A(new_n9044), .Y(new_n9068));
  INVx1_ASAP7_75t_L         g08812(.A(new_n9024), .Y(new_n9069));
  A2O1A1O1Ixp25_ASAP7_75t_L g08813(.A1(new_n8696), .A2(new_n8699), .B(new_n9029), .C(new_n9020), .D(new_n9069), .Y(new_n9070));
  NAND2xp33_ASAP7_75t_L     g08814(.A(new_n9005), .B(new_n9002), .Y(new_n9071));
  INVx1_ASAP7_75t_L         g08815(.A(new_n9071), .Y(new_n9072));
  A2O1A1Ixp33_ASAP7_75t_L   g08816(.A1(\a[14] ), .A2(new_n9009), .B(new_n9010), .C(new_n9072), .Y(new_n9073));
  NAND2xp33_ASAP7_75t_L     g08817(.A(new_n8949), .B(new_n8946), .Y(new_n9074));
  MAJIxp5_ASAP7_75t_L       g08818(.A(new_n8804), .B(new_n9074), .C(new_n8955), .Y(new_n9075));
  A2O1A1O1Ixp25_ASAP7_75t_L g08819(.A1(new_n8624), .A2(new_n8596), .B(new_n8607), .C(new_n8938), .D(new_n8948), .Y(new_n9076));
  NOR3xp33_ASAP7_75t_L      g08820(.A(new_n8923), .B(new_n8921), .C(new_n8924), .Y(new_n9077));
  NOR2xp33_ASAP7_75t_L      g08821(.A(new_n1895), .B(new_n3509), .Y(new_n9078));
  AOI221xp5_ASAP7_75t_L     g08822(.A1(\b[20] ), .A2(new_n3708), .B1(\b[22] ), .B2(new_n3503), .C(new_n9078), .Y(new_n9079));
  O2A1O1Ixp33_ASAP7_75t_L   g08823(.A1(new_n3513), .A2(new_n2522), .B(new_n9079), .C(new_n3493), .Y(new_n9080));
  INVx1_ASAP7_75t_L         g08824(.A(new_n9080), .Y(new_n9081));
  O2A1O1Ixp33_ASAP7_75t_L   g08825(.A1(new_n3513), .A2(new_n2522), .B(new_n9079), .C(\a[32] ), .Y(new_n9082));
  AOI21xp33_ASAP7_75t_L     g08826(.A1(new_n9081), .A2(\a[32] ), .B(new_n9082), .Y(new_n9083));
  A2O1A1O1Ixp25_ASAP7_75t_L g08827(.A1(new_n8465), .A2(new_n8806), .B(new_n8565), .C(new_n8916), .D(new_n8910), .Y(new_n9084));
  NAND2xp33_ASAP7_75t_L     g08828(.A(new_n8892), .B(new_n8891), .Y(new_n9085));
  O2A1O1Ixp33_ASAP7_75t_L   g08829(.A1(new_n5626), .A2(new_n8824), .B(new_n8826), .C(new_n9085), .Y(new_n9086));
  NAND3xp33_ASAP7_75t_L     g08830(.A(new_n8850), .B(new_n8856), .C(new_n8862), .Y(new_n9087));
  MAJIxp5_ASAP7_75t_L       g08831(.A(new_n8495), .B(new_n8839), .C(new_n8855), .Y(new_n9088));
  NAND2xp33_ASAP7_75t_L     g08832(.A(\b[3] ), .B(new_n8169), .Y(new_n9089));
  OAI221xp5_ASAP7_75t_L     g08833(.A1(new_n8483), .A2(new_n289), .B1(new_n332), .B2(new_n8843), .C(new_n9089), .Y(new_n9090));
  A2O1A1Ixp33_ASAP7_75t_L   g08834(.A1(new_n342), .A2(new_n8490), .B(new_n9090), .C(\a[50] ), .Y(new_n9091));
  AOI211xp5_ASAP7_75t_L     g08835(.A1(new_n342), .A2(new_n8490), .B(new_n8172), .C(new_n9090), .Y(new_n9092));
  A2O1A1O1Ixp25_ASAP7_75t_L g08836(.A1(new_n8490), .A2(new_n342), .B(new_n9090), .C(new_n9091), .D(new_n9092), .Y(new_n9093));
  NAND2xp33_ASAP7_75t_L     g08837(.A(new_n8836), .B(new_n8835), .Y(new_n9094));
  XNOR2x2_ASAP7_75t_L       g08838(.A(\a[52] ), .B(\a[51] ), .Y(new_n9095));
  NOR2xp33_ASAP7_75t_L      g08839(.A(new_n9095), .B(new_n9094), .Y(new_n9096));
  INVx1_ASAP7_75t_L         g08840(.A(\a[52] ), .Y(new_n9097));
  NAND2xp33_ASAP7_75t_L     g08841(.A(\a[53] ), .B(new_n9097), .Y(new_n9098));
  INVx1_ASAP7_75t_L         g08842(.A(\a[53] ), .Y(new_n9099));
  NAND2xp33_ASAP7_75t_L     g08843(.A(\a[52] ), .B(new_n9099), .Y(new_n9100));
  NAND2xp33_ASAP7_75t_L     g08844(.A(new_n9100), .B(new_n9098), .Y(new_n9101));
  NOR2xp33_ASAP7_75t_L      g08845(.A(new_n9101), .B(new_n8837), .Y(new_n9102));
  AOI22xp33_ASAP7_75t_L     g08846(.A1(new_n9096), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n9102), .Y(new_n9103));
  NAND2xp33_ASAP7_75t_L     g08847(.A(new_n9101), .B(new_n9094), .Y(new_n9104));
  OA21x2_ASAP7_75t_L        g08848(.A1(new_n9104), .A2(new_n274), .B(new_n9103), .Y(new_n9105));
  NAND3xp33_ASAP7_75t_L     g08849(.A(new_n9105), .B(new_n8839), .C(\a[53] ), .Y(new_n9106));
  INVx1_ASAP7_75t_L         g08850(.A(new_n9106), .Y(new_n9107));
  O2A1O1Ixp33_ASAP7_75t_L   g08851(.A1(new_n9104), .A2(new_n274), .B(new_n9103), .C(new_n9099), .Y(new_n9108));
  INVx1_ASAP7_75t_L         g08852(.A(new_n9108), .Y(new_n9109));
  O2A1O1Ixp33_ASAP7_75t_L   g08853(.A1(new_n9104), .A2(new_n274), .B(new_n9103), .C(\a[53] ), .Y(new_n9110));
  O2A1O1Ixp33_ASAP7_75t_L   g08854(.A1(new_n8839), .A2(new_n9109), .B(\a[53] ), .C(new_n9110), .Y(new_n9111));
  OAI21xp33_ASAP7_75t_L     g08855(.A1(new_n9107), .A2(new_n9111), .B(new_n9093), .Y(new_n9112));
  INVx1_ASAP7_75t_L         g08856(.A(new_n9092), .Y(new_n9113));
  A2O1A1Ixp33_ASAP7_75t_L   g08857(.A1(new_n342), .A2(new_n8490), .B(new_n9090), .C(new_n8172), .Y(new_n9114));
  NAND2xp33_ASAP7_75t_L     g08858(.A(new_n9114), .B(new_n9113), .Y(new_n9115));
  INVx1_ASAP7_75t_L         g08859(.A(new_n9110), .Y(new_n9116));
  A2O1A1Ixp33_ASAP7_75t_L   g08860(.A1(new_n8838), .A2(new_n9108), .B(new_n9099), .C(new_n9116), .Y(new_n9117));
  NAND3xp33_ASAP7_75t_L     g08861(.A(new_n9115), .B(new_n9106), .C(new_n9117), .Y(new_n9118));
  NAND3xp33_ASAP7_75t_L     g08862(.A(new_n9088), .B(new_n9118), .C(new_n9112), .Y(new_n9119));
  MAJIxp5_ASAP7_75t_L       g08863(.A(new_n8849), .B(new_n8838), .C(new_n8833), .Y(new_n9120));
  AOI21xp33_ASAP7_75t_L     g08864(.A1(new_n9117), .A2(new_n9106), .B(new_n9115), .Y(new_n9121));
  NOR3xp33_ASAP7_75t_L      g08865(.A(new_n9111), .B(new_n9093), .C(new_n9107), .Y(new_n9122));
  OAI21xp33_ASAP7_75t_L     g08866(.A1(new_n9122), .A2(new_n9121), .B(new_n9120), .Y(new_n9123));
  NOR2xp33_ASAP7_75t_L      g08867(.A(new_n448), .B(new_n7318), .Y(new_n9124));
  AOI221xp5_ASAP7_75t_L     g08868(.A1(new_n7333), .A2(\b[6] ), .B1(new_n7609), .B2(\b[5] ), .C(new_n9124), .Y(new_n9125));
  O2A1O1Ixp33_ASAP7_75t_L   g08869(.A1(new_n7321), .A2(new_n456), .B(new_n9125), .C(new_n7316), .Y(new_n9126));
  OAI21xp33_ASAP7_75t_L     g08870(.A1(new_n7321), .A2(new_n456), .B(new_n9125), .Y(new_n9127));
  NAND2xp33_ASAP7_75t_L     g08871(.A(new_n7316), .B(new_n9127), .Y(new_n9128));
  OA21x2_ASAP7_75t_L        g08872(.A1(new_n7316), .A2(new_n9126), .B(new_n9128), .Y(new_n9129));
  NAND3xp33_ASAP7_75t_L     g08873(.A(new_n9119), .B(new_n9123), .C(new_n9129), .Y(new_n9130));
  NOR3xp33_ASAP7_75t_L      g08874(.A(new_n9121), .B(new_n9122), .C(new_n9120), .Y(new_n9131));
  AOI21xp33_ASAP7_75t_L     g08875(.A1(new_n9118), .A2(new_n9112), .B(new_n9088), .Y(new_n9132));
  NOR2xp33_ASAP7_75t_L      g08876(.A(new_n7316), .B(new_n9127), .Y(new_n9133));
  O2A1O1Ixp33_ASAP7_75t_L   g08877(.A1(new_n7321), .A2(new_n456), .B(new_n9125), .C(\a[47] ), .Y(new_n9134));
  OAI22xp33_ASAP7_75t_L     g08878(.A1(new_n9132), .A2(new_n9131), .B1(new_n9134), .B2(new_n9133), .Y(new_n9135));
  NAND4xp25_ASAP7_75t_L     g08879(.A(new_n8878), .B(new_n9130), .C(new_n9135), .D(new_n9087), .Y(new_n9136));
  NAND2xp33_ASAP7_75t_L     g08880(.A(new_n9130), .B(new_n9135), .Y(new_n9137));
  A2O1A1Ixp33_ASAP7_75t_L   g08881(.A1(new_n8863), .A2(new_n8864), .B(new_n8869), .C(new_n9087), .Y(new_n9138));
  NAND2xp33_ASAP7_75t_L     g08882(.A(new_n9138), .B(new_n9137), .Y(new_n9139));
  OAI22xp33_ASAP7_75t_L     g08883(.A1(new_n7304), .A2(new_n590), .B1(new_n534), .B2(new_n6741), .Y(new_n9140));
  AOI221xp5_ASAP7_75t_L     g08884(.A1(new_n6442), .A2(\b[10] ), .B1(new_n6450), .B2(new_n690), .C(new_n9140), .Y(new_n9141));
  XNOR2x2_ASAP7_75t_L       g08885(.A(new_n6439), .B(new_n9141), .Y(new_n9142));
  INVx1_ASAP7_75t_L         g08886(.A(new_n9142), .Y(new_n9143));
  NAND3xp33_ASAP7_75t_L     g08887(.A(new_n9143), .B(new_n9139), .C(new_n9136), .Y(new_n9144));
  NOR2xp33_ASAP7_75t_L      g08888(.A(new_n9138), .B(new_n9137), .Y(new_n9145));
  AND2x2_ASAP7_75t_L        g08889(.A(new_n9138), .B(new_n9137), .Y(new_n9146));
  OAI21xp33_ASAP7_75t_L     g08890(.A1(new_n9145), .A2(new_n9146), .B(new_n9142), .Y(new_n9147));
  A2O1A1Ixp33_ASAP7_75t_L   g08891(.A1(new_n8528), .A2(new_n8480), .B(new_n8515), .C(new_n8517), .Y(new_n9148));
  A2O1A1Ixp33_ASAP7_75t_L   g08892(.A1(new_n9148), .A2(new_n8876), .B(new_n8889), .C(new_n9147), .Y(new_n9149));
  A2O1A1O1Ixp25_ASAP7_75t_L g08893(.A1(new_n8529), .A2(new_n8534), .B(new_n8536), .C(new_n8876), .D(new_n8889), .Y(new_n9150));
  AOI21xp33_ASAP7_75t_L     g08894(.A1(new_n9147), .A2(new_n9144), .B(new_n9150), .Y(new_n9151));
  NAND2xp33_ASAP7_75t_L     g08895(.A(\b[12] ), .B(new_n5623), .Y(new_n9152));
  OAI221xp5_ASAP7_75t_L     g08896(.A1(new_n5641), .A2(new_n936), .B1(new_n748), .B2(new_n5925), .C(new_n9152), .Y(new_n9153));
  AOI211xp5_ASAP7_75t_L     g08897(.A1(new_n1166), .A2(new_n5637), .B(new_n9153), .C(new_n5626), .Y(new_n9154));
  INVx1_ASAP7_75t_L         g08898(.A(new_n9154), .Y(new_n9155));
  A2O1A1Ixp33_ASAP7_75t_L   g08899(.A1(new_n1166), .A2(new_n5637), .B(new_n9153), .C(new_n5626), .Y(new_n9156));
  NAND2xp33_ASAP7_75t_L     g08900(.A(new_n9156), .B(new_n9155), .Y(new_n9157));
  AOI311xp33_ASAP7_75t_L    g08901(.A1(new_n9149), .A2(new_n9144), .A3(new_n9147), .B(new_n9157), .C(new_n9151), .Y(new_n9158));
  AOI21xp33_ASAP7_75t_L     g08902(.A1(new_n9136), .A2(new_n9139), .B(new_n9143), .Y(new_n9159));
  O2A1O1Ixp33_ASAP7_75t_L   g08903(.A1(new_n8888), .A2(new_n8828), .B(new_n8882), .C(new_n9159), .Y(new_n9160));
  NAND3xp33_ASAP7_75t_L     g08904(.A(new_n9150), .B(new_n9144), .C(new_n9147), .Y(new_n9161));
  A2O1A1Ixp33_ASAP7_75t_L   g08905(.A1(new_n1166), .A2(new_n5637), .B(new_n9153), .C(\a[41] ), .Y(new_n9162));
  A2O1A1O1Ixp25_ASAP7_75t_L g08906(.A1(new_n5637), .A2(new_n1166), .B(new_n9153), .C(new_n9162), .D(new_n9154), .Y(new_n9163));
  A2O1A1O1Ixp25_ASAP7_75t_L g08907(.A1(new_n9144), .A2(new_n9160), .B(new_n9150), .C(new_n9161), .D(new_n9163), .Y(new_n9164));
  NOR2xp33_ASAP7_75t_L      g08908(.A(new_n9158), .B(new_n9164), .Y(new_n9165));
  A2O1A1Ixp33_ASAP7_75t_L   g08909(.A1(new_n8894), .A2(new_n8821), .B(new_n9086), .C(new_n9165), .Y(new_n9166));
  NOR2xp33_ASAP7_75t_L      g08910(.A(new_n8885), .B(new_n8884), .Y(new_n9167));
  MAJIxp5_ASAP7_75t_L       g08911(.A(new_n8821), .B(new_n8827), .C(new_n9167), .Y(new_n9168));
  OAI21xp33_ASAP7_75t_L     g08912(.A1(new_n9158), .A2(new_n9164), .B(new_n9168), .Y(new_n9169));
  OAI22xp33_ASAP7_75t_L     g08913(.A1(new_n5144), .A2(new_n960), .B1(new_n1043), .B2(new_n4903), .Y(new_n9170));
  AOI221xp5_ASAP7_75t_L     g08914(.A1(new_n4917), .A2(\b[16] ), .B1(new_n4912), .B2(new_n1156), .C(new_n9170), .Y(new_n9171));
  XNOR2x2_ASAP7_75t_L       g08915(.A(new_n4906), .B(new_n9171), .Y(new_n9172));
  NAND3xp33_ASAP7_75t_L     g08916(.A(new_n9166), .B(new_n9169), .C(new_n9172), .Y(new_n9173));
  NOR3xp33_ASAP7_75t_L      g08917(.A(new_n9168), .B(new_n9158), .C(new_n9164), .Y(new_n9174));
  A2O1A1O1Ixp25_ASAP7_75t_L g08918(.A1(new_n8220), .A2(new_n8242), .B(new_n8243), .C(new_n8526), .D(new_n8540), .Y(new_n9175));
  AOI21xp33_ASAP7_75t_L     g08919(.A1(new_n8893), .A2(new_n8886), .B(new_n9175), .Y(new_n9176));
  NOR3xp33_ASAP7_75t_L      g08920(.A(new_n9165), .B(new_n9176), .C(new_n9086), .Y(new_n9177));
  XNOR2x2_ASAP7_75t_L       g08921(.A(\a[38] ), .B(new_n9171), .Y(new_n9178));
  OAI21xp33_ASAP7_75t_L     g08922(.A1(new_n9174), .A2(new_n9177), .B(new_n9178), .Y(new_n9179));
  A2O1A1Ixp33_ASAP7_75t_L   g08923(.A1(new_n8896), .A2(new_n8886), .B(new_n9176), .C(new_n8820), .Y(new_n9180));
  A2O1A1O1Ixp25_ASAP7_75t_L g08924(.A1(new_n8471), .A2(new_n8553), .B(new_n8814), .C(new_n9180), .D(new_n8897), .Y(new_n9181));
  NAND3xp33_ASAP7_75t_L     g08925(.A(new_n9181), .B(new_n9179), .C(new_n9173), .Y(new_n9182));
  AO21x2_ASAP7_75t_L        g08926(.A1(new_n9173), .A2(new_n9179), .B(new_n9181), .Y(new_n9183));
  NAND2xp33_ASAP7_75t_L     g08927(.A(\b[18] ), .B(new_n4155), .Y(new_n9184));
  OAI221xp5_ASAP7_75t_L     g08928(.A1(new_n4147), .A2(new_n1599), .B1(new_n1349), .B2(new_n4397), .C(new_n9184), .Y(new_n9185));
  A2O1A1Ixp33_ASAP7_75t_L   g08929(.A1(new_n1607), .A2(new_n4151), .B(new_n9185), .C(\a[35] ), .Y(new_n9186));
  NAND2xp33_ASAP7_75t_L     g08930(.A(\a[35] ), .B(new_n9186), .Y(new_n9187));
  A2O1A1Ixp33_ASAP7_75t_L   g08931(.A1(new_n1607), .A2(new_n4151), .B(new_n9185), .C(new_n4145), .Y(new_n9188));
  NAND2xp33_ASAP7_75t_L     g08932(.A(new_n9188), .B(new_n9187), .Y(new_n9189));
  NAND3xp33_ASAP7_75t_L     g08933(.A(new_n9189), .B(new_n9183), .C(new_n9182), .Y(new_n9190));
  AOI21xp33_ASAP7_75t_L     g08934(.A1(new_n9183), .A2(new_n9182), .B(new_n9189), .Y(new_n9191));
  O2A1O1Ixp33_ASAP7_75t_L   g08935(.A1(new_n8911), .A2(new_n8914), .B(new_n8915), .C(new_n9191), .Y(new_n9192));
  AO21x2_ASAP7_75t_L        g08936(.A1(new_n9182), .A2(new_n9183), .B(new_n9189), .Y(new_n9193));
  NAND3xp33_ASAP7_75t_L     g08937(.A(new_n9084), .B(new_n9190), .C(new_n9193), .Y(new_n9194));
  A2O1A1O1Ixp25_ASAP7_75t_L g08938(.A1(new_n9190), .A2(new_n9192), .B(new_n9084), .C(new_n9194), .D(new_n9083), .Y(new_n9195));
  AOI21xp33_ASAP7_75t_L     g08939(.A1(new_n9193), .A2(new_n9190), .B(new_n9084), .Y(new_n9196));
  AND3x1_ASAP7_75t_L        g08940(.A(new_n9084), .B(new_n9193), .C(new_n9190), .Y(new_n9197));
  OAI21xp33_ASAP7_75t_L     g08941(.A1(new_n9196), .A2(new_n9197), .B(new_n9083), .Y(new_n9198));
  OAI21xp33_ASAP7_75t_L     g08942(.A1(new_n9083), .A2(new_n9195), .B(new_n9198), .Y(new_n9199));
  AOI211xp5_ASAP7_75t_L     g08943(.A1(new_n8927), .A2(new_n8930), .B(new_n9077), .C(new_n9199), .Y(new_n9200));
  INVx1_ASAP7_75t_L         g08944(.A(new_n9077), .Y(new_n9201));
  INVx1_ASAP7_75t_L         g08945(.A(new_n9082), .Y(new_n9202));
  OAI21xp33_ASAP7_75t_L     g08946(.A1(new_n3493), .A2(new_n9080), .B(new_n9202), .Y(new_n9203));
  A2O1A1O1Ixp25_ASAP7_75t_L g08947(.A1(new_n9190), .A2(new_n9192), .B(new_n9084), .C(new_n9194), .D(new_n9203), .Y(new_n9204));
  NOR3xp33_ASAP7_75t_L      g08948(.A(new_n9197), .B(new_n9083), .C(new_n9196), .Y(new_n9205));
  NOR2xp33_ASAP7_75t_L      g08949(.A(new_n9204), .B(new_n9205), .Y(new_n9206));
  O2A1O1Ixp33_ASAP7_75t_L   g08950(.A1(new_n8941), .A2(new_n8933), .B(new_n9201), .C(new_n9206), .Y(new_n9207));
  OAI22xp33_ASAP7_75t_L     g08951(.A1(new_n3133), .A2(new_n2188), .B1(new_n2205), .B2(new_n2925), .Y(new_n9208));
  AOI221xp5_ASAP7_75t_L     g08952(.A1(new_n2938), .A2(\b[25] ), .B1(new_n2932), .B2(new_n5001), .C(new_n9208), .Y(new_n9209));
  XNOR2x2_ASAP7_75t_L       g08953(.A(\a[29] ), .B(new_n9209), .Y(new_n9210));
  NOR3xp33_ASAP7_75t_L      g08954(.A(new_n9200), .B(new_n9207), .C(new_n9210), .Y(new_n9211));
  OAI211xp5_ASAP7_75t_L     g08955(.A1(new_n8941), .A2(new_n8933), .B(new_n9206), .C(new_n9201), .Y(new_n9212));
  A2O1A1Ixp33_ASAP7_75t_L   g08956(.A1(new_n8927), .A2(new_n8930), .B(new_n9077), .C(new_n9199), .Y(new_n9213));
  XNOR2x2_ASAP7_75t_L       g08957(.A(new_n2928), .B(new_n9209), .Y(new_n9214));
  AOI21xp33_ASAP7_75t_L     g08958(.A1(new_n9212), .A2(new_n9213), .B(new_n9214), .Y(new_n9215));
  NOR3xp33_ASAP7_75t_L      g08959(.A(new_n9076), .B(new_n9211), .C(new_n9215), .Y(new_n9216));
  A2O1A1Ixp33_ASAP7_75t_L   g08960(.A1(new_n8606), .A2(new_n8294), .B(new_n8597), .C(new_n8596), .Y(new_n9217));
  A2O1A1Ixp33_ASAP7_75t_L   g08961(.A1(new_n9217), .A2(new_n8604), .B(new_n8947), .C(new_n8945), .Y(new_n9218));
  NAND3xp33_ASAP7_75t_L     g08962(.A(new_n9212), .B(new_n9213), .C(new_n9214), .Y(new_n9219));
  OAI21xp33_ASAP7_75t_L     g08963(.A1(new_n9207), .A2(new_n9200), .B(new_n9210), .Y(new_n9220));
  AOI21xp33_ASAP7_75t_L     g08964(.A1(new_n9220), .A2(new_n9219), .B(new_n9218), .Y(new_n9221));
  NOR2xp33_ASAP7_75t_L      g08965(.A(new_n3079), .B(new_n2415), .Y(new_n9222));
  AOI221xp5_ASAP7_75t_L     g08966(.A1(\b[26] ), .A2(new_n2577), .B1(\b[27] ), .B2(new_n2421), .C(new_n9222), .Y(new_n9223));
  O2A1O1Ixp33_ASAP7_75t_L   g08967(.A1(new_n2425), .A2(new_n3087), .B(new_n9223), .C(new_n2413), .Y(new_n9224));
  O2A1O1Ixp33_ASAP7_75t_L   g08968(.A1(new_n2425), .A2(new_n3087), .B(new_n9223), .C(\a[26] ), .Y(new_n9225));
  INVx1_ASAP7_75t_L         g08969(.A(new_n9225), .Y(new_n9226));
  OAI21xp33_ASAP7_75t_L     g08970(.A1(new_n2413), .A2(new_n9224), .B(new_n9226), .Y(new_n9227));
  OAI21xp33_ASAP7_75t_L     g08971(.A1(new_n9221), .A2(new_n9216), .B(new_n9227), .Y(new_n9228));
  NAND3xp33_ASAP7_75t_L     g08972(.A(new_n9218), .B(new_n9219), .C(new_n9220), .Y(new_n9229));
  OAI21xp33_ASAP7_75t_L     g08973(.A1(new_n9211), .A2(new_n9215), .B(new_n9076), .Y(new_n9230));
  OAI21xp33_ASAP7_75t_L     g08974(.A1(new_n2425), .A2(new_n3087), .B(new_n9223), .Y(new_n9231));
  NOR2xp33_ASAP7_75t_L      g08975(.A(new_n2413), .B(new_n9231), .Y(new_n9232));
  NOR2xp33_ASAP7_75t_L      g08976(.A(new_n9225), .B(new_n9232), .Y(new_n9233));
  NAND3xp33_ASAP7_75t_L     g08977(.A(new_n9229), .B(new_n9230), .C(new_n9233), .Y(new_n9234));
  AOI21xp33_ASAP7_75t_L     g08978(.A1(new_n9234), .A2(new_n9228), .B(new_n9075), .Y(new_n9235));
  O2A1O1Ixp33_ASAP7_75t_L   g08979(.A1(new_n8952), .A2(new_n2413), .B(new_n8959), .C(new_n9074), .Y(new_n9236));
  INVx1_ASAP7_75t_L         g08980(.A(new_n9236), .Y(new_n9237));
  NAND2xp33_ASAP7_75t_L     g08981(.A(new_n8965), .B(new_n8962), .Y(new_n9238));
  NAND2xp33_ASAP7_75t_L     g08982(.A(new_n9234), .B(new_n9228), .Y(new_n9239));
  AOI21xp33_ASAP7_75t_L     g08983(.A1(new_n9238), .A2(new_n9237), .B(new_n9239), .Y(new_n9240));
  NOR2xp33_ASAP7_75t_L      g08984(.A(new_n3456), .B(new_n1962), .Y(new_n9241));
  AOI221xp5_ASAP7_75t_L     g08985(.A1(new_n1955), .A2(\b[31] ), .B1(new_n2093), .B2(\b[29] ), .C(new_n9241), .Y(new_n9242));
  O2A1O1Ixp33_ASAP7_75t_L   g08986(.A1(new_n1956), .A2(new_n3681), .B(new_n9242), .C(new_n1952), .Y(new_n9243));
  O2A1O1Ixp33_ASAP7_75t_L   g08987(.A1(new_n1956), .A2(new_n3681), .B(new_n9242), .C(\a[23] ), .Y(new_n9244));
  INVx1_ASAP7_75t_L         g08988(.A(new_n9244), .Y(new_n9245));
  OAI21xp33_ASAP7_75t_L     g08989(.A1(new_n1952), .A2(new_n9243), .B(new_n9245), .Y(new_n9246));
  NOR3xp33_ASAP7_75t_L      g08990(.A(new_n9240), .B(new_n9246), .C(new_n9235), .Y(new_n9247));
  AO221x2_ASAP7_75t_L       g08991(.A1(new_n8962), .A2(new_n8965), .B1(new_n9228), .B2(new_n9234), .C(new_n9236), .Y(new_n9248));
  NAND3xp33_ASAP7_75t_L     g08992(.A(new_n9075), .B(new_n9228), .C(new_n9234), .Y(new_n9249));
  INVx1_ASAP7_75t_L         g08993(.A(new_n9243), .Y(new_n9250));
  AOI21xp33_ASAP7_75t_L     g08994(.A1(new_n9250), .A2(\a[23] ), .B(new_n9244), .Y(new_n9251));
  AOI21xp33_ASAP7_75t_L     g08995(.A1(new_n9248), .A2(new_n9249), .B(new_n9251), .Y(new_n9252));
  NOR3xp33_ASAP7_75t_L      g08996(.A(new_n8972), .B(new_n8966), .C(new_n8963), .Y(new_n9253));
  OAI21xp33_ASAP7_75t_L     g08997(.A1(new_n9253), .A2(new_n8802), .B(new_n8973), .Y(new_n9254));
  NOR3xp33_ASAP7_75t_L      g08998(.A(new_n9254), .B(new_n9252), .C(new_n9247), .Y(new_n9255));
  NAND3xp33_ASAP7_75t_L     g08999(.A(new_n9248), .B(new_n9249), .C(new_n9251), .Y(new_n9256));
  OAI21xp33_ASAP7_75t_L     g09000(.A1(new_n9235), .A2(new_n9240), .B(new_n9246), .Y(new_n9257));
  AOI21xp33_ASAP7_75t_L     g09001(.A1(new_n8974), .A2(new_n8975), .B(new_n8971), .Y(new_n9258));
  A2O1A1O1Ixp25_ASAP7_75t_L g09002(.A1(new_n8629), .A2(new_n8642), .B(new_n8801), .C(new_n8976), .D(new_n9258), .Y(new_n9259));
  AOI21xp33_ASAP7_75t_L     g09003(.A1(new_n9257), .A2(new_n9256), .B(new_n9259), .Y(new_n9260));
  NOR2xp33_ASAP7_75t_L      g09004(.A(new_n4101), .B(new_n1517), .Y(new_n9261));
  AOI221xp5_ASAP7_75t_L     g09005(.A1(\b[32] ), .A2(new_n1659), .B1(\b[34] ), .B2(new_n1511), .C(new_n9261), .Y(new_n9262));
  O2A1O1Ixp33_ASAP7_75t_L   g09006(.A1(new_n1521), .A2(new_n4352), .B(new_n9262), .C(new_n1501), .Y(new_n9263));
  INVx1_ASAP7_75t_L         g09007(.A(new_n9262), .Y(new_n9264));
  A2O1A1Ixp33_ASAP7_75t_L   g09008(.A1(new_n5599), .A2(new_n1513), .B(new_n9264), .C(new_n1501), .Y(new_n9265));
  OAI21xp33_ASAP7_75t_L     g09009(.A1(new_n1501), .A2(new_n9263), .B(new_n9265), .Y(new_n9266));
  NOR3xp33_ASAP7_75t_L      g09010(.A(new_n9255), .B(new_n9260), .C(new_n9266), .Y(new_n9267));
  NAND3xp33_ASAP7_75t_L     g09011(.A(new_n9259), .B(new_n9257), .C(new_n9256), .Y(new_n9268));
  OAI21xp33_ASAP7_75t_L     g09012(.A1(new_n9247), .A2(new_n9252), .B(new_n9254), .Y(new_n9269));
  INVx1_ASAP7_75t_L         g09013(.A(new_n9266), .Y(new_n9270));
  AOI21xp33_ASAP7_75t_L     g09014(.A1(new_n9268), .A2(new_n9269), .B(new_n9270), .Y(new_n9271));
  NOR2xp33_ASAP7_75t_L      g09015(.A(new_n9271), .B(new_n9267), .Y(new_n9272));
  NOR2xp33_ASAP7_75t_L      g09016(.A(new_n8979), .B(new_n8978), .Y(new_n9273));
  MAJIxp5_ASAP7_75t_L       g09017(.A(new_n8800), .B(new_n9273), .C(new_n8985), .Y(new_n9274));
  NAND2xp33_ASAP7_75t_L     g09018(.A(new_n9272), .B(new_n9274), .Y(new_n9275));
  XNOR2x2_ASAP7_75t_L       g09019(.A(new_n8802), .B(new_n8977), .Y(new_n9276));
  INVx1_ASAP7_75t_L         g09020(.A(new_n8985), .Y(new_n9277));
  MAJIxp5_ASAP7_75t_L       g09021(.A(new_n8991), .B(new_n9277), .C(new_n9276), .Y(new_n9278));
  OAI21xp33_ASAP7_75t_L     g09022(.A1(new_n9267), .A2(new_n9271), .B(new_n9278), .Y(new_n9279));
  NOR2xp33_ASAP7_75t_L      g09023(.A(new_n4613), .B(new_n2118), .Y(new_n9280));
  AOI221xp5_ASAP7_75t_L     g09024(.A1(\b[35] ), .A2(new_n1290), .B1(\b[37] ), .B2(new_n1209), .C(new_n9280), .Y(new_n9281));
  O2A1O1Ixp33_ASAP7_75t_L   g09025(.A1(new_n1210), .A2(new_n5083), .B(new_n9281), .C(new_n1206), .Y(new_n9282));
  INVx1_ASAP7_75t_L         g09026(.A(new_n9282), .Y(new_n9283));
  O2A1O1Ixp33_ASAP7_75t_L   g09027(.A1(new_n1210), .A2(new_n5083), .B(new_n9281), .C(\a[17] ), .Y(new_n9284));
  AOI21xp33_ASAP7_75t_L     g09028(.A1(new_n9283), .A2(\a[17] ), .B(new_n9284), .Y(new_n9285));
  NAND3xp33_ASAP7_75t_L     g09029(.A(new_n9275), .B(new_n9279), .C(new_n9285), .Y(new_n9286));
  AO21x2_ASAP7_75t_L        g09030(.A1(new_n9279), .A2(new_n9275), .B(new_n9285), .Y(new_n9287));
  NAND3xp33_ASAP7_75t_L     g09031(.A(new_n8989), .B(new_n8997), .C(new_n8993), .Y(new_n9288));
  A2O1A1O1Ixp25_ASAP7_75t_L g09032(.A1(new_n8668), .A2(new_n8669), .B(new_n8677), .C(new_n9288), .D(new_n8998), .Y(new_n9289));
  AND3x1_ASAP7_75t_L        g09033(.A(new_n9289), .B(new_n9287), .C(new_n9286), .Y(new_n9290));
  AOI21xp33_ASAP7_75t_L     g09034(.A1(new_n9287), .A2(new_n9286), .B(new_n9289), .Y(new_n9291));
  NOR2xp33_ASAP7_75t_L      g09035(.A(new_n5570), .B(new_n864), .Y(new_n9292));
  AOI221xp5_ASAP7_75t_L     g09036(.A1(\b[38] ), .A2(new_n985), .B1(\b[40] ), .B2(new_n886), .C(new_n9292), .Y(new_n9293));
  O2A1O1Ixp33_ASAP7_75t_L   g09037(.A1(new_n872), .A2(new_n5862), .B(new_n9293), .C(new_n867), .Y(new_n9294));
  INVx1_ASAP7_75t_L         g09038(.A(new_n9294), .Y(new_n9295));
  O2A1O1Ixp33_ASAP7_75t_L   g09039(.A1(new_n872), .A2(new_n5862), .B(new_n9293), .C(\a[14] ), .Y(new_n9296));
  AOI21xp33_ASAP7_75t_L     g09040(.A1(new_n9295), .A2(\a[14] ), .B(new_n9296), .Y(new_n9297));
  INVx1_ASAP7_75t_L         g09041(.A(new_n9297), .Y(new_n9298));
  NOR3xp33_ASAP7_75t_L      g09042(.A(new_n9290), .B(new_n9291), .C(new_n9298), .Y(new_n9299));
  NAND3xp33_ASAP7_75t_L     g09043(.A(new_n9289), .B(new_n9287), .C(new_n9286), .Y(new_n9300));
  AO21x2_ASAP7_75t_L        g09044(.A1(new_n9286), .A2(new_n9287), .B(new_n9289), .Y(new_n9301));
  AOI21xp33_ASAP7_75t_L     g09045(.A1(new_n9301), .A2(new_n9300), .B(new_n9297), .Y(new_n9302));
  NOR2xp33_ASAP7_75t_L      g09046(.A(new_n9302), .B(new_n9299), .Y(new_n9303));
  NAND3xp33_ASAP7_75t_L     g09047(.A(new_n9303), .B(new_n9022), .C(new_n9073), .Y(new_n9304));
  MAJIxp5_ASAP7_75t_L       g09048(.A(new_n9015), .B(new_n9071), .C(new_n9011), .Y(new_n9305));
  OAI21xp33_ASAP7_75t_L     g09049(.A1(new_n9299), .A2(new_n9302), .B(new_n9305), .Y(new_n9306));
  OAI22xp33_ASAP7_75t_L     g09050(.A1(new_n1550), .A2(new_n6378), .B1(new_n6110), .B2(new_n712), .Y(new_n9307));
  AOI221xp5_ASAP7_75t_L     g09051(.A1(new_n640), .A2(\b[43] ), .B1(new_n718), .B2(new_n6682), .C(new_n9307), .Y(new_n9308));
  XNOR2x2_ASAP7_75t_L       g09052(.A(new_n637), .B(new_n9308), .Y(new_n9309));
  INVx1_ASAP7_75t_L         g09053(.A(new_n9309), .Y(new_n9310));
  NAND3xp33_ASAP7_75t_L     g09054(.A(new_n9310), .B(new_n9306), .C(new_n9304), .Y(new_n9311));
  AOI21xp33_ASAP7_75t_L     g09055(.A1(new_n9304), .A2(new_n9306), .B(new_n9310), .Y(new_n9312));
  O2A1O1Ixp33_ASAP7_75t_L   g09056(.A1(new_n9028), .A2(new_n9030), .B(new_n9024), .C(new_n9312), .Y(new_n9313));
  NAND3xp33_ASAP7_75t_L     g09057(.A(new_n9301), .B(new_n9300), .C(new_n9297), .Y(new_n9314));
  OAI21xp33_ASAP7_75t_L     g09058(.A1(new_n9291), .A2(new_n9290), .B(new_n9298), .Y(new_n9315));
  NAND2xp33_ASAP7_75t_L     g09059(.A(new_n9314), .B(new_n9315), .Y(new_n9316));
  NOR2xp33_ASAP7_75t_L      g09060(.A(new_n9305), .B(new_n9316), .Y(new_n9317));
  AOI21xp33_ASAP7_75t_L     g09061(.A1(new_n9022), .A2(new_n9073), .B(new_n9303), .Y(new_n9318));
  OAI21xp33_ASAP7_75t_L     g09062(.A1(new_n9317), .A2(new_n9318), .B(new_n9309), .Y(new_n9319));
  NAND3xp33_ASAP7_75t_L     g09063(.A(new_n9070), .B(new_n9311), .C(new_n9319), .Y(new_n9320));
  OAI22xp33_ASAP7_75t_L     g09064(.A1(new_n513), .A2(new_n7249), .B1(new_n6944), .B2(new_n506), .Y(new_n9321));
  AOI221xp5_ASAP7_75t_L     g09065(.A1(new_n475), .A2(\b[46] ), .B1(new_n483), .B2(new_n7278), .C(new_n9321), .Y(new_n9322));
  XNOR2x2_ASAP7_75t_L       g09066(.A(new_n466), .B(new_n9322), .Y(new_n9323));
  INVx1_ASAP7_75t_L         g09067(.A(new_n9323), .Y(new_n9324));
  A2O1A1O1Ixp25_ASAP7_75t_L g09068(.A1(new_n9311), .A2(new_n9313), .B(new_n9070), .C(new_n9320), .D(new_n9324), .Y(new_n9325));
  AOI21xp33_ASAP7_75t_L     g09069(.A1(new_n9311), .A2(new_n9319), .B(new_n9070), .Y(new_n9326));
  NOR3xp33_ASAP7_75t_L      g09070(.A(new_n9318), .B(new_n9309), .C(new_n9317), .Y(new_n9327));
  A2O1A1O1Ixp25_ASAP7_75t_L g09071(.A1(new_n9020), .A2(new_n9026), .B(new_n9069), .C(new_n9319), .D(new_n9327), .Y(new_n9328));
  AOI211xp5_ASAP7_75t_L     g09072(.A1(new_n9328), .A2(new_n9319), .B(new_n9323), .C(new_n9326), .Y(new_n9329));
  A2O1A1Ixp33_ASAP7_75t_L   g09073(.A1(new_n8721), .A2(new_n8416), .B(new_n8720), .C(new_n8710), .Y(new_n9330));
  AOI22xp33_ASAP7_75t_L     g09074(.A1(new_n9042), .A2(new_n9039), .B1(new_n8716), .B2(new_n9330), .Y(new_n9331));
  NOR4xp25_ASAP7_75t_L      g09075(.A(new_n9331), .B(new_n9325), .C(new_n9329), .D(new_n9068), .Y(new_n9332));
  A2O1A1Ixp33_ASAP7_75t_L   g09076(.A1(new_n9328), .A2(new_n9319), .B(new_n9326), .C(new_n9323), .Y(new_n9333));
  A2O1A1Ixp33_ASAP7_75t_L   g09077(.A1(new_n8715), .A2(new_n9025), .B(new_n9028), .C(new_n9024), .Y(new_n9334));
  OAI21xp33_ASAP7_75t_L     g09078(.A1(new_n9327), .A2(new_n9312), .B(new_n9334), .Y(new_n9335));
  NAND3xp33_ASAP7_75t_L     g09079(.A(new_n9335), .B(new_n9320), .C(new_n9324), .Y(new_n9336));
  AOI21xp33_ASAP7_75t_L     g09080(.A1(new_n9031), .A2(new_n9027), .B(new_n9038), .Y(new_n9337));
  OAI22xp33_ASAP7_75t_L     g09081(.A1(new_n8744), .A2(new_n8722), .B1(new_n9337), .B2(new_n9045), .Y(new_n9338));
  AOI22xp33_ASAP7_75t_L     g09082(.A1(new_n9333), .A2(new_n9336), .B1(new_n9044), .B2(new_n9338), .Y(new_n9339));
  OAI22xp33_ASAP7_75t_L     g09083(.A1(new_n350), .A2(new_n7860), .B1(new_n7552), .B2(new_n375), .Y(new_n9340));
  AOI221xp5_ASAP7_75t_L     g09084(.A1(new_n361), .A2(\b[49] ), .B1(new_n359), .B2(new_n8438), .C(new_n9340), .Y(new_n9341));
  XNOR2x2_ASAP7_75t_L       g09085(.A(new_n346), .B(new_n9341), .Y(new_n9342));
  INVx1_ASAP7_75t_L         g09086(.A(new_n9342), .Y(new_n9343));
  NOR3xp33_ASAP7_75t_L      g09087(.A(new_n9343), .B(new_n9332), .C(new_n9339), .Y(new_n9344));
  NAND4xp25_ASAP7_75t_L     g09088(.A(new_n9338), .B(new_n9333), .C(new_n9044), .D(new_n9336), .Y(new_n9345));
  A2O1A1Ixp33_ASAP7_75t_L   g09089(.A1(new_n9313), .A2(new_n9311), .B(new_n9070), .C(new_n9320), .Y(new_n9346));
  A2O1A1Ixp33_ASAP7_75t_L   g09090(.A1(new_n9328), .A2(new_n9319), .B(new_n9326), .C(new_n9324), .Y(new_n9347));
  A2O1A1Ixp33_ASAP7_75t_L   g09091(.A1(new_n9039), .A2(new_n9038), .B(new_n8723), .C(new_n9044), .Y(new_n9348));
  A2O1A1Ixp33_ASAP7_75t_L   g09092(.A1(new_n9347), .A2(new_n9346), .B(new_n9329), .C(new_n9348), .Y(new_n9349));
  AOI21xp33_ASAP7_75t_L     g09093(.A1(new_n9349), .A2(new_n9345), .B(new_n9342), .Y(new_n9350));
  NOR3xp33_ASAP7_75t_L      g09094(.A(new_n9067), .B(new_n9344), .C(new_n9350), .Y(new_n9351));
  NAND3xp33_ASAP7_75t_L     g09095(.A(new_n9349), .B(new_n9345), .C(new_n9342), .Y(new_n9352));
  OAI21xp33_ASAP7_75t_L     g09096(.A1(new_n9339), .A2(new_n9332), .B(new_n9343), .Y(new_n9353));
  AOI221xp5_ASAP7_75t_L     g09097(.A1(new_n9057), .A2(new_n9053), .B1(new_n9352), .B2(new_n9353), .C(new_n9066), .Y(new_n9354));
  INVx1_ASAP7_75t_L         g09098(.A(\b[52] ), .Y(new_n9355));
  NAND2xp33_ASAP7_75t_L     g09099(.A(\b[50] ), .B(new_n286), .Y(new_n9356));
  OAI221xp5_ASAP7_75t_L     g09100(.A1(new_n285), .A2(new_n8779), .B1(new_n9355), .B2(new_n269), .C(new_n9356), .Y(new_n9357));
  A2O1A1Ixp33_ASAP7_75t_L   g09101(.A1(new_n8433), .A2(new_n8753), .B(new_n8758), .C(new_n8786), .Y(new_n9358));
  NOR2xp33_ASAP7_75t_L      g09102(.A(\b[51] ), .B(\b[52] ), .Y(new_n9359));
  NOR2xp33_ASAP7_75t_L      g09103(.A(new_n8779), .B(new_n9355), .Y(new_n9360));
  NOR2xp33_ASAP7_75t_L      g09104(.A(new_n9359), .B(new_n9360), .Y(new_n9361));
  A2O1A1Ixp33_ASAP7_75t_L   g09105(.A1(new_n9358), .A2(new_n8784), .B(new_n8783), .C(new_n9361), .Y(new_n9362));
  INVx1_ASAP7_75t_L         g09106(.A(new_n9362), .Y(new_n9363));
  INVx1_ASAP7_75t_L         g09107(.A(new_n8783), .Y(new_n9364));
  A2O1A1Ixp33_ASAP7_75t_L   g09108(.A1(new_n8787), .A2(new_n8786), .B(new_n8782), .C(new_n9364), .Y(new_n9365));
  NOR2xp33_ASAP7_75t_L      g09109(.A(new_n9361), .B(new_n9365), .Y(new_n9366));
  NOR2xp33_ASAP7_75t_L      g09110(.A(new_n9363), .B(new_n9366), .Y(new_n9367));
  A2O1A1Ixp33_ASAP7_75t_L   g09111(.A1(new_n9367), .A2(new_n273), .B(new_n9357), .C(\a[2] ), .Y(new_n9368));
  NAND2xp33_ASAP7_75t_L     g09112(.A(\a[2] ), .B(new_n9368), .Y(new_n9369));
  A2O1A1Ixp33_ASAP7_75t_L   g09113(.A1(new_n9367), .A2(new_n273), .B(new_n9357), .C(new_n257), .Y(new_n9370));
  NAND2xp33_ASAP7_75t_L     g09114(.A(new_n9370), .B(new_n9369), .Y(new_n9371));
  OA21x2_ASAP7_75t_L        g09115(.A1(new_n9354), .A2(new_n9351), .B(new_n9371), .Y(new_n9372));
  INVx1_ASAP7_75t_L         g09116(.A(new_n9372), .Y(new_n9373));
  INVx1_ASAP7_75t_L         g09117(.A(new_n9053), .Y(new_n9374));
  A2O1A1Ixp33_ASAP7_75t_L   g09118(.A1(new_n8749), .A2(new_n8795), .B(new_n9374), .C(new_n9054), .Y(new_n9375));
  NAND3xp33_ASAP7_75t_L     g09119(.A(new_n9375), .B(new_n9352), .C(new_n9353), .Y(new_n9376));
  NAND2xp33_ASAP7_75t_L     g09120(.A(new_n9352), .B(new_n9353), .Y(new_n9377));
  NAND2xp33_ASAP7_75t_L     g09121(.A(new_n9067), .B(new_n9377), .Y(new_n9378));
  INVx1_ASAP7_75t_L         g09122(.A(new_n9371), .Y(new_n9379));
  NAND3xp33_ASAP7_75t_L     g09123(.A(new_n9376), .B(new_n9378), .C(new_n9379), .Y(new_n9380));
  NAND2xp33_ASAP7_75t_L     g09124(.A(new_n9380), .B(new_n9373), .Y(new_n9381));
  XOR2x2_ASAP7_75t_L        g09125(.A(new_n9064), .B(new_n9381), .Y(\f[52] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g09126(.A1(new_n9061), .A2(new_n8778), .B(new_n9059), .C(new_n9380), .D(new_n9372), .Y(new_n9383));
  NAND2xp33_ASAP7_75t_L     g09127(.A(new_n9345), .B(new_n9349), .Y(new_n9384));
  NAND3xp33_ASAP7_75t_L     g09128(.A(new_n9349), .B(new_n9345), .C(new_n9343), .Y(new_n9385));
  A2O1A1Ixp33_ASAP7_75t_L   g09129(.A1(new_n9353), .A2(new_n9384), .B(new_n9067), .C(new_n9385), .Y(new_n9386));
  NOR2xp33_ASAP7_75t_L      g09130(.A(new_n9291), .B(new_n9290), .Y(new_n9387));
  A2O1A1Ixp33_ASAP7_75t_L   g09131(.A1(\a[14] ), .A2(new_n9295), .B(new_n9296), .C(new_n9387), .Y(new_n9388));
  NAND2xp33_ASAP7_75t_L     g09132(.A(new_n9279), .B(new_n9275), .Y(new_n9389));
  INVx1_ASAP7_75t_L         g09133(.A(new_n9389), .Y(new_n9390));
  A2O1A1Ixp33_ASAP7_75t_L   g09134(.A1(\a[17] ), .A2(new_n9283), .B(new_n9284), .C(new_n9390), .Y(new_n9391));
  NAND2xp33_ASAP7_75t_L     g09135(.A(new_n9249), .B(new_n9248), .Y(new_n9392));
  MAJIxp5_ASAP7_75t_L       g09136(.A(new_n9259), .B(new_n9392), .C(new_n9251), .Y(new_n9393));
  NOR2xp33_ASAP7_75t_L      g09137(.A(new_n3674), .B(new_n1962), .Y(new_n9394));
  AOI221xp5_ASAP7_75t_L     g09138(.A1(new_n1955), .A2(\b[32] ), .B1(new_n2093), .B2(\b[30] ), .C(new_n9394), .Y(new_n9395));
  INVx1_ASAP7_75t_L         g09139(.A(new_n9395), .Y(new_n9396));
  A2O1A1Ixp33_ASAP7_75t_L   g09140(.A1(new_n3900), .A2(new_n1964), .B(new_n9396), .C(\a[23] ), .Y(new_n9397));
  O2A1O1Ixp33_ASAP7_75t_L   g09141(.A1(new_n1956), .A2(new_n3897), .B(new_n9395), .C(new_n1952), .Y(new_n9398));
  NOR2xp33_ASAP7_75t_L      g09142(.A(new_n1952), .B(new_n9398), .Y(new_n9399));
  A2O1A1O1Ixp25_ASAP7_75t_L g09143(.A1(new_n3900), .A2(new_n1964), .B(new_n9396), .C(new_n9397), .D(new_n9399), .Y(new_n9400));
  AOI21xp33_ASAP7_75t_L     g09144(.A1(new_n9229), .A2(new_n9230), .B(new_n9233), .Y(new_n9401));
  A2O1A1O1Ixp25_ASAP7_75t_L g09145(.A1(new_n8965), .A2(new_n8962), .B(new_n9236), .C(new_n9234), .D(new_n9401), .Y(new_n9402));
  OAI22xp33_ASAP7_75t_L     g09146(.A1(new_n2572), .A2(new_n2879), .B1(new_n3079), .B2(new_n2410), .Y(new_n9403));
  AOI221xp5_ASAP7_75t_L     g09147(.A1(new_n2423), .A2(\b[29] ), .B1(new_n2417), .B2(new_n3873), .C(new_n9403), .Y(new_n9404));
  XNOR2x2_ASAP7_75t_L       g09148(.A(new_n2413), .B(new_n9404), .Y(new_n9405));
  INVx1_ASAP7_75t_L         g09149(.A(new_n9405), .Y(new_n9406));
  NAND2xp33_ASAP7_75t_L     g09150(.A(new_n9213), .B(new_n9212), .Y(new_n9407));
  MAJIxp5_ASAP7_75t_L       g09151(.A(new_n9076), .B(new_n9214), .C(new_n9407), .Y(new_n9408));
  A2O1A1Ixp33_ASAP7_75t_L   g09152(.A1(new_n8922), .A2(new_n8926), .B(new_n8933), .C(new_n9201), .Y(new_n9409));
  NOR2xp33_ASAP7_75t_L      g09153(.A(new_n2045), .B(new_n3509), .Y(new_n9410));
  AOI221xp5_ASAP7_75t_L     g09154(.A1(\b[21] ), .A2(new_n3708), .B1(\b[23] ), .B2(new_n3503), .C(new_n9410), .Y(new_n9411));
  INVx1_ASAP7_75t_L         g09155(.A(new_n9411), .Y(new_n9412));
  A2O1A1Ixp33_ASAP7_75t_L   g09156(.A1(new_n2679), .A2(new_n3505), .B(new_n9412), .C(\a[32] ), .Y(new_n9413));
  O2A1O1Ixp33_ASAP7_75t_L   g09157(.A1(new_n3513), .A2(new_n2194), .B(new_n9411), .C(\a[32] ), .Y(new_n9414));
  AOI21xp33_ASAP7_75t_L     g09158(.A1(new_n9413), .A2(\a[32] ), .B(new_n9414), .Y(new_n9415));
  INVx1_ASAP7_75t_L         g09159(.A(new_n9190), .Y(new_n9416));
  NAND3xp33_ASAP7_75t_L     g09160(.A(new_n9166), .B(new_n9169), .C(new_n9178), .Y(new_n9417));
  A2O1A1Ixp33_ASAP7_75t_L   g09161(.A1(new_n9172), .A2(new_n9173), .B(new_n9181), .C(new_n9417), .Y(new_n9418));
  OAI22xp33_ASAP7_75t_L     g09162(.A1(new_n5144), .A2(new_n1043), .B1(new_n1150), .B2(new_n4903), .Y(new_n9419));
  AOI221xp5_ASAP7_75t_L     g09163(.A1(new_n4917), .A2(\b[17] ), .B1(new_n4912), .B2(new_n1633), .C(new_n9419), .Y(new_n9420));
  XNOR2x2_ASAP7_75t_L       g09164(.A(\a[38] ), .B(new_n9420), .Y(new_n9421));
  INVx1_ASAP7_75t_L         g09165(.A(new_n9151), .Y(new_n9422));
  NAND3xp33_ASAP7_75t_L     g09166(.A(new_n9422), .B(new_n9161), .C(new_n9163), .Y(new_n9423));
  A2O1A1O1Ixp25_ASAP7_75t_L g09167(.A1(new_n8821), .A2(new_n8894), .B(new_n9086), .C(new_n9423), .D(new_n9164), .Y(new_n9424));
  OAI22xp33_ASAP7_75t_L     g09168(.A1(new_n5640), .A2(new_n936), .B1(new_n833), .B2(new_n5925), .Y(new_n9425));
  AOI221xp5_ASAP7_75t_L     g09169(.A1(new_n5629), .A2(\b[14] ), .B1(new_n5637), .B2(new_n971), .C(new_n9425), .Y(new_n9426));
  XNOR2x2_ASAP7_75t_L       g09170(.A(new_n5626), .B(new_n9426), .Y(new_n9427));
  NOR3xp33_ASAP7_75t_L      g09171(.A(new_n9146), .B(new_n9142), .C(new_n9145), .Y(new_n9428));
  A2O1A1O1Ixp25_ASAP7_75t_L g09172(.A1(new_n8876), .A2(new_n9148), .B(new_n8889), .C(new_n9147), .D(new_n9428), .Y(new_n9429));
  OAI22xp33_ASAP7_75t_L     g09173(.A1(new_n7304), .A2(new_n680), .B1(new_n590), .B2(new_n6741), .Y(new_n9430));
  AOI221xp5_ASAP7_75t_L     g09174(.A1(new_n6442), .A2(\b[11] ), .B1(new_n6450), .B2(new_n976), .C(new_n9430), .Y(new_n9431));
  XNOR2x2_ASAP7_75t_L       g09175(.A(new_n6439), .B(new_n9431), .Y(new_n9432));
  INVx1_ASAP7_75t_L         g09176(.A(new_n9432), .Y(new_n9433));
  NAND2xp33_ASAP7_75t_L     g09177(.A(new_n9123), .B(new_n9119), .Y(new_n9434));
  O2A1O1Ixp33_ASAP7_75t_L   g09178(.A1(new_n9126), .A2(new_n7316), .B(new_n9128), .C(new_n9434), .Y(new_n9435));
  OAI21xp33_ASAP7_75t_L     g09179(.A1(new_n9120), .A2(new_n9121), .B(new_n9118), .Y(new_n9436));
  INVx1_ASAP7_75t_L         g09180(.A(new_n9104), .Y(new_n9437));
  INVx1_ASAP7_75t_L         g09181(.A(new_n9101), .Y(new_n9438));
  NAND2xp33_ASAP7_75t_L     g09182(.A(new_n9094), .B(new_n9438), .Y(new_n9439));
  NAND3xp33_ASAP7_75t_L     g09183(.A(new_n8837), .B(new_n9095), .C(new_n9101), .Y(new_n9440));
  NAND2xp33_ASAP7_75t_L     g09184(.A(\b[1] ), .B(new_n9096), .Y(new_n9441));
  OAI221xp5_ASAP7_75t_L     g09185(.A1(new_n9440), .A2(new_n284), .B1(new_n289), .B2(new_n9439), .C(new_n9441), .Y(new_n9442));
  A2O1A1Ixp33_ASAP7_75t_L   g09186(.A1(new_n294), .A2(new_n9437), .B(new_n9442), .C(\a[53] ), .Y(new_n9443));
  A2O1A1Ixp33_ASAP7_75t_L   g09187(.A1(new_n294), .A2(new_n9437), .B(new_n9442), .C(new_n9099), .Y(new_n9444));
  INVx1_ASAP7_75t_L         g09188(.A(new_n9444), .Y(new_n9445));
  A2O1A1O1Ixp25_ASAP7_75t_L g09189(.A1(new_n9105), .A2(new_n8839), .B(new_n9443), .C(\a[53] ), .D(new_n9445), .Y(new_n9446));
  OAI21xp33_ASAP7_75t_L     g09190(.A1(new_n9104), .A2(new_n274), .B(new_n9103), .Y(new_n9447));
  NOR2xp33_ASAP7_75t_L      g09191(.A(new_n9104), .B(new_n509), .Y(new_n9448));
  NOR5xp2_ASAP7_75t_L       g09192(.A(new_n9447), .B(new_n9442), .C(new_n9448), .D(new_n8838), .E(new_n9099), .Y(new_n9449));
  NAND2xp33_ASAP7_75t_L     g09193(.A(\b[4] ), .B(new_n8169), .Y(new_n9450));
  OAI221xp5_ASAP7_75t_L     g09194(.A1(new_n8483), .A2(new_n301), .B1(new_n384), .B2(new_n8843), .C(new_n9450), .Y(new_n9451));
  A2O1A1Ixp33_ASAP7_75t_L   g09195(.A1(new_n394), .A2(new_n8490), .B(new_n9451), .C(\a[50] ), .Y(new_n9452));
  INVx1_ASAP7_75t_L         g09196(.A(new_n9451), .Y(new_n9453));
  O2A1O1Ixp33_ASAP7_75t_L   g09197(.A1(new_n728), .A2(new_n8176), .B(new_n9453), .C(\a[50] ), .Y(new_n9454));
  AOI21xp33_ASAP7_75t_L     g09198(.A1(new_n9452), .A2(\a[50] ), .B(new_n9454), .Y(new_n9455));
  NOR3xp33_ASAP7_75t_L      g09199(.A(new_n9446), .B(new_n9449), .C(new_n9455), .Y(new_n9456));
  NOR2xp33_ASAP7_75t_L      g09200(.A(new_n9448), .B(new_n9442), .Y(new_n9457));
  NAND2xp33_ASAP7_75t_L     g09201(.A(\a[53] ), .B(new_n9457), .Y(new_n9458));
  NAND3xp33_ASAP7_75t_L     g09202(.A(new_n9458), .B(new_n9106), .C(new_n9444), .Y(new_n9459));
  NAND4xp25_ASAP7_75t_L     g09203(.A(new_n9457), .B(\a[53] ), .C(new_n8839), .D(new_n9105), .Y(new_n9460));
  AOI221xp5_ASAP7_75t_L     g09204(.A1(new_n9452), .A2(\a[50] ), .B1(new_n9460), .B2(new_n9459), .C(new_n9454), .Y(new_n9461));
  OAI21xp33_ASAP7_75t_L     g09205(.A1(new_n9456), .A2(new_n9461), .B(new_n9436), .Y(new_n9462));
  AOI21xp33_ASAP7_75t_L     g09206(.A1(new_n9088), .A2(new_n9112), .B(new_n9122), .Y(new_n9463));
  INVx1_ASAP7_75t_L         g09207(.A(new_n9456), .Y(new_n9464));
  OAI21xp33_ASAP7_75t_L     g09208(.A1(new_n9449), .A2(new_n9446), .B(new_n9455), .Y(new_n9465));
  NAND3xp33_ASAP7_75t_L     g09209(.A(new_n9463), .B(new_n9464), .C(new_n9465), .Y(new_n9466));
  NOR2xp33_ASAP7_75t_L      g09210(.A(new_n534), .B(new_n7318), .Y(new_n9467));
  AOI221xp5_ASAP7_75t_L     g09211(.A1(new_n7333), .A2(\b[7] ), .B1(new_n7609), .B2(\b[6] ), .C(new_n9467), .Y(new_n9468));
  O2A1O1Ixp33_ASAP7_75t_L   g09212(.A1(new_n7321), .A2(new_n540), .B(new_n9468), .C(new_n7316), .Y(new_n9469));
  OAI21xp33_ASAP7_75t_L     g09213(.A1(new_n7321), .A2(new_n540), .B(new_n9468), .Y(new_n9470));
  NAND2xp33_ASAP7_75t_L     g09214(.A(new_n7316), .B(new_n9470), .Y(new_n9471));
  OA21x2_ASAP7_75t_L        g09215(.A1(new_n7316), .A2(new_n9469), .B(new_n9471), .Y(new_n9472));
  NAND3xp33_ASAP7_75t_L     g09216(.A(new_n9466), .B(new_n9462), .C(new_n9472), .Y(new_n9473));
  AOI21xp33_ASAP7_75t_L     g09217(.A1(new_n9464), .A2(new_n9465), .B(new_n9463), .Y(new_n9474));
  A2O1A1O1Ixp25_ASAP7_75t_L g09218(.A1(new_n9112), .A2(new_n9088), .B(new_n9122), .C(new_n9465), .D(new_n9456), .Y(new_n9475));
  OAI21xp33_ASAP7_75t_L     g09219(.A1(new_n7316), .A2(new_n9469), .B(new_n9471), .Y(new_n9476));
  A2O1A1Ixp33_ASAP7_75t_L   g09220(.A1(new_n9475), .A2(new_n9465), .B(new_n9474), .C(new_n9476), .Y(new_n9477));
  AND2x2_ASAP7_75t_L        g09221(.A(new_n9473), .B(new_n9477), .Y(new_n9478));
  A2O1A1Ixp33_ASAP7_75t_L   g09222(.A1(new_n9137), .A2(new_n9138), .B(new_n9435), .C(new_n9478), .Y(new_n9479));
  NAND2xp33_ASAP7_75t_L     g09223(.A(new_n9473), .B(new_n9477), .Y(new_n9480));
  OAI211xp5_ASAP7_75t_L     g09224(.A1(new_n9434), .A2(new_n9129), .B(new_n9480), .C(new_n9139), .Y(new_n9481));
  AOI21xp33_ASAP7_75t_L     g09225(.A1(new_n9479), .A2(new_n9481), .B(new_n9433), .Y(new_n9482));
  O2A1O1Ixp33_ASAP7_75t_L   g09226(.A1(new_n9434), .A2(new_n9129), .B(new_n9139), .C(new_n9480), .Y(new_n9483));
  NOR3xp33_ASAP7_75t_L      g09227(.A(new_n9478), .B(new_n9146), .C(new_n9435), .Y(new_n9484));
  NOR3xp33_ASAP7_75t_L      g09228(.A(new_n9484), .B(new_n9432), .C(new_n9483), .Y(new_n9485));
  NOR3xp33_ASAP7_75t_L      g09229(.A(new_n9429), .B(new_n9482), .C(new_n9485), .Y(new_n9486));
  OAI21xp33_ASAP7_75t_L     g09230(.A1(new_n9159), .A2(new_n9150), .B(new_n9144), .Y(new_n9487));
  OAI21xp33_ASAP7_75t_L     g09231(.A1(new_n9483), .A2(new_n9484), .B(new_n9432), .Y(new_n9488));
  NAND3xp33_ASAP7_75t_L     g09232(.A(new_n9433), .B(new_n9479), .C(new_n9481), .Y(new_n9489));
  AOI21xp33_ASAP7_75t_L     g09233(.A1(new_n9489), .A2(new_n9488), .B(new_n9487), .Y(new_n9490));
  NOR3xp33_ASAP7_75t_L      g09234(.A(new_n9427), .B(new_n9486), .C(new_n9490), .Y(new_n9491));
  NAND3xp33_ASAP7_75t_L     g09235(.A(new_n9487), .B(new_n9488), .C(new_n9489), .Y(new_n9492));
  OAI21xp33_ASAP7_75t_L     g09236(.A1(new_n9485), .A2(new_n9482), .B(new_n9429), .Y(new_n9493));
  NAND3xp33_ASAP7_75t_L     g09237(.A(new_n9427), .B(new_n9492), .C(new_n9493), .Y(new_n9494));
  O2A1O1Ixp33_ASAP7_75t_L   g09238(.A1(new_n9427), .A2(new_n9491), .B(new_n9494), .C(new_n9424), .Y(new_n9495));
  NAND2xp33_ASAP7_75t_L     g09239(.A(new_n8827), .B(new_n9167), .Y(new_n9496));
  INVx1_ASAP7_75t_L         g09240(.A(new_n9164), .Y(new_n9497));
  A2O1A1Ixp33_ASAP7_75t_L   g09241(.A1(new_n8902), .A2(new_n9496), .B(new_n9158), .C(new_n9497), .Y(new_n9498));
  XNOR2x2_ASAP7_75t_L       g09242(.A(\a[41] ), .B(new_n9426), .Y(new_n9499));
  OAI21xp33_ASAP7_75t_L     g09243(.A1(new_n9490), .A2(new_n9486), .B(new_n9499), .Y(new_n9500));
  NAND2xp33_ASAP7_75t_L     g09244(.A(new_n9500), .B(new_n9494), .Y(new_n9501));
  NOR2xp33_ASAP7_75t_L      g09245(.A(new_n9498), .B(new_n9501), .Y(new_n9502));
  OAI21xp33_ASAP7_75t_L     g09246(.A1(new_n9495), .A2(new_n9502), .B(new_n9421), .Y(new_n9503));
  XNOR2x2_ASAP7_75t_L       g09247(.A(new_n4906), .B(new_n9420), .Y(new_n9504));
  A2O1A1Ixp33_ASAP7_75t_L   g09248(.A1(new_n9144), .A2(new_n9160), .B(new_n9150), .C(new_n9161), .Y(new_n9505));
  A2O1A1Ixp33_ASAP7_75t_L   g09249(.A1(new_n9157), .A2(new_n9505), .B(new_n9174), .C(new_n9501), .Y(new_n9506));
  NAND3xp33_ASAP7_75t_L     g09250(.A(new_n9424), .B(new_n9494), .C(new_n9500), .Y(new_n9507));
  NAND3xp33_ASAP7_75t_L     g09251(.A(new_n9506), .B(new_n9504), .C(new_n9507), .Y(new_n9508));
  NAND3xp33_ASAP7_75t_L     g09252(.A(new_n9418), .B(new_n9503), .C(new_n9508), .Y(new_n9509));
  NOR3xp33_ASAP7_75t_L      g09253(.A(new_n9177), .B(new_n9178), .C(new_n9174), .Y(new_n9510));
  AOI21xp33_ASAP7_75t_L     g09254(.A1(new_n9417), .A2(new_n9178), .B(new_n9510), .Y(new_n9511));
  AOI21xp33_ASAP7_75t_L     g09255(.A1(new_n9506), .A2(new_n9507), .B(new_n9504), .Y(new_n9512));
  NOR3xp33_ASAP7_75t_L      g09256(.A(new_n9502), .B(new_n9495), .C(new_n9421), .Y(new_n9513));
  OAI221xp5_ASAP7_75t_L     g09257(.A1(new_n9512), .A2(new_n9513), .B1(new_n9181), .B2(new_n9511), .C(new_n9417), .Y(new_n9514));
  NOR2xp33_ASAP7_75t_L      g09258(.A(new_n1745), .B(new_n4147), .Y(new_n9515));
  AOI221xp5_ASAP7_75t_L     g09259(.A1(\b[18] ), .A2(new_n4402), .B1(\b[19] ), .B2(new_n4155), .C(new_n9515), .Y(new_n9516));
  O2A1O1Ixp33_ASAP7_75t_L   g09260(.A1(new_n4150), .A2(new_n1754), .B(new_n9516), .C(new_n4145), .Y(new_n9517));
  OAI21xp33_ASAP7_75t_L     g09261(.A1(new_n4150), .A2(new_n1754), .B(new_n9516), .Y(new_n9518));
  NAND2xp33_ASAP7_75t_L     g09262(.A(new_n4145), .B(new_n9518), .Y(new_n9519));
  OAI21xp33_ASAP7_75t_L     g09263(.A1(new_n4145), .A2(new_n9517), .B(new_n9519), .Y(new_n9520));
  AOI21xp33_ASAP7_75t_L     g09264(.A1(new_n9514), .A2(new_n9509), .B(new_n9520), .Y(new_n9521));
  OAI21xp33_ASAP7_75t_L     g09265(.A1(new_n9512), .A2(new_n9513), .B(new_n9418), .Y(new_n9522));
  NOR3xp33_ASAP7_75t_L      g09266(.A(new_n9502), .B(new_n9495), .C(new_n9504), .Y(new_n9523));
  O2A1O1Ixp33_ASAP7_75t_L   g09267(.A1(new_n9504), .A2(new_n9523), .B(new_n9508), .C(new_n9418), .Y(new_n9524));
  OA21x2_ASAP7_75t_L        g09268(.A1(new_n4145), .A2(new_n9517), .B(new_n9519), .Y(new_n9525));
  AOI211xp5_ASAP7_75t_L     g09269(.A1(new_n9522), .A2(new_n9418), .B(new_n9524), .C(new_n9525), .Y(new_n9526));
  OAI22xp33_ASAP7_75t_L     g09270(.A1(new_n9192), .A2(new_n9416), .B1(new_n9521), .B2(new_n9526), .Y(new_n9527));
  INVx1_ASAP7_75t_L         g09271(.A(new_n8565), .Y(new_n9528));
  A2O1A1Ixp33_ASAP7_75t_L   g09272(.A1(new_n8266), .A2(new_n8464), .B(new_n8575), .C(new_n9528), .Y(new_n9529));
  A2O1A1Ixp33_ASAP7_75t_L   g09273(.A1(new_n9529), .A2(new_n8912), .B(new_n8910), .C(new_n9193), .Y(new_n9530));
  A2O1A1Ixp33_ASAP7_75t_L   g09274(.A1(new_n9522), .A2(new_n9418), .B(new_n9524), .C(new_n9525), .Y(new_n9531));
  NAND3xp33_ASAP7_75t_L     g09275(.A(new_n9514), .B(new_n9509), .C(new_n9520), .Y(new_n9532));
  NAND4xp25_ASAP7_75t_L     g09276(.A(new_n9530), .B(new_n9531), .C(new_n9532), .D(new_n9190), .Y(new_n9533));
  AOI21xp33_ASAP7_75t_L     g09277(.A1(new_n9533), .A2(new_n9527), .B(new_n9415), .Y(new_n9534));
  O2A1O1Ixp33_ASAP7_75t_L   g09278(.A1(new_n3513), .A2(new_n2194), .B(new_n9411), .C(new_n3493), .Y(new_n9535));
  INVx1_ASAP7_75t_L         g09279(.A(new_n9414), .Y(new_n9536));
  OAI21xp33_ASAP7_75t_L     g09280(.A1(new_n3493), .A2(new_n9535), .B(new_n9536), .Y(new_n9537));
  AOI22xp33_ASAP7_75t_L     g09281(.A1(new_n9531), .A2(new_n9532), .B1(new_n9190), .B2(new_n9530), .Y(new_n9538));
  NOR4xp25_ASAP7_75t_L      g09282(.A(new_n9192), .B(new_n9526), .C(new_n9416), .D(new_n9521), .Y(new_n9539));
  NOR3xp33_ASAP7_75t_L      g09283(.A(new_n9538), .B(new_n9539), .C(new_n9537), .Y(new_n9540));
  NOR2xp33_ASAP7_75t_L      g09284(.A(new_n9534), .B(new_n9540), .Y(new_n9541));
  A2O1A1Ixp33_ASAP7_75t_L   g09285(.A1(new_n9199), .A2(new_n9409), .B(new_n9195), .C(new_n9541), .Y(new_n9542));
  INVx1_ASAP7_75t_L         g09286(.A(new_n9195), .Y(new_n9543));
  AOI21xp33_ASAP7_75t_L     g09287(.A1(new_n8930), .A2(new_n8927), .B(new_n9077), .Y(new_n9544));
  OAI221xp5_ASAP7_75t_L     g09288(.A1(new_n9534), .A2(new_n9540), .B1(new_n9206), .B2(new_n9544), .C(new_n9543), .Y(new_n9545));
  NOR2xp33_ASAP7_75t_L      g09289(.A(new_n2377), .B(new_n2925), .Y(new_n9546));
  AOI221xp5_ASAP7_75t_L     g09290(.A1(\b[24] ), .A2(new_n3129), .B1(\b[26] ), .B2(new_n2938), .C(new_n9546), .Y(new_n9547));
  O2A1O1Ixp33_ASAP7_75t_L   g09291(.A1(new_n2940), .A2(new_n2708), .B(new_n9547), .C(new_n2928), .Y(new_n9548));
  INVx1_ASAP7_75t_L         g09292(.A(new_n9548), .Y(new_n9549));
  O2A1O1Ixp33_ASAP7_75t_L   g09293(.A1(new_n2940), .A2(new_n2708), .B(new_n9547), .C(\a[29] ), .Y(new_n9550));
  AOI21xp33_ASAP7_75t_L     g09294(.A1(new_n9549), .A2(\a[29] ), .B(new_n9550), .Y(new_n9551));
  NAND3xp33_ASAP7_75t_L     g09295(.A(new_n9542), .B(new_n9545), .C(new_n9551), .Y(new_n9552));
  OAI21xp33_ASAP7_75t_L     g09296(.A1(new_n9539), .A2(new_n9538), .B(new_n9537), .Y(new_n9553));
  NAND3xp33_ASAP7_75t_L     g09297(.A(new_n9533), .B(new_n9415), .C(new_n9527), .Y(new_n9554));
  NAND2xp33_ASAP7_75t_L     g09298(.A(new_n9554), .B(new_n9553), .Y(new_n9555));
  O2A1O1Ixp33_ASAP7_75t_L   g09299(.A1(new_n9206), .A2(new_n9544), .B(new_n9543), .C(new_n9555), .Y(new_n9556));
  AOI221xp5_ASAP7_75t_L     g09300(.A1(new_n9554), .A2(new_n9553), .B1(new_n9199), .B2(new_n9409), .C(new_n9195), .Y(new_n9557));
  INVx1_ASAP7_75t_L         g09301(.A(new_n9551), .Y(new_n9558));
  OAI21xp33_ASAP7_75t_L     g09302(.A1(new_n9557), .A2(new_n9556), .B(new_n9558), .Y(new_n9559));
  NAND3xp33_ASAP7_75t_L     g09303(.A(new_n9408), .B(new_n9552), .C(new_n9559), .Y(new_n9560));
  NOR2xp33_ASAP7_75t_L      g09304(.A(new_n9207), .B(new_n9200), .Y(new_n9561));
  MAJIxp5_ASAP7_75t_L       g09305(.A(new_n9218), .B(new_n9210), .C(new_n9561), .Y(new_n9562));
  NAND2xp33_ASAP7_75t_L     g09306(.A(new_n9559), .B(new_n9552), .Y(new_n9563));
  NAND2xp33_ASAP7_75t_L     g09307(.A(new_n9562), .B(new_n9563), .Y(new_n9564));
  AOI21xp33_ASAP7_75t_L     g09308(.A1(new_n9560), .A2(new_n9564), .B(new_n9406), .Y(new_n9565));
  NOR2xp33_ASAP7_75t_L      g09309(.A(new_n9562), .B(new_n9563), .Y(new_n9566));
  NOR2xp33_ASAP7_75t_L      g09310(.A(new_n9214), .B(new_n9407), .Y(new_n9567));
  NAND2xp33_ASAP7_75t_L     g09311(.A(new_n9219), .B(new_n9220), .Y(new_n9568));
  AOI221xp5_ASAP7_75t_L     g09312(.A1(new_n9552), .A2(new_n9559), .B1(new_n9218), .B2(new_n9568), .C(new_n9567), .Y(new_n9569));
  NOR3xp33_ASAP7_75t_L      g09313(.A(new_n9566), .B(new_n9569), .C(new_n9405), .Y(new_n9570));
  NOR3xp33_ASAP7_75t_L      g09314(.A(new_n9402), .B(new_n9565), .C(new_n9570), .Y(new_n9571));
  AO21x2_ASAP7_75t_L        g09315(.A1(new_n9234), .A2(new_n9075), .B(new_n9401), .Y(new_n9572));
  OAI21xp33_ASAP7_75t_L     g09316(.A1(new_n9569), .A2(new_n9566), .B(new_n9405), .Y(new_n9573));
  NAND3xp33_ASAP7_75t_L     g09317(.A(new_n9406), .B(new_n9560), .C(new_n9564), .Y(new_n9574));
  AOI21xp33_ASAP7_75t_L     g09318(.A1(new_n9574), .A2(new_n9573), .B(new_n9572), .Y(new_n9575));
  OAI21xp33_ASAP7_75t_L     g09319(.A1(new_n9571), .A2(new_n9575), .B(new_n9400), .Y(new_n9576));
  OR3x1_ASAP7_75t_L         g09320(.A(new_n9575), .B(new_n9400), .C(new_n9571), .Y(new_n9577));
  NAND3xp33_ASAP7_75t_L     g09321(.A(new_n9393), .B(new_n9576), .C(new_n9577), .Y(new_n9578));
  NOR2xp33_ASAP7_75t_L      g09322(.A(new_n9235), .B(new_n9240), .Y(new_n9579));
  MAJIxp5_ASAP7_75t_L       g09323(.A(new_n9254), .B(new_n9246), .C(new_n9579), .Y(new_n9580));
  OA21x2_ASAP7_75t_L        g09324(.A1(new_n9571), .A2(new_n9575), .B(new_n9400), .Y(new_n9581));
  NOR3xp33_ASAP7_75t_L      g09325(.A(new_n9575), .B(new_n9571), .C(new_n9400), .Y(new_n9582));
  OAI21xp33_ASAP7_75t_L     g09326(.A1(new_n9581), .A2(new_n9582), .B(new_n9580), .Y(new_n9583));
  NOR2xp33_ASAP7_75t_L      g09327(.A(new_n4344), .B(new_n1517), .Y(new_n9584));
  AOI221xp5_ASAP7_75t_L     g09328(.A1(\b[33] ), .A2(new_n1659), .B1(\b[35] ), .B2(new_n1511), .C(new_n9584), .Y(new_n9585));
  INVx1_ASAP7_75t_L         g09329(.A(new_n9585), .Y(new_n9586));
  O2A1O1Ixp33_ASAP7_75t_L   g09330(.A1(new_n1521), .A2(new_n4589), .B(new_n9585), .C(new_n1501), .Y(new_n9587));
  INVx1_ASAP7_75t_L         g09331(.A(new_n9587), .Y(new_n9588));
  NOR2xp33_ASAP7_75t_L      g09332(.A(new_n1501), .B(new_n9587), .Y(new_n9589));
  A2O1A1O1Ixp25_ASAP7_75t_L g09333(.A1(new_n7773), .A2(new_n1513), .B(new_n9586), .C(new_n9588), .D(new_n9589), .Y(new_n9590));
  NAND3xp33_ASAP7_75t_L     g09334(.A(new_n9578), .B(new_n9583), .C(new_n9590), .Y(new_n9591));
  NOR3xp33_ASAP7_75t_L      g09335(.A(new_n9580), .B(new_n9581), .C(new_n9582), .Y(new_n9592));
  AOI21xp33_ASAP7_75t_L     g09336(.A1(new_n9577), .A2(new_n9576), .B(new_n9393), .Y(new_n9593));
  O2A1O1Ixp33_ASAP7_75t_L   g09337(.A1(new_n1521), .A2(new_n4589), .B(new_n9585), .C(\a[20] ), .Y(new_n9594));
  OAI22xp33_ASAP7_75t_L     g09338(.A1(new_n9592), .A2(new_n9593), .B1(new_n9594), .B2(new_n9589), .Y(new_n9595));
  AND2x2_ASAP7_75t_L        g09339(.A(new_n9591), .B(new_n9595), .Y(new_n9596));
  NAND3xp33_ASAP7_75t_L     g09340(.A(new_n9268), .B(new_n9269), .C(new_n9266), .Y(new_n9597));
  INVx1_ASAP7_75t_L         g09341(.A(new_n9597), .Y(new_n9598));
  O2A1O1Ixp33_ASAP7_75t_L   g09342(.A1(new_n9267), .A2(new_n9271), .B(new_n9278), .C(new_n9598), .Y(new_n9599));
  NAND2xp33_ASAP7_75t_L     g09343(.A(new_n9599), .B(new_n9596), .Y(new_n9600));
  NAND2xp33_ASAP7_75t_L     g09344(.A(new_n9591), .B(new_n9595), .Y(new_n9601));
  OAI21xp33_ASAP7_75t_L     g09345(.A1(new_n9272), .A2(new_n9274), .B(new_n9597), .Y(new_n9602));
  NAND2xp33_ASAP7_75t_L     g09346(.A(new_n9601), .B(new_n9602), .Y(new_n9603));
  OAI22xp33_ASAP7_75t_L     g09347(.A1(new_n1285), .A2(new_n4613), .B1(new_n5074), .B2(new_n2118), .Y(new_n9604));
  AOI221xp5_ASAP7_75t_L     g09348(.A1(new_n1209), .A2(\b[38] ), .B1(new_n1216), .B2(new_n6083), .C(new_n9604), .Y(new_n9605));
  XNOR2x2_ASAP7_75t_L       g09349(.A(\a[17] ), .B(new_n9605), .Y(new_n9606));
  INVx1_ASAP7_75t_L         g09350(.A(new_n9606), .Y(new_n9607));
  NAND3xp33_ASAP7_75t_L     g09351(.A(new_n9607), .B(new_n9603), .C(new_n9600), .Y(new_n9608));
  NOR2xp33_ASAP7_75t_L      g09352(.A(new_n9601), .B(new_n9602), .Y(new_n9609));
  AOI22xp33_ASAP7_75t_L     g09353(.A1(new_n9591), .A2(new_n9595), .B1(new_n9597), .B2(new_n9279), .Y(new_n9610));
  OAI21xp33_ASAP7_75t_L     g09354(.A1(new_n9610), .A2(new_n9609), .B(new_n9606), .Y(new_n9611));
  NAND4xp25_ASAP7_75t_L     g09355(.A(new_n9301), .B(new_n9608), .C(new_n9611), .D(new_n9391), .Y(new_n9612));
  NOR3xp33_ASAP7_75t_L      g09356(.A(new_n9609), .B(new_n9610), .C(new_n9606), .Y(new_n9613));
  AOI21xp33_ASAP7_75t_L     g09357(.A1(new_n9600), .A2(new_n9603), .B(new_n9607), .Y(new_n9614));
  MAJIxp5_ASAP7_75t_L       g09358(.A(new_n9289), .B(new_n9389), .C(new_n9285), .Y(new_n9615));
  OAI21xp33_ASAP7_75t_L     g09359(.A1(new_n9613), .A2(new_n9614), .B(new_n9615), .Y(new_n9616));
  NOR2xp33_ASAP7_75t_L      g09360(.A(new_n6110), .B(new_n869), .Y(new_n9617));
  AOI221xp5_ASAP7_75t_L     g09361(.A1(\b[39] ), .A2(new_n985), .B1(\b[40] ), .B2(new_n885), .C(new_n9617), .Y(new_n9618));
  O2A1O1Ixp33_ASAP7_75t_L   g09362(.A1(new_n872), .A2(new_n6117), .B(new_n9618), .C(new_n867), .Y(new_n9619));
  OAI21xp33_ASAP7_75t_L     g09363(.A1(new_n872), .A2(new_n6117), .B(new_n9618), .Y(new_n9620));
  NAND2xp33_ASAP7_75t_L     g09364(.A(new_n867), .B(new_n9620), .Y(new_n9621));
  OAI21xp33_ASAP7_75t_L     g09365(.A1(new_n867), .A2(new_n9619), .B(new_n9621), .Y(new_n9622));
  INVx1_ASAP7_75t_L         g09366(.A(new_n9622), .Y(new_n9623));
  NAND3xp33_ASAP7_75t_L     g09367(.A(new_n9612), .B(new_n9623), .C(new_n9616), .Y(new_n9624));
  NOR3xp33_ASAP7_75t_L      g09368(.A(new_n9615), .B(new_n9614), .C(new_n9613), .Y(new_n9625));
  OA21x2_ASAP7_75t_L        g09369(.A1(new_n9613), .A2(new_n9614), .B(new_n9615), .Y(new_n9626));
  OAI21xp33_ASAP7_75t_L     g09370(.A1(new_n9625), .A2(new_n9626), .B(new_n9622), .Y(new_n9627));
  AND4x1_ASAP7_75t_L        g09371(.A(new_n9306), .B(new_n9388), .C(new_n9627), .D(new_n9624), .Y(new_n9628));
  MAJIxp5_ASAP7_75t_L       g09372(.A(new_n9305), .B(new_n9298), .C(new_n9387), .Y(new_n9629));
  AOI21xp33_ASAP7_75t_L     g09373(.A1(new_n9627), .A2(new_n9624), .B(new_n9629), .Y(new_n9630));
  NOR2xp33_ASAP7_75t_L      g09374(.A(new_n6944), .B(new_n710), .Y(new_n9631));
  AOI221xp5_ASAP7_75t_L     g09375(.A1(\b[43] ), .A2(new_n635), .B1(\b[42] ), .B2(new_n713), .C(new_n9631), .Y(new_n9632));
  O2A1O1Ixp33_ASAP7_75t_L   g09376(.A1(new_n641), .A2(new_n6951), .B(new_n9632), .C(new_n637), .Y(new_n9633));
  OAI21xp33_ASAP7_75t_L     g09377(.A1(new_n641), .A2(new_n6951), .B(new_n9632), .Y(new_n9634));
  NAND2xp33_ASAP7_75t_L     g09378(.A(new_n637), .B(new_n9634), .Y(new_n9635));
  OAI21xp33_ASAP7_75t_L     g09379(.A1(new_n637), .A2(new_n9633), .B(new_n9635), .Y(new_n9636));
  INVx1_ASAP7_75t_L         g09380(.A(new_n9636), .Y(new_n9637));
  NOR3xp33_ASAP7_75t_L      g09381(.A(new_n9628), .B(new_n9630), .C(new_n9637), .Y(new_n9638));
  AND2x2_ASAP7_75t_L        g09382(.A(new_n9624), .B(new_n9627), .Y(new_n9639));
  NAND2xp33_ASAP7_75t_L     g09383(.A(new_n9629), .B(new_n9639), .Y(new_n9640));
  INVx1_ASAP7_75t_L         g09384(.A(new_n9388), .Y(new_n9641));
  NAND2xp33_ASAP7_75t_L     g09385(.A(new_n9624), .B(new_n9627), .Y(new_n9642));
  A2O1A1Ixp33_ASAP7_75t_L   g09386(.A1(new_n9316), .A2(new_n9305), .B(new_n9641), .C(new_n9642), .Y(new_n9643));
  AOI21xp33_ASAP7_75t_L     g09387(.A1(new_n9640), .A2(new_n9643), .B(new_n9636), .Y(new_n9644));
  OAI22xp33_ASAP7_75t_L     g09388(.A1(new_n9313), .A2(new_n9327), .B1(new_n9644), .B2(new_n9638), .Y(new_n9645));
  NAND3xp33_ASAP7_75t_L     g09389(.A(new_n9640), .B(new_n9643), .C(new_n9636), .Y(new_n9646));
  OAI21xp33_ASAP7_75t_L     g09390(.A1(new_n9630), .A2(new_n9628), .B(new_n9637), .Y(new_n9647));
  NAND3xp33_ASAP7_75t_L     g09391(.A(new_n9328), .B(new_n9646), .C(new_n9647), .Y(new_n9648));
  NOR2xp33_ASAP7_75t_L      g09392(.A(new_n7249), .B(new_n506), .Y(new_n9649));
  AOI221xp5_ASAP7_75t_L     g09393(.A1(\b[47] ), .A2(new_n475), .B1(new_n470), .B2(\b[46] ), .C(new_n9649), .Y(new_n9650));
  O2A1O1Ixp33_ASAP7_75t_L   g09394(.A1(new_n477), .A2(new_n7560), .B(new_n9650), .C(new_n466), .Y(new_n9651));
  OAI21xp33_ASAP7_75t_L     g09395(.A1(new_n477), .A2(new_n7560), .B(new_n9650), .Y(new_n9652));
  NAND2xp33_ASAP7_75t_L     g09396(.A(new_n466), .B(new_n9652), .Y(new_n9653));
  OAI21xp33_ASAP7_75t_L     g09397(.A1(new_n466), .A2(new_n9651), .B(new_n9653), .Y(new_n9654));
  AOI21xp33_ASAP7_75t_L     g09398(.A1(new_n9645), .A2(new_n9648), .B(new_n9654), .Y(new_n9655));
  AOI21xp33_ASAP7_75t_L     g09399(.A1(new_n9647), .A2(new_n9646), .B(new_n9328), .Y(new_n9656));
  NOR4xp25_ASAP7_75t_L      g09400(.A(new_n9313), .B(new_n9644), .C(new_n9327), .D(new_n9638), .Y(new_n9657));
  INVx1_ASAP7_75t_L         g09401(.A(new_n9654), .Y(new_n9658));
  NOR3xp33_ASAP7_75t_L      g09402(.A(new_n9657), .B(new_n9658), .C(new_n9656), .Y(new_n9659));
  NOR2xp33_ASAP7_75t_L      g09403(.A(new_n9655), .B(new_n9659), .Y(new_n9660));
  A2O1A1O1Ixp25_ASAP7_75t_L g09404(.A1(new_n9311), .A2(new_n9313), .B(new_n9070), .C(new_n9320), .D(new_n9323), .Y(new_n9661));
  O2A1O1Ixp33_ASAP7_75t_L   g09405(.A1(new_n9325), .A2(new_n9329), .B(new_n9348), .C(new_n9661), .Y(new_n9662));
  NAND2xp33_ASAP7_75t_L     g09406(.A(new_n9662), .B(new_n9660), .Y(new_n9663));
  OAI21xp33_ASAP7_75t_L     g09407(.A1(new_n9656), .A2(new_n9657), .B(new_n9658), .Y(new_n9664));
  NAND3xp33_ASAP7_75t_L     g09408(.A(new_n9645), .B(new_n9648), .C(new_n9654), .Y(new_n9665));
  NAND2xp33_ASAP7_75t_L     g09409(.A(new_n9665), .B(new_n9664), .Y(new_n9666));
  OAI21xp33_ASAP7_75t_L     g09410(.A1(new_n9661), .A2(new_n9339), .B(new_n9666), .Y(new_n9667));
  OAI22xp33_ASAP7_75t_L     g09411(.A1(new_n350), .A2(new_n8427), .B1(new_n7860), .B2(new_n375), .Y(new_n9668));
  AOI221xp5_ASAP7_75t_L     g09412(.A1(new_n361), .A2(\b[50] ), .B1(new_n359), .B2(new_n8763), .C(new_n9668), .Y(new_n9669));
  XNOR2x2_ASAP7_75t_L       g09413(.A(new_n346), .B(new_n9669), .Y(new_n9670));
  INVx1_ASAP7_75t_L         g09414(.A(new_n9670), .Y(new_n9671));
  NAND3xp33_ASAP7_75t_L     g09415(.A(new_n9663), .B(new_n9667), .C(new_n9671), .Y(new_n9672));
  NOR3xp33_ASAP7_75t_L      g09416(.A(new_n9666), .B(new_n9339), .C(new_n9661), .Y(new_n9673));
  NOR2xp33_ASAP7_75t_L      g09417(.A(new_n9662), .B(new_n9660), .Y(new_n9674));
  OAI21xp33_ASAP7_75t_L     g09418(.A1(new_n9674), .A2(new_n9673), .B(new_n9670), .Y(new_n9675));
  NAND3xp33_ASAP7_75t_L     g09419(.A(new_n9386), .B(new_n9672), .C(new_n9675), .Y(new_n9676));
  NOR3xp33_ASAP7_75t_L      g09420(.A(new_n9673), .B(new_n9674), .C(new_n9670), .Y(new_n9677));
  AOI21xp33_ASAP7_75t_L     g09421(.A1(new_n9663), .A2(new_n9667), .B(new_n9671), .Y(new_n9678));
  NOR3xp33_ASAP7_75t_L      g09422(.A(new_n9386), .B(new_n9677), .C(new_n9678), .Y(new_n9679));
  NOR2xp33_ASAP7_75t_L      g09423(.A(new_n8779), .B(new_n287), .Y(new_n9680));
  AOI221xp5_ASAP7_75t_L     g09424(.A1(\b[52] ), .A2(new_n264), .B1(\b[53] ), .B2(new_n283), .C(new_n9680), .Y(new_n9681));
  NOR2xp33_ASAP7_75t_L      g09425(.A(\b[52] ), .B(\b[53] ), .Y(new_n9682));
  INVx1_ASAP7_75t_L         g09426(.A(\b[53] ), .Y(new_n9683));
  NOR2xp33_ASAP7_75t_L      g09427(.A(new_n9355), .B(new_n9683), .Y(new_n9684));
  NOR2xp33_ASAP7_75t_L      g09428(.A(new_n9682), .B(new_n9684), .Y(new_n9685));
  A2O1A1Ixp33_ASAP7_75t_L   g09429(.A1(new_n9365), .A2(new_n9361), .B(new_n9360), .C(new_n9685), .Y(new_n9686));
  A2O1A1O1Ixp25_ASAP7_75t_L g09430(.A1(new_n8784), .A2(new_n9358), .B(new_n8783), .C(new_n9361), .D(new_n9360), .Y(new_n9687));
  INVx1_ASAP7_75t_L         g09431(.A(new_n9685), .Y(new_n9688));
  NAND2xp33_ASAP7_75t_L     g09432(.A(new_n9688), .B(new_n9687), .Y(new_n9689));
  AND2x2_ASAP7_75t_L        g09433(.A(new_n9689), .B(new_n9686), .Y(new_n9690));
  INVx1_ASAP7_75t_L         g09434(.A(new_n9690), .Y(new_n9691));
  O2A1O1Ixp33_ASAP7_75t_L   g09435(.A1(new_n279), .A2(new_n9691), .B(new_n9681), .C(new_n257), .Y(new_n9692));
  OAI21xp33_ASAP7_75t_L     g09436(.A1(new_n279), .A2(new_n9691), .B(new_n9681), .Y(new_n9693));
  NAND2xp33_ASAP7_75t_L     g09437(.A(new_n257), .B(new_n9693), .Y(new_n9694));
  OA21x2_ASAP7_75t_L        g09438(.A1(new_n257), .A2(new_n9692), .B(new_n9694), .Y(new_n9695));
  A2O1A1Ixp33_ASAP7_75t_L   g09439(.A1(new_n9676), .A2(new_n9386), .B(new_n9679), .C(new_n9695), .Y(new_n9696));
  AOI21xp33_ASAP7_75t_L     g09440(.A1(new_n9676), .A2(new_n9386), .B(new_n9679), .Y(new_n9697));
  INVx1_ASAP7_75t_L         g09441(.A(new_n9695), .Y(new_n9698));
  NAND2xp33_ASAP7_75t_L     g09442(.A(new_n9698), .B(new_n9697), .Y(new_n9699));
  AOI21xp33_ASAP7_75t_L     g09443(.A1(new_n9699), .A2(new_n9696), .B(new_n9383), .Y(new_n9700));
  AND3x1_ASAP7_75t_L        g09444(.A(new_n9699), .B(new_n9696), .C(new_n9383), .Y(new_n9701));
  NOR2xp33_ASAP7_75t_L      g09445(.A(new_n9700), .B(new_n9701), .Y(\f[53] ));
  A2O1A1Ixp33_ASAP7_75t_L   g09446(.A1(new_n9676), .A2(new_n9386), .B(new_n9679), .C(new_n9698), .Y(new_n9703));
  NOR2xp33_ASAP7_75t_L      g09447(.A(new_n9355), .B(new_n287), .Y(new_n9704));
  AOI221xp5_ASAP7_75t_L     g09448(.A1(\b[53] ), .A2(new_n264), .B1(\b[54] ), .B2(new_n283), .C(new_n9704), .Y(new_n9705));
  INVx1_ASAP7_75t_L         g09449(.A(new_n9360), .Y(new_n9706));
  A2O1A1O1Ixp25_ASAP7_75t_L g09450(.A1(new_n9364), .A2(new_n8785), .B(new_n9359), .C(new_n9706), .D(new_n9688), .Y(new_n9707));
  NOR2xp33_ASAP7_75t_L      g09451(.A(\b[53] ), .B(\b[54] ), .Y(new_n9708));
  INVx1_ASAP7_75t_L         g09452(.A(\b[54] ), .Y(new_n9709));
  NOR2xp33_ASAP7_75t_L      g09453(.A(new_n9683), .B(new_n9709), .Y(new_n9710));
  NOR2xp33_ASAP7_75t_L      g09454(.A(new_n9708), .B(new_n9710), .Y(new_n9711));
  A2O1A1Ixp33_ASAP7_75t_L   g09455(.A1(\b[53] ), .A2(\b[52] ), .B(new_n9707), .C(new_n9711), .Y(new_n9712));
  INVx1_ASAP7_75t_L         g09456(.A(new_n9712), .Y(new_n9713));
  INVx1_ASAP7_75t_L         g09457(.A(new_n9684), .Y(new_n9714));
  A2O1A1Ixp33_ASAP7_75t_L   g09458(.A1(new_n9362), .A2(new_n9706), .B(new_n9688), .C(new_n9714), .Y(new_n9715));
  NOR2xp33_ASAP7_75t_L      g09459(.A(new_n9711), .B(new_n9715), .Y(new_n9716));
  NOR2xp33_ASAP7_75t_L      g09460(.A(new_n9716), .B(new_n9713), .Y(new_n9717));
  INVx1_ASAP7_75t_L         g09461(.A(new_n9717), .Y(new_n9718));
  O2A1O1Ixp33_ASAP7_75t_L   g09462(.A1(new_n279), .A2(new_n9718), .B(new_n9705), .C(new_n257), .Y(new_n9719));
  NOR2xp33_ASAP7_75t_L      g09463(.A(new_n257), .B(new_n9719), .Y(new_n9720));
  O2A1O1Ixp33_ASAP7_75t_L   g09464(.A1(new_n279), .A2(new_n9718), .B(new_n9705), .C(\a[2] ), .Y(new_n9721));
  NOR2xp33_ASAP7_75t_L      g09465(.A(new_n9721), .B(new_n9720), .Y(new_n9722));
  NOR2xp33_ASAP7_75t_L      g09466(.A(new_n9342), .B(new_n9384), .Y(new_n9723));
  A2O1A1O1Ixp25_ASAP7_75t_L g09467(.A1(new_n9375), .A2(new_n9377), .B(new_n9723), .C(new_n9675), .D(new_n9677), .Y(new_n9724));
  NOR2xp33_ASAP7_75t_L      g09468(.A(new_n7270), .B(new_n506), .Y(new_n9725));
  AOI221xp5_ASAP7_75t_L     g09469(.A1(\b[48] ), .A2(new_n475), .B1(new_n470), .B2(\b[47] ), .C(new_n9725), .Y(new_n9726));
  O2A1O1Ixp33_ASAP7_75t_L   g09470(.A1(new_n477), .A2(new_n7868), .B(new_n9726), .C(new_n466), .Y(new_n9727));
  OAI21xp33_ASAP7_75t_L     g09471(.A1(new_n477), .A2(new_n7868), .B(new_n9726), .Y(new_n9728));
  NAND2xp33_ASAP7_75t_L     g09472(.A(new_n466), .B(new_n9728), .Y(new_n9729));
  OAI21xp33_ASAP7_75t_L     g09473(.A1(new_n466), .A2(new_n9727), .B(new_n9729), .Y(new_n9730));
  A2O1A1Ixp33_ASAP7_75t_L   g09474(.A1(new_n9026), .A2(new_n9020), .B(new_n9069), .C(new_n9319), .Y(new_n9731));
  A2O1A1Ixp33_ASAP7_75t_L   g09475(.A1(new_n9731), .A2(new_n9311), .B(new_n9644), .C(new_n9646), .Y(new_n9732));
  NOR2xp33_ASAP7_75t_L      g09476(.A(new_n7249), .B(new_n710), .Y(new_n9733));
  AOI221xp5_ASAP7_75t_L     g09477(.A1(\b[44] ), .A2(new_n635), .B1(\b[43] ), .B2(new_n713), .C(new_n9733), .Y(new_n9734));
  O2A1O1Ixp33_ASAP7_75t_L   g09478(.A1(new_n641), .A2(new_n7255), .B(new_n9734), .C(new_n637), .Y(new_n9735));
  OAI21xp33_ASAP7_75t_L     g09479(.A1(new_n641), .A2(new_n7255), .B(new_n9734), .Y(new_n9736));
  NAND2xp33_ASAP7_75t_L     g09480(.A(new_n637), .B(new_n9736), .Y(new_n9737));
  OAI21xp33_ASAP7_75t_L     g09481(.A1(new_n637), .A2(new_n9735), .B(new_n9737), .Y(new_n9738));
  INVx1_ASAP7_75t_L         g09482(.A(new_n9738), .Y(new_n9739));
  NAND3xp33_ASAP7_75t_L     g09483(.A(new_n9612), .B(new_n9616), .C(new_n9622), .Y(new_n9740));
  A2O1A1Ixp33_ASAP7_75t_L   g09484(.A1(new_n9623), .A2(new_n9624), .B(new_n9629), .C(new_n9740), .Y(new_n9741));
  NAND2xp33_ASAP7_75t_L     g09485(.A(new_n9583), .B(new_n9578), .Y(new_n9742));
  INVx1_ASAP7_75t_L         g09486(.A(new_n9742), .Y(new_n9743));
  A2O1A1Ixp33_ASAP7_75t_L   g09487(.A1(\a[20] ), .A2(new_n9588), .B(new_n9594), .C(new_n9743), .Y(new_n9744));
  A2O1A1Ixp33_ASAP7_75t_L   g09488(.A1(\a[23] ), .A2(new_n9250), .B(new_n9244), .C(new_n9579), .Y(new_n9745));
  A2O1A1Ixp33_ASAP7_75t_L   g09489(.A1(new_n9269), .A2(new_n9745), .B(new_n9581), .C(new_n9577), .Y(new_n9746));
  A2O1A1O1Ixp25_ASAP7_75t_L g09490(.A1(new_n9075), .A2(new_n9234), .B(new_n9401), .C(new_n9573), .D(new_n9570), .Y(new_n9747));
  OAI22xp33_ASAP7_75t_L     g09491(.A1(new_n2572), .A2(new_n3079), .B1(new_n3098), .B2(new_n2410), .Y(new_n9748));
  AOI221xp5_ASAP7_75t_L     g09492(.A1(new_n2423), .A2(\b[30] ), .B1(new_n2417), .B2(new_n4813), .C(new_n9748), .Y(new_n9749));
  XNOR2x2_ASAP7_75t_L       g09493(.A(new_n2413), .B(new_n9749), .Y(new_n9750));
  O2A1O1Ixp33_ASAP7_75t_L   g09494(.A1(new_n9206), .A2(new_n9544), .B(new_n9543), .C(new_n9541), .Y(new_n9751));
  O2A1O1Ixp33_ASAP7_75t_L   g09495(.A1(new_n9541), .A2(new_n9751), .B(new_n9542), .C(new_n9551), .Y(new_n9752));
  A2O1A1O1Ixp25_ASAP7_75t_L g09496(.A1(new_n9218), .A2(new_n9568), .B(new_n9567), .C(new_n9552), .D(new_n9752), .Y(new_n9753));
  NOR2xp33_ASAP7_75t_L      g09497(.A(new_n2703), .B(new_n2925), .Y(new_n9754));
  AOI221xp5_ASAP7_75t_L     g09498(.A1(\b[25] ), .A2(new_n3129), .B1(\b[27] ), .B2(new_n2938), .C(new_n9754), .Y(new_n9755));
  O2A1O1Ixp33_ASAP7_75t_L   g09499(.A1(new_n2940), .A2(new_n2889), .B(new_n9755), .C(new_n2928), .Y(new_n9756));
  INVx1_ASAP7_75t_L         g09500(.A(new_n9756), .Y(new_n9757));
  O2A1O1Ixp33_ASAP7_75t_L   g09501(.A1(new_n2940), .A2(new_n2889), .B(new_n9755), .C(\a[29] ), .Y(new_n9758));
  AOI21xp33_ASAP7_75t_L     g09502(.A1(new_n9757), .A2(\a[29] ), .B(new_n9758), .Y(new_n9759));
  NAND2xp33_ASAP7_75t_L     g09503(.A(new_n9527), .B(new_n9533), .Y(new_n9760));
  O2A1O1Ixp33_ASAP7_75t_L   g09504(.A1(new_n3493), .A2(new_n9535), .B(new_n9536), .C(new_n9760), .Y(new_n9761));
  A2O1A1O1Ixp25_ASAP7_75t_L g09505(.A1(new_n9199), .A2(new_n9409), .B(new_n9195), .C(new_n9555), .D(new_n9761), .Y(new_n9762));
  OAI22xp33_ASAP7_75t_L     g09506(.A1(new_n3703), .A2(new_n2045), .B1(new_n2188), .B2(new_n3509), .Y(new_n9763));
  AOI221xp5_ASAP7_75t_L     g09507(.A1(new_n3503), .A2(\b[24] ), .B1(new_n3505), .B2(new_n2216), .C(new_n9763), .Y(new_n9764));
  XNOR2x2_ASAP7_75t_L       g09508(.A(\a[32] ), .B(new_n9764), .Y(new_n9765));
  A2O1A1Ixp33_ASAP7_75t_L   g09509(.A1(new_n9522), .A2(new_n9418), .B(new_n9524), .C(new_n9520), .Y(new_n9766));
  INVx1_ASAP7_75t_L         g09510(.A(new_n9766), .Y(new_n9767));
  NAND2xp33_ASAP7_75t_L     g09511(.A(\b[20] ), .B(new_n4155), .Y(new_n9768));
  OAI221xp5_ASAP7_75t_L     g09512(.A1(new_n4147), .A2(new_n1895), .B1(new_n1599), .B2(new_n4397), .C(new_n9768), .Y(new_n9769));
  A2O1A1Ixp33_ASAP7_75t_L   g09513(.A1(new_n2836), .A2(new_n4151), .B(new_n9769), .C(\a[35] ), .Y(new_n9770));
  AOI211xp5_ASAP7_75t_L     g09514(.A1(new_n2836), .A2(new_n4151), .B(new_n9769), .C(new_n4145), .Y(new_n9771));
  A2O1A1O1Ixp25_ASAP7_75t_L g09515(.A1(new_n4151), .A2(new_n2836), .B(new_n9769), .C(new_n9770), .D(new_n9771), .Y(new_n9772));
  INVx1_ASAP7_75t_L         g09516(.A(new_n9772), .Y(new_n9773));
  NAND2xp33_ASAP7_75t_L     g09517(.A(new_n9503), .B(new_n9508), .Y(new_n9774));
  NOR2xp33_ASAP7_75t_L      g09518(.A(new_n1458), .B(new_n4908), .Y(new_n9775));
  AOI221xp5_ASAP7_75t_L     g09519(.A1(\b[16] ), .A2(new_n5139), .B1(\b[17] ), .B2(new_n4916), .C(new_n9775), .Y(new_n9776));
  O2A1O1Ixp33_ASAP7_75t_L   g09520(.A1(new_n4911), .A2(new_n1464), .B(new_n9776), .C(new_n4906), .Y(new_n9777));
  OAI21xp33_ASAP7_75t_L     g09521(.A1(new_n4911), .A2(new_n1464), .B(new_n9776), .Y(new_n9778));
  NAND2xp33_ASAP7_75t_L     g09522(.A(new_n4906), .B(new_n9778), .Y(new_n9779));
  OA21x2_ASAP7_75t_L        g09523(.A1(new_n4906), .A2(new_n9777), .B(new_n9779), .Y(new_n9780));
  NOR2xp33_ASAP7_75t_L      g09524(.A(new_n960), .B(new_n5640), .Y(new_n9781));
  AOI221xp5_ASAP7_75t_L     g09525(.A1(\b[13] ), .A2(new_n5920), .B1(\b[15] ), .B2(new_n5629), .C(new_n9781), .Y(new_n9782));
  INVx1_ASAP7_75t_L         g09526(.A(new_n9782), .Y(new_n9783));
  A2O1A1Ixp33_ASAP7_75t_L   g09527(.A1(new_n1052), .A2(new_n5637), .B(new_n9783), .C(\a[41] ), .Y(new_n9784));
  O2A1O1Ixp33_ASAP7_75t_L   g09528(.A1(new_n5630), .A2(new_n1774), .B(new_n9782), .C(\a[41] ), .Y(new_n9785));
  AOI21xp33_ASAP7_75t_L     g09529(.A1(new_n9784), .A2(\a[41] ), .B(new_n9785), .Y(new_n9786));
  A2O1A1Ixp33_ASAP7_75t_L   g09530(.A1(new_n9149), .A2(new_n9144), .B(new_n9482), .C(new_n9489), .Y(new_n9787));
  NOR2xp33_ASAP7_75t_L      g09531(.A(new_n680), .B(new_n6741), .Y(new_n9788));
  AOI221xp5_ASAP7_75t_L     g09532(.A1(\b[12] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[11] ), .C(new_n9788), .Y(new_n9789));
  OA211x2_ASAP7_75t_L       g09533(.A1(new_n6443), .A2(new_n841), .B(\a[44] ), .C(new_n9789), .Y(new_n9790));
  O2A1O1Ixp33_ASAP7_75t_L   g09534(.A1(new_n6443), .A2(new_n841), .B(new_n9789), .C(\a[44] ), .Y(new_n9791));
  NOR2xp33_ASAP7_75t_L      g09535(.A(new_n9791), .B(new_n9790), .Y(new_n9792));
  INVx1_ASAP7_75t_L         g09536(.A(new_n9792), .Y(new_n9793));
  NOR2xp33_ASAP7_75t_L      g09537(.A(new_n534), .B(new_n7312), .Y(new_n9794));
  AOI221xp5_ASAP7_75t_L     g09538(.A1(\b[7] ), .A2(new_n7609), .B1(\b[9] ), .B2(new_n7334), .C(new_n9794), .Y(new_n9795));
  O2A1O1Ixp33_ASAP7_75t_L   g09539(.A1(new_n7321), .A2(new_n1066), .B(new_n9795), .C(new_n7316), .Y(new_n9796));
  INVx1_ASAP7_75t_L         g09540(.A(new_n9796), .Y(new_n9797));
  O2A1O1Ixp33_ASAP7_75t_L   g09541(.A1(new_n7321), .A2(new_n1066), .B(new_n9795), .C(\a[47] ), .Y(new_n9798));
  AOI21xp33_ASAP7_75t_L     g09542(.A1(new_n9797), .A2(\a[47] ), .B(new_n9798), .Y(new_n9799));
  O2A1O1Ixp33_ASAP7_75t_L   g09543(.A1(new_n9120), .A2(new_n9121), .B(new_n9118), .C(new_n9461), .Y(new_n9800));
  INVx1_ASAP7_75t_L         g09544(.A(\a[54] ), .Y(new_n9801));
  NAND2xp33_ASAP7_75t_L     g09545(.A(\a[53] ), .B(new_n9801), .Y(new_n9802));
  NAND2xp33_ASAP7_75t_L     g09546(.A(\a[54] ), .B(new_n9099), .Y(new_n9803));
  AND2x2_ASAP7_75t_L        g09547(.A(new_n9802), .B(new_n9803), .Y(new_n9804));
  NOR2xp33_ASAP7_75t_L      g09548(.A(new_n284), .B(new_n9804), .Y(new_n9805));
  A2O1A1Ixp33_ASAP7_75t_L   g09549(.A1(new_n9458), .A2(new_n9444), .B(new_n9106), .C(new_n9805), .Y(new_n9806));
  A2O1A1Ixp33_ASAP7_75t_L   g09550(.A1(new_n9802), .A2(new_n9803), .B(new_n284), .C(new_n9449), .Y(new_n9807));
  NAND2xp33_ASAP7_75t_L     g09551(.A(\b[2] ), .B(new_n9096), .Y(new_n9808));
  OAI221xp5_ASAP7_75t_L     g09552(.A1(new_n9440), .A2(new_n262), .B1(new_n301), .B2(new_n9439), .C(new_n9808), .Y(new_n9809));
  NOR2xp33_ASAP7_75t_L      g09553(.A(new_n9104), .B(new_n319), .Y(new_n9810));
  A2O1A1Ixp33_ASAP7_75t_L   g09554(.A1(new_n312), .A2(new_n9437), .B(new_n9809), .C(\a[53] ), .Y(new_n9811));
  NOR3xp33_ASAP7_75t_L      g09555(.A(new_n9809), .B(new_n9810), .C(new_n9099), .Y(new_n9812));
  O2A1O1Ixp33_ASAP7_75t_L   g09556(.A1(new_n9809), .A2(new_n9810), .B(new_n9811), .C(new_n9812), .Y(new_n9813));
  AOI21xp33_ASAP7_75t_L     g09557(.A1(new_n9806), .A2(new_n9807), .B(new_n9813), .Y(new_n9814));
  INVx1_ASAP7_75t_L         g09558(.A(new_n9805), .Y(new_n9815));
  NOR2xp33_ASAP7_75t_L      g09559(.A(new_n9815), .B(new_n9449), .Y(new_n9816));
  NOR2xp33_ASAP7_75t_L      g09560(.A(new_n9805), .B(new_n9460), .Y(new_n9817));
  INVx1_ASAP7_75t_L         g09561(.A(new_n9813), .Y(new_n9818));
  NOR3xp33_ASAP7_75t_L      g09562(.A(new_n9818), .B(new_n9817), .C(new_n9816), .Y(new_n9819));
  NAND2xp33_ASAP7_75t_L     g09563(.A(\b[5] ), .B(new_n8169), .Y(new_n9820));
  OAI221xp5_ASAP7_75t_L     g09564(.A1(new_n8483), .A2(new_n332), .B1(new_n427), .B2(new_n8843), .C(new_n9820), .Y(new_n9821));
  A2O1A1Ixp33_ASAP7_75t_L   g09565(.A1(new_n5363), .A2(new_n8490), .B(new_n9821), .C(\a[50] ), .Y(new_n9822));
  NAND2xp33_ASAP7_75t_L     g09566(.A(\a[50] ), .B(new_n9822), .Y(new_n9823));
  A2O1A1Ixp33_ASAP7_75t_L   g09567(.A1(new_n5363), .A2(new_n8490), .B(new_n9821), .C(new_n8172), .Y(new_n9824));
  NAND2xp33_ASAP7_75t_L     g09568(.A(new_n9824), .B(new_n9823), .Y(new_n9825));
  NOR3xp33_ASAP7_75t_L      g09569(.A(new_n9814), .B(new_n9819), .C(new_n9825), .Y(new_n9826));
  OAI21xp33_ASAP7_75t_L     g09570(.A1(new_n9816), .A2(new_n9817), .B(new_n9818), .Y(new_n9827));
  NAND3xp33_ASAP7_75t_L     g09571(.A(new_n9806), .B(new_n9807), .C(new_n9813), .Y(new_n9828));
  INVx1_ASAP7_75t_L         g09572(.A(new_n9825), .Y(new_n9829));
  AOI21xp33_ASAP7_75t_L     g09573(.A1(new_n9828), .A2(new_n9827), .B(new_n9829), .Y(new_n9830));
  OAI22xp33_ASAP7_75t_L     g09574(.A1(new_n9830), .A2(new_n9826), .B1(new_n9456), .B2(new_n9800), .Y(new_n9831));
  NOR2xp33_ASAP7_75t_L      g09575(.A(new_n9826), .B(new_n9830), .Y(new_n9832));
  NAND2xp33_ASAP7_75t_L     g09576(.A(new_n9475), .B(new_n9832), .Y(new_n9833));
  AO21x2_ASAP7_75t_L        g09577(.A1(new_n9831), .A2(new_n9833), .B(new_n9799), .Y(new_n9834));
  A2O1A1O1Ixp25_ASAP7_75t_L g09578(.A1(new_n9464), .A2(new_n9800), .B(new_n9463), .C(new_n9466), .D(new_n9472), .Y(new_n9835));
  A2O1A1O1Ixp25_ASAP7_75t_L g09579(.A1(new_n9138), .A2(new_n9137), .B(new_n9435), .C(new_n9473), .D(new_n9835), .Y(new_n9836));
  NAND3xp33_ASAP7_75t_L     g09580(.A(new_n9833), .B(new_n9831), .C(new_n9799), .Y(new_n9837));
  AOI21xp33_ASAP7_75t_L     g09581(.A1(new_n9834), .A2(new_n9837), .B(new_n9836), .Y(new_n9838));
  AND2x2_ASAP7_75t_L        g09582(.A(new_n9837), .B(new_n9836), .Y(new_n9839));
  A2O1A1Ixp33_ASAP7_75t_L   g09583(.A1(new_n9839), .A2(new_n9834), .B(new_n9838), .C(new_n9793), .Y(new_n9840));
  AO21x2_ASAP7_75t_L        g09584(.A1(new_n9837), .A2(new_n9834), .B(new_n9836), .Y(new_n9841));
  NAND3xp33_ASAP7_75t_L     g09585(.A(new_n9836), .B(new_n9834), .C(new_n9837), .Y(new_n9842));
  NAND3xp33_ASAP7_75t_L     g09586(.A(new_n9841), .B(new_n9792), .C(new_n9842), .Y(new_n9843));
  NAND2xp33_ASAP7_75t_L     g09587(.A(new_n9843), .B(new_n9840), .Y(new_n9844));
  AND3x1_ASAP7_75t_L        g09588(.A(new_n9841), .B(new_n9842), .C(new_n9792), .Y(new_n9845));
  AOI211xp5_ASAP7_75t_L     g09589(.A1(new_n9487), .A2(new_n9488), .B(new_n9485), .C(new_n9845), .Y(new_n9846));
  AOI221xp5_ASAP7_75t_L     g09590(.A1(new_n9787), .A2(new_n9844), .B1(new_n9840), .B2(new_n9846), .C(new_n9786), .Y(new_n9847));
  AO21x2_ASAP7_75t_L        g09591(.A1(\a[41] ), .A2(new_n9784), .B(new_n9785), .Y(new_n9848));
  INVx1_ASAP7_75t_L         g09592(.A(new_n9798), .Y(new_n9849));
  NAND2xp33_ASAP7_75t_L     g09593(.A(new_n9831), .B(new_n9833), .Y(new_n9850));
  INVx1_ASAP7_75t_L         g09594(.A(new_n9850), .Y(new_n9851));
  O2A1O1Ixp33_ASAP7_75t_L   g09595(.A1(new_n7316), .A2(new_n9796), .B(new_n9849), .C(new_n9851), .Y(new_n9852));
  NAND2xp33_ASAP7_75t_L     g09596(.A(new_n9837), .B(new_n9836), .Y(new_n9853));
  O2A1O1Ixp33_ASAP7_75t_L   g09597(.A1(new_n9853), .A2(new_n9852), .B(new_n9841), .C(new_n9792), .Y(new_n9854));
  OAI21xp33_ASAP7_75t_L     g09598(.A1(new_n9854), .A2(new_n9845), .B(new_n9787), .Y(new_n9855));
  OAI211xp5_ASAP7_75t_L     g09599(.A1(new_n9482), .A2(new_n9429), .B(new_n9489), .C(new_n9843), .Y(new_n9856));
  O2A1O1Ixp33_ASAP7_75t_L   g09600(.A1(new_n9854), .A2(new_n9856), .B(new_n9855), .C(new_n9848), .Y(new_n9857));
  NOR2xp33_ASAP7_75t_L      g09601(.A(new_n9847), .B(new_n9857), .Y(new_n9858));
  A2O1A1Ixp33_ASAP7_75t_L   g09602(.A1(new_n9501), .A2(new_n9498), .B(new_n9491), .C(new_n9858), .Y(new_n9859));
  INVx1_ASAP7_75t_L         g09603(.A(new_n9491), .Y(new_n9860));
  AND2x2_ASAP7_75t_L        g09604(.A(new_n9500), .B(new_n9494), .Y(new_n9861));
  OAI221xp5_ASAP7_75t_L     g09605(.A1(new_n9847), .A2(new_n9857), .B1(new_n9424), .B2(new_n9861), .C(new_n9860), .Y(new_n9862));
  AO21x2_ASAP7_75t_L        g09606(.A1(new_n9862), .A2(new_n9859), .B(new_n9780), .Y(new_n9863));
  NAND3xp33_ASAP7_75t_L     g09607(.A(new_n9859), .B(new_n9780), .C(new_n9862), .Y(new_n9864));
  NAND2xp33_ASAP7_75t_L     g09608(.A(new_n9864), .B(new_n9863), .Y(new_n9865));
  A2O1A1Ixp33_ASAP7_75t_L   g09609(.A1(new_n9774), .A2(new_n9418), .B(new_n9523), .C(new_n9865), .Y(new_n9866));
  O2A1O1Ixp33_ASAP7_75t_L   g09610(.A1(new_n9512), .A2(new_n9513), .B(new_n9418), .C(new_n9523), .Y(new_n9867));
  NAND3xp33_ASAP7_75t_L     g09611(.A(new_n9867), .B(new_n9863), .C(new_n9864), .Y(new_n9868));
  NAND3xp33_ASAP7_75t_L     g09612(.A(new_n9866), .B(new_n9773), .C(new_n9868), .Y(new_n9869));
  AOI21xp33_ASAP7_75t_L     g09613(.A1(new_n9864), .A2(new_n9863), .B(new_n9867), .Y(new_n9870));
  AND3x1_ASAP7_75t_L        g09614(.A(new_n9859), .B(new_n9780), .C(new_n9862), .Y(new_n9871));
  AOI211xp5_ASAP7_75t_L     g09615(.A1(new_n9774), .A2(new_n9418), .B(new_n9523), .C(new_n9871), .Y(new_n9872));
  A2O1A1Ixp33_ASAP7_75t_L   g09616(.A1(new_n9872), .A2(new_n9863), .B(new_n9870), .C(new_n9772), .Y(new_n9873));
  OAI211xp5_ASAP7_75t_L     g09617(.A1(new_n9767), .A2(new_n9538), .B(new_n9869), .C(new_n9873), .Y(new_n9874));
  OAI21xp33_ASAP7_75t_L     g09618(.A1(new_n9191), .A2(new_n9084), .B(new_n9190), .Y(new_n9875));
  O2A1O1Ixp33_ASAP7_75t_L   g09619(.A1(new_n9521), .A2(new_n9526), .B(new_n9875), .C(new_n9767), .Y(new_n9876));
  AOI211xp5_ASAP7_75t_L     g09620(.A1(new_n9863), .A2(new_n9872), .B(new_n9772), .C(new_n9870), .Y(new_n9877));
  INVx1_ASAP7_75t_L         g09621(.A(new_n9865), .Y(new_n9878));
  O2A1O1Ixp33_ASAP7_75t_L   g09622(.A1(new_n9867), .A2(new_n9878), .B(new_n9868), .C(new_n9773), .Y(new_n9879));
  OAI21xp33_ASAP7_75t_L     g09623(.A1(new_n9877), .A2(new_n9879), .B(new_n9876), .Y(new_n9880));
  NAND3xp33_ASAP7_75t_L     g09624(.A(new_n9874), .B(new_n9765), .C(new_n9880), .Y(new_n9881));
  XNOR2x2_ASAP7_75t_L       g09625(.A(new_n3493), .B(new_n9764), .Y(new_n9882));
  AOI211xp5_ASAP7_75t_L     g09626(.A1(new_n9527), .A2(new_n9766), .B(new_n9877), .C(new_n9879), .Y(new_n9883));
  AOI211xp5_ASAP7_75t_L     g09627(.A1(new_n9873), .A2(new_n9869), .B(new_n9767), .C(new_n9538), .Y(new_n9884));
  OAI21xp33_ASAP7_75t_L     g09628(.A1(new_n9883), .A2(new_n9884), .B(new_n9882), .Y(new_n9885));
  NAND2xp33_ASAP7_75t_L     g09629(.A(new_n9885), .B(new_n9881), .Y(new_n9886));
  NOR2xp33_ASAP7_75t_L      g09630(.A(new_n9762), .B(new_n9886), .Y(new_n9887));
  OAI21xp33_ASAP7_75t_L     g09631(.A1(new_n9206), .A2(new_n9544), .B(new_n9543), .Y(new_n9888));
  AOI221xp5_ASAP7_75t_L     g09632(.A1(new_n9885), .A2(new_n9881), .B1(new_n9555), .B2(new_n9888), .C(new_n9761), .Y(new_n9889));
  NOR3xp33_ASAP7_75t_L      g09633(.A(new_n9887), .B(new_n9889), .C(new_n9759), .Y(new_n9890));
  INVx1_ASAP7_75t_L         g09634(.A(new_n9759), .Y(new_n9891));
  INVx1_ASAP7_75t_L         g09635(.A(new_n9761), .Y(new_n9892));
  A2O1A1Ixp33_ASAP7_75t_L   g09636(.A1(new_n9213), .A2(new_n9543), .B(new_n9541), .C(new_n9892), .Y(new_n9893));
  AND2x2_ASAP7_75t_L        g09637(.A(new_n9885), .B(new_n9881), .Y(new_n9894));
  NAND2xp33_ASAP7_75t_L     g09638(.A(new_n9894), .B(new_n9893), .Y(new_n9895));
  NAND2xp33_ASAP7_75t_L     g09639(.A(new_n9762), .B(new_n9886), .Y(new_n9896));
  AOI21xp33_ASAP7_75t_L     g09640(.A1(new_n9895), .A2(new_n9896), .B(new_n9891), .Y(new_n9897));
  NOR3xp33_ASAP7_75t_L      g09641(.A(new_n9753), .B(new_n9890), .C(new_n9897), .Y(new_n9898));
  NAND3xp33_ASAP7_75t_L     g09642(.A(new_n9895), .B(new_n9891), .C(new_n9896), .Y(new_n9899));
  OAI21xp33_ASAP7_75t_L     g09643(.A1(new_n9889), .A2(new_n9887), .B(new_n9759), .Y(new_n9900));
  AOI221xp5_ASAP7_75t_L     g09644(.A1(new_n9408), .A2(new_n9552), .B1(new_n9900), .B2(new_n9899), .C(new_n9752), .Y(new_n9901));
  NOR3xp33_ASAP7_75t_L      g09645(.A(new_n9898), .B(new_n9901), .C(new_n9750), .Y(new_n9902));
  XNOR2x2_ASAP7_75t_L       g09646(.A(\a[26] ), .B(new_n9749), .Y(new_n9903));
  INVx1_ASAP7_75t_L         g09647(.A(new_n9552), .Y(new_n9904));
  OAI21xp33_ASAP7_75t_L     g09648(.A1(new_n9904), .A2(new_n9562), .B(new_n9559), .Y(new_n9905));
  NAND3xp33_ASAP7_75t_L     g09649(.A(new_n9905), .B(new_n9899), .C(new_n9900), .Y(new_n9906));
  OAI21xp33_ASAP7_75t_L     g09650(.A1(new_n9890), .A2(new_n9897), .B(new_n9753), .Y(new_n9907));
  AOI21xp33_ASAP7_75t_L     g09651(.A1(new_n9906), .A2(new_n9907), .B(new_n9903), .Y(new_n9908));
  NOR3xp33_ASAP7_75t_L      g09652(.A(new_n9747), .B(new_n9902), .C(new_n9908), .Y(new_n9909));
  NAND3xp33_ASAP7_75t_L     g09653(.A(new_n9906), .B(new_n9903), .C(new_n9907), .Y(new_n9910));
  OAI21xp33_ASAP7_75t_L     g09654(.A1(new_n9901), .A2(new_n9898), .B(new_n9750), .Y(new_n9911));
  AOI221xp5_ASAP7_75t_L     g09655(.A1(new_n9572), .A2(new_n9573), .B1(new_n9910), .B2(new_n9911), .C(new_n9570), .Y(new_n9912));
  NOR2xp33_ASAP7_75t_L      g09656(.A(new_n3891), .B(new_n1962), .Y(new_n9913));
  AOI221xp5_ASAP7_75t_L     g09657(.A1(new_n1955), .A2(\b[33] ), .B1(new_n2093), .B2(\b[31] ), .C(new_n9913), .Y(new_n9914));
  O2A1O1Ixp33_ASAP7_75t_L   g09658(.A1(new_n1956), .A2(new_n4108), .B(new_n9914), .C(new_n1952), .Y(new_n9915));
  INVx1_ASAP7_75t_L         g09659(.A(new_n9914), .Y(new_n9916));
  A2O1A1Ixp33_ASAP7_75t_L   g09660(.A1(new_n4831), .A2(new_n1964), .B(new_n9916), .C(new_n1952), .Y(new_n9917));
  OAI21xp33_ASAP7_75t_L     g09661(.A1(new_n1952), .A2(new_n9915), .B(new_n9917), .Y(new_n9918));
  NOR3xp33_ASAP7_75t_L      g09662(.A(new_n9912), .B(new_n9909), .C(new_n9918), .Y(new_n9919));
  OAI21xp33_ASAP7_75t_L     g09663(.A1(new_n9565), .A2(new_n9402), .B(new_n9574), .Y(new_n9920));
  NAND3xp33_ASAP7_75t_L     g09664(.A(new_n9920), .B(new_n9910), .C(new_n9911), .Y(new_n9921));
  OAI21xp33_ASAP7_75t_L     g09665(.A1(new_n9908), .A2(new_n9902), .B(new_n9747), .Y(new_n9922));
  INVx1_ASAP7_75t_L         g09666(.A(new_n9915), .Y(new_n9923));
  NOR2xp33_ASAP7_75t_L      g09667(.A(new_n1952), .B(new_n9915), .Y(new_n9924));
  A2O1A1O1Ixp25_ASAP7_75t_L g09668(.A1(new_n4831), .A2(new_n1964), .B(new_n9916), .C(new_n9923), .D(new_n9924), .Y(new_n9925));
  AOI21xp33_ASAP7_75t_L     g09669(.A1(new_n9921), .A2(new_n9922), .B(new_n9925), .Y(new_n9926));
  NOR2xp33_ASAP7_75t_L      g09670(.A(new_n9919), .B(new_n9926), .Y(new_n9927));
  NAND2xp33_ASAP7_75t_L     g09671(.A(new_n9746), .B(new_n9927), .Y(new_n9928));
  O2A1O1Ixp33_ASAP7_75t_L   g09672(.A1(new_n9243), .A2(new_n1952), .B(new_n9245), .C(new_n9392), .Y(new_n9929));
  NAND2xp33_ASAP7_75t_L     g09673(.A(new_n9256), .B(new_n9257), .Y(new_n9930));
  A2O1A1O1Ixp25_ASAP7_75t_L g09674(.A1(new_n9254), .A2(new_n9930), .B(new_n9929), .C(new_n9576), .D(new_n9582), .Y(new_n9931));
  NAND3xp33_ASAP7_75t_L     g09675(.A(new_n9921), .B(new_n9922), .C(new_n9925), .Y(new_n9932));
  OAI21xp33_ASAP7_75t_L     g09676(.A1(new_n9909), .A2(new_n9912), .B(new_n9918), .Y(new_n9933));
  NAND2xp33_ASAP7_75t_L     g09677(.A(new_n9933), .B(new_n9932), .Y(new_n9934));
  NAND2xp33_ASAP7_75t_L     g09678(.A(new_n9931), .B(new_n9934), .Y(new_n9935));
  OAI22xp33_ASAP7_75t_L     g09679(.A1(new_n1654), .A2(new_n4344), .B1(new_n4581), .B2(new_n1517), .Y(new_n9936));
  AOI221xp5_ASAP7_75t_L     g09680(.A1(new_n1511), .A2(\b[36] ), .B1(new_n1513), .B2(new_n4621), .C(new_n9936), .Y(new_n9937));
  XNOR2x2_ASAP7_75t_L       g09681(.A(new_n1501), .B(new_n9937), .Y(new_n9938));
  AOI21xp33_ASAP7_75t_L     g09682(.A1(new_n9928), .A2(new_n9935), .B(new_n9938), .Y(new_n9939));
  NOR2xp33_ASAP7_75t_L      g09683(.A(new_n9931), .B(new_n9934), .Y(new_n9940));
  AOI221xp5_ASAP7_75t_L     g09684(.A1(new_n9932), .A2(new_n9933), .B1(new_n9393), .B2(new_n9576), .C(new_n9582), .Y(new_n9941));
  XNOR2x2_ASAP7_75t_L       g09685(.A(\a[20] ), .B(new_n9937), .Y(new_n9942));
  NOR3xp33_ASAP7_75t_L      g09686(.A(new_n9940), .B(new_n9941), .C(new_n9942), .Y(new_n9943));
  OAI221xp5_ASAP7_75t_L     g09687(.A1(new_n9939), .A2(new_n9943), .B1(new_n9599), .B2(new_n9596), .C(new_n9744), .Y(new_n9944));
  INVx1_ASAP7_75t_L         g09688(.A(new_n9594), .Y(new_n9945));
  O2A1O1Ixp33_ASAP7_75t_L   g09689(.A1(new_n9587), .A2(new_n1501), .B(new_n9945), .C(new_n9742), .Y(new_n9946));
  NOR2xp33_ASAP7_75t_L      g09690(.A(new_n9943), .B(new_n9939), .Y(new_n9947));
  OAI21xp33_ASAP7_75t_L     g09691(.A1(new_n9946), .A2(new_n9610), .B(new_n9947), .Y(new_n9948));
  NOR2xp33_ASAP7_75t_L      g09692(.A(new_n5311), .B(new_n2118), .Y(new_n9949));
  AOI221xp5_ASAP7_75t_L     g09693(.A1(\b[37] ), .A2(new_n1290), .B1(\b[39] ), .B2(new_n1209), .C(new_n9949), .Y(new_n9950));
  O2A1O1Ixp33_ASAP7_75t_L   g09694(.A1(new_n1210), .A2(new_n5578), .B(new_n9950), .C(new_n1206), .Y(new_n9951));
  INVx1_ASAP7_75t_L         g09695(.A(new_n9951), .Y(new_n9952));
  O2A1O1Ixp33_ASAP7_75t_L   g09696(.A1(new_n1210), .A2(new_n5578), .B(new_n9950), .C(\a[17] ), .Y(new_n9953));
  AOI21xp33_ASAP7_75t_L     g09697(.A1(new_n9952), .A2(\a[17] ), .B(new_n9953), .Y(new_n9954));
  NAND3xp33_ASAP7_75t_L     g09698(.A(new_n9948), .B(new_n9944), .C(new_n9954), .Y(new_n9955));
  OAI21xp33_ASAP7_75t_L     g09699(.A1(new_n9941), .A2(new_n9940), .B(new_n9942), .Y(new_n9956));
  NAND3xp33_ASAP7_75t_L     g09700(.A(new_n9928), .B(new_n9935), .C(new_n9938), .Y(new_n9957));
  AOI221xp5_ASAP7_75t_L     g09701(.A1(new_n9957), .A2(new_n9956), .B1(new_n9601), .B2(new_n9602), .C(new_n9946), .Y(new_n9958));
  NAND2xp33_ASAP7_75t_L     g09702(.A(new_n9956), .B(new_n9957), .Y(new_n9959));
  O2A1O1Ixp33_ASAP7_75t_L   g09703(.A1(new_n9596), .A2(new_n9599), .B(new_n9744), .C(new_n9959), .Y(new_n9960));
  INVx1_ASAP7_75t_L         g09704(.A(new_n9954), .Y(new_n9961));
  OAI21xp33_ASAP7_75t_L     g09705(.A1(new_n9958), .A2(new_n9960), .B(new_n9961), .Y(new_n9962));
  NOR2xp33_ASAP7_75t_L      g09706(.A(new_n9610), .B(new_n9609), .Y(new_n9963));
  MAJIxp5_ASAP7_75t_L       g09707(.A(new_n9615), .B(new_n9963), .C(new_n9606), .Y(new_n9964));
  NAND3xp33_ASAP7_75t_L     g09708(.A(new_n9964), .B(new_n9962), .C(new_n9955), .Y(new_n9965));
  NAND2xp33_ASAP7_75t_L     g09709(.A(new_n9606), .B(new_n9963), .Y(new_n9966));
  INVx1_ASAP7_75t_L         g09710(.A(new_n9966), .Y(new_n9967));
  NAND2xp33_ASAP7_75t_L     g09711(.A(new_n9611), .B(new_n9608), .Y(new_n9968));
  NAND2xp33_ASAP7_75t_L     g09712(.A(new_n9955), .B(new_n9962), .Y(new_n9969));
  A2O1A1Ixp33_ASAP7_75t_L   g09713(.A1(new_n9968), .A2(new_n9615), .B(new_n9967), .C(new_n9969), .Y(new_n9970));
  OAI22xp33_ASAP7_75t_L     g09714(.A1(new_n980), .A2(new_n5855), .B1(new_n6110), .B2(new_n864), .Y(new_n9971));
  AOI221xp5_ASAP7_75t_L     g09715(.A1(new_n886), .A2(\b[42] ), .B1(new_n873), .B2(new_n6389), .C(new_n9971), .Y(new_n9972));
  XNOR2x2_ASAP7_75t_L       g09716(.A(\a[14] ), .B(new_n9972), .Y(new_n9973));
  AOI21xp33_ASAP7_75t_L     g09717(.A1(new_n9970), .A2(new_n9965), .B(new_n9973), .Y(new_n9974));
  AND4x1_ASAP7_75t_L        g09718(.A(new_n9616), .B(new_n9966), .C(new_n9962), .D(new_n9955), .Y(new_n9975));
  AOI21xp33_ASAP7_75t_L     g09719(.A1(new_n9962), .A2(new_n9955), .B(new_n9964), .Y(new_n9976));
  XNOR2x2_ASAP7_75t_L       g09720(.A(new_n867), .B(new_n9972), .Y(new_n9977));
  NOR3xp33_ASAP7_75t_L      g09721(.A(new_n9975), .B(new_n9976), .C(new_n9977), .Y(new_n9978));
  NOR2xp33_ASAP7_75t_L      g09722(.A(new_n9974), .B(new_n9978), .Y(new_n9979));
  NAND2xp33_ASAP7_75t_L     g09723(.A(new_n9979), .B(new_n9741), .Y(new_n9980));
  OAI221xp5_ASAP7_75t_L     g09724(.A1(new_n9974), .A2(new_n9978), .B1(new_n9629), .B2(new_n9639), .C(new_n9740), .Y(new_n9981));
  AOI21xp33_ASAP7_75t_L     g09725(.A1(new_n9980), .A2(new_n9981), .B(new_n9739), .Y(new_n9982));
  OAI21xp33_ASAP7_75t_L     g09726(.A1(new_n9976), .A2(new_n9975), .B(new_n9977), .Y(new_n9983));
  NAND3xp33_ASAP7_75t_L     g09727(.A(new_n9970), .B(new_n9965), .C(new_n9973), .Y(new_n9984));
  NAND2xp33_ASAP7_75t_L     g09728(.A(new_n9984), .B(new_n9983), .Y(new_n9985));
  O2A1O1Ixp33_ASAP7_75t_L   g09729(.A1(new_n9639), .A2(new_n9629), .B(new_n9740), .C(new_n9985), .Y(new_n9986));
  INVx1_ASAP7_75t_L         g09730(.A(new_n9740), .Y(new_n9987));
  A2O1A1Ixp33_ASAP7_75t_L   g09731(.A1(new_n9022), .A2(new_n9073), .B(new_n9303), .C(new_n9388), .Y(new_n9988));
  AOI221xp5_ASAP7_75t_L     g09732(.A1(new_n9983), .A2(new_n9984), .B1(new_n9642), .B2(new_n9988), .C(new_n9987), .Y(new_n9989));
  NOR3xp33_ASAP7_75t_L      g09733(.A(new_n9986), .B(new_n9989), .C(new_n9738), .Y(new_n9990));
  OAI21xp33_ASAP7_75t_L     g09734(.A1(new_n9982), .A2(new_n9990), .B(new_n9732), .Y(new_n9991));
  OAI21xp33_ASAP7_75t_L     g09735(.A1(new_n9989), .A2(new_n9986), .B(new_n9738), .Y(new_n9992));
  NAND3xp33_ASAP7_75t_L     g09736(.A(new_n9980), .B(new_n9739), .C(new_n9981), .Y(new_n9993));
  AOI21xp33_ASAP7_75t_L     g09737(.A1(new_n9993), .A2(new_n9992), .B(new_n9732), .Y(new_n9994));
  A2O1A1Ixp33_ASAP7_75t_L   g09738(.A1(new_n9991), .A2(new_n9732), .B(new_n9994), .C(new_n9730), .Y(new_n9995));
  NAND3xp33_ASAP7_75t_L     g09739(.A(new_n9732), .B(new_n9992), .C(new_n9993), .Y(new_n9996));
  A2O1A1O1Ixp25_ASAP7_75t_L g09740(.A1(new_n9319), .A2(new_n9334), .B(new_n9327), .C(new_n9647), .D(new_n9638), .Y(new_n9997));
  OAI21xp33_ASAP7_75t_L     g09741(.A1(new_n9982), .A2(new_n9990), .B(new_n9997), .Y(new_n9998));
  AOI21xp33_ASAP7_75t_L     g09742(.A1(new_n9998), .A2(new_n9996), .B(new_n9730), .Y(new_n9999));
  AOI21xp33_ASAP7_75t_L     g09743(.A1(new_n9995), .A2(new_n9730), .B(new_n9999), .Y(new_n10000));
  O2A1O1Ixp33_ASAP7_75t_L   g09744(.A1(new_n9644), .A2(new_n9732), .B(new_n9645), .C(new_n9658), .Y(new_n10001));
  O2A1O1Ixp33_ASAP7_75t_L   g09745(.A1(new_n9661), .A2(new_n9339), .B(new_n9666), .C(new_n10001), .Y(new_n10002));
  NAND2xp33_ASAP7_75t_L     g09746(.A(new_n10000), .B(new_n10002), .Y(new_n10003));
  MAJx2_ASAP7_75t_L         g09747(.A(new_n9348), .B(new_n9324), .C(new_n9346), .Y(new_n10004));
  INVx1_ASAP7_75t_L         g09748(.A(new_n9730), .Y(new_n10005));
  A2O1A1Ixp33_ASAP7_75t_L   g09749(.A1(new_n9991), .A2(new_n9732), .B(new_n9994), .C(new_n10005), .Y(new_n10006));
  NAND3xp33_ASAP7_75t_L     g09750(.A(new_n9998), .B(new_n9996), .C(new_n9730), .Y(new_n10007));
  NAND2xp33_ASAP7_75t_L     g09751(.A(new_n10007), .B(new_n10006), .Y(new_n10008));
  A2O1A1Ixp33_ASAP7_75t_L   g09752(.A1(new_n9666), .A2(new_n10004), .B(new_n10001), .C(new_n10008), .Y(new_n10009));
  OAI22xp33_ASAP7_75t_L     g09753(.A1(new_n350), .A2(new_n8755), .B1(new_n8427), .B2(new_n375), .Y(new_n10010));
  AOI221xp5_ASAP7_75t_L     g09754(.A1(new_n361), .A2(\b[51] ), .B1(new_n359), .B2(new_n8790), .C(new_n10010), .Y(new_n10011));
  XNOR2x2_ASAP7_75t_L       g09755(.A(new_n346), .B(new_n10011), .Y(new_n10012));
  INVx1_ASAP7_75t_L         g09756(.A(new_n10012), .Y(new_n10013));
  AOI21xp33_ASAP7_75t_L     g09757(.A1(new_n10003), .A2(new_n10009), .B(new_n10013), .Y(new_n10014));
  A2O1A1Ixp33_ASAP7_75t_L   g09758(.A1(new_n9027), .A2(new_n9024), .B(new_n9312), .C(new_n9311), .Y(new_n10015));
  A2O1A1Ixp33_ASAP7_75t_L   g09759(.A1(new_n9334), .A2(new_n9319), .B(new_n9327), .C(new_n9647), .Y(new_n10016));
  O2A1O1Ixp33_ASAP7_75t_L   g09760(.A1(new_n9638), .A2(new_n10016), .B(new_n10015), .C(new_n9657), .Y(new_n10017));
  INVx1_ASAP7_75t_L         g09761(.A(new_n10001), .Y(new_n10018));
  A2O1A1Ixp33_ASAP7_75t_L   g09762(.A1(new_n10017), .A2(new_n9665), .B(new_n9662), .C(new_n10018), .Y(new_n10019));
  NOR2xp33_ASAP7_75t_L      g09763(.A(new_n10008), .B(new_n10019), .Y(new_n10020));
  AOI21xp33_ASAP7_75t_L     g09764(.A1(new_n9667), .A2(new_n10018), .B(new_n10000), .Y(new_n10021));
  NOR3xp33_ASAP7_75t_L      g09765(.A(new_n10020), .B(new_n10021), .C(new_n10012), .Y(new_n10022));
  NOR3xp33_ASAP7_75t_L      g09766(.A(new_n9724), .B(new_n10014), .C(new_n10022), .Y(new_n10023));
  OAI21xp33_ASAP7_75t_L     g09767(.A1(new_n10021), .A2(new_n10020), .B(new_n10012), .Y(new_n10024));
  NAND3xp33_ASAP7_75t_L     g09768(.A(new_n10013), .B(new_n10003), .C(new_n10009), .Y(new_n10025));
  AOI221xp5_ASAP7_75t_L     g09769(.A1(new_n9386), .A2(new_n9675), .B1(new_n10024), .B2(new_n10025), .C(new_n9677), .Y(new_n10026));
  NOR3xp33_ASAP7_75t_L      g09770(.A(new_n10026), .B(new_n10023), .C(new_n9722), .Y(new_n10027));
  INVx1_ASAP7_75t_L         g09771(.A(new_n10027), .Y(new_n10028));
  OAI21xp33_ASAP7_75t_L     g09772(.A1(new_n10023), .A2(new_n10026), .B(new_n9722), .Y(new_n10029));
  NAND2xp33_ASAP7_75t_L     g09773(.A(new_n10029), .B(new_n10028), .Y(new_n10030));
  A2O1A1O1Ixp25_ASAP7_75t_L g09774(.A1(new_n9696), .A2(new_n9699), .B(new_n9383), .C(new_n9703), .D(new_n10030), .Y(new_n10031));
  MAJIxp5_ASAP7_75t_L       g09775(.A(new_n9383), .B(new_n9695), .C(new_n9697), .Y(new_n10032));
  AOI21xp33_ASAP7_75t_L     g09776(.A1(new_n10028), .A2(new_n10029), .B(new_n10032), .Y(new_n10033));
  NOR2xp33_ASAP7_75t_L      g09777(.A(new_n10033), .B(new_n10031), .Y(\f[54] ));
  O2A1O1Ixp33_ASAP7_75t_L   g09778(.A1(new_n9692), .A2(new_n257), .B(new_n9694), .C(new_n9697), .Y(new_n10035));
  O2A1O1Ixp33_ASAP7_75t_L   g09779(.A1(new_n10035), .A2(new_n9700), .B(new_n10029), .C(new_n10027), .Y(new_n10036));
  A2O1A1Ixp33_ASAP7_75t_L   g09780(.A1(new_n9377), .A2(new_n9375), .B(new_n9723), .C(new_n9675), .Y(new_n10037));
  A2O1A1Ixp33_ASAP7_75t_L   g09781(.A1(new_n10037), .A2(new_n9672), .B(new_n10014), .C(new_n10025), .Y(new_n10038));
  INVx1_ASAP7_75t_L         g09782(.A(new_n9995), .Y(new_n10039));
  OAI22xp33_ASAP7_75t_L     g09783(.A1(new_n513), .A2(new_n7860), .B1(new_n7552), .B2(new_n506), .Y(new_n10040));
  AOI221xp5_ASAP7_75t_L     g09784(.A1(new_n475), .A2(\b[49] ), .B1(new_n483), .B2(new_n8438), .C(new_n10040), .Y(new_n10041));
  XNOR2x2_ASAP7_75t_L       g09785(.A(new_n466), .B(new_n10041), .Y(new_n10042));
  INVx1_ASAP7_75t_L         g09786(.A(new_n10042), .Y(new_n10043));
  NAND2xp33_ASAP7_75t_L     g09787(.A(new_n9981), .B(new_n9980), .Y(new_n10044));
  MAJIxp5_ASAP7_75t_L       g09788(.A(new_n9997), .B(new_n9739), .C(new_n10044), .Y(new_n10045));
  A2O1A1Ixp33_ASAP7_75t_L   g09789(.A1(new_n9643), .A2(new_n9740), .B(new_n9974), .C(new_n9984), .Y(new_n10046));
  OAI22xp33_ASAP7_75t_L     g09790(.A1(new_n3703), .A2(new_n2188), .B1(new_n2205), .B2(new_n3509), .Y(new_n10047));
  AOI221xp5_ASAP7_75t_L     g09791(.A1(new_n3503), .A2(\b[25] ), .B1(new_n3505), .B2(new_n5001), .C(new_n10047), .Y(new_n10048));
  XNOR2x2_ASAP7_75t_L       g09792(.A(\a[32] ), .B(new_n10048), .Y(new_n10049));
  A2O1A1Ixp33_ASAP7_75t_L   g09793(.A1(new_n8530), .A2(new_n8517), .B(new_n8888), .C(new_n8882), .Y(new_n10050));
  A2O1A1O1Ixp25_ASAP7_75t_L g09794(.A1(new_n10050), .A2(new_n9147), .B(new_n9428), .C(new_n9488), .D(new_n9485), .Y(new_n10051));
  NAND2xp33_ASAP7_75t_L     g09795(.A(new_n9842), .B(new_n9841), .Y(new_n10052));
  NAND3xp33_ASAP7_75t_L     g09796(.A(new_n9841), .B(new_n9793), .C(new_n9842), .Y(new_n10053));
  A2O1A1Ixp33_ASAP7_75t_L   g09797(.A1(new_n9840), .A2(new_n10052), .B(new_n10051), .C(new_n10053), .Y(new_n10054));
  OAI22xp33_ASAP7_75t_L     g09798(.A1(new_n7304), .A2(new_n833), .B1(new_n748), .B2(new_n6741), .Y(new_n10055));
  AOI221xp5_ASAP7_75t_L     g09799(.A1(new_n6442), .A2(\b[13] ), .B1(new_n6450), .B2(new_n1166), .C(new_n10055), .Y(new_n10056));
  XNOR2x2_ASAP7_75t_L       g09800(.A(new_n6439), .B(new_n10056), .Y(new_n10057));
  AOI22xp33_ASAP7_75t_L     g09801(.A1(new_n7333), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n7609), .Y(new_n10058));
  OAI221xp5_ASAP7_75t_L     g09802(.A1(new_n680), .A2(new_n7318), .B1(new_n7321), .B2(new_n1175), .C(new_n10058), .Y(new_n10059));
  XNOR2x2_ASAP7_75t_L       g09803(.A(new_n7316), .B(new_n10059), .Y(new_n10060));
  NAND3xp33_ASAP7_75t_L     g09804(.A(new_n9828), .B(new_n9827), .C(new_n9825), .Y(new_n10061));
  NAND3xp33_ASAP7_75t_L     g09805(.A(new_n9829), .B(new_n9828), .C(new_n9827), .Y(new_n10062));
  A2O1A1Ixp33_ASAP7_75t_L   g09806(.A1(new_n10062), .A2(new_n9829), .B(new_n9475), .C(new_n10061), .Y(new_n10063));
  INVx1_ASAP7_75t_L         g09807(.A(new_n8168), .Y(new_n10064));
  NAND2xp33_ASAP7_75t_L     g09808(.A(new_n10064), .B(new_n7906), .Y(new_n10065));
  NOR2xp33_ASAP7_75t_L      g09809(.A(new_n427), .B(new_n10065), .Y(new_n10066));
  AOI221xp5_ASAP7_75t_L     g09810(.A1(new_n8175), .A2(\b[7] ), .B1(new_n8484), .B2(\b[5] ), .C(new_n10066), .Y(new_n10067));
  NAND2xp33_ASAP7_75t_L     g09811(.A(new_n8490), .B(new_n1188), .Y(new_n10068));
  O2A1O1Ixp33_ASAP7_75t_L   g09812(.A1(new_n8176), .A2(new_n456), .B(new_n10067), .C(new_n8172), .Y(new_n10069));
  OAI211xp5_ASAP7_75t_L     g09813(.A1(new_n8176), .A2(new_n456), .B(\a[50] ), .C(new_n10067), .Y(new_n10070));
  A2O1A1Ixp33_ASAP7_75t_L   g09814(.A1(new_n10068), .A2(new_n10067), .B(new_n10069), .C(new_n10070), .Y(new_n10071));
  MAJIxp5_ASAP7_75t_L       g09815(.A(new_n9813), .B(new_n9815), .C(new_n9460), .Y(new_n10072));
  NAND2xp33_ASAP7_75t_L     g09816(.A(\b[3] ), .B(new_n9096), .Y(new_n10073));
  OAI221xp5_ASAP7_75t_L     g09817(.A1(new_n9440), .A2(new_n289), .B1(new_n332), .B2(new_n9439), .C(new_n10073), .Y(new_n10074));
  A2O1A1Ixp33_ASAP7_75t_L   g09818(.A1(new_n342), .A2(new_n9437), .B(new_n10074), .C(\a[53] ), .Y(new_n10075));
  AOI211xp5_ASAP7_75t_L     g09819(.A1(new_n342), .A2(new_n9437), .B(new_n9099), .C(new_n10074), .Y(new_n10076));
  A2O1A1O1Ixp25_ASAP7_75t_L g09820(.A1(new_n9437), .A2(new_n342), .B(new_n10074), .C(new_n10075), .D(new_n10076), .Y(new_n10077));
  NAND2xp33_ASAP7_75t_L     g09821(.A(new_n9803), .B(new_n9802), .Y(new_n10078));
  XNOR2x2_ASAP7_75t_L       g09822(.A(\a[55] ), .B(\a[54] ), .Y(new_n10079));
  NOR2xp33_ASAP7_75t_L      g09823(.A(new_n10079), .B(new_n10078), .Y(new_n10080));
  INVx1_ASAP7_75t_L         g09824(.A(\a[55] ), .Y(new_n10081));
  NAND2xp33_ASAP7_75t_L     g09825(.A(\a[56] ), .B(new_n10081), .Y(new_n10082));
  INVx1_ASAP7_75t_L         g09826(.A(\a[56] ), .Y(new_n10083));
  NAND2xp33_ASAP7_75t_L     g09827(.A(\a[55] ), .B(new_n10083), .Y(new_n10084));
  NAND2xp33_ASAP7_75t_L     g09828(.A(new_n10084), .B(new_n10082), .Y(new_n10085));
  NOR2xp33_ASAP7_75t_L      g09829(.A(new_n10085), .B(new_n9804), .Y(new_n10086));
  AOI22xp33_ASAP7_75t_L     g09830(.A1(new_n10080), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n10086), .Y(new_n10087));
  NAND2xp33_ASAP7_75t_L     g09831(.A(new_n10085), .B(new_n10078), .Y(new_n10088));
  OAI21xp33_ASAP7_75t_L     g09832(.A1(new_n10088), .A2(new_n274), .B(new_n10087), .Y(new_n10089));
  INVx1_ASAP7_75t_L         g09833(.A(new_n10089), .Y(new_n10090));
  NAND3xp33_ASAP7_75t_L     g09834(.A(new_n10090), .B(new_n9815), .C(\a[56] ), .Y(new_n10091));
  O2A1O1Ixp33_ASAP7_75t_L   g09835(.A1(new_n10088), .A2(new_n274), .B(new_n10087), .C(new_n10083), .Y(new_n10092));
  NAND2xp33_ASAP7_75t_L     g09836(.A(new_n10083), .B(new_n10089), .Y(new_n10093));
  A2O1A1Ixp33_ASAP7_75t_L   g09837(.A1(new_n9805), .A2(new_n10092), .B(new_n10083), .C(new_n10093), .Y(new_n10094));
  NAND2xp33_ASAP7_75t_L     g09838(.A(new_n10091), .B(new_n10094), .Y(new_n10095));
  NAND2xp33_ASAP7_75t_L     g09839(.A(new_n10077), .B(new_n10095), .Y(new_n10096));
  INVx1_ASAP7_75t_L         g09840(.A(new_n10076), .Y(new_n10097));
  A2O1A1Ixp33_ASAP7_75t_L   g09841(.A1(new_n342), .A2(new_n9437), .B(new_n10074), .C(new_n9099), .Y(new_n10098));
  NAND2xp33_ASAP7_75t_L     g09842(.A(new_n10098), .B(new_n10097), .Y(new_n10099));
  NAND3xp33_ASAP7_75t_L     g09843(.A(new_n10099), .B(new_n10091), .C(new_n10094), .Y(new_n10100));
  NAND3xp33_ASAP7_75t_L     g09844(.A(new_n10096), .B(new_n10072), .C(new_n10100), .Y(new_n10101));
  MAJIxp5_ASAP7_75t_L       g09845(.A(new_n9818), .B(new_n9449), .C(new_n9805), .Y(new_n10102));
  AOI21xp33_ASAP7_75t_L     g09846(.A1(new_n10094), .A2(new_n10091), .B(new_n10099), .Y(new_n10103));
  NOR2xp33_ASAP7_75t_L      g09847(.A(new_n10077), .B(new_n10095), .Y(new_n10104));
  OAI21xp33_ASAP7_75t_L     g09848(.A1(new_n10103), .A2(new_n10104), .B(new_n10102), .Y(new_n10105));
  AO21x2_ASAP7_75t_L        g09849(.A1(new_n10101), .A2(new_n10105), .B(new_n10071), .Y(new_n10106));
  NAND3xp33_ASAP7_75t_L     g09850(.A(new_n10105), .B(new_n10101), .C(new_n10071), .Y(new_n10107));
  NAND3xp33_ASAP7_75t_L     g09851(.A(new_n10063), .B(new_n10106), .C(new_n10107), .Y(new_n10108));
  AOI21xp33_ASAP7_75t_L     g09852(.A1(new_n10105), .A2(new_n10101), .B(new_n10071), .Y(new_n10109));
  AND3x1_ASAP7_75t_L        g09853(.A(new_n10105), .B(new_n10101), .C(new_n10071), .Y(new_n10110));
  OAI211xp5_ASAP7_75t_L     g09854(.A1(new_n10109), .A2(new_n10110), .B(new_n9831), .C(new_n10061), .Y(new_n10111));
  AO21x2_ASAP7_75t_L        g09855(.A1(new_n10108), .A2(new_n10111), .B(new_n10060), .Y(new_n10112));
  NAND3xp33_ASAP7_75t_L     g09856(.A(new_n10111), .B(new_n10108), .C(new_n10060), .Y(new_n10113));
  NAND2xp33_ASAP7_75t_L     g09857(.A(new_n10113), .B(new_n10112), .Y(new_n10114));
  O2A1O1Ixp33_ASAP7_75t_L   g09858(.A1(new_n9799), .A2(new_n9850), .B(new_n9841), .C(new_n10114), .Y(new_n10115));
  MAJIxp5_ASAP7_75t_L       g09859(.A(new_n9836), .B(new_n9799), .C(new_n9850), .Y(new_n10116));
  AOI21xp33_ASAP7_75t_L     g09860(.A1(new_n10113), .A2(new_n10112), .B(new_n10116), .Y(new_n10117));
  OAI21xp33_ASAP7_75t_L     g09861(.A1(new_n10117), .A2(new_n10115), .B(new_n10057), .Y(new_n10118));
  AND2x2_ASAP7_75t_L        g09862(.A(\a[44] ), .B(new_n10056), .Y(new_n10119));
  NOR2xp33_ASAP7_75t_L      g09863(.A(\a[44] ), .B(new_n10056), .Y(new_n10120));
  NAND3xp33_ASAP7_75t_L     g09864(.A(new_n10116), .B(new_n10112), .C(new_n10113), .Y(new_n10121));
  MAJx2_ASAP7_75t_L         g09865(.A(new_n9836), .B(new_n9799), .C(new_n9850), .Y(new_n10122));
  NAND2xp33_ASAP7_75t_L     g09866(.A(new_n10114), .B(new_n10122), .Y(new_n10123));
  OAI211xp5_ASAP7_75t_L     g09867(.A1(new_n10119), .A2(new_n10120), .B(new_n10123), .C(new_n10121), .Y(new_n10124));
  NAND3xp33_ASAP7_75t_L     g09868(.A(new_n10054), .B(new_n10118), .C(new_n10124), .Y(new_n10125));
  INVx1_ASAP7_75t_L         g09869(.A(new_n10053), .Y(new_n10126));
  O2A1O1Ixp33_ASAP7_75t_L   g09870(.A1(new_n9845), .A2(new_n9793), .B(new_n9787), .C(new_n10126), .Y(new_n10127));
  NAND2xp33_ASAP7_75t_L     g09871(.A(new_n10118), .B(new_n10124), .Y(new_n10128));
  NAND2xp33_ASAP7_75t_L     g09872(.A(new_n10127), .B(new_n10128), .Y(new_n10129));
  OAI22xp33_ASAP7_75t_L     g09873(.A1(new_n5640), .A2(new_n1043), .B1(new_n960), .B2(new_n5925), .Y(new_n10130));
  AOI221xp5_ASAP7_75t_L     g09874(.A1(new_n5629), .A2(\b[16] ), .B1(new_n5637), .B2(new_n1156), .C(new_n10130), .Y(new_n10131));
  XNOR2x2_ASAP7_75t_L       g09875(.A(new_n5626), .B(new_n10131), .Y(new_n10132));
  NAND3xp33_ASAP7_75t_L     g09876(.A(new_n10129), .B(new_n10125), .C(new_n10132), .Y(new_n10133));
  AO21x2_ASAP7_75t_L        g09877(.A1(new_n10125), .A2(new_n10129), .B(new_n10132), .Y(new_n10134));
  O2A1O1Ixp33_ASAP7_75t_L   g09878(.A1(new_n9792), .A2(new_n10126), .B(new_n9843), .C(new_n10051), .Y(new_n10135));
  A2O1A1Ixp33_ASAP7_75t_L   g09879(.A1(new_n9846), .A2(new_n9840), .B(new_n10135), .C(new_n9786), .Y(new_n10136));
  A2O1A1O1Ixp25_ASAP7_75t_L g09880(.A1(new_n9498), .A2(new_n9501), .B(new_n9491), .C(new_n10136), .D(new_n9847), .Y(new_n10137));
  NAND3xp33_ASAP7_75t_L     g09881(.A(new_n10137), .B(new_n10134), .C(new_n10133), .Y(new_n10138));
  INVx1_ASAP7_75t_L         g09882(.A(new_n10138), .Y(new_n10139));
  AO21x2_ASAP7_75t_L        g09883(.A1(new_n10133), .A2(new_n10134), .B(new_n10137), .Y(new_n10140));
  INVx1_ASAP7_75t_L         g09884(.A(new_n10140), .Y(new_n10141));
  OAI22xp33_ASAP7_75t_L     g09885(.A1(new_n5144), .A2(new_n1349), .B1(new_n1458), .B2(new_n4903), .Y(new_n10142));
  AOI221xp5_ASAP7_75t_L     g09886(.A1(new_n4917), .A2(\b[19] ), .B1(new_n4912), .B2(new_n1607), .C(new_n10142), .Y(new_n10143));
  XNOR2x2_ASAP7_75t_L       g09887(.A(new_n4906), .B(new_n10143), .Y(new_n10144));
  OAI21xp33_ASAP7_75t_L     g09888(.A1(new_n10139), .A2(new_n10141), .B(new_n10144), .Y(new_n10145));
  INVx1_ASAP7_75t_L         g09889(.A(new_n9780), .Y(new_n10146));
  NAND3xp33_ASAP7_75t_L     g09890(.A(new_n10146), .B(new_n9859), .C(new_n9862), .Y(new_n10147));
  A2O1A1Ixp33_ASAP7_75t_L   g09891(.A1(new_n9864), .A2(new_n9780), .B(new_n9867), .C(new_n10147), .Y(new_n10148));
  NOR3xp33_ASAP7_75t_L      g09892(.A(new_n10141), .B(new_n10144), .C(new_n10139), .Y(new_n10149));
  XNOR2x2_ASAP7_75t_L       g09893(.A(\a[38] ), .B(new_n10143), .Y(new_n10150));
  AOI21xp33_ASAP7_75t_L     g09894(.A1(new_n10140), .A2(new_n10138), .B(new_n10150), .Y(new_n10151));
  OA21x2_ASAP7_75t_L        g09895(.A1(new_n10149), .A2(new_n10151), .B(new_n10148), .Y(new_n10152));
  INVx1_ASAP7_75t_L         g09896(.A(new_n9523), .Y(new_n10153));
  NOR2xp33_ASAP7_75t_L      g09897(.A(new_n9513), .B(new_n9512), .Y(new_n10154));
  A2O1A1Ixp33_ASAP7_75t_L   g09898(.A1(new_n9417), .A2(new_n9183), .B(new_n10154), .C(new_n10153), .Y(new_n10155));
  INVx1_ASAP7_75t_L         g09899(.A(new_n10147), .Y(new_n10156));
  A2O1A1O1Ixp25_ASAP7_75t_L g09900(.A1(new_n9865), .A2(new_n10155), .B(new_n10156), .C(new_n10145), .D(new_n10149), .Y(new_n10157));
  OAI22xp33_ASAP7_75t_L     g09901(.A1(new_n4397), .A2(new_n1745), .B1(new_n1895), .B2(new_n4142), .Y(new_n10158));
  AOI221xp5_ASAP7_75t_L     g09902(.A1(new_n4156), .A2(\b[22] ), .B1(new_n4151), .B2(new_n2056), .C(new_n10158), .Y(new_n10159));
  XNOR2x2_ASAP7_75t_L       g09903(.A(new_n4145), .B(new_n10159), .Y(new_n10160));
  A2O1A1Ixp33_ASAP7_75t_L   g09904(.A1(new_n10157), .A2(new_n10145), .B(new_n10152), .C(new_n10160), .Y(new_n10161));
  A2O1A1O1Ixp25_ASAP7_75t_L g09905(.A1(new_n9864), .A2(new_n9780), .B(new_n9867), .C(new_n10147), .D(new_n10151), .Y(new_n10162));
  OAI21xp33_ASAP7_75t_L     g09906(.A1(new_n10149), .A2(new_n10151), .B(new_n10148), .Y(new_n10163));
  XNOR2x2_ASAP7_75t_L       g09907(.A(\a[35] ), .B(new_n10159), .Y(new_n10164));
  OAI311xp33_ASAP7_75t_L    g09908(.A1(new_n10149), .A2(new_n10162), .A3(new_n10151), .B1(new_n10163), .C1(new_n10164), .Y(new_n10165));
  NAND2xp33_ASAP7_75t_L     g09909(.A(new_n9532), .B(new_n9531), .Y(new_n10166));
  A2O1A1O1Ixp25_ASAP7_75t_L g09910(.A1(new_n9875), .A2(new_n10166), .B(new_n9767), .C(new_n9873), .D(new_n9877), .Y(new_n10167));
  NAND3xp33_ASAP7_75t_L     g09911(.A(new_n10167), .B(new_n10161), .C(new_n10165), .Y(new_n10168));
  AO21x2_ASAP7_75t_L        g09912(.A1(new_n10165), .A2(new_n10161), .B(new_n10167), .Y(new_n10169));
  NAND3xp33_ASAP7_75t_L     g09913(.A(new_n10169), .B(new_n10049), .C(new_n10168), .Y(new_n10170));
  AND3x1_ASAP7_75t_L        g09914(.A(new_n10167), .B(new_n10161), .C(new_n10165), .Y(new_n10171));
  AOI21xp33_ASAP7_75t_L     g09915(.A1(new_n10161), .A2(new_n10165), .B(new_n10167), .Y(new_n10172));
  NOR3xp33_ASAP7_75t_L      g09916(.A(new_n10171), .B(new_n10049), .C(new_n10172), .Y(new_n10173));
  AOI21xp33_ASAP7_75t_L     g09917(.A1(new_n10170), .A2(new_n10049), .B(new_n10173), .Y(new_n10174));
  INVx1_ASAP7_75t_L         g09918(.A(new_n9881), .Y(new_n10175));
  A2O1A1O1Ixp25_ASAP7_75t_L g09919(.A1(new_n9555), .A2(new_n9888), .B(new_n9761), .C(new_n9885), .D(new_n10175), .Y(new_n10176));
  NAND2xp33_ASAP7_75t_L     g09920(.A(new_n10174), .B(new_n10176), .Y(new_n10177));
  XNOR2x2_ASAP7_75t_L       g09921(.A(new_n3493), .B(new_n10048), .Y(new_n10178));
  NAND3xp33_ASAP7_75t_L     g09922(.A(new_n10169), .B(new_n10178), .C(new_n10168), .Y(new_n10179));
  OAI21xp33_ASAP7_75t_L     g09923(.A1(new_n10172), .A2(new_n10171), .B(new_n10049), .Y(new_n10180));
  NAND2xp33_ASAP7_75t_L     g09924(.A(new_n10179), .B(new_n10180), .Y(new_n10181));
  A2O1A1Ixp33_ASAP7_75t_L   g09925(.A1(new_n9894), .A2(new_n9893), .B(new_n10175), .C(new_n10181), .Y(new_n10182));
  NOR2xp33_ASAP7_75t_L      g09926(.A(new_n3079), .B(new_n2930), .Y(new_n10183));
  AOI221xp5_ASAP7_75t_L     g09927(.A1(\b[26] ), .A2(new_n3129), .B1(\b[27] ), .B2(new_n2936), .C(new_n10183), .Y(new_n10184));
  O2A1O1Ixp33_ASAP7_75t_L   g09928(.A1(new_n2940), .A2(new_n3087), .B(new_n10184), .C(new_n2928), .Y(new_n10185));
  OAI21xp33_ASAP7_75t_L     g09929(.A1(new_n2940), .A2(new_n3087), .B(new_n10184), .Y(new_n10186));
  NAND2xp33_ASAP7_75t_L     g09930(.A(new_n2928), .B(new_n10186), .Y(new_n10187));
  OA21x2_ASAP7_75t_L        g09931(.A1(new_n2928), .A2(new_n10185), .B(new_n10187), .Y(new_n10188));
  NAND3xp33_ASAP7_75t_L     g09932(.A(new_n10177), .B(new_n10182), .C(new_n10188), .Y(new_n10189));
  AO21x2_ASAP7_75t_L        g09933(.A1(new_n10182), .A2(new_n10177), .B(new_n10188), .Y(new_n10190));
  A2O1A1O1Ixp25_ASAP7_75t_L g09934(.A1(new_n9552), .A2(new_n9408), .B(new_n9752), .C(new_n9900), .D(new_n9890), .Y(new_n10191));
  NAND3xp33_ASAP7_75t_L     g09935(.A(new_n10191), .B(new_n10190), .C(new_n10189), .Y(new_n10192));
  AO21x2_ASAP7_75t_L        g09936(.A1(new_n10189), .A2(new_n10190), .B(new_n10191), .Y(new_n10193));
  NOR2xp33_ASAP7_75t_L      g09937(.A(new_n3456), .B(new_n2410), .Y(new_n10194));
  AOI221xp5_ASAP7_75t_L     g09938(.A1(\b[29] ), .A2(new_n2577), .B1(\b[31] ), .B2(new_n2423), .C(new_n10194), .Y(new_n10195));
  O2A1O1Ixp33_ASAP7_75t_L   g09939(.A1(new_n2425), .A2(new_n3681), .B(new_n10195), .C(new_n2413), .Y(new_n10196));
  INVx1_ASAP7_75t_L         g09940(.A(new_n10196), .Y(new_n10197));
  O2A1O1Ixp33_ASAP7_75t_L   g09941(.A1(new_n2425), .A2(new_n3681), .B(new_n10195), .C(\a[26] ), .Y(new_n10198));
  AOI21xp33_ASAP7_75t_L     g09942(.A1(new_n10197), .A2(\a[26] ), .B(new_n10198), .Y(new_n10199));
  NAND3xp33_ASAP7_75t_L     g09943(.A(new_n10193), .B(new_n10192), .C(new_n10199), .Y(new_n10200));
  AND3x1_ASAP7_75t_L        g09944(.A(new_n10191), .B(new_n10190), .C(new_n10189), .Y(new_n10201));
  AOI21xp33_ASAP7_75t_L     g09945(.A1(new_n10190), .A2(new_n10189), .B(new_n10191), .Y(new_n10202));
  INVx1_ASAP7_75t_L         g09946(.A(new_n10198), .Y(new_n10203));
  OAI21xp33_ASAP7_75t_L     g09947(.A1(new_n2413), .A2(new_n10196), .B(new_n10203), .Y(new_n10204));
  OAI21xp33_ASAP7_75t_L     g09948(.A1(new_n10202), .A2(new_n10201), .B(new_n10204), .Y(new_n10205));
  A2O1A1O1Ixp25_ASAP7_75t_L g09949(.A1(new_n9573), .A2(new_n9572), .B(new_n9570), .C(new_n9911), .D(new_n9902), .Y(new_n10206));
  NAND3xp33_ASAP7_75t_L     g09950(.A(new_n10206), .B(new_n10205), .C(new_n10200), .Y(new_n10207));
  NOR3xp33_ASAP7_75t_L      g09951(.A(new_n10201), .B(new_n10202), .C(new_n10204), .Y(new_n10208));
  AOI21xp33_ASAP7_75t_L     g09952(.A1(new_n10193), .A2(new_n10192), .B(new_n10199), .Y(new_n10209));
  OAI21xp33_ASAP7_75t_L     g09953(.A1(new_n9908), .A2(new_n9747), .B(new_n9910), .Y(new_n10210));
  OAI21xp33_ASAP7_75t_L     g09954(.A1(new_n10208), .A2(new_n10209), .B(new_n10210), .Y(new_n10211));
  NOR2xp33_ASAP7_75t_L      g09955(.A(new_n4101), .B(new_n1962), .Y(new_n10212));
  AOI221xp5_ASAP7_75t_L     g09956(.A1(new_n1955), .A2(\b[34] ), .B1(new_n2093), .B2(\b[32] ), .C(new_n10212), .Y(new_n10213));
  O2A1O1Ixp33_ASAP7_75t_L   g09957(.A1(new_n1956), .A2(new_n4352), .B(new_n10213), .C(new_n1952), .Y(new_n10214));
  O2A1O1Ixp33_ASAP7_75t_L   g09958(.A1(new_n1956), .A2(new_n4352), .B(new_n10213), .C(\a[23] ), .Y(new_n10215));
  INVx1_ASAP7_75t_L         g09959(.A(new_n10215), .Y(new_n10216));
  OA21x2_ASAP7_75t_L        g09960(.A1(new_n1952), .A2(new_n10214), .B(new_n10216), .Y(new_n10217));
  NAND3xp33_ASAP7_75t_L     g09961(.A(new_n10207), .B(new_n10211), .C(new_n10217), .Y(new_n10218));
  NOR3xp33_ASAP7_75t_L      g09962(.A(new_n10210), .B(new_n10209), .C(new_n10208), .Y(new_n10219));
  AOI21xp33_ASAP7_75t_L     g09963(.A1(new_n10205), .A2(new_n10200), .B(new_n10206), .Y(new_n10220));
  NOR2xp33_ASAP7_75t_L      g09964(.A(new_n1952), .B(new_n10214), .Y(new_n10221));
  OAI22xp33_ASAP7_75t_L     g09965(.A1(new_n10220), .A2(new_n10219), .B1(new_n10215), .B2(new_n10221), .Y(new_n10222));
  NAND2xp33_ASAP7_75t_L     g09966(.A(new_n9922), .B(new_n9921), .Y(new_n10223));
  O2A1O1Ixp33_ASAP7_75t_L   g09967(.A1(new_n9915), .A2(new_n1952), .B(new_n9917), .C(new_n10223), .Y(new_n10224));
  AOI21xp33_ASAP7_75t_L     g09968(.A1(new_n9746), .A2(new_n9934), .B(new_n10224), .Y(new_n10225));
  NAND3xp33_ASAP7_75t_L     g09969(.A(new_n10225), .B(new_n10222), .C(new_n10218), .Y(new_n10226));
  NAND2xp33_ASAP7_75t_L     g09970(.A(new_n10218), .B(new_n10222), .Y(new_n10227));
  A2O1A1Ixp33_ASAP7_75t_L   g09971(.A1(new_n9934), .A2(new_n9746), .B(new_n10224), .C(new_n10227), .Y(new_n10228));
  INVx1_ASAP7_75t_L         g09972(.A(new_n5083), .Y(new_n10229));
  OAI22xp33_ASAP7_75t_L     g09973(.A1(new_n1654), .A2(new_n4581), .B1(new_n4613), .B2(new_n1517), .Y(new_n10230));
  AOI221xp5_ASAP7_75t_L     g09974(.A1(new_n1511), .A2(\b[37] ), .B1(new_n1513), .B2(new_n10229), .C(new_n10230), .Y(new_n10231));
  XNOR2x2_ASAP7_75t_L       g09975(.A(new_n1501), .B(new_n10231), .Y(new_n10232));
  NAND3xp33_ASAP7_75t_L     g09976(.A(new_n10226), .B(new_n10228), .C(new_n10232), .Y(new_n10233));
  AO21x2_ASAP7_75t_L        g09977(.A1(new_n10228), .A2(new_n10226), .B(new_n10232), .Y(new_n10234));
  A2O1A1O1Ixp25_ASAP7_75t_L g09978(.A1(new_n9601), .A2(new_n9602), .B(new_n9946), .C(new_n9957), .D(new_n9939), .Y(new_n10235));
  NAND3xp33_ASAP7_75t_L     g09979(.A(new_n10235), .B(new_n10234), .C(new_n10233), .Y(new_n10236));
  AO21x2_ASAP7_75t_L        g09980(.A1(new_n10233), .A2(new_n10234), .B(new_n10235), .Y(new_n10237));
  NOR2xp33_ASAP7_75t_L      g09981(.A(new_n5570), .B(new_n2118), .Y(new_n10238));
  AOI221xp5_ASAP7_75t_L     g09982(.A1(\b[38] ), .A2(new_n1290), .B1(\b[40] ), .B2(new_n1209), .C(new_n10238), .Y(new_n10239));
  O2A1O1Ixp33_ASAP7_75t_L   g09983(.A1(new_n1210), .A2(new_n5862), .B(new_n10239), .C(new_n1206), .Y(new_n10240));
  INVx1_ASAP7_75t_L         g09984(.A(new_n10239), .Y(new_n10241));
  A2O1A1Ixp33_ASAP7_75t_L   g09985(.A1(new_n6651), .A2(new_n1216), .B(new_n10241), .C(new_n1206), .Y(new_n10242));
  OAI21xp33_ASAP7_75t_L     g09986(.A1(new_n1206), .A2(new_n10240), .B(new_n10242), .Y(new_n10243));
  INVx1_ASAP7_75t_L         g09987(.A(new_n10243), .Y(new_n10244));
  NAND3xp33_ASAP7_75t_L     g09988(.A(new_n10237), .B(new_n10236), .C(new_n10244), .Y(new_n10245));
  AND3x1_ASAP7_75t_L        g09989(.A(new_n10235), .B(new_n10234), .C(new_n10233), .Y(new_n10246));
  AOI21xp33_ASAP7_75t_L     g09990(.A1(new_n10234), .A2(new_n10233), .B(new_n10235), .Y(new_n10247));
  OAI21xp33_ASAP7_75t_L     g09991(.A1(new_n10247), .A2(new_n10246), .B(new_n10243), .Y(new_n10248));
  NAND2xp33_ASAP7_75t_L     g09992(.A(new_n10245), .B(new_n10248), .Y(new_n10249));
  NOR2xp33_ASAP7_75t_L      g09993(.A(new_n9958), .B(new_n9960), .Y(new_n10250));
  A2O1A1Ixp33_ASAP7_75t_L   g09994(.A1(\a[17] ), .A2(new_n9952), .B(new_n9953), .C(new_n10250), .Y(new_n10251));
  A2O1A1Ixp33_ASAP7_75t_L   g09995(.A1(new_n9955), .A2(new_n9962), .B(new_n9964), .C(new_n10251), .Y(new_n10252));
  NOR2xp33_ASAP7_75t_L      g09996(.A(new_n10249), .B(new_n10252), .Y(new_n10253));
  INVx1_ASAP7_75t_L         g09997(.A(new_n10250), .Y(new_n10254));
  NAND3xp33_ASAP7_75t_L     g09998(.A(new_n10237), .B(new_n10236), .C(new_n10243), .Y(new_n10255));
  NOR3xp33_ASAP7_75t_L      g09999(.A(new_n10246), .B(new_n10247), .C(new_n10243), .Y(new_n10256));
  AOI21xp33_ASAP7_75t_L     g10000(.A1(new_n10255), .A2(new_n10243), .B(new_n10256), .Y(new_n10257));
  O2A1O1Ixp33_ASAP7_75t_L   g10001(.A1(new_n10254), .A2(new_n9954), .B(new_n9970), .C(new_n10257), .Y(new_n10258));
  OAI22xp33_ASAP7_75t_L     g10002(.A1(new_n980), .A2(new_n6110), .B1(new_n6378), .B2(new_n864), .Y(new_n10259));
  AOI221xp5_ASAP7_75t_L     g10003(.A1(new_n886), .A2(\b[43] ), .B1(new_n873), .B2(new_n6682), .C(new_n10259), .Y(new_n10260));
  XNOR2x2_ASAP7_75t_L       g10004(.A(new_n867), .B(new_n10260), .Y(new_n10261));
  NOR3xp33_ASAP7_75t_L      g10005(.A(new_n10258), .B(new_n10261), .C(new_n10253), .Y(new_n10262));
  OAI21xp33_ASAP7_75t_L     g10006(.A1(new_n10253), .A2(new_n10258), .B(new_n10261), .Y(new_n10263));
  INVx1_ASAP7_75t_L         g10007(.A(new_n10263), .Y(new_n10264));
  OAI21xp33_ASAP7_75t_L     g10008(.A1(new_n10262), .A2(new_n10264), .B(new_n10046), .Y(new_n10265));
  A2O1A1O1Ixp25_ASAP7_75t_L g10009(.A1(new_n9642), .A2(new_n9988), .B(new_n9987), .C(new_n9983), .D(new_n9978), .Y(new_n10266));
  INVx1_ASAP7_75t_L         g10010(.A(new_n10262), .Y(new_n10267));
  NAND3xp33_ASAP7_75t_L     g10011(.A(new_n10267), .B(new_n10266), .C(new_n10263), .Y(new_n10268));
  OAI22xp33_ASAP7_75t_L     g10012(.A1(new_n1550), .A2(new_n7249), .B1(new_n6944), .B2(new_n712), .Y(new_n10269));
  AOI221xp5_ASAP7_75t_L     g10013(.A1(new_n640), .A2(\b[46] ), .B1(new_n718), .B2(new_n7278), .C(new_n10269), .Y(new_n10270));
  XNOR2x2_ASAP7_75t_L       g10014(.A(new_n637), .B(new_n10270), .Y(new_n10271));
  NAND3xp33_ASAP7_75t_L     g10015(.A(new_n10265), .B(new_n10268), .C(new_n10271), .Y(new_n10272));
  AOI21xp33_ASAP7_75t_L     g10016(.A1(new_n10267), .A2(new_n10263), .B(new_n10266), .Y(new_n10273));
  A2O1A1O1Ixp25_ASAP7_75t_L g10017(.A1(new_n9983), .A2(new_n9741), .B(new_n9978), .C(new_n10263), .D(new_n10262), .Y(new_n10274));
  INVx1_ASAP7_75t_L         g10018(.A(new_n10271), .Y(new_n10275));
  A2O1A1Ixp33_ASAP7_75t_L   g10019(.A1(new_n10274), .A2(new_n10263), .B(new_n10273), .C(new_n10275), .Y(new_n10276));
  NAND3xp33_ASAP7_75t_L     g10020(.A(new_n10045), .B(new_n10272), .C(new_n10276), .Y(new_n10277));
  NOR2xp33_ASAP7_75t_L      g10021(.A(new_n9989), .B(new_n9986), .Y(new_n10278));
  MAJIxp5_ASAP7_75t_L       g10022(.A(new_n9732), .B(new_n9738), .C(new_n10278), .Y(new_n10279));
  AOI211xp5_ASAP7_75t_L     g10023(.A1(new_n10274), .A2(new_n10263), .B(new_n10275), .C(new_n10273), .Y(new_n10280));
  AOI21xp33_ASAP7_75t_L     g10024(.A1(new_n10265), .A2(new_n10268), .B(new_n10271), .Y(new_n10281));
  OAI21xp33_ASAP7_75t_L     g10025(.A1(new_n10281), .A2(new_n10280), .B(new_n10279), .Y(new_n10282));
  AOI21xp33_ASAP7_75t_L     g10026(.A1(new_n10277), .A2(new_n10282), .B(new_n10043), .Y(new_n10283));
  NOR3xp33_ASAP7_75t_L      g10027(.A(new_n10279), .B(new_n10280), .C(new_n10281), .Y(new_n10284));
  O2A1O1Ixp33_ASAP7_75t_L   g10028(.A1(new_n637), .A2(new_n9735), .B(new_n9737), .C(new_n10044), .Y(new_n10285));
  NAND2xp33_ASAP7_75t_L     g10029(.A(new_n9993), .B(new_n9992), .Y(new_n10286));
  AOI221xp5_ASAP7_75t_L     g10030(.A1(new_n9732), .A2(new_n10286), .B1(new_n10272), .B2(new_n10276), .C(new_n10285), .Y(new_n10287));
  NOR3xp33_ASAP7_75t_L      g10031(.A(new_n10284), .B(new_n10287), .C(new_n10042), .Y(new_n10288));
  NOR2xp33_ASAP7_75t_L      g10032(.A(new_n10288), .B(new_n10283), .Y(new_n10289));
  OAI21xp33_ASAP7_75t_L     g10033(.A1(new_n10039), .A2(new_n10021), .B(new_n10289), .Y(new_n10290));
  OAI221xp5_ASAP7_75t_L     g10034(.A1(new_n10002), .A2(new_n10000), .B1(new_n10283), .B2(new_n10288), .C(new_n9995), .Y(new_n10291));
  OAI22xp33_ASAP7_75t_L     g10035(.A1(new_n350), .A2(new_n8779), .B1(new_n8755), .B2(new_n375), .Y(new_n10292));
  AOI221xp5_ASAP7_75t_L     g10036(.A1(new_n361), .A2(\b[52] ), .B1(new_n359), .B2(new_n9367), .C(new_n10292), .Y(new_n10293));
  XNOR2x2_ASAP7_75t_L       g10037(.A(new_n346), .B(new_n10293), .Y(new_n10294));
  NAND3xp33_ASAP7_75t_L     g10038(.A(new_n10290), .B(new_n10291), .C(new_n10294), .Y(new_n10295));
  A2O1A1O1Ixp25_ASAP7_75t_L g10039(.A1(new_n9666), .A2(new_n10004), .B(new_n10001), .C(new_n10008), .D(new_n10039), .Y(new_n10296));
  OAI21xp33_ASAP7_75t_L     g10040(.A1(new_n10287), .A2(new_n10284), .B(new_n10042), .Y(new_n10297));
  NAND3xp33_ASAP7_75t_L     g10041(.A(new_n10277), .B(new_n10043), .C(new_n10282), .Y(new_n10298));
  NAND2xp33_ASAP7_75t_L     g10042(.A(new_n10297), .B(new_n10298), .Y(new_n10299));
  NOR2xp33_ASAP7_75t_L      g10043(.A(new_n10299), .B(new_n10296), .Y(new_n10300));
  AOI221xp5_ASAP7_75t_L     g10044(.A1(new_n10019), .A2(new_n10008), .B1(new_n10297), .B2(new_n10298), .C(new_n10039), .Y(new_n10301));
  INVx1_ASAP7_75t_L         g10045(.A(new_n10294), .Y(new_n10302));
  OAI21xp33_ASAP7_75t_L     g10046(.A1(new_n10301), .A2(new_n10300), .B(new_n10302), .Y(new_n10303));
  NAND3xp33_ASAP7_75t_L     g10047(.A(new_n10038), .B(new_n10295), .C(new_n10303), .Y(new_n10304));
  A2O1A1O1Ixp25_ASAP7_75t_L g10048(.A1(new_n9386), .A2(new_n9675), .B(new_n9677), .C(new_n10024), .D(new_n10022), .Y(new_n10305));
  NOR3xp33_ASAP7_75t_L      g10049(.A(new_n10300), .B(new_n10301), .C(new_n10302), .Y(new_n10306));
  AOI21xp33_ASAP7_75t_L     g10050(.A1(new_n10290), .A2(new_n10291), .B(new_n10294), .Y(new_n10307));
  OAI21xp33_ASAP7_75t_L     g10051(.A1(new_n10306), .A2(new_n10307), .B(new_n10305), .Y(new_n10308));
  INVx1_ASAP7_75t_L         g10052(.A(\b[55] ), .Y(new_n10309));
  NAND2xp33_ASAP7_75t_L     g10053(.A(\b[53] ), .B(new_n286), .Y(new_n10310));
  OAI221xp5_ASAP7_75t_L     g10054(.A1(new_n285), .A2(new_n9709), .B1(new_n10309), .B2(new_n269), .C(new_n10310), .Y(new_n10311));
  NOR2xp33_ASAP7_75t_L      g10055(.A(\b[54] ), .B(\b[55] ), .Y(new_n10312));
  NOR2xp33_ASAP7_75t_L      g10056(.A(new_n9709), .B(new_n10309), .Y(new_n10313));
  NOR2xp33_ASAP7_75t_L      g10057(.A(new_n10312), .B(new_n10313), .Y(new_n10314));
  A2O1A1Ixp33_ASAP7_75t_L   g10058(.A1(new_n9715), .A2(new_n9711), .B(new_n9710), .C(new_n10314), .Y(new_n10315));
  INVx1_ASAP7_75t_L         g10059(.A(new_n10315), .Y(new_n10316));
  INVx1_ASAP7_75t_L         g10060(.A(new_n9710), .Y(new_n10317));
  A2O1A1Ixp33_ASAP7_75t_L   g10061(.A1(new_n9686), .A2(new_n9714), .B(new_n9708), .C(new_n10317), .Y(new_n10318));
  NOR2xp33_ASAP7_75t_L      g10062(.A(new_n10314), .B(new_n10318), .Y(new_n10319));
  NOR2xp33_ASAP7_75t_L      g10063(.A(new_n10316), .B(new_n10319), .Y(new_n10320));
  A2O1A1Ixp33_ASAP7_75t_L   g10064(.A1(new_n10320), .A2(new_n273), .B(new_n10311), .C(\a[2] ), .Y(new_n10321));
  AOI211xp5_ASAP7_75t_L     g10065(.A1(new_n10320), .A2(new_n273), .B(new_n10311), .C(new_n257), .Y(new_n10322));
  A2O1A1O1Ixp25_ASAP7_75t_L g10066(.A1(new_n273), .A2(new_n10320), .B(new_n10311), .C(new_n10321), .D(new_n10322), .Y(new_n10323));
  AOI21xp33_ASAP7_75t_L     g10067(.A1(new_n10304), .A2(new_n10308), .B(new_n10323), .Y(new_n10324));
  INVx1_ASAP7_75t_L         g10068(.A(new_n10324), .Y(new_n10325));
  NAND3xp33_ASAP7_75t_L     g10069(.A(new_n10304), .B(new_n10308), .C(new_n10323), .Y(new_n10326));
  NAND2xp33_ASAP7_75t_L     g10070(.A(new_n10326), .B(new_n10325), .Y(new_n10327));
  XOR2x2_ASAP7_75t_L        g10071(.A(new_n10036), .B(new_n10327), .Y(\f[55] ));
  NOR2xp33_ASAP7_75t_L      g10072(.A(new_n9709), .B(new_n287), .Y(new_n10329));
  AOI221xp5_ASAP7_75t_L     g10073(.A1(\b[55] ), .A2(new_n264), .B1(\b[56] ), .B2(new_n283), .C(new_n10329), .Y(new_n10330));
  NOR2xp33_ASAP7_75t_L      g10074(.A(\b[55] ), .B(\b[56] ), .Y(new_n10331));
  INVx1_ASAP7_75t_L         g10075(.A(\b[56] ), .Y(new_n10332));
  NOR2xp33_ASAP7_75t_L      g10076(.A(new_n10309), .B(new_n10332), .Y(new_n10333));
  NOR2xp33_ASAP7_75t_L      g10077(.A(new_n10331), .B(new_n10333), .Y(new_n10334));
  A2O1A1Ixp33_ASAP7_75t_L   g10078(.A1(new_n10318), .A2(new_n10314), .B(new_n10313), .C(new_n10334), .Y(new_n10335));
  A2O1A1O1Ixp25_ASAP7_75t_L g10079(.A1(new_n9711), .A2(new_n9715), .B(new_n9710), .C(new_n10314), .D(new_n10313), .Y(new_n10336));
  INVx1_ASAP7_75t_L         g10080(.A(new_n10334), .Y(new_n10337));
  NAND2xp33_ASAP7_75t_L     g10081(.A(new_n10337), .B(new_n10336), .Y(new_n10338));
  NAND2xp33_ASAP7_75t_L     g10082(.A(new_n10338), .B(new_n10335), .Y(new_n10339));
  O2A1O1Ixp33_ASAP7_75t_L   g10083(.A1(new_n279), .A2(new_n10339), .B(new_n10330), .C(new_n257), .Y(new_n10340));
  OAI21xp33_ASAP7_75t_L     g10084(.A1(new_n279), .A2(new_n10339), .B(new_n10330), .Y(new_n10341));
  NAND2xp33_ASAP7_75t_L     g10085(.A(new_n257), .B(new_n10341), .Y(new_n10342));
  OAI21xp33_ASAP7_75t_L     g10086(.A1(new_n257), .A2(new_n10340), .B(new_n10342), .Y(new_n10343));
  INVx1_ASAP7_75t_L         g10087(.A(new_n10343), .Y(new_n10344));
  NAND2xp33_ASAP7_75t_L     g10088(.A(new_n10291), .B(new_n10290), .Y(new_n10345));
  MAJIxp5_ASAP7_75t_L       g10089(.A(new_n10305), .B(new_n10294), .C(new_n10345), .Y(new_n10346));
  A2O1A1O1Ixp25_ASAP7_75t_L g10090(.A1(new_n10008), .A2(new_n10019), .B(new_n10039), .C(new_n10297), .D(new_n10288), .Y(new_n10347));
  OAI22xp33_ASAP7_75t_L     g10091(.A1(new_n513), .A2(new_n8427), .B1(new_n7860), .B2(new_n506), .Y(new_n10348));
  AOI221xp5_ASAP7_75t_L     g10092(.A1(new_n475), .A2(\b[50] ), .B1(new_n483), .B2(new_n8763), .C(new_n10348), .Y(new_n10349));
  XNOR2x2_ASAP7_75t_L       g10093(.A(new_n466), .B(new_n10349), .Y(new_n10350));
  INVx1_ASAP7_75t_L         g10094(.A(new_n10350), .Y(new_n10351));
  A2O1A1O1Ixp25_ASAP7_75t_L g10095(.A1(new_n9732), .A2(new_n10286), .B(new_n10285), .C(new_n10272), .D(new_n10281), .Y(new_n10352));
  NAND2xp33_ASAP7_75t_L     g10096(.A(new_n10192), .B(new_n10193), .Y(new_n10353));
  MAJIxp5_ASAP7_75t_L       g10097(.A(new_n10206), .B(new_n10353), .C(new_n10199), .Y(new_n10354));
  NOR2xp33_ASAP7_75t_L      g10098(.A(new_n3674), .B(new_n2410), .Y(new_n10355));
  AOI221xp5_ASAP7_75t_L     g10099(.A1(\b[30] ), .A2(new_n2577), .B1(\b[32] ), .B2(new_n2423), .C(new_n10355), .Y(new_n10356));
  O2A1O1Ixp33_ASAP7_75t_L   g10100(.A1(new_n2425), .A2(new_n3897), .B(new_n10356), .C(new_n2413), .Y(new_n10357));
  INVx1_ASAP7_75t_L         g10101(.A(new_n10356), .Y(new_n10358));
  A2O1A1Ixp33_ASAP7_75t_L   g10102(.A1(new_n3900), .A2(new_n2417), .B(new_n10358), .C(new_n2413), .Y(new_n10359));
  OAI21xp33_ASAP7_75t_L     g10103(.A1(new_n2413), .A2(new_n10357), .B(new_n10359), .Y(new_n10360));
  INVx1_ASAP7_75t_L         g10104(.A(new_n10360), .Y(new_n10361));
  NOR2xp33_ASAP7_75t_L      g10105(.A(new_n2928), .B(new_n10186), .Y(new_n10362));
  O2A1O1Ixp33_ASAP7_75t_L   g10106(.A1(new_n2940), .A2(new_n3087), .B(new_n10184), .C(\a[29] ), .Y(new_n10363));
  OAI211xp5_ASAP7_75t_L     g10107(.A1(new_n10362), .A2(new_n10363), .B(new_n10177), .C(new_n10182), .Y(new_n10364));
  A2O1A1Ixp33_ASAP7_75t_L   g10108(.A1(new_n10188), .A2(new_n10189), .B(new_n10191), .C(new_n10364), .Y(new_n10365));
  A2O1A1Ixp33_ASAP7_75t_L   g10109(.A1(new_n10179), .A2(new_n10180), .B(new_n10176), .C(new_n10170), .Y(new_n10366));
  A2O1A1Ixp33_ASAP7_75t_L   g10110(.A1(new_n10157), .A2(new_n10145), .B(new_n10152), .C(new_n10164), .Y(new_n10367));
  A2O1A1Ixp33_ASAP7_75t_L   g10111(.A1(new_n10161), .A2(new_n10165), .B(new_n10167), .C(new_n10367), .Y(new_n10368));
  NAND2xp33_ASAP7_75t_L     g10112(.A(new_n10125), .B(new_n10129), .Y(new_n10369));
  MAJIxp5_ASAP7_75t_L       g10113(.A(new_n10137), .B(new_n10132), .C(new_n10369), .Y(new_n10370));
  OAI22xp33_ASAP7_75t_L     g10114(.A1(new_n5640), .A2(new_n1150), .B1(new_n1043), .B2(new_n5925), .Y(new_n10371));
  AOI221xp5_ASAP7_75t_L     g10115(.A1(new_n5629), .A2(\b[17] ), .B1(new_n5637), .B2(new_n1633), .C(new_n10371), .Y(new_n10372));
  XNOR2x2_ASAP7_75t_L       g10116(.A(\a[41] ), .B(new_n10372), .Y(new_n10373));
  NOR3xp33_ASAP7_75t_L      g10117(.A(new_n10115), .B(new_n10117), .C(new_n10057), .Y(new_n10374));
  A2O1A1O1Ixp25_ASAP7_75t_L g10118(.A1(new_n9787), .A2(new_n9844), .B(new_n10126), .C(new_n10118), .D(new_n10374), .Y(new_n10375));
  INVx1_ASAP7_75t_L         g10119(.A(new_n10113), .Y(new_n10376));
  NOR2xp33_ASAP7_75t_L      g10120(.A(new_n680), .B(new_n7312), .Y(new_n10377));
  AOI221xp5_ASAP7_75t_L     g10121(.A1(\b[9] ), .A2(new_n7609), .B1(\b[11] ), .B2(new_n7334), .C(new_n10377), .Y(new_n10378));
  O2A1O1Ixp33_ASAP7_75t_L   g10122(.A1(new_n7321), .A2(new_n754), .B(new_n10378), .C(new_n7316), .Y(new_n10379));
  INVx1_ASAP7_75t_L         g10123(.A(new_n10378), .Y(new_n10380));
  A2O1A1Ixp33_ASAP7_75t_L   g10124(.A1(new_n976), .A2(new_n7322), .B(new_n10380), .C(new_n7316), .Y(new_n10381));
  OAI21xp33_ASAP7_75t_L     g10125(.A1(new_n7316), .A2(new_n10379), .B(new_n10381), .Y(new_n10382));
  A2O1A1Ixp33_ASAP7_75t_L   g10126(.A1(new_n9831), .A2(new_n10061), .B(new_n10109), .C(new_n10107), .Y(new_n10383));
  NAND2xp33_ASAP7_75t_L     g10127(.A(new_n9805), .B(new_n9449), .Y(new_n10384));
  A2O1A1Ixp33_ASAP7_75t_L   g10128(.A1(new_n9827), .A2(new_n10384), .B(new_n10103), .C(new_n10100), .Y(new_n10385));
  INVx1_ASAP7_75t_L         g10129(.A(new_n10088), .Y(new_n10386));
  INVx1_ASAP7_75t_L         g10130(.A(new_n10079), .Y(new_n10387));
  NAND2xp33_ASAP7_75t_L     g10131(.A(new_n10387), .B(new_n9804), .Y(new_n10388));
  NAND2xp33_ASAP7_75t_L     g10132(.A(\b[2] ), .B(new_n10086), .Y(new_n10389));
  NAND3xp33_ASAP7_75t_L     g10133(.A(new_n9804), .B(new_n10079), .C(new_n10085), .Y(new_n10390));
  OAI221xp5_ASAP7_75t_L     g10134(.A1(new_n10388), .A2(new_n262), .B1(new_n10390), .B2(new_n284), .C(new_n10389), .Y(new_n10391));
  A2O1A1Ixp33_ASAP7_75t_L   g10135(.A1(new_n294), .A2(new_n10386), .B(new_n10391), .C(\a[56] ), .Y(new_n10392));
  A2O1A1Ixp33_ASAP7_75t_L   g10136(.A1(new_n294), .A2(new_n10386), .B(new_n10391), .C(new_n10083), .Y(new_n10393));
  INVx1_ASAP7_75t_L         g10137(.A(new_n10393), .Y(new_n10394));
  A2O1A1O1Ixp25_ASAP7_75t_L g10138(.A1(new_n10090), .A2(new_n9815), .B(new_n10392), .C(\a[56] ), .D(new_n10394), .Y(new_n10395));
  NOR2xp33_ASAP7_75t_L      g10139(.A(new_n10088), .B(new_n509), .Y(new_n10396));
  NOR5xp2_ASAP7_75t_L       g10140(.A(new_n10089), .B(new_n10391), .C(new_n10396), .D(new_n9805), .E(new_n10083), .Y(new_n10397));
  INVx1_ASAP7_75t_L         g10141(.A(new_n9440), .Y(new_n10398));
  INVx1_ASAP7_75t_L         g10142(.A(new_n9095), .Y(new_n10399));
  NAND2xp33_ASAP7_75t_L     g10143(.A(new_n10399), .B(new_n8837), .Y(new_n10400));
  NOR2xp33_ASAP7_75t_L      g10144(.A(new_n332), .B(new_n10400), .Y(new_n10401));
  AOI221xp5_ASAP7_75t_L     g10145(.A1(new_n9102), .A2(\b[5] ), .B1(new_n10398), .B2(\b[3] ), .C(new_n10401), .Y(new_n10402));
  O2A1O1Ixp33_ASAP7_75t_L   g10146(.A1(new_n728), .A2(new_n9104), .B(new_n10402), .C(new_n9099), .Y(new_n10403));
  NOR2xp33_ASAP7_75t_L      g10147(.A(new_n9099), .B(new_n10403), .Y(new_n10404));
  O2A1O1Ixp33_ASAP7_75t_L   g10148(.A1(new_n728), .A2(new_n9104), .B(new_n10402), .C(\a[53] ), .Y(new_n10405));
  NOR2xp33_ASAP7_75t_L      g10149(.A(new_n10405), .B(new_n10404), .Y(new_n10406));
  NOR3xp33_ASAP7_75t_L      g10150(.A(new_n10406), .B(new_n10395), .C(new_n10397), .Y(new_n10407));
  NOR2xp33_ASAP7_75t_L      g10151(.A(new_n10396), .B(new_n10391), .Y(new_n10408));
  NAND2xp33_ASAP7_75t_L     g10152(.A(\a[56] ), .B(new_n10408), .Y(new_n10409));
  NAND3xp33_ASAP7_75t_L     g10153(.A(new_n10409), .B(new_n10091), .C(new_n10393), .Y(new_n10410));
  INVx1_ASAP7_75t_L         g10154(.A(new_n10397), .Y(new_n10411));
  INVx1_ASAP7_75t_L         g10155(.A(new_n10405), .Y(new_n10412));
  OAI21xp33_ASAP7_75t_L     g10156(.A1(new_n9099), .A2(new_n10403), .B(new_n10412), .Y(new_n10413));
  AOI21xp33_ASAP7_75t_L     g10157(.A1(new_n10410), .A2(new_n10411), .B(new_n10413), .Y(new_n10414));
  OAI21xp33_ASAP7_75t_L     g10158(.A1(new_n10407), .A2(new_n10414), .B(new_n10385), .Y(new_n10415));
  AOI21xp33_ASAP7_75t_L     g10159(.A1(new_n10096), .A2(new_n10072), .B(new_n10104), .Y(new_n10416));
  NAND3xp33_ASAP7_75t_L     g10160(.A(new_n10413), .B(new_n10410), .C(new_n10411), .Y(new_n10417));
  OAI21xp33_ASAP7_75t_L     g10161(.A1(new_n10397), .A2(new_n10395), .B(new_n10406), .Y(new_n10418));
  NAND3xp33_ASAP7_75t_L     g10162(.A(new_n10416), .B(new_n10417), .C(new_n10418), .Y(new_n10419));
  NOR2xp33_ASAP7_75t_L      g10163(.A(new_n448), .B(new_n10065), .Y(new_n10420));
  AOI221xp5_ASAP7_75t_L     g10164(.A1(new_n8175), .A2(\b[8] ), .B1(new_n8484), .B2(\b[6] ), .C(new_n10420), .Y(new_n10421));
  O2A1O1Ixp33_ASAP7_75t_L   g10165(.A1(new_n8176), .A2(new_n540), .B(new_n10421), .C(new_n8172), .Y(new_n10422));
  INVx1_ASAP7_75t_L         g10166(.A(new_n10422), .Y(new_n10423));
  O2A1O1Ixp33_ASAP7_75t_L   g10167(.A1(new_n8176), .A2(new_n540), .B(new_n10421), .C(\a[50] ), .Y(new_n10424));
  AOI21xp33_ASAP7_75t_L     g10168(.A1(new_n10423), .A2(\a[50] ), .B(new_n10424), .Y(new_n10425));
  NAND3xp33_ASAP7_75t_L     g10169(.A(new_n10419), .B(new_n10415), .C(new_n10425), .Y(new_n10426));
  AO21x2_ASAP7_75t_L        g10170(.A1(new_n10415), .A2(new_n10419), .B(new_n10425), .Y(new_n10427));
  NAND3xp33_ASAP7_75t_L     g10171(.A(new_n10383), .B(new_n10426), .C(new_n10427), .Y(new_n10428));
  AOI21xp33_ASAP7_75t_L     g10172(.A1(new_n10063), .A2(new_n10106), .B(new_n10110), .Y(new_n10429));
  AND3x1_ASAP7_75t_L        g10173(.A(new_n10419), .B(new_n10425), .C(new_n10415), .Y(new_n10430));
  AOI21xp33_ASAP7_75t_L     g10174(.A1(new_n10419), .A2(new_n10415), .B(new_n10425), .Y(new_n10431));
  OAI21xp33_ASAP7_75t_L     g10175(.A1(new_n10430), .A2(new_n10431), .B(new_n10429), .Y(new_n10432));
  AOI21xp33_ASAP7_75t_L     g10176(.A1(new_n10428), .A2(new_n10432), .B(new_n10382), .Y(new_n10433));
  INVx1_ASAP7_75t_L         g10177(.A(new_n10382), .Y(new_n10434));
  NOR3xp33_ASAP7_75t_L      g10178(.A(new_n10429), .B(new_n10430), .C(new_n10431), .Y(new_n10435));
  AOI21xp33_ASAP7_75t_L     g10179(.A1(new_n10427), .A2(new_n10426), .B(new_n10383), .Y(new_n10436));
  NOR3xp33_ASAP7_75t_L      g10180(.A(new_n10435), .B(new_n10436), .C(new_n10434), .Y(new_n10437));
  NOR2xp33_ASAP7_75t_L      g10181(.A(new_n10433), .B(new_n10437), .Y(new_n10438));
  A2O1A1Ixp33_ASAP7_75t_L   g10182(.A1(new_n10112), .A2(new_n10116), .B(new_n10376), .C(new_n10438), .Y(new_n10439));
  O2A1O1Ixp33_ASAP7_75t_L   g10183(.A1(new_n7316), .A2(new_n9796), .B(new_n9849), .C(new_n9850), .Y(new_n10440));
  O2A1O1Ixp33_ASAP7_75t_L   g10184(.A1(new_n10440), .A2(new_n9838), .B(new_n10112), .C(new_n10376), .Y(new_n10441));
  OAI21xp33_ASAP7_75t_L     g10185(.A1(new_n10436), .A2(new_n10435), .B(new_n10434), .Y(new_n10442));
  NAND3xp33_ASAP7_75t_L     g10186(.A(new_n10428), .B(new_n10382), .C(new_n10432), .Y(new_n10443));
  NAND2xp33_ASAP7_75t_L     g10187(.A(new_n10443), .B(new_n10442), .Y(new_n10444));
  NAND2xp33_ASAP7_75t_L     g10188(.A(new_n10444), .B(new_n10441), .Y(new_n10445));
  OAI22xp33_ASAP7_75t_L     g10189(.A1(new_n7304), .A2(new_n936), .B1(new_n833), .B2(new_n6741), .Y(new_n10446));
  AOI221xp5_ASAP7_75t_L     g10190(.A1(new_n6442), .A2(\b[14] ), .B1(new_n6450), .B2(new_n971), .C(new_n10446), .Y(new_n10447));
  XNOR2x2_ASAP7_75t_L       g10191(.A(new_n6439), .B(new_n10447), .Y(new_n10448));
  NAND3xp33_ASAP7_75t_L     g10192(.A(new_n10439), .B(new_n10448), .C(new_n10445), .Y(new_n10449));
  O2A1O1Ixp33_ASAP7_75t_L   g10193(.A1(new_n10122), .A2(new_n10114), .B(new_n10113), .C(new_n10444), .Y(new_n10450));
  A2O1A1Ixp33_ASAP7_75t_L   g10194(.A1(new_n9797), .A2(\a[47] ), .B(new_n9798), .C(new_n9851), .Y(new_n10451));
  A2O1A1Ixp33_ASAP7_75t_L   g10195(.A1(new_n10451), .A2(new_n9841), .B(new_n10114), .C(new_n10113), .Y(new_n10452));
  NOR2xp33_ASAP7_75t_L      g10196(.A(new_n10438), .B(new_n10452), .Y(new_n10453));
  XNOR2x2_ASAP7_75t_L       g10197(.A(\a[44] ), .B(new_n10447), .Y(new_n10454));
  OAI21xp33_ASAP7_75t_L     g10198(.A1(new_n10450), .A2(new_n10453), .B(new_n10454), .Y(new_n10455));
  AOI21xp33_ASAP7_75t_L     g10199(.A1(new_n10455), .A2(new_n10449), .B(new_n10375), .Y(new_n10456));
  AND3x1_ASAP7_75t_L        g10200(.A(new_n10375), .B(new_n10455), .C(new_n10449), .Y(new_n10457));
  OAI21xp33_ASAP7_75t_L     g10201(.A1(new_n10456), .A2(new_n10457), .B(new_n10373), .Y(new_n10458));
  XNOR2x2_ASAP7_75t_L       g10202(.A(new_n5626), .B(new_n10372), .Y(new_n10459));
  AO21x2_ASAP7_75t_L        g10203(.A1(new_n10455), .A2(new_n10449), .B(new_n10375), .Y(new_n10460));
  NAND3xp33_ASAP7_75t_L     g10204(.A(new_n10375), .B(new_n10449), .C(new_n10455), .Y(new_n10461));
  NAND3xp33_ASAP7_75t_L     g10205(.A(new_n10460), .B(new_n10459), .C(new_n10461), .Y(new_n10462));
  NAND2xp33_ASAP7_75t_L     g10206(.A(new_n10462), .B(new_n10458), .Y(new_n10463));
  NAND2xp33_ASAP7_75t_L     g10207(.A(new_n10370), .B(new_n10463), .Y(new_n10464));
  NOR3xp33_ASAP7_75t_L      g10208(.A(new_n10457), .B(new_n10456), .C(new_n10459), .Y(new_n10465));
  O2A1O1Ixp33_ASAP7_75t_L   g10209(.A1(new_n10459), .A2(new_n10465), .B(new_n10462), .C(new_n10370), .Y(new_n10466));
  NOR2xp33_ASAP7_75t_L      g10210(.A(new_n1745), .B(new_n4908), .Y(new_n10467));
  AOI221xp5_ASAP7_75t_L     g10211(.A1(\b[18] ), .A2(new_n5139), .B1(\b[19] ), .B2(new_n4916), .C(new_n10467), .Y(new_n10468));
  O2A1O1Ixp33_ASAP7_75t_L   g10212(.A1(new_n4911), .A2(new_n1754), .B(new_n10468), .C(new_n4906), .Y(new_n10469));
  OAI21xp33_ASAP7_75t_L     g10213(.A1(new_n4911), .A2(new_n1754), .B(new_n10468), .Y(new_n10470));
  NAND2xp33_ASAP7_75t_L     g10214(.A(new_n4906), .B(new_n10470), .Y(new_n10471));
  OA21x2_ASAP7_75t_L        g10215(.A1(new_n4906), .A2(new_n10469), .B(new_n10471), .Y(new_n10472));
  A2O1A1Ixp33_ASAP7_75t_L   g10216(.A1(new_n10464), .A2(new_n10370), .B(new_n10466), .C(new_n10472), .Y(new_n10473));
  AOI21xp33_ASAP7_75t_L     g10217(.A1(new_n10460), .A2(new_n10461), .B(new_n10459), .Y(new_n10474));
  NOR3xp33_ASAP7_75t_L      g10218(.A(new_n10457), .B(new_n10456), .C(new_n10373), .Y(new_n10475));
  NOR2xp33_ASAP7_75t_L      g10219(.A(new_n10474), .B(new_n10475), .Y(new_n10476));
  NAND2xp33_ASAP7_75t_L     g10220(.A(new_n10370), .B(new_n10476), .Y(new_n10477));
  OAI211xp5_ASAP7_75t_L     g10221(.A1(new_n10369), .A2(new_n10132), .B(new_n10463), .C(new_n10140), .Y(new_n10478));
  OAI21xp33_ASAP7_75t_L     g10222(.A1(new_n4906), .A2(new_n10469), .B(new_n10471), .Y(new_n10479));
  NAND3xp33_ASAP7_75t_L     g10223(.A(new_n10478), .B(new_n10477), .C(new_n10479), .Y(new_n10480));
  NAND2xp33_ASAP7_75t_L     g10224(.A(new_n10480), .B(new_n10473), .Y(new_n10481));
  NOR2xp33_ASAP7_75t_L      g10225(.A(new_n10157), .B(new_n10481), .Y(new_n10482));
  AOI211xp5_ASAP7_75t_L     g10226(.A1(new_n10473), .A2(new_n10480), .B(new_n10162), .C(new_n10149), .Y(new_n10483));
  NAND2xp33_ASAP7_75t_L     g10227(.A(\b[22] ), .B(new_n4155), .Y(new_n10484));
  OAI221xp5_ASAP7_75t_L     g10228(.A1(new_n4147), .A2(new_n2188), .B1(new_n1895), .B2(new_n4397), .C(new_n10484), .Y(new_n10485));
  A2O1A1Ixp33_ASAP7_75t_L   g10229(.A1(new_n2679), .A2(new_n4151), .B(new_n10485), .C(\a[35] ), .Y(new_n10486));
  AOI211xp5_ASAP7_75t_L     g10230(.A1(new_n2679), .A2(new_n4151), .B(new_n10485), .C(new_n4145), .Y(new_n10487));
  A2O1A1O1Ixp25_ASAP7_75t_L g10231(.A1(new_n4151), .A2(new_n2679), .B(new_n10485), .C(new_n10486), .D(new_n10487), .Y(new_n10488));
  INVx1_ASAP7_75t_L         g10232(.A(new_n10488), .Y(new_n10489));
  OAI21xp33_ASAP7_75t_L     g10233(.A1(new_n10483), .A2(new_n10482), .B(new_n10489), .Y(new_n10490));
  OAI211xp5_ASAP7_75t_L     g10234(.A1(new_n10149), .A2(new_n10162), .B(new_n10473), .C(new_n10480), .Y(new_n10491));
  A2O1A1Ixp33_ASAP7_75t_L   g10235(.A1(new_n10464), .A2(new_n10370), .B(new_n10466), .C(new_n10479), .Y(new_n10492));
  AOI21xp33_ASAP7_75t_L     g10236(.A1(new_n10478), .A2(new_n10477), .B(new_n10479), .Y(new_n10493));
  A2O1A1Ixp33_ASAP7_75t_L   g10237(.A1(new_n10479), .A2(new_n10492), .B(new_n10493), .C(new_n10157), .Y(new_n10494));
  NAND3xp33_ASAP7_75t_L     g10238(.A(new_n10494), .B(new_n10491), .C(new_n10488), .Y(new_n10495));
  AOI21xp33_ASAP7_75t_L     g10239(.A1(new_n10495), .A2(new_n10490), .B(new_n10368), .Y(new_n10496));
  A2O1A1O1Ixp25_ASAP7_75t_L g10240(.A1(new_n10140), .A2(new_n10138), .B(new_n10150), .C(new_n10157), .D(new_n10152), .Y(new_n10497));
  NAND2xp33_ASAP7_75t_L     g10241(.A(new_n10495), .B(new_n10490), .Y(new_n10498));
  O2A1O1Ixp33_ASAP7_75t_L   g10242(.A1(new_n10497), .A2(new_n10160), .B(new_n10169), .C(new_n10498), .Y(new_n10499));
  OAI22xp33_ASAP7_75t_L     g10243(.A1(new_n3703), .A2(new_n2205), .B1(new_n2377), .B2(new_n3509), .Y(new_n10500));
  AOI221xp5_ASAP7_75t_L     g10244(.A1(new_n3503), .A2(\b[26] ), .B1(new_n3505), .B2(new_n2709), .C(new_n10500), .Y(new_n10501));
  XNOR2x2_ASAP7_75t_L       g10245(.A(new_n3493), .B(new_n10501), .Y(new_n10502));
  NOR3xp33_ASAP7_75t_L      g10246(.A(new_n10499), .B(new_n10502), .C(new_n10496), .Y(new_n10503));
  NAND3xp33_ASAP7_75t_L     g10247(.A(new_n10498), .B(new_n10169), .C(new_n10367), .Y(new_n10504));
  NAND3xp33_ASAP7_75t_L     g10248(.A(new_n10368), .B(new_n10490), .C(new_n10495), .Y(new_n10505));
  XNOR2x2_ASAP7_75t_L       g10249(.A(\a[32] ), .B(new_n10501), .Y(new_n10506));
  AOI21xp33_ASAP7_75t_L     g10250(.A1(new_n10504), .A2(new_n10505), .B(new_n10506), .Y(new_n10507));
  OAI21xp33_ASAP7_75t_L     g10251(.A1(new_n10503), .A2(new_n10507), .B(new_n10366), .Y(new_n10508));
  INVx1_ASAP7_75t_L         g10252(.A(new_n10170), .Y(new_n10509));
  A2O1A1O1Ixp25_ASAP7_75t_L g10253(.A1(new_n9893), .A2(new_n9885), .B(new_n10175), .C(new_n10181), .D(new_n10509), .Y(new_n10510));
  NAND3xp33_ASAP7_75t_L     g10254(.A(new_n10504), .B(new_n10505), .C(new_n10506), .Y(new_n10511));
  OAI21xp33_ASAP7_75t_L     g10255(.A1(new_n10496), .A2(new_n10499), .B(new_n10502), .Y(new_n10512));
  NAND3xp33_ASAP7_75t_L     g10256(.A(new_n10510), .B(new_n10511), .C(new_n10512), .Y(new_n10513));
  OAI22xp33_ASAP7_75t_L     g10257(.A1(new_n3133), .A2(new_n2879), .B1(new_n3079), .B2(new_n2925), .Y(new_n10514));
  AOI221xp5_ASAP7_75t_L     g10258(.A1(new_n2938), .A2(\b[29] ), .B1(new_n2932), .B2(new_n3873), .C(new_n10514), .Y(new_n10515));
  XNOR2x2_ASAP7_75t_L       g10259(.A(new_n2928), .B(new_n10515), .Y(new_n10516));
  NAND3xp33_ASAP7_75t_L     g10260(.A(new_n10513), .B(new_n10508), .C(new_n10516), .Y(new_n10517));
  AO21x2_ASAP7_75t_L        g10261(.A1(new_n10508), .A2(new_n10513), .B(new_n10516), .Y(new_n10518));
  AND3x1_ASAP7_75t_L        g10262(.A(new_n10365), .B(new_n10518), .C(new_n10517), .Y(new_n10519));
  AOI21xp33_ASAP7_75t_L     g10263(.A1(new_n10518), .A2(new_n10517), .B(new_n10365), .Y(new_n10520));
  OAI21xp33_ASAP7_75t_L     g10264(.A1(new_n10520), .A2(new_n10519), .B(new_n10361), .Y(new_n10521));
  NAND3xp33_ASAP7_75t_L     g10265(.A(new_n10365), .B(new_n10518), .C(new_n10517), .Y(new_n10522));
  AO21x2_ASAP7_75t_L        g10266(.A1(new_n10517), .A2(new_n10518), .B(new_n10365), .Y(new_n10523));
  NAND3xp33_ASAP7_75t_L     g10267(.A(new_n10523), .B(new_n10522), .C(new_n10360), .Y(new_n10524));
  NAND3xp33_ASAP7_75t_L     g10268(.A(new_n10354), .B(new_n10521), .C(new_n10524), .Y(new_n10525));
  NOR2xp33_ASAP7_75t_L      g10269(.A(new_n10202), .B(new_n10201), .Y(new_n10526));
  MAJIxp5_ASAP7_75t_L       g10270(.A(new_n10210), .B(new_n10204), .C(new_n10526), .Y(new_n10527));
  AOI21xp33_ASAP7_75t_L     g10271(.A1(new_n10523), .A2(new_n10522), .B(new_n10360), .Y(new_n10528));
  NOR3xp33_ASAP7_75t_L      g10272(.A(new_n10519), .B(new_n10520), .C(new_n10361), .Y(new_n10529));
  OAI21xp33_ASAP7_75t_L     g10273(.A1(new_n10528), .A2(new_n10529), .B(new_n10527), .Y(new_n10530));
  OAI22xp33_ASAP7_75t_L     g10274(.A1(new_n2089), .A2(new_n4101), .B1(new_n4344), .B2(new_n1962), .Y(new_n10531));
  AOI221xp5_ASAP7_75t_L     g10275(.A1(new_n1955), .A2(\b[35] ), .B1(new_n1964), .B2(new_n7773), .C(new_n10531), .Y(new_n10532));
  XNOR2x2_ASAP7_75t_L       g10276(.A(new_n1952), .B(new_n10532), .Y(new_n10533));
  NAND3xp33_ASAP7_75t_L     g10277(.A(new_n10525), .B(new_n10530), .C(new_n10533), .Y(new_n10534));
  NOR3xp33_ASAP7_75t_L      g10278(.A(new_n10527), .B(new_n10528), .C(new_n10529), .Y(new_n10535));
  AOI21xp33_ASAP7_75t_L     g10279(.A1(new_n10524), .A2(new_n10521), .B(new_n10354), .Y(new_n10536));
  AND2x2_ASAP7_75t_L        g10280(.A(\a[23] ), .B(new_n10532), .Y(new_n10537));
  NOR2xp33_ASAP7_75t_L      g10281(.A(\a[23] ), .B(new_n10532), .Y(new_n10538));
  OAI22xp33_ASAP7_75t_L     g10282(.A1(new_n10536), .A2(new_n10535), .B1(new_n10538), .B2(new_n10537), .Y(new_n10539));
  NAND2xp33_ASAP7_75t_L     g10283(.A(new_n10534), .B(new_n10539), .Y(new_n10540));
  NAND2xp33_ASAP7_75t_L     g10284(.A(new_n10211), .B(new_n10207), .Y(new_n10541));
  MAJIxp5_ASAP7_75t_L       g10285(.A(new_n10225), .B(new_n10541), .C(new_n10217), .Y(new_n10542));
  NOR2xp33_ASAP7_75t_L      g10286(.A(new_n10540), .B(new_n10542), .Y(new_n10543));
  NOR3xp33_ASAP7_75t_L      g10287(.A(new_n10536), .B(new_n10535), .C(new_n10533), .Y(new_n10544));
  O2A1O1Ixp33_ASAP7_75t_L   g10288(.A1(new_n10214), .A2(new_n1952), .B(new_n10216), .C(new_n10541), .Y(new_n10545));
  A2O1A1O1Ixp25_ASAP7_75t_L g10289(.A1(new_n9746), .A2(new_n9934), .B(new_n10224), .C(new_n10227), .D(new_n10545), .Y(new_n10546));
  O2A1O1Ixp33_ASAP7_75t_L   g10290(.A1(new_n10533), .A2(new_n10544), .B(new_n10534), .C(new_n10546), .Y(new_n10547));
  OAI22xp33_ASAP7_75t_L     g10291(.A1(new_n1654), .A2(new_n4613), .B1(new_n5074), .B2(new_n1517), .Y(new_n10548));
  AOI221xp5_ASAP7_75t_L     g10292(.A1(new_n1511), .A2(\b[38] ), .B1(new_n1513), .B2(new_n6083), .C(new_n10548), .Y(new_n10549));
  XNOR2x2_ASAP7_75t_L       g10293(.A(\a[20] ), .B(new_n10549), .Y(new_n10550));
  NOR3xp33_ASAP7_75t_L      g10294(.A(new_n10547), .B(new_n10550), .C(new_n10543), .Y(new_n10551));
  AND2x2_ASAP7_75t_L        g10295(.A(new_n10534), .B(new_n10539), .Y(new_n10552));
  NAND2xp33_ASAP7_75t_L     g10296(.A(new_n10546), .B(new_n10552), .Y(new_n10553));
  NAND2xp33_ASAP7_75t_L     g10297(.A(new_n10540), .B(new_n10542), .Y(new_n10554));
  INVx1_ASAP7_75t_L         g10298(.A(new_n10550), .Y(new_n10555));
  AOI21xp33_ASAP7_75t_L     g10299(.A1(new_n10553), .A2(new_n10554), .B(new_n10555), .Y(new_n10556));
  NAND2xp33_ASAP7_75t_L     g10300(.A(new_n10228), .B(new_n10226), .Y(new_n10557));
  MAJIxp5_ASAP7_75t_L       g10301(.A(new_n10235), .B(new_n10557), .C(new_n10232), .Y(new_n10558));
  NOR3xp33_ASAP7_75t_L      g10302(.A(new_n10558), .B(new_n10556), .C(new_n10551), .Y(new_n10559));
  OA21x2_ASAP7_75t_L        g10303(.A1(new_n10551), .A2(new_n10556), .B(new_n10558), .Y(new_n10560));
  NOR2xp33_ASAP7_75t_L      g10304(.A(new_n6110), .B(new_n1284), .Y(new_n10561));
  AOI221xp5_ASAP7_75t_L     g10305(.A1(\b[39] ), .A2(new_n1290), .B1(\b[40] ), .B2(new_n1204), .C(new_n10561), .Y(new_n10562));
  O2A1O1Ixp33_ASAP7_75t_L   g10306(.A1(new_n1210), .A2(new_n6117), .B(new_n10562), .C(new_n1206), .Y(new_n10563));
  OAI21xp33_ASAP7_75t_L     g10307(.A1(new_n1210), .A2(new_n6117), .B(new_n10562), .Y(new_n10564));
  NAND2xp33_ASAP7_75t_L     g10308(.A(new_n1206), .B(new_n10564), .Y(new_n10565));
  OAI21xp33_ASAP7_75t_L     g10309(.A1(new_n1206), .A2(new_n10563), .B(new_n10565), .Y(new_n10566));
  NOR3xp33_ASAP7_75t_L      g10310(.A(new_n10560), .B(new_n10566), .C(new_n10559), .Y(new_n10567));
  OR2x4_ASAP7_75t_L         g10311(.A(new_n10232), .B(new_n10557), .Y(new_n10568));
  NAND3xp33_ASAP7_75t_L     g10312(.A(new_n10555), .B(new_n10553), .C(new_n10554), .Y(new_n10569));
  OAI21xp33_ASAP7_75t_L     g10313(.A1(new_n10543), .A2(new_n10547), .B(new_n10550), .Y(new_n10570));
  NAND4xp25_ASAP7_75t_L     g10314(.A(new_n10237), .B(new_n10569), .C(new_n10570), .D(new_n10568), .Y(new_n10571));
  OAI21xp33_ASAP7_75t_L     g10315(.A1(new_n10551), .A2(new_n10556), .B(new_n10558), .Y(new_n10572));
  INVx1_ASAP7_75t_L         g10316(.A(new_n10566), .Y(new_n10573));
  AOI21xp33_ASAP7_75t_L     g10317(.A1(new_n10571), .A2(new_n10572), .B(new_n10573), .Y(new_n10574));
  NOR2xp33_ASAP7_75t_L      g10318(.A(new_n10574), .B(new_n10567), .Y(new_n10575));
  INVx1_ASAP7_75t_L         g10319(.A(new_n10255), .Y(new_n10576));
  AOI21xp33_ASAP7_75t_L     g10320(.A1(new_n10252), .A2(new_n10249), .B(new_n10576), .Y(new_n10577));
  NAND2xp33_ASAP7_75t_L     g10321(.A(new_n10577), .B(new_n10575), .Y(new_n10578));
  NAND3xp33_ASAP7_75t_L     g10322(.A(new_n10571), .B(new_n10572), .C(new_n10573), .Y(new_n10579));
  OAI21xp33_ASAP7_75t_L     g10323(.A1(new_n10559), .A2(new_n10560), .B(new_n10566), .Y(new_n10580));
  NAND2xp33_ASAP7_75t_L     g10324(.A(new_n10579), .B(new_n10580), .Y(new_n10581));
  A2O1A1Ixp33_ASAP7_75t_L   g10325(.A1(new_n10249), .A2(new_n10252), .B(new_n10576), .C(new_n10581), .Y(new_n10582));
  NOR2xp33_ASAP7_75t_L      g10326(.A(new_n6944), .B(new_n869), .Y(new_n10583));
  AOI221xp5_ASAP7_75t_L     g10327(.A1(\b[42] ), .A2(new_n985), .B1(\b[43] ), .B2(new_n885), .C(new_n10583), .Y(new_n10584));
  O2A1O1Ixp33_ASAP7_75t_L   g10328(.A1(new_n872), .A2(new_n6951), .B(new_n10584), .C(new_n867), .Y(new_n10585));
  OAI21xp33_ASAP7_75t_L     g10329(.A1(new_n872), .A2(new_n6951), .B(new_n10584), .Y(new_n10586));
  NAND2xp33_ASAP7_75t_L     g10330(.A(new_n867), .B(new_n10586), .Y(new_n10587));
  OAI21xp33_ASAP7_75t_L     g10331(.A1(new_n867), .A2(new_n10585), .B(new_n10587), .Y(new_n10588));
  NAND3xp33_ASAP7_75t_L     g10332(.A(new_n10582), .B(new_n10578), .C(new_n10588), .Y(new_n10589));
  A2O1A1Ixp33_ASAP7_75t_L   g10333(.A1(new_n9970), .A2(new_n10251), .B(new_n10257), .C(new_n10255), .Y(new_n10590));
  NOR2xp33_ASAP7_75t_L      g10334(.A(new_n10581), .B(new_n10590), .Y(new_n10591));
  NAND3xp33_ASAP7_75t_L     g10335(.A(new_n10571), .B(new_n10572), .C(new_n10566), .Y(new_n10592));
  INVx1_ASAP7_75t_L         g10336(.A(new_n10592), .Y(new_n10593));
  O2A1O1Ixp33_ASAP7_75t_L   g10337(.A1(new_n10573), .A2(new_n10593), .B(new_n10579), .C(new_n10577), .Y(new_n10594));
  INVx1_ASAP7_75t_L         g10338(.A(new_n10588), .Y(new_n10595));
  OAI21xp33_ASAP7_75t_L     g10339(.A1(new_n10594), .A2(new_n10591), .B(new_n10595), .Y(new_n10596));
  AOI21xp33_ASAP7_75t_L     g10340(.A1(new_n10596), .A2(new_n10589), .B(new_n10274), .Y(new_n10597));
  AND3x1_ASAP7_75t_L        g10341(.A(new_n10274), .B(new_n10596), .C(new_n10589), .Y(new_n10598));
  NOR2xp33_ASAP7_75t_L      g10342(.A(new_n10597), .B(new_n10598), .Y(new_n10599));
  AOI21xp33_ASAP7_75t_L     g10343(.A1(new_n10582), .A2(new_n10578), .B(new_n10588), .Y(new_n10600));
  O2A1O1Ixp33_ASAP7_75t_L   g10344(.A1(new_n10266), .A2(new_n10264), .B(new_n10267), .C(new_n10600), .Y(new_n10601));
  NAND3xp33_ASAP7_75t_L     g10345(.A(new_n10274), .B(new_n10589), .C(new_n10596), .Y(new_n10602));
  OAI22xp33_ASAP7_75t_L     g10346(.A1(new_n1550), .A2(new_n7270), .B1(new_n7249), .B2(new_n712), .Y(new_n10603));
  AOI221xp5_ASAP7_75t_L     g10347(.A1(new_n640), .A2(\b[47] ), .B1(new_n718), .B2(new_n8726), .C(new_n10603), .Y(new_n10604));
  XNOR2x2_ASAP7_75t_L       g10348(.A(\a[11] ), .B(new_n10604), .Y(new_n10605));
  INVx1_ASAP7_75t_L         g10349(.A(new_n10605), .Y(new_n10606));
  A2O1A1O1Ixp25_ASAP7_75t_L g10350(.A1(new_n10589), .A2(new_n10601), .B(new_n10274), .C(new_n10602), .D(new_n10606), .Y(new_n10607));
  O2A1O1Ixp33_ASAP7_75t_L   g10351(.A1(new_n10253), .A2(new_n10258), .B(new_n10261), .C(new_n10266), .Y(new_n10608));
  NOR3xp33_ASAP7_75t_L      g10352(.A(new_n10591), .B(new_n10594), .C(new_n10595), .Y(new_n10609));
  OAI22xp33_ASAP7_75t_L     g10353(.A1(new_n10608), .A2(new_n10262), .B1(new_n10600), .B2(new_n10609), .Y(new_n10610));
  NAND3xp33_ASAP7_75t_L     g10354(.A(new_n10610), .B(new_n10602), .C(new_n10605), .Y(new_n10611));
  O2A1O1Ixp33_ASAP7_75t_L   g10355(.A1(new_n10599), .A2(new_n10607), .B(new_n10611), .C(new_n10352), .Y(new_n10612));
  NAND2xp33_ASAP7_75t_L     g10356(.A(new_n9738), .B(new_n10278), .Y(new_n10613));
  A2O1A1Ixp33_ASAP7_75t_L   g10357(.A1(new_n9991), .A2(new_n10613), .B(new_n10280), .C(new_n10276), .Y(new_n10614));
  OAI21xp33_ASAP7_75t_L     g10358(.A1(new_n10597), .A2(new_n10598), .B(new_n10606), .Y(new_n10615));
  NAND2xp33_ASAP7_75t_L     g10359(.A(new_n10615), .B(new_n10611), .Y(new_n10616));
  NOR2xp33_ASAP7_75t_L      g10360(.A(new_n10614), .B(new_n10616), .Y(new_n10617));
  OAI21xp33_ASAP7_75t_L     g10361(.A1(new_n10612), .A2(new_n10617), .B(new_n10351), .Y(new_n10618));
  A2O1A1Ixp33_ASAP7_75t_L   g10362(.A1(new_n10589), .A2(new_n10601), .B(new_n10274), .C(new_n10602), .Y(new_n10619));
  A2O1A1O1Ixp25_ASAP7_75t_L g10363(.A1(new_n10263), .A2(new_n10046), .B(new_n10262), .C(new_n10596), .D(new_n10609), .Y(new_n10620));
  A2O1A1Ixp33_ASAP7_75t_L   g10364(.A1(new_n10620), .A2(new_n10596), .B(new_n10597), .C(new_n10605), .Y(new_n10621));
  NOR3xp33_ASAP7_75t_L      g10365(.A(new_n10598), .B(new_n10606), .C(new_n10597), .Y(new_n10622));
  A2O1A1Ixp33_ASAP7_75t_L   g10366(.A1(new_n10619), .A2(new_n10621), .B(new_n10622), .C(new_n10614), .Y(new_n10623));
  A2O1A1O1Ixp25_ASAP7_75t_L g10367(.A1(new_n10589), .A2(new_n10601), .B(new_n10274), .C(new_n10602), .D(new_n10605), .Y(new_n10624));
  NOR2xp33_ASAP7_75t_L      g10368(.A(new_n10624), .B(new_n10622), .Y(new_n10625));
  NAND2xp33_ASAP7_75t_L     g10369(.A(new_n10352), .B(new_n10625), .Y(new_n10626));
  NAND3xp33_ASAP7_75t_L     g10370(.A(new_n10626), .B(new_n10623), .C(new_n10350), .Y(new_n10627));
  AOI21xp33_ASAP7_75t_L     g10371(.A1(new_n10627), .A2(new_n10618), .B(new_n10347), .Y(new_n10628));
  NAND3xp33_ASAP7_75t_L     g10372(.A(new_n10626), .B(new_n10623), .C(new_n10351), .Y(new_n10629));
  NOR3xp33_ASAP7_75t_L      g10373(.A(new_n10617), .B(new_n10612), .C(new_n10351), .Y(new_n10630));
  A2O1A1Ixp33_ASAP7_75t_L   g10374(.A1(new_n10351), .A2(new_n10629), .B(new_n10630), .C(new_n10347), .Y(new_n10631));
  OAI22xp33_ASAP7_75t_L     g10375(.A1(new_n350), .A2(new_n9355), .B1(new_n8779), .B2(new_n375), .Y(new_n10632));
  AOI221xp5_ASAP7_75t_L     g10376(.A1(new_n361), .A2(\b[53] ), .B1(new_n359), .B2(new_n9690), .C(new_n10632), .Y(new_n10633));
  XNOR2x2_ASAP7_75t_L       g10377(.A(new_n346), .B(new_n10633), .Y(new_n10634));
  OAI211xp5_ASAP7_75t_L     g10378(.A1(new_n10347), .A2(new_n10628), .B(new_n10631), .C(new_n10634), .Y(new_n10635));
  NAND2xp33_ASAP7_75t_L     g10379(.A(new_n10618), .B(new_n10627), .Y(new_n10636));
  AO21x2_ASAP7_75t_L        g10380(.A1(new_n10627), .A2(new_n10618), .B(new_n10347), .Y(new_n10637));
  NOR2xp33_ASAP7_75t_L      g10381(.A(new_n10347), .B(new_n10636), .Y(new_n10638));
  INVx1_ASAP7_75t_L         g10382(.A(new_n10634), .Y(new_n10639));
  A2O1A1Ixp33_ASAP7_75t_L   g10383(.A1(new_n10637), .A2(new_n10636), .B(new_n10638), .C(new_n10639), .Y(new_n10640));
  NAND3xp33_ASAP7_75t_L     g10384(.A(new_n10346), .B(new_n10635), .C(new_n10640), .Y(new_n10641));
  NOR2xp33_ASAP7_75t_L      g10385(.A(new_n10301), .B(new_n10300), .Y(new_n10642));
  MAJIxp5_ASAP7_75t_L       g10386(.A(new_n10038), .B(new_n10302), .C(new_n10642), .Y(new_n10643));
  AOI211xp5_ASAP7_75t_L     g10387(.A1(new_n10637), .A2(new_n10636), .B(new_n10639), .C(new_n10638), .Y(new_n10644));
  O2A1O1Ixp33_ASAP7_75t_L   g10388(.A1(new_n10347), .A2(new_n10628), .B(new_n10631), .C(new_n10634), .Y(new_n10645));
  OAI21xp33_ASAP7_75t_L     g10389(.A1(new_n10645), .A2(new_n10644), .B(new_n10643), .Y(new_n10646));
  NAND3xp33_ASAP7_75t_L     g10390(.A(new_n10641), .B(new_n10646), .C(new_n10343), .Y(new_n10647));
  INVx1_ASAP7_75t_L         g10391(.A(new_n10647), .Y(new_n10648));
  NAND3xp33_ASAP7_75t_L     g10392(.A(new_n10641), .B(new_n10646), .C(new_n10344), .Y(new_n10649));
  A2O1A1O1Ixp25_ASAP7_75t_L g10393(.A1(new_n10029), .A2(new_n10032), .B(new_n10027), .C(new_n10326), .D(new_n10324), .Y(new_n10650));
  O2A1O1Ixp33_ASAP7_75t_L   g10394(.A1(new_n10344), .A2(new_n10648), .B(new_n10649), .C(new_n10650), .Y(new_n10651));
  OAI21xp33_ASAP7_75t_L     g10395(.A1(new_n10344), .A2(new_n10648), .B(new_n10649), .Y(new_n10652));
  INVx1_ASAP7_75t_L         g10396(.A(new_n10650), .Y(new_n10653));
  NOR2xp33_ASAP7_75t_L      g10397(.A(new_n10653), .B(new_n10652), .Y(new_n10654));
  NOR2xp33_ASAP7_75t_L      g10398(.A(new_n10651), .B(new_n10654), .Y(\f[56] ));
  NAND2xp33_ASAP7_75t_L     g10399(.A(new_n10302), .B(new_n10642), .Y(new_n10656));
  OAI21xp33_ASAP7_75t_L     g10400(.A1(new_n10306), .A2(new_n10307), .B(new_n10038), .Y(new_n10657));
  A2O1A1Ixp33_ASAP7_75t_L   g10401(.A1(new_n10657), .A2(new_n10656), .B(new_n10644), .C(new_n10640), .Y(new_n10658));
  OAI22xp33_ASAP7_75t_L     g10402(.A1(new_n350), .A2(new_n9683), .B1(new_n9355), .B2(new_n375), .Y(new_n10659));
  AOI221xp5_ASAP7_75t_L     g10403(.A1(new_n361), .A2(\b[54] ), .B1(new_n359), .B2(new_n9717), .C(new_n10659), .Y(new_n10660));
  XNOR2x2_ASAP7_75t_L       g10404(.A(new_n346), .B(new_n10660), .Y(new_n10661));
  INVx1_ASAP7_75t_L         g10405(.A(new_n10661), .Y(new_n10662));
  NOR2xp33_ASAP7_75t_L      g10406(.A(new_n8427), .B(new_n506), .Y(new_n10663));
  AOI221xp5_ASAP7_75t_L     g10407(.A1(\b[51] ), .A2(new_n475), .B1(new_n470), .B2(\b[50] ), .C(new_n10663), .Y(new_n10664));
  O2A1O1Ixp33_ASAP7_75t_L   g10408(.A1(new_n477), .A2(new_n8789), .B(new_n10664), .C(new_n466), .Y(new_n10665));
  OAI21xp33_ASAP7_75t_L     g10409(.A1(new_n477), .A2(new_n8789), .B(new_n10664), .Y(new_n10666));
  NAND2xp33_ASAP7_75t_L     g10410(.A(new_n466), .B(new_n10666), .Y(new_n10667));
  OAI21xp33_ASAP7_75t_L     g10411(.A1(new_n466), .A2(new_n10665), .B(new_n10667), .Y(new_n10668));
  INVx1_ASAP7_75t_L         g10412(.A(new_n10668), .Y(new_n10669));
  A2O1A1Ixp33_ASAP7_75t_L   g10413(.A1(new_n9741), .A2(new_n9983), .B(new_n9978), .C(new_n10263), .Y(new_n10670));
  A2O1A1Ixp33_ASAP7_75t_L   g10414(.A1(new_n10670), .A2(new_n10267), .B(new_n10600), .C(new_n10589), .Y(new_n10671));
  NOR2xp33_ASAP7_75t_L      g10415(.A(new_n7860), .B(new_n710), .Y(new_n10672));
  AOI221xp5_ASAP7_75t_L     g10416(.A1(\b[47] ), .A2(new_n635), .B1(\b[46] ), .B2(new_n713), .C(new_n10672), .Y(new_n10673));
  O2A1O1Ixp33_ASAP7_75t_L   g10417(.A1(new_n641), .A2(new_n7868), .B(new_n10673), .C(new_n637), .Y(new_n10674));
  OAI21xp33_ASAP7_75t_L     g10418(.A1(new_n641), .A2(new_n7868), .B(new_n10673), .Y(new_n10675));
  NAND2xp33_ASAP7_75t_L     g10419(.A(new_n637), .B(new_n10675), .Y(new_n10676));
  OAI21xp33_ASAP7_75t_L     g10420(.A1(new_n637), .A2(new_n10674), .B(new_n10676), .Y(new_n10677));
  NOR2xp33_ASAP7_75t_L      g10421(.A(new_n7249), .B(new_n869), .Y(new_n10678));
  AOI221xp5_ASAP7_75t_L     g10422(.A1(\b[43] ), .A2(new_n985), .B1(\b[44] ), .B2(new_n885), .C(new_n10678), .Y(new_n10679));
  O2A1O1Ixp33_ASAP7_75t_L   g10423(.A1(new_n872), .A2(new_n7255), .B(new_n10679), .C(new_n867), .Y(new_n10680));
  OAI21xp33_ASAP7_75t_L     g10424(.A1(new_n872), .A2(new_n7255), .B(new_n10679), .Y(new_n10681));
  NAND2xp33_ASAP7_75t_L     g10425(.A(new_n867), .B(new_n10681), .Y(new_n10682));
  OAI21xp33_ASAP7_75t_L     g10426(.A1(new_n867), .A2(new_n10680), .B(new_n10682), .Y(new_n10683));
  NOR2xp33_ASAP7_75t_L      g10427(.A(new_n10543), .B(new_n10547), .Y(new_n10684));
  NAND2xp33_ASAP7_75t_L     g10428(.A(new_n10550), .B(new_n10684), .Y(new_n10685));
  INVx1_ASAP7_75t_L         g10429(.A(new_n10544), .Y(new_n10686));
  A2O1A1Ixp33_ASAP7_75t_L   g10430(.A1(\a[26] ), .A2(new_n10197), .B(new_n10198), .C(new_n10526), .Y(new_n10687));
  A2O1A1Ixp33_ASAP7_75t_L   g10431(.A1(new_n10211), .A2(new_n10687), .B(new_n10528), .C(new_n10524), .Y(new_n10688));
  O2A1O1Ixp33_ASAP7_75t_L   g10432(.A1(new_n10174), .A2(new_n10176), .B(new_n10170), .C(new_n10507), .Y(new_n10689));
  A2O1A1O1Ixp25_ASAP7_75t_L g10433(.A1(new_n10511), .A2(new_n10689), .B(new_n10510), .C(new_n10513), .D(new_n10516), .Y(new_n10690));
  AO21x2_ASAP7_75t_L        g10434(.A1(new_n10517), .A2(new_n10365), .B(new_n10690), .Y(new_n10691));
  OAI22xp33_ASAP7_75t_L     g10435(.A1(new_n3133), .A2(new_n3079), .B1(new_n3098), .B2(new_n2925), .Y(new_n10692));
  AOI221xp5_ASAP7_75t_L     g10436(.A1(new_n2938), .A2(\b[30] ), .B1(new_n2932), .B2(new_n4813), .C(new_n10692), .Y(new_n10693));
  XNOR2x2_ASAP7_75t_L       g10437(.A(new_n2928), .B(new_n10693), .Y(new_n10694));
  A2O1A1Ixp33_ASAP7_75t_L   g10438(.A1(new_n9199), .A2(new_n9409), .B(new_n9195), .C(new_n9555), .Y(new_n10695));
  A2O1A1Ixp33_ASAP7_75t_L   g10439(.A1(new_n9892), .A2(new_n10695), .B(new_n9886), .C(new_n9881), .Y(new_n10696));
  A2O1A1O1Ixp25_ASAP7_75t_L g10440(.A1(new_n10181), .A2(new_n10696), .B(new_n10509), .C(new_n10512), .D(new_n10503), .Y(new_n10697));
  INVx1_ASAP7_75t_L         g10441(.A(new_n10149), .Y(new_n10698));
  A2O1A1Ixp33_ASAP7_75t_L   g10442(.A1(new_n9866), .A2(new_n10147), .B(new_n10151), .C(new_n10698), .Y(new_n10699));
  INVx1_ASAP7_75t_L         g10443(.A(new_n10492), .Y(new_n10700));
  NAND2xp33_ASAP7_75t_L     g10444(.A(\b[20] ), .B(new_n4916), .Y(new_n10701));
  OAI221xp5_ASAP7_75t_L     g10445(.A1(new_n4908), .A2(new_n1895), .B1(new_n1599), .B2(new_n5144), .C(new_n10701), .Y(new_n10702));
  A2O1A1Ixp33_ASAP7_75t_L   g10446(.A1(new_n2836), .A2(new_n4912), .B(new_n10702), .C(\a[38] ), .Y(new_n10703));
  AOI211xp5_ASAP7_75t_L     g10447(.A1(new_n2836), .A2(new_n4912), .B(new_n10702), .C(new_n4906), .Y(new_n10704));
  A2O1A1O1Ixp25_ASAP7_75t_L g10448(.A1(new_n4912), .A2(new_n2836), .B(new_n10702), .C(new_n10703), .D(new_n10704), .Y(new_n10705));
  AO21x2_ASAP7_75t_L        g10449(.A1(new_n10370), .A2(new_n10463), .B(new_n10465), .Y(new_n10706));
  NOR2xp33_ASAP7_75t_L      g10450(.A(new_n1458), .B(new_n5641), .Y(new_n10707));
  AOI221xp5_ASAP7_75t_L     g10451(.A1(\b[16] ), .A2(new_n5920), .B1(\b[17] ), .B2(new_n5623), .C(new_n10707), .Y(new_n10708));
  O2A1O1Ixp33_ASAP7_75t_L   g10452(.A1(new_n5630), .A2(new_n1464), .B(new_n10708), .C(new_n5626), .Y(new_n10709));
  OAI21xp33_ASAP7_75t_L     g10453(.A1(new_n5630), .A2(new_n1464), .B(new_n10708), .Y(new_n10710));
  NAND2xp33_ASAP7_75t_L     g10454(.A(new_n5626), .B(new_n10710), .Y(new_n10711));
  OA21x2_ASAP7_75t_L        g10455(.A1(new_n5626), .A2(new_n10709), .B(new_n10711), .Y(new_n10712));
  NAND3xp33_ASAP7_75t_L     g10456(.A(new_n10439), .B(new_n10454), .C(new_n10445), .Y(new_n10713));
  A2O1A1Ixp33_ASAP7_75t_L   g10457(.A1(new_n10449), .A2(new_n10455), .B(new_n10375), .C(new_n10713), .Y(new_n10714));
  NOR2xp33_ASAP7_75t_L      g10458(.A(new_n960), .B(new_n7304), .Y(new_n10715));
  AOI221xp5_ASAP7_75t_L     g10459(.A1(\b[13] ), .A2(new_n6742), .B1(\b[15] ), .B2(new_n6442), .C(new_n10715), .Y(new_n10716));
  O2A1O1Ixp33_ASAP7_75t_L   g10460(.A1(new_n6443), .A2(new_n1774), .B(new_n10716), .C(new_n6439), .Y(new_n10717));
  O2A1O1Ixp33_ASAP7_75t_L   g10461(.A1(new_n6443), .A2(new_n1774), .B(new_n10716), .C(\a[44] ), .Y(new_n10718));
  INVx1_ASAP7_75t_L         g10462(.A(new_n10718), .Y(new_n10719));
  OAI21xp33_ASAP7_75t_L     g10463(.A1(new_n6439), .A2(new_n10717), .B(new_n10719), .Y(new_n10720));
  NOR2xp33_ASAP7_75t_L      g10464(.A(new_n748), .B(new_n7312), .Y(new_n10721));
  AOI221xp5_ASAP7_75t_L     g10465(.A1(\b[10] ), .A2(new_n7609), .B1(\b[12] ), .B2(new_n7334), .C(new_n10721), .Y(new_n10722));
  O2A1O1Ixp33_ASAP7_75t_L   g10466(.A1(new_n7321), .A2(new_n841), .B(new_n10722), .C(new_n7316), .Y(new_n10723));
  NOR2xp33_ASAP7_75t_L      g10467(.A(new_n7316), .B(new_n10723), .Y(new_n10724));
  O2A1O1Ixp33_ASAP7_75t_L   g10468(.A1(new_n7321), .A2(new_n841), .B(new_n10722), .C(\a[47] ), .Y(new_n10725));
  NOR2xp33_ASAP7_75t_L      g10469(.A(new_n10725), .B(new_n10724), .Y(new_n10726));
  A2O1A1O1Ixp25_ASAP7_75t_L g10470(.A1(new_n10106), .A2(new_n10063), .B(new_n10110), .C(new_n10426), .D(new_n10431), .Y(new_n10727));
  O2A1O1Ixp33_ASAP7_75t_L   g10471(.A1(new_n10103), .A2(new_n10102), .B(new_n10100), .C(new_n10414), .Y(new_n10728));
  INVx1_ASAP7_75t_L         g10472(.A(\a[57] ), .Y(new_n10729));
  NAND2xp33_ASAP7_75t_L     g10473(.A(\a[56] ), .B(new_n10729), .Y(new_n10730));
  NAND2xp33_ASAP7_75t_L     g10474(.A(\a[57] ), .B(new_n10083), .Y(new_n10731));
  AND2x2_ASAP7_75t_L        g10475(.A(new_n10730), .B(new_n10731), .Y(new_n10732));
  NOR2xp33_ASAP7_75t_L      g10476(.A(new_n284), .B(new_n10732), .Y(new_n10733));
  INVx1_ASAP7_75t_L         g10477(.A(new_n10733), .Y(new_n10734));
  NOR2xp33_ASAP7_75t_L      g10478(.A(new_n10734), .B(new_n10397), .Y(new_n10735));
  NOR2xp33_ASAP7_75t_L      g10479(.A(new_n10733), .B(new_n10411), .Y(new_n10736));
  NAND2xp33_ASAP7_75t_L     g10480(.A(\b[3] ), .B(new_n10086), .Y(new_n10737));
  OAI221xp5_ASAP7_75t_L     g10481(.A1(new_n10388), .A2(new_n289), .B1(new_n262), .B2(new_n10390), .C(new_n10737), .Y(new_n10738));
  NOR2xp33_ASAP7_75t_L      g10482(.A(new_n10088), .B(new_n319), .Y(new_n10739));
  OR3x1_ASAP7_75t_L         g10483(.A(new_n10738), .B(new_n10083), .C(new_n10739), .Y(new_n10740));
  A2O1A1Ixp33_ASAP7_75t_L   g10484(.A1(new_n312), .A2(new_n10386), .B(new_n10738), .C(new_n10083), .Y(new_n10741));
  NAND2xp33_ASAP7_75t_L     g10485(.A(new_n10741), .B(new_n10740), .Y(new_n10742));
  OAI21xp33_ASAP7_75t_L     g10486(.A1(new_n10735), .A2(new_n10736), .B(new_n10742), .Y(new_n10743));
  A2O1A1Ixp33_ASAP7_75t_L   g10487(.A1(new_n10409), .A2(new_n10393), .B(new_n10091), .C(new_n10733), .Y(new_n10744));
  A2O1A1Ixp33_ASAP7_75t_L   g10488(.A1(new_n10730), .A2(new_n10731), .B(new_n284), .C(new_n10397), .Y(new_n10745));
  A2O1A1Ixp33_ASAP7_75t_L   g10489(.A1(new_n312), .A2(new_n10386), .B(new_n10738), .C(\a[56] ), .Y(new_n10746));
  NOR3xp33_ASAP7_75t_L      g10490(.A(new_n10738), .B(new_n10739), .C(new_n10083), .Y(new_n10747));
  O2A1O1Ixp33_ASAP7_75t_L   g10491(.A1(new_n10738), .A2(new_n10739), .B(new_n10746), .C(new_n10747), .Y(new_n10748));
  NAND3xp33_ASAP7_75t_L     g10492(.A(new_n10744), .B(new_n10748), .C(new_n10745), .Y(new_n10749));
  NAND2xp33_ASAP7_75t_L     g10493(.A(\b[5] ), .B(new_n9096), .Y(new_n10750));
  OAI221xp5_ASAP7_75t_L     g10494(.A1(new_n9440), .A2(new_n332), .B1(new_n427), .B2(new_n9439), .C(new_n10750), .Y(new_n10751));
  A2O1A1Ixp33_ASAP7_75t_L   g10495(.A1(new_n5363), .A2(new_n9437), .B(new_n10751), .C(\a[53] ), .Y(new_n10752));
  NAND2xp33_ASAP7_75t_L     g10496(.A(\a[53] ), .B(new_n10752), .Y(new_n10753));
  A2O1A1Ixp33_ASAP7_75t_L   g10497(.A1(new_n5363), .A2(new_n9437), .B(new_n10751), .C(new_n9099), .Y(new_n10754));
  NAND2xp33_ASAP7_75t_L     g10498(.A(new_n10754), .B(new_n10753), .Y(new_n10755));
  INVx1_ASAP7_75t_L         g10499(.A(new_n10755), .Y(new_n10756));
  NAND3xp33_ASAP7_75t_L     g10500(.A(new_n10743), .B(new_n10749), .C(new_n10756), .Y(new_n10757));
  AOI21xp33_ASAP7_75t_L     g10501(.A1(new_n10744), .A2(new_n10745), .B(new_n10748), .Y(new_n10758));
  NOR3xp33_ASAP7_75t_L      g10502(.A(new_n10736), .B(new_n10742), .C(new_n10735), .Y(new_n10759));
  OAI21xp33_ASAP7_75t_L     g10503(.A1(new_n10758), .A2(new_n10759), .B(new_n10755), .Y(new_n10760));
  OAI211xp5_ASAP7_75t_L     g10504(.A1(new_n10407), .A2(new_n10728), .B(new_n10760), .C(new_n10757), .Y(new_n10761));
  A2O1A1O1Ixp25_ASAP7_75t_L g10505(.A1(new_n10096), .A2(new_n10072), .B(new_n10104), .C(new_n10418), .D(new_n10407), .Y(new_n10762));
  NAND3xp33_ASAP7_75t_L     g10506(.A(new_n10743), .B(new_n10749), .C(new_n10755), .Y(new_n10763));
  NOR3xp33_ASAP7_75t_L      g10507(.A(new_n10759), .B(new_n10758), .C(new_n10755), .Y(new_n10764));
  A2O1A1Ixp33_ASAP7_75t_L   g10508(.A1(new_n10763), .A2(new_n10755), .B(new_n10764), .C(new_n10762), .Y(new_n10765));
  NAND2xp33_ASAP7_75t_L     g10509(.A(\b[8] ), .B(new_n8169), .Y(new_n10766));
  OAI221xp5_ASAP7_75t_L     g10510(.A1(new_n8483), .A2(new_n448), .B1(new_n590), .B2(new_n8843), .C(new_n10766), .Y(new_n10767));
  A2O1A1Ixp33_ASAP7_75t_L   g10511(.A1(new_n602), .A2(new_n8490), .B(new_n10767), .C(\a[50] ), .Y(new_n10768));
  NAND2xp33_ASAP7_75t_L     g10512(.A(\a[50] ), .B(new_n10768), .Y(new_n10769));
  A2O1A1Ixp33_ASAP7_75t_L   g10513(.A1(new_n602), .A2(new_n8490), .B(new_n10767), .C(new_n8172), .Y(new_n10770));
  AOI22xp33_ASAP7_75t_L     g10514(.A1(new_n10769), .A2(new_n10770), .B1(new_n10761), .B2(new_n10765), .Y(new_n10771));
  AOI21xp33_ASAP7_75t_L     g10515(.A1(new_n10743), .A2(new_n10749), .B(new_n10756), .Y(new_n10772));
  NOR3xp33_ASAP7_75t_L      g10516(.A(new_n10762), .B(new_n10764), .C(new_n10772), .Y(new_n10773));
  AOI211xp5_ASAP7_75t_L     g10517(.A1(new_n10760), .A2(new_n10757), .B(new_n10407), .C(new_n10728), .Y(new_n10774));
  NAND2xp33_ASAP7_75t_L     g10518(.A(new_n10770), .B(new_n10769), .Y(new_n10775));
  NOR3xp33_ASAP7_75t_L      g10519(.A(new_n10774), .B(new_n10775), .C(new_n10773), .Y(new_n10776));
  NOR3xp33_ASAP7_75t_L      g10520(.A(new_n10727), .B(new_n10771), .C(new_n10776), .Y(new_n10777));
  OAI21xp33_ASAP7_75t_L     g10521(.A1(new_n10773), .A2(new_n10774), .B(new_n10775), .Y(new_n10778));
  NAND4xp25_ASAP7_75t_L     g10522(.A(new_n10765), .B(new_n10761), .C(new_n10769), .D(new_n10770), .Y(new_n10779));
  AOI221xp5_ASAP7_75t_L     g10523(.A1(new_n10383), .A2(new_n10426), .B1(new_n10779), .B2(new_n10778), .C(new_n10431), .Y(new_n10780));
  OA21x2_ASAP7_75t_L        g10524(.A1(new_n10780), .A2(new_n10777), .B(new_n10726), .Y(new_n10781));
  NOR3xp33_ASAP7_75t_L      g10525(.A(new_n10777), .B(new_n10726), .C(new_n10780), .Y(new_n10782));
  NOR2xp33_ASAP7_75t_L      g10526(.A(new_n10782), .B(new_n10781), .Y(new_n10783));
  A2O1A1Ixp33_ASAP7_75t_L   g10527(.A1(new_n10438), .A2(new_n10452), .B(new_n10437), .C(new_n10783), .Y(new_n10784));
  A2O1A1O1Ixp25_ASAP7_75t_L g10528(.A1(new_n10112), .A2(new_n10116), .B(new_n10376), .C(new_n10442), .D(new_n10437), .Y(new_n10785));
  OAI21xp33_ASAP7_75t_L     g10529(.A1(new_n10781), .A2(new_n10782), .B(new_n10785), .Y(new_n10786));
  NAND3xp33_ASAP7_75t_L     g10530(.A(new_n10784), .B(new_n10720), .C(new_n10786), .Y(new_n10787));
  INVx1_ASAP7_75t_L         g10531(.A(new_n10717), .Y(new_n10788));
  AOI21xp33_ASAP7_75t_L     g10532(.A1(new_n10788), .A2(\a[44] ), .B(new_n10718), .Y(new_n10789));
  NOR3xp33_ASAP7_75t_L      g10533(.A(new_n10785), .B(new_n10781), .C(new_n10782), .Y(new_n10790));
  INVx1_ASAP7_75t_L         g10534(.A(new_n10786), .Y(new_n10791));
  OAI21xp33_ASAP7_75t_L     g10535(.A1(new_n10790), .A2(new_n10791), .B(new_n10789), .Y(new_n10792));
  NAND3xp33_ASAP7_75t_L     g10536(.A(new_n10714), .B(new_n10787), .C(new_n10792), .Y(new_n10793));
  NOR3xp33_ASAP7_75t_L      g10537(.A(new_n10453), .B(new_n10454), .C(new_n10450), .Y(new_n10794));
  AOI21xp33_ASAP7_75t_L     g10538(.A1(new_n10713), .A2(new_n10454), .B(new_n10794), .Y(new_n10795));
  NOR3xp33_ASAP7_75t_L      g10539(.A(new_n10789), .B(new_n10791), .C(new_n10790), .Y(new_n10796));
  AOI21xp33_ASAP7_75t_L     g10540(.A1(new_n10784), .A2(new_n10786), .B(new_n10720), .Y(new_n10797));
  OAI221xp5_ASAP7_75t_L     g10541(.A1(new_n10797), .A2(new_n10796), .B1(new_n10795), .B2(new_n10375), .C(new_n10713), .Y(new_n10798));
  AO21x2_ASAP7_75t_L        g10542(.A1(new_n10798), .A2(new_n10793), .B(new_n10712), .Y(new_n10799));
  NAND3xp33_ASAP7_75t_L     g10543(.A(new_n10793), .B(new_n10712), .C(new_n10798), .Y(new_n10800));
  NAND2xp33_ASAP7_75t_L     g10544(.A(new_n10800), .B(new_n10799), .Y(new_n10801));
  NAND2xp33_ASAP7_75t_L     g10545(.A(new_n10792), .B(new_n10787), .Y(new_n10802));
  XNOR2x2_ASAP7_75t_L       g10546(.A(new_n10714), .B(new_n10802), .Y(new_n10803));
  AOI221xp5_ASAP7_75t_L     g10547(.A1(new_n10803), .A2(new_n10712), .B1(new_n10370), .B2(new_n10463), .C(new_n10465), .Y(new_n10804));
  AOI221xp5_ASAP7_75t_L     g10548(.A1(new_n10706), .A2(new_n10801), .B1(new_n10799), .B2(new_n10804), .C(new_n10705), .Y(new_n10805));
  INVx1_ASAP7_75t_L         g10549(.A(new_n10705), .Y(new_n10806));
  O2A1O1Ixp33_ASAP7_75t_L   g10550(.A1(new_n10474), .A2(new_n10475), .B(new_n10370), .C(new_n10465), .Y(new_n10807));
  OAI21xp33_ASAP7_75t_L     g10551(.A1(new_n5626), .A2(new_n10709), .B(new_n10711), .Y(new_n10808));
  NAND3xp33_ASAP7_75t_L     g10552(.A(new_n10793), .B(new_n10808), .C(new_n10798), .Y(new_n10809));
  AOI21xp33_ASAP7_75t_L     g10553(.A1(new_n10793), .A2(new_n10798), .B(new_n10712), .Y(new_n10810));
  AOI21xp33_ASAP7_75t_L     g10554(.A1(new_n10803), .A2(new_n10809), .B(new_n10810), .Y(new_n10811));
  NAND3xp33_ASAP7_75t_L     g10555(.A(new_n10807), .B(new_n10799), .C(new_n10800), .Y(new_n10812));
  O2A1O1Ixp33_ASAP7_75t_L   g10556(.A1(new_n10807), .A2(new_n10811), .B(new_n10812), .C(new_n10806), .Y(new_n10813));
  NOR2xp33_ASAP7_75t_L      g10557(.A(new_n10805), .B(new_n10813), .Y(new_n10814));
  A2O1A1Ixp33_ASAP7_75t_L   g10558(.A1(new_n10481), .A2(new_n10699), .B(new_n10700), .C(new_n10814), .Y(new_n10815));
  O2A1O1Ixp33_ASAP7_75t_L   g10559(.A1(new_n10369), .A2(new_n10132), .B(new_n10140), .C(new_n10463), .Y(new_n10816));
  NOR3xp33_ASAP7_75t_L      g10560(.A(new_n10816), .B(new_n10466), .C(new_n10472), .Y(new_n10817));
  OAI22xp33_ASAP7_75t_L     g10561(.A1(new_n10162), .A2(new_n10149), .B1(new_n10817), .B2(new_n10493), .Y(new_n10818));
  OAI211xp5_ASAP7_75t_L     g10562(.A1(new_n10807), .A2(new_n10811), .B(new_n10806), .C(new_n10812), .Y(new_n10819));
  INVx1_ASAP7_75t_L         g10563(.A(new_n10809), .Y(new_n10820));
  O2A1O1Ixp33_ASAP7_75t_L   g10564(.A1(new_n10712), .A2(new_n10820), .B(new_n10800), .C(new_n10807), .Y(new_n10821));
  A2O1A1Ixp33_ASAP7_75t_L   g10565(.A1(new_n10804), .A2(new_n10799), .B(new_n10821), .C(new_n10705), .Y(new_n10822));
  NAND2xp33_ASAP7_75t_L     g10566(.A(new_n10819), .B(new_n10822), .Y(new_n10823));
  NAND3xp33_ASAP7_75t_L     g10567(.A(new_n10823), .B(new_n10818), .C(new_n10492), .Y(new_n10824));
  OAI22xp33_ASAP7_75t_L     g10568(.A1(new_n4397), .A2(new_n2045), .B1(new_n2188), .B2(new_n4142), .Y(new_n10825));
  AOI221xp5_ASAP7_75t_L     g10569(.A1(new_n4156), .A2(\b[24] ), .B1(new_n4151), .B2(new_n2216), .C(new_n10825), .Y(new_n10826));
  XNOR2x2_ASAP7_75t_L       g10570(.A(new_n4145), .B(new_n10826), .Y(new_n10827));
  NAND3xp33_ASAP7_75t_L     g10571(.A(new_n10815), .B(new_n10824), .C(new_n10827), .Y(new_n10828));
  O2A1O1Ixp33_ASAP7_75t_L   g10572(.A1(new_n10474), .A2(new_n10475), .B(new_n10464), .C(new_n10816), .Y(new_n10829));
  O2A1O1Ixp33_ASAP7_75t_L   g10573(.A1(new_n10829), .A2(new_n10472), .B(new_n10818), .C(new_n10823), .Y(new_n10830));
  A2O1A1Ixp33_ASAP7_75t_L   g10574(.A1(new_n10473), .A2(new_n10480), .B(new_n10157), .C(new_n10492), .Y(new_n10831));
  NOR2xp33_ASAP7_75t_L      g10575(.A(new_n10814), .B(new_n10831), .Y(new_n10832));
  INVx1_ASAP7_75t_L         g10576(.A(new_n10827), .Y(new_n10833));
  OAI21xp33_ASAP7_75t_L     g10577(.A1(new_n10832), .A2(new_n10830), .B(new_n10833), .Y(new_n10834));
  INVx1_ASAP7_75t_L         g10578(.A(new_n10367), .Y(new_n10835));
  INVx1_ASAP7_75t_L         g10579(.A(new_n10490), .Y(new_n10836));
  O2A1O1Ixp33_ASAP7_75t_L   g10580(.A1(new_n10835), .A2(new_n10172), .B(new_n10495), .C(new_n10836), .Y(new_n10837));
  NAND3xp33_ASAP7_75t_L     g10581(.A(new_n10837), .B(new_n10834), .C(new_n10828), .Y(new_n10838));
  NAND2xp33_ASAP7_75t_L     g10582(.A(new_n10828), .B(new_n10834), .Y(new_n10839));
  INVx1_ASAP7_75t_L         g10583(.A(new_n10495), .Y(new_n10840));
  A2O1A1Ixp33_ASAP7_75t_L   g10584(.A1(new_n10169), .A2(new_n10367), .B(new_n10840), .C(new_n10490), .Y(new_n10841));
  NAND2xp33_ASAP7_75t_L     g10585(.A(new_n10841), .B(new_n10839), .Y(new_n10842));
  OAI22xp33_ASAP7_75t_L     g10586(.A1(new_n3703), .A2(new_n2377), .B1(new_n2703), .B2(new_n3509), .Y(new_n10843));
  AOI221xp5_ASAP7_75t_L     g10587(.A1(new_n3503), .A2(\b[27] ), .B1(new_n3505), .B2(new_n2887), .C(new_n10843), .Y(new_n10844));
  XNOR2x2_ASAP7_75t_L       g10588(.A(\a[32] ), .B(new_n10844), .Y(new_n10845));
  AOI21xp33_ASAP7_75t_L     g10589(.A1(new_n10842), .A2(new_n10838), .B(new_n10845), .Y(new_n10846));
  NOR2xp33_ASAP7_75t_L      g10590(.A(new_n10841), .B(new_n10839), .Y(new_n10847));
  AOI21xp33_ASAP7_75t_L     g10591(.A1(new_n10834), .A2(new_n10828), .B(new_n10837), .Y(new_n10848));
  XNOR2x2_ASAP7_75t_L       g10592(.A(new_n3493), .B(new_n10844), .Y(new_n10849));
  NOR3xp33_ASAP7_75t_L      g10593(.A(new_n10847), .B(new_n10848), .C(new_n10849), .Y(new_n10850));
  NOR3xp33_ASAP7_75t_L      g10594(.A(new_n10697), .B(new_n10846), .C(new_n10850), .Y(new_n10851));
  OAI21xp33_ASAP7_75t_L     g10595(.A1(new_n10848), .A2(new_n10847), .B(new_n10849), .Y(new_n10852));
  NAND3xp33_ASAP7_75t_L     g10596(.A(new_n10842), .B(new_n10838), .C(new_n10845), .Y(new_n10853));
  AOI211xp5_ASAP7_75t_L     g10597(.A1(new_n10852), .A2(new_n10853), .B(new_n10689), .C(new_n10503), .Y(new_n10854));
  NOR3xp33_ASAP7_75t_L      g10598(.A(new_n10851), .B(new_n10854), .C(new_n10694), .Y(new_n10855));
  XNOR2x2_ASAP7_75t_L       g10599(.A(\a[29] ), .B(new_n10693), .Y(new_n10856));
  OAI211xp5_ASAP7_75t_L     g10600(.A1(new_n10503), .A2(new_n10689), .B(new_n10852), .C(new_n10853), .Y(new_n10857));
  OAI21xp33_ASAP7_75t_L     g10601(.A1(new_n10846), .A2(new_n10850), .B(new_n10697), .Y(new_n10858));
  AOI21xp33_ASAP7_75t_L     g10602(.A1(new_n10857), .A2(new_n10858), .B(new_n10856), .Y(new_n10859));
  NOR2xp33_ASAP7_75t_L      g10603(.A(new_n10859), .B(new_n10855), .Y(new_n10860));
  NAND2xp33_ASAP7_75t_L     g10604(.A(new_n10691), .B(new_n10860), .Y(new_n10861));
  AOI21xp33_ASAP7_75t_L     g10605(.A1(new_n10365), .A2(new_n10517), .B(new_n10690), .Y(new_n10862));
  NAND3xp33_ASAP7_75t_L     g10606(.A(new_n10857), .B(new_n10856), .C(new_n10858), .Y(new_n10863));
  OAI21xp33_ASAP7_75t_L     g10607(.A1(new_n10854), .A2(new_n10851), .B(new_n10694), .Y(new_n10864));
  NAND2xp33_ASAP7_75t_L     g10608(.A(new_n10863), .B(new_n10864), .Y(new_n10865));
  NAND2xp33_ASAP7_75t_L     g10609(.A(new_n10862), .B(new_n10865), .Y(new_n10866));
  NOR2xp33_ASAP7_75t_L      g10610(.A(new_n4101), .B(new_n2415), .Y(new_n10867));
  AOI221xp5_ASAP7_75t_L     g10611(.A1(\b[31] ), .A2(new_n2577), .B1(\b[32] ), .B2(new_n2421), .C(new_n10867), .Y(new_n10868));
  O2A1O1Ixp33_ASAP7_75t_L   g10612(.A1(new_n2425), .A2(new_n4108), .B(new_n10868), .C(new_n2413), .Y(new_n10869));
  OAI21xp33_ASAP7_75t_L     g10613(.A1(new_n2425), .A2(new_n4108), .B(new_n10868), .Y(new_n10870));
  NAND2xp33_ASAP7_75t_L     g10614(.A(new_n2413), .B(new_n10870), .Y(new_n10871));
  OAI21xp33_ASAP7_75t_L     g10615(.A1(new_n2413), .A2(new_n10869), .B(new_n10871), .Y(new_n10872));
  INVx1_ASAP7_75t_L         g10616(.A(new_n10872), .Y(new_n10873));
  NAND3xp33_ASAP7_75t_L     g10617(.A(new_n10861), .B(new_n10866), .C(new_n10873), .Y(new_n10874));
  NOR2xp33_ASAP7_75t_L      g10618(.A(new_n10862), .B(new_n10865), .Y(new_n10875));
  AOI221xp5_ASAP7_75t_L     g10619(.A1(new_n10365), .A2(new_n10517), .B1(new_n10863), .B2(new_n10864), .C(new_n10690), .Y(new_n10876));
  OAI21xp33_ASAP7_75t_L     g10620(.A1(new_n10876), .A2(new_n10875), .B(new_n10872), .Y(new_n10877));
  NAND3xp33_ASAP7_75t_L     g10621(.A(new_n10688), .B(new_n10874), .C(new_n10877), .Y(new_n10878));
  O2A1O1Ixp33_ASAP7_75t_L   g10622(.A1(new_n10196), .A2(new_n2413), .B(new_n10203), .C(new_n10353), .Y(new_n10879));
  NAND2xp33_ASAP7_75t_L     g10623(.A(new_n10200), .B(new_n10205), .Y(new_n10880));
  A2O1A1O1Ixp25_ASAP7_75t_L g10624(.A1(new_n10210), .A2(new_n10880), .B(new_n10879), .C(new_n10521), .D(new_n10529), .Y(new_n10881));
  NOR3xp33_ASAP7_75t_L      g10625(.A(new_n10875), .B(new_n10876), .C(new_n10872), .Y(new_n10882));
  AOI21xp33_ASAP7_75t_L     g10626(.A1(new_n10861), .A2(new_n10866), .B(new_n10873), .Y(new_n10883));
  OAI21xp33_ASAP7_75t_L     g10627(.A1(new_n10883), .A2(new_n10882), .B(new_n10881), .Y(new_n10884));
  OAI22xp33_ASAP7_75t_L     g10628(.A1(new_n2089), .A2(new_n4344), .B1(new_n4581), .B2(new_n1962), .Y(new_n10885));
  AOI221xp5_ASAP7_75t_L     g10629(.A1(new_n1955), .A2(\b[36] ), .B1(new_n1964), .B2(new_n4621), .C(new_n10885), .Y(new_n10886));
  XNOR2x2_ASAP7_75t_L       g10630(.A(new_n1952), .B(new_n10886), .Y(new_n10887));
  AOI21xp33_ASAP7_75t_L     g10631(.A1(new_n10878), .A2(new_n10884), .B(new_n10887), .Y(new_n10888));
  NOR3xp33_ASAP7_75t_L      g10632(.A(new_n10881), .B(new_n10882), .C(new_n10883), .Y(new_n10889));
  AOI221xp5_ASAP7_75t_L     g10633(.A1(new_n10354), .A2(new_n10521), .B1(new_n10877), .B2(new_n10874), .C(new_n10529), .Y(new_n10890));
  XNOR2x2_ASAP7_75t_L       g10634(.A(\a[23] ), .B(new_n10886), .Y(new_n10891));
  NOR3xp33_ASAP7_75t_L      g10635(.A(new_n10889), .B(new_n10890), .C(new_n10891), .Y(new_n10892));
  OAI221xp5_ASAP7_75t_L     g10636(.A1(new_n10888), .A2(new_n10892), .B1(new_n10546), .B2(new_n10552), .C(new_n10686), .Y(new_n10893));
  NOR2xp33_ASAP7_75t_L      g10637(.A(new_n10892), .B(new_n10888), .Y(new_n10894));
  A2O1A1Ixp33_ASAP7_75t_L   g10638(.A1(new_n10540), .A2(new_n10542), .B(new_n10544), .C(new_n10894), .Y(new_n10895));
  NOR2xp33_ASAP7_75t_L      g10639(.A(new_n5311), .B(new_n1517), .Y(new_n10896));
  AOI221xp5_ASAP7_75t_L     g10640(.A1(\b[37] ), .A2(new_n1659), .B1(\b[39] ), .B2(new_n1511), .C(new_n10896), .Y(new_n10897));
  O2A1O1Ixp33_ASAP7_75t_L   g10641(.A1(new_n1521), .A2(new_n5578), .B(new_n10897), .C(new_n1501), .Y(new_n10898));
  INVx1_ASAP7_75t_L         g10642(.A(new_n10898), .Y(new_n10899));
  O2A1O1Ixp33_ASAP7_75t_L   g10643(.A1(new_n1521), .A2(new_n5578), .B(new_n10897), .C(\a[20] ), .Y(new_n10900));
  AOI21xp33_ASAP7_75t_L     g10644(.A1(new_n10899), .A2(\a[20] ), .B(new_n10900), .Y(new_n10901));
  NAND3xp33_ASAP7_75t_L     g10645(.A(new_n10895), .B(new_n10893), .C(new_n10901), .Y(new_n10902));
  OAI21xp33_ASAP7_75t_L     g10646(.A1(new_n10890), .A2(new_n10889), .B(new_n10891), .Y(new_n10903));
  NAND3xp33_ASAP7_75t_L     g10647(.A(new_n10878), .B(new_n10884), .C(new_n10887), .Y(new_n10904));
  AOI221xp5_ASAP7_75t_L     g10648(.A1(new_n10904), .A2(new_n10903), .B1(new_n10540), .B2(new_n10542), .C(new_n10544), .Y(new_n10905));
  NAND2xp33_ASAP7_75t_L     g10649(.A(new_n10903), .B(new_n10904), .Y(new_n10906));
  O2A1O1Ixp33_ASAP7_75t_L   g10650(.A1(new_n10552), .A2(new_n10546), .B(new_n10686), .C(new_n10906), .Y(new_n10907));
  INVx1_ASAP7_75t_L         g10651(.A(new_n10901), .Y(new_n10908));
  OAI21xp33_ASAP7_75t_L     g10652(.A1(new_n10905), .A2(new_n10907), .B(new_n10908), .Y(new_n10909));
  AND4x1_ASAP7_75t_L        g10653(.A(new_n10572), .B(new_n10685), .C(new_n10909), .D(new_n10902), .Y(new_n10910));
  MAJIxp5_ASAP7_75t_L       g10654(.A(new_n10558), .B(new_n10550), .C(new_n10684), .Y(new_n10911));
  AOI21xp33_ASAP7_75t_L     g10655(.A1(new_n10909), .A2(new_n10902), .B(new_n10911), .Y(new_n10912));
  OAI22xp33_ASAP7_75t_L     g10656(.A1(new_n1285), .A2(new_n5855), .B1(new_n6110), .B2(new_n2118), .Y(new_n10913));
  AOI221xp5_ASAP7_75t_L     g10657(.A1(new_n1209), .A2(\b[42] ), .B1(new_n1216), .B2(new_n6389), .C(new_n10913), .Y(new_n10914));
  XNOR2x2_ASAP7_75t_L       g10658(.A(new_n1206), .B(new_n10914), .Y(new_n10915));
  OAI21xp33_ASAP7_75t_L     g10659(.A1(new_n10912), .A2(new_n10910), .B(new_n10915), .Y(new_n10916));
  NAND3xp33_ASAP7_75t_L     g10660(.A(new_n10911), .B(new_n10909), .C(new_n10902), .Y(new_n10917));
  INVx1_ASAP7_75t_L         g10661(.A(new_n10685), .Y(new_n10918));
  NAND2xp33_ASAP7_75t_L     g10662(.A(new_n10570), .B(new_n10569), .Y(new_n10919));
  NAND2xp33_ASAP7_75t_L     g10663(.A(new_n10909), .B(new_n10902), .Y(new_n10920));
  A2O1A1Ixp33_ASAP7_75t_L   g10664(.A1(new_n10919), .A2(new_n10558), .B(new_n10918), .C(new_n10920), .Y(new_n10921));
  XNOR2x2_ASAP7_75t_L       g10665(.A(\a[17] ), .B(new_n10914), .Y(new_n10922));
  NAND3xp33_ASAP7_75t_L     g10666(.A(new_n10921), .B(new_n10917), .C(new_n10922), .Y(new_n10923));
  NAND2xp33_ASAP7_75t_L     g10667(.A(new_n10923), .B(new_n10916), .Y(new_n10924));
  O2A1O1Ixp33_ASAP7_75t_L   g10668(.A1(new_n10575), .A2(new_n10577), .B(new_n10592), .C(new_n10924), .Y(new_n10925));
  AOI221xp5_ASAP7_75t_L     g10669(.A1(new_n10916), .A2(new_n10923), .B1(new_n10581), .B2(new_n10590), .C(new_n10593), .Y(new_n10926));
  OAI21xp33_ASAP7_75t_L     g10670(.A1(new_n10926), .A2(new_n10925), .B(new_n10683), .Y(new_n10927));
  INVx1_ASAP7_75t_L         g10671(.A(new_n10683), .Y(new_n10928));
  OAI21xp33_ASAP7_75t_L     g10672(.A1(new_n10577), .A2(new_n10575), .B(new_n10592), .Y(new_n10929));
  AOI21xp33_ASAP7_75t_L     g10673(.A1(new_n10921), .A2(new_n10917), .B(new_n10922), .Y(new_n10930));
  NOR3xp33_ASAP7_75t_L      g10674(.A(new_n10910), .B(new_n10912), .C(new_n10915), .Y(new_n10931));
  NOR2xp33_ASAP7_75t_L      g10675(.A(new_n10930), .B(new_n10931), .Y(new_n10932));
  NAND2xp33_ASAP7_75t_L     g10676(.A(new_n10932), .B(new_n10929), .Y(new_n10933));
  OAI221xp5_ASAP7_75t_L     g10677(.A1(new_n10575), .A2(new_n10577), .B1(new_n10930), .B2(new_n10931), .C(new_n10592), .Y(new_n10934));
  NAND3xp33_ASAP7_75t_L     g10678(.A(new_n10933), .B(new_n10928), .C(new_n10934), .Y(new_n10935));
  NAND2xp33_ASAP7_75t_L     g10679(.A(new_n10935), .B(new_n10927), .Y(new_n10936));
  AOI21xp33_ASAP7_75t_L     g10680(.A1(new_n10933), .A2(new_n10934), .B(new_n10928), .Y(new_n10937));
  NOR3xp33_ASAP7_75t_L      g10681(.A(new_n10925), .B(new_n10926), .C(new_n10683), .Y(new_n10938));
  NOR4xp25_ASAP7_75t_L      g10682(.A(new_n10601), .B(new_n10938), .C(new_n10937), .D(new_n10609), .Y(new_n10939));
  A2O1A1Ixp33_ASAP7_75t_L   g10683(.A1(new_n10671), .A2(new_n10936), .B(new_n10939), .C(new_n10677), .Y(new_n10940));
  INVx1_ASAP7_75t_L         g10684(.A(new_n10940), .Y(new_n10941));
  INVx1_ASAP7_75t_L         g10685(.A(new_n10677), .Y(new_n10942));
  OAI22xp33_ASAP7_75t_L     g10686(.A1(new_n10601), .A2(new_n10609), .B1(new_n10938), .B2(new_n10937), .Y(new_n10943));
  OAI211xp5_ASAP7_75t_L     g10687(.A1(new_n10274), .A2(new_n10600), .B(new_n10935), .C(new_n10589), .Y(new_n10944));
  OAI211xp5_ASAP7_75t_L     g10688(.A1(new_n10937), .A2(new_n10944), .B(new_n10943), .C(new_n10942), .Y(new_n10945));
  NAND2xp33_ASAP7_75t_L     g10689(.A(new_n10945), .B(new_n10940), .Y(new_n10946));
  A2O1A1Ixp33_ASAP7_75t_L   g10690(.A1(new_n10616), .A2(new_n10614), .B(new_n10607), .C(new_n10946), .Y(new_n10947));
  OAI211xp5_ASAP7_75t_L     g10691(.A1(new_n10352), .A2(new_n10625), .B(new_n10945), .C(new_n10621), .Y(new_n10948));
  O2A1O1Ixp33_ASAP7_75t_L   g10692(.A1(new_n10948), .A2(new_n10941), .B(new_n10947), .C(new_n10669), .Y(new_n10949));
  INVx1_ASAP7_75t_L         g10693(.A(new_n10949), .Y(new_n10950));
  AOI21xp33_ASAP7_75t_L     g10694(.A1(new_n10629), .A2(new_n10351), .B(new_n10630), .Y(new_n10951));
  MAJIxp5_ASAP7_75t_L       g10695(.A(new_n10352), .B(new_n10599), .C(new_n10606), .Y(new_n10952));
  O2A1O1Ixp33_ASAP7_75t_L   g10696(.A1(new_n10609), .A2(new_n10601), .B(new_n10936), .C(new_n10939), .Y(new_n10953));
  AOI221xp5_ASAP7_75t_L     g10697(.A1(new_n10942), .A2(new_n10953), .B1(new_n10614), .B2(new_n10616), .C(new_n10607), .Y(new_n10954));
  AOI221xp5_ASAP7_75t_L     g10698(.A1(new_n10952), .A2(new_n10946), .B1(new_n10940), .B2(new_n10954), .C(new_n10668), .Y(new_n10955));
  NOR2xp33_ASAP7_75t_L      g10699(.A(new_n10955), .B(new_n10949), .Y(new_n10956));
  O2A1O1Ixp33_ASAP7_75t_L   g10700(.A1(new_n10347), .A2(new_n10951), .B(new_n10629), .C(new_n10956), .Y(new_n10957));
  A2O1A1Ixp33_ASAP7_75t_L   g10701(.A1(new_n10618), .A2(new_n10627), .B(new_n10347), .C(new_n10629), .Y(new_n10958));
  NOR2xp33_ASAP7_75t_L      g10702(.A(new_n10955), .B(new_n10958), .Y(new_n10959));
  A2O1A1Ixp33_ASAP7_75t_L   g10703(.A1(new_n10959), .A2(new_n10950), .B(new_n10957), .C(new_n10662), .Y(new_n10960));
  OAI211xp5_ASAP7_75t_L     g10704(.A1(new_n10941), .A2(new_n10948), .B(new_n10947), .C(new_n10668), .Y(new_n10961));
  A2O1A1Ixp33_ASAP7_75t_L   g10705(.A1(new_n10668), .A2(new_n10961), .B(new_n10955), .C(new_n10958), .Y(new_n10962));
  OAI211xp5_ASAP7_75t_L     g10706(.A1(new_n10941), .A2(new_n10948), .B(new_n10947), .C(new_n10669), .Y(new_n10963));
  OAI211xp5_ASAP7_75t_L     g10707(.A1(new_n10347), .A2(new_n10951), .B(new_n10963), .C(new_n10629), .Y(new_n10964));
  OAI211xp5_ASAP7_75t_L     g10708(.A1(new_n10949), .A2(new_n10964), .B(new_n10962), .C(new_n10661), .Y(new_n10965));
  NAND3xp33_ASAP7_75t_L     g10709(.A(new_n10658), .B(new_n10960), .C(new_n10965), .Y(new_n10966));
  NOR2xp33_ASAP7_75t_L      g10710(.A(new_n10294), .B(new_n10345), .Y(new_n10967));
  NAND2xp33_ASAP7_75t_L     g10711(.A(new_n10295), .B(new_n10303), .Y(new_n10968));
  A2O1A1O1Ixp25_ASAP7_75t_L g10712(.A1(new_n10038), .A2(new_n10968), .B(new_n10967), .C(new_n10635), .D(new_n10645), .Y(new_n10969));
  O2A1O1Ixp33_ASAP7_75t_L   g10713(.A1(new_n10949), .A2(new_n10964), .B(new_n10962), .C(new_n10661), .Y(new_n10970));
  AOI221xp5_ASAP7_75t_L     g10714(.A1(new_n10952), .A2(new_n10946), .B1(new_n10940), .B2(new_n10954), .C(new_n10669), .Y(new_n10971));
  OAI21xp33_ASAP7_75t_L     g10715(.A1(new_n10669), .A2(new_n10971), .B(new_n10963), .Y(new_n10972));
  AOI221xp5_ASAP7_75t_L     g10716(.A1(new_n10958), .A2(new_n10972), .B1(new_n10950), .B2(new_n10959), .C(new_n10662), .Y(new_n10973));
  OAI21xp33_ASAP7_75t_L     g10717(.A1(new_n10970), .A2(new_n10973), .B(new_n10969), .Y(new_n10974));
  OAI211xp5_ASAP7_75t_L     g10718(.A1(new_n10949), .A2(new_n10964), .B(new_n10962), .C(new_n10662), .Y(new_n10975));
  A2O1A1Ixp33_ASAP7_75t_L   g10719(.A1(new_n10662), .A2(new_n10975), .B(new_n10973), .C(new_n10658), .Y(new_n10976));
  INVx1_ASAP7_75t_L         g10720(.A(new_n10976), .Y(new_n10977));
  INVx1_ASAP7_75t_L         g10721(.A(\b[57] ), .Y(new_n10978));
  NAND2xp33_ASAP7_75t_L     g10722(.A(\b[55] ), .B(new_n286), .Y(new_n10979));
  OAI221xp5_ASAP7_75t_L     g10723(.A1(new_n285), .A2(new_n10332), .B1(new_n10978), .B2(new_n269), .C(new_n10979), .Y(new_n10980));
  O2A1O1Ixp33_ASAP7_75t_L   g10724(.A1(new_n9709), .A2(new_n10309), .B(new_n10315), .C(new_n10337), .Y(new_n10981));
  NOR2xp33_ASAP7_75t_L      g10725(.A(\b[56] ), .B(\b[57] ), .Y(new_n10982));
  NOR2xp33_ASAP7_75t_L      g10726(.A(new_n10332), .B(new_n10978), .Y(new_n10983));
  NOR2xp33_ASAP7_75t_L      g10727(.A(new_n10982), .B(new_n10983), .Y(new_n10984));
  A2O1A1Ixp33_ASAP7_75t_L   g10728(.A1(\b[56] ), .A2(\b[55] ), .B(new_n10981), .C(new_n10984), .Y(new_n10985));
  INVx1_ASAP7_75t_L         g10729(.A(new_n10985), .Y(new_n10986));
  INVx1_ASAP7_75t_L         g10730(.A(new_n10313), .Y(new_n10987));
  INVx1_ASAP7_75t_L         g10731(.A(new_n10333), .Y(new_n10988));
  A2O1A1Ixp33_ASAP7_75t_L   g10732(.A1(new_n10315), .A2(new_n10987), .B(new_n10337), .C(new_n10988), .Y(new_n10989));
  NOR2xp33_ASAP7_75t_L      g10733(.A(new_n10984), .B(new_n10989), .Y(new_n10990));
  NOR2xp33_ASAP7_75t_L      g10734(.A(new_n10990), .B(new_n10986), .Y(new_n10991));
  A2O1A1Ixp33_ASAP7_75t_L   g10735(.A1(new_n10991), .A2(new_n273), .B(new_n10980), .C(\a[2] ), .Y(new_n10992));
  AOI211xp5_ASAP7_75t_L     g10736(.A1(new_n10991), .A2(new_n273), .B(new_n10980), .C(new_n257), .Y(new_n10993));
  A2O1A1O1Ixp25_ASAP7_75t_L g10737(.A1(new_n273), .A2(new_n10991), .B(new_n10980), .C(new_n10992), .D(new_n10993), .Y(new_n10994));
  O2A1O1Ixp33_ASAP7_75t_L   g10738(.A1(new_n10969), .A2(new_n10977), .B(new_n10974), .C(new_n10994), .Y(new_n10995));
  NAND2xp33_ASAP7_75t_L     g10739(.A(new_n10974), .B(new_n10966), .Y(new_n10996));
  INVx1_ASAP7_75t_L         g10740(.A(new_n10996), .Y(new_n10997));
  INVx1_ASAP7_75t_L         g10741(.A(new_n10994), .Y(new_n10998));
  NAND2xp33_ASAP7_75t_L     g10742(.A(new_n10998), .B(new_n10997), .Y(new_n10999));
  A2O1A1Ixp33_ASAP7_75t_L   g10743(.A1(new_n10974), .A2(new_n10966), .B(new_n10995), .C(new_n10999), .Y(new_n11000));
  A2O1A1Ixp33_ASAP7_75t_L   g10744(.A1(new_n10653), .A2(new_n10652), .B(new_n10648), .C(new_n11000), .Y(new_n11001));
  INVx1_ASAP7_75t_L         g10745(.A(new_n11001), .Y(new_n11002));
  A2O1A1Ixp33_ASAP7_75t_L   g10746(.A1(new_n10344), .A2(new_n10649), .B(new_n10650), .C(new_n10647), .Y(new_n11003));
  NOR2xp33_ASAP7_75t_L      g10747(.A(new_n11003), .B(new_n11000), .Y(new_n11004));
  NOR2xp33_ASAP7_75t_L      g10748(.A(new_n11004), .B(new_n11002), .Y(\f[57] ));
  A2O1A1Ixp33_ASAP7_75t_L   g10749(.A1(new_n10668), .A2(new_n10961), .B(new_n10964), .C(new_n10962), .Y(new_n11006));
  MAJIxp5_ASAP7_75t_L       g10750(.A(new_n10969), .B(new_n10661), .C(new_n11006), .Y(new_n11007));
  OAI22xp33_ASAP7_75t_L     g10751(.A1(new_n350), .A2(new_n9709), .B1(new_n9683), .B2(new_n375), .Y(new_n11008));
  AOI221xp5_ASAP7_75t_L     g10752(.A1(new_n361), .A2(\b[55] ), .B1(new_n359), .B2(new_n10320), .C(new_n11008), .Y(new_n11009));
  XNOR2x2_ASAP7_75t_L       g10753(.A(new_n346), .B(new_n11009), .Y(new_n11010));
  O2A1O1Ixp33_ASAP7_75t_L   g10754(.A1(new_n10955), .A2(new_n10668), .B(new_n10958), .C(new_n10971), .Y(new_n11011));
  OAI22xp33_ASAP7_75t_L     g10755(.A1(new_n513), .A2(new_n8779), .B1(new_n8755), .B2(new_n506), .Y(new_n11012));
  AOI221xp5_ASAP7_75t_L     g10756(.A1(new_n475), .A2(\b[52] ), .B1(new_n483), .B2(new_n9367), .C(new_n11012), .Y(new_n11013));
  XNOR2x2_ASAP7_75t_L       g10757(.A(new_n466), .B(new_n11013), .Y(new_n11014));
  INVx1_ASAP7_75t_L         g10758(.A(new_n11014), .Y(new_n11015));
  O2A1O1Ixp33_ASAP7_75t_L   g10759(.A1(new_n10622), .A2(new_n10619), .B(new_n10614), .C(new_n10607), .Y(new_n11016));
  NAND2xp33_ASAP7_75t_L     g10760(.A(new_n10677), .B(new_n10953), .Y(new_n11017));
  A2O1A1Ixp33_ASAP7_75t_L   g10761(.A1(new_n10945), .A2(new_n10942), .B(new_n11016), .C(new_n11017), .Y(new_n11018));
  OAI22xp33_ASAP7_75t_L     g10762(.A1(new_n1550), .A2(new_n7860), .B1(new_n7552), .B2(new_n712), .Y(new_n11019));
  AOI221xp5_ASAP7_75t_L     g10763(.A1(new_n640), .A2(\b[49] ), .B1(new_n718), .B2(new_n8438), .C(new_n11019), .Y(new_n11020));
  XNOR2x2_ASAP7_75t_L       g10764(.A(new_n637), .B(new_n11020), .Y(new_n11021));
  NAND3xp33_ASAP7_75t_L     g10765(.A(new_n10933), .B(new_n10683), .C(new_n10934), .Y(new_n11022));
  A2O1A1O1Ixp25_ASAP7_75t_L g10766(.A1(new_n10512), .A2(new_n10366), .B(new_n10503), .C(new_n10852), .D(new_n10850), .Y(new_n11023));
  OAI22xp33_ASAP7_75t_L     g10767(.A1(new_n7304), .A2(new_n1043), .B1(new_n960), .B2(new_n6741), .Y(new_n11024));
  AOI221xp5_ASAP7_75t_L     g10768(.A1(new_n6442), .A2(\b[16] ), .B1(new_n6450), .B2(new_n1156), .C(new_n11024), .Y(new_n11025));
  XNOR2x2_ASAP7_75t_L       g10769(.A(new_n6439), .B(new_n11025), .Y(new_n11026));
  OAI21xp33_ASAP7_75t_L     g10770(.A1(new_n10780), .A2(new_n10777), .B(new_n10726), .Y(new_n11027));
  A2O1A1O1Ixp25_ASAP7_75t_L g10771(.A1(new_n10442), .A2(new_n10452), .B(new_n10437), .C(new_n11027), .D(new_n10782), .Y(new_n11028));
  A2O1A1Ixp33_ASAP7_75t_L   g10772(.A1(new_n10757), .A2(new_n10756), .B(new_n10762), .C(new_n10763), .Y(new_n11029));
  NOR2xp33_ASAP7_75t_L      g10773(.A(new_n427), .B(new_n10400), .Y(new_n11030));
  AOI221xp5_ASAP7_75t_L     g10774(.A1(new_n9102), .A2(\b[7] ), .B1(new_n10398), .B2(\b[5] ), .C(new_n11030), .Y(new_n11031));
  O2A1O1Ixp33_ASAP7_75t_L   g10775(.A1(new_n9104), .A2(new_n456), .B(new_n11031), .C(new_n9099), .Y(new_n11032));
  OAI21xp33_ASAP7_75t_L     g10776(.A1(new_n9104), .A2(new_n456), .B(new_n11031), .Y(new_n11033));
  NAND2xp33_ASAP7_75t_L     g10777(.A(new_n9099), .B(new_n11033), .Y(new_n11034));
  OAI21xp33_ASAP7_75t_L     g10778(.A1(new_n9099), .A2(new_n11032), .B(new_n11034), .Y(new_n11035));
  INVx1_ASAP7_75t_L         g10779(.A(new_n11035), .Y(new_n11036));
  MAJIxp5_ASAP7_75t_L       g10780(.A(new_n10742), .B(new_n10397), .C(new_n10733), .Y(new_n11037));
  NAND2xp33_ASAP7_75t_L     g10781(.A(\b[4] ), .B(new_n10086), .Y(new_n11038));
  OAI221xp5_ASAP7_75t_L     g10782(.A1(new_n10388), .A2(new_n301), .B1(new_n289), .B2(new_n10390), .C(new_n11038), .Y(new_n11039));
  AOI211xp5_ASAP7_75t_L     g10783(.A1(new_n342), .A2(new_n10386), .B(new_n10083), .C(new_n11039), .Y(new_n11040));
  AOI21xp33_ASAP7_75t_L     g10784(.A1(new_n342), .A2(new_n10386), .B(new_n11039), .Y(new_n11041));
  NOR2xp33_ASAP7_75t_L      g10785(.A(\a[56] ), .B(new_n11041), .Y(new_n11042));
  NAND2xp33_ASAP7_75t_L     g10786(.A(new_n10731), .B(new_n10730), .Y(new_n11043));
  XNOR2x2_ASAP7_75t_L       g10787(.A(\a[58] ), .B(\a[57] ), .Y(new_n11044));
  NOR2xp33_ASAP7_75t_L      g10788(.A(new_n11044), .B(new_n11043), .Y(new_n11045));
  INVx1_ASAP7_75t_L         g10789(.A(\a[58] ), .Y(new_n11046));
  NAND2xp33_ASAP7_75t_L     g10790(.A(\a[59] ), .B(new_n11046), .Y(new_n11047));
  INVx1_ASAP7_75t_L         g10791(.A(\a[59] ), .Y(new_n11048));
  NAND2xp33_ASAP7_75t_L     g10792(.A(\a[58] ), .B(new_n11048), .Y(new_n11049));
  NAND2xp33_ASAP7_75t_L     g10793(.A(new_n11049), .B(new_n11047), .Y(new_n11050));
  NOR2xp33_ASAP7_75t_L      g10794(.A(new_n11050), .B(new_n10732), .Y(new_n11051));
  AOI22xp33_ASAP7_75t_L     g10795(.A1(new_n11045), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n11051), .Y(new_n11052));
  NAND2xp33_ASAP7_75t_L     g10796(.A(new_n11050), .B(new_n11043), .Y(new_n11053));
  OAI21xp33_ASAP7_75t_L     g10797(.A1(new_n11053), .A2(new_n274), .B(new_n11052), .Y(new_n11054));
  INVx1_ASAP7_75t_L         g10798(.A(new_n11054), .Y(new_n11055));
  NAND3xp33_ASAP7_75t_L     g10799(.A(new_n11055), .B(new_n10734), .C(\a[59] ), .Y(new_n11056));
  O2A1O1Ixp33_ASAP7_75t_L   g10800(.A1(new_n11053), .A2(new_n274), .B(new_n11052), .C(new_n11048), .Y(new_n11057));
  NAND2xp33_ASAP7_75t_L     g10801(.A(new_n11048), .B(new_n11054), .Y(new_n11058));
  A2O1A1Ixp33_ASAP7_75t_L   g10802(.A1(new_n10733), .A2(new_n11057), .B(new_n11048), .C(new_n11058), .Y(new_n11059));
  AOI211xp5_ASAP7_75t_L     g10803(.A1(new_n11059), .A2(new_n11056), .B(new_n11040), .C(new_n11042), .Y(new_n11060));
  OAI211xp5_ASAP7_75t_L     g10804(.A1(new_n11040), .A2(new_n11042), .B(new_n11056), .C(new_n11059), .Y(new_n11061));
  INVx1_ASAP7_75t_L         g10805(.A(new_n11061), .Y(new_n11062));
  NOR3xp33_ASAP7_75t_L      g10806(.A(new_n11062), .B(new_n11060), .C(new_n11037), .Y(new_n11063));
  MAJIxp5_ASAP7_75t_L       g10807(.A(new_n10748), .B(new_n10734), .C(new_n10411), .Y(new_n11064));
  A2O1A1Ixp33_ASAP7_75t_L   g10808(.A1(new_n342), .A2(new_n10386), .B(new_n11039), .C(\a[56] ), .Y(new_n11065));
  A2O1A1O1Ixp25_ASAP7_75t_L g10809(.A1(new_n10386), .A2(new_n342), .B(new_n11039), .C(new_n11065), .D(new_n11040), .Y(new_n11066));
  NAND2xp33_ASAP7_75t_L     g10810(.A(new_n11056), .B(new_n11059), .Y(new_n11067));
  NAND2xp33_ASAP7_75t_L     g10811(.A(new_n11066), .B(new_n11067), .Y(new_n11068));
  AOI21xp33_ASAP7_75t_L     g10812(.A1(new_n11068), .A2(new_n11061), .B(new_n11064), .Y(new_n11069));
  OAI21xp33_ASAP7_75t_L     g10813(.A1(new_n11069), .A2(new_n11063), .B(new_n11036), .Y(new_n11070));
  NAND3xp33_ASAP7_75t_L     g10814(.A(new_n11064), .B(new_n11068), .C(new_n11061), .Y(new_n11071));
  OAI21xp33_ASAP7_75t_L     g10815(.A1(new_n11060), .A2(new_n11062), .B(new_n11037), .Y(new_n11072));
  NAND3xp33_ASAP7_75t_L     g10816(.A(new_n11072), .B(new_n11071), .C(new_n11035), .Y(new_n11073));
  NAND3xp33_ASAP7_75t_L     g10817(.A(new_n11029), .B(new_n11070), .C(new_n11073), .Y(new_n11074));
  NOR2xp33_ASAP7_75t_L      g10818(.A(new_n10772), .B(new_n10764), .Y(new_n11075));
  AOI21xp33_ASAP7_75t_L     g10819(.A1(new_n11072), .A2(new_n11071), .B(new_n11035), .Y(new_n11076));
  NOR3xp33_ASAP7_75t_L      g10820(.A(new_n11063), .B(new_n11069), .C(new_n11036), .Y(new_n11077));
  OAI221xp5_ASAP7_75t_L     g10821(.A1(new_n11076), .A2(new_n11077), .B1(new_n10762), .B2(new_n11075), .C(new_n10763), .Y(new_n11078));
  OAI22xp33_ASAP7_75t_L     g10822(.A1(new_n8483), .A2(new_n534), .B1(new_n590), .B2(new_n10065), .Y(new_n11079));
  AOI221xp5_ASAP7_75t_L     g10823(.A1(new_n8175), .A2(\b[10] ), .B1(new_n8490), .B2(new_n690), .C(new_n11079), .Y(new_n11080));
  XNOR2x2_ASAP7_75t_L       g10824(.A(new_n8172), .B(new_n11080), .Y(new_n11081));
  NAND3xp33_ASAP7_75t_L     g10825(.A(new_n11078), .B(new_n11074), .C(new_n11081), .Y(new_n11082));
  AO21x2_ASAP7_75t_L        g10826(.A1(new_n11074), .A2(new_n11078), .B(new_n11081), .Y(new_n11083));
  A2O1A1O1Ixp25_ASAP7_75t_L g10827(.A1(new_n10426), .A2(new_n10383), .B(new_n10431), .C(new_n10779), .D(new_n10771), .Y(new_n11084));
  NAND3xp33_ASAP7_75t_L     g10828(.A(new_n11084), .B(new_n11083), .C(new_n11082), .Y(new_n11085));
  XNOR2x2_ASAP7_75t_L       g10829(.A(\a[50] ), .B(new_n11080), .Y(new_n11086));
  NAND3xp33_ASAP7_75t_L     g10830(.A(new_n11078), .B(new_n11074), .C(new_n11086), .Y(new_n11087));
  AND3x1_ASAP7_75t_L        g10831(.A(new_n11078), .B(new_n11074), .C(new_n11081), .Y(new_n11088));
  OAI21xp33_ASAP7_75t_L     g10832(.A1(new_n10776), .A2(new_n10727), .B(new_n10778), .Y(new_n11089));
  A2O1A1Ixp33_ASAP7_75t_L   g10833(.A1(new_n11087), .A2(new_n11086), .B(new_n11088), .C(new_n11089), .Y(new_n11090));
  OAI22xp33_ASAP7_75t_L     g10834(.A1(new_n7614), .A2(new_n748), .B1(new_n833), .B2(new_n7312), .Y(new_n11091));
  AOI221xp5_ASAP7_75t_L     g10835(.A1(new_n7334), .A2(\b[13] ), .B1(new_n7322), .B2(new_n1166), .C(new_n11091), .Y(new_n11092));
  XNOR2x2_ASAP7_75t_L       g10836(.A(\a[47] ), .B(new_n11092), .Y(new_n11093));
  NAND3xp33_ASAP7_75t_L     g10837(.A(new_n11093), .B(new_n11090), .C(new_n11085), .Y(new_n11094));
  INVx1_ASAP7_75t_L         g10838(.A(new_n10782), .Y(new_n11095));
  AOI21xp33_ASAP7_75t_L     g10839(.A1(new_n11090), .A2(new_n11085), .B(new_n11093), .Y(new_n11096));
  O2A1O1Ixp33_ASAP7_75t_L   g10840(.A1(new_n10781), .A2(new_n10785), .B(new_n11095), .C(new_n11096), .Y(new_n11097));
  AO21x2_ASAP7_75t_L        g10841(.A1(new_n11085), .A2(new_n11090), .B(new_n11093), .Y(new_n11098));
  NAND3xp33_ASAP7_75t_L     g10842(.A(new_n11028), .B(new_n11094), .C(new_n11098), .Y(new_n11099));
  A2O1A1O1Ixp25_ASAP7_75t_L g10843(.A1(new_n11094), .A2(new_n11097), .B(new_n11028), .C(new_n11099), .D(new_n11026), .Y(new_n11100));
  AOI21xp33_ASAP7_75t_L     g10844(.A1(new_n11098), .A2(new_n11094), .B(new_n11028), .Y(new_n11101));
  INVx1_ASAP7_75t_L         g10845(.A(new_n11094), .Y(new_n11102));
  O2A1O1Ixp33_ASAP7_75t_L   g10846(.A1(new_n10782), .A2(new_n10790), .B(new_n11098), .C(new_n11102), .Y(new_n11103));
  A2O1A1Ixp33_ASAP7_75t_L   g10847(.A1(new_n11103), .A2(new_n11098), .B(new_n11101), .C(new_n11026), .Y(new_n11104));
  OAI21xp33_ASAP7_75t_L     g10848(.A1(new_n11026), .A2(new_n11100), .B(new_n11104), .Y(new_n11105));
  A2O1A1Ixp33_ASAP7_75t_L   g10849(.A1(new_n10460), .A2(new_n10713), .B(new_n10802), .C(new_n10787), .Y(new_n11106));
  NOR2xp33_ASAP7_75t_L      g10850(.A(new_n11105), .B(new_n11106), .Y(new_n11107));
  AOI21xp33_ASAP7_75t_L     g10851(.A1(new_n10714), .A2(new_n10792), .B(new_n10796), .Y(new_n11108));
  O2A1O1Ixp33_ASAP7_75t_L   g10852(.A1(new_n11026), .A2(new_n11100), .B(new_n11104), .C(new_n11108), .Y(new_n11109));
  OAI22xp33_ASAP7_75t_L     g10853(.A1(new_n5640), .A2(new_n1458), .B1(new_n1349), .B2(new_n5925), .Y(new_n11110));
  AOI221xp5_ASAP7_75t_L     g10854(.A1(new_n5629), .A2(\b[19] ), .B1(new_n5637), .B2(new_n1607), .C(new_n11110), .Y(new_n11111));
  XNOR2x2_ASAP7_75t_L       g10855(.A(new_n5626), .B(new_n11111), .Y(new_n11112));
  OAI21xp33_ASAP7_75t_L     g10856(.A1(new_n11109), .A2(new_n11107), .B(new_n11112), .Y(new_n11113));
  A2O1A1O1Ixp25_ASAP7_75t_L g10857(.A1(new_n10370), .A2(new_n10463), .B(new_n10465), .C(new_n10801), .D(new_n10820), .Y(new_n11114));
  NOR3xp33_ASAP7_75t_L      g10858(.A(new_n11107), .B(new_n11109), .C(new_n11112), .Y(new_n11115));
  INVx1_ASAP7_75t_L         g10859(.A(new_n11115), .Y(new_n11116));
  AOI21xp33_ASAP7_75t_L     g10860(.A1(new_n11113), .A2(new_n11116), .B(new_n11114), .Y(new_n11117));
  A2O1A1O1Ixp25_ASAP7_75t_L g10861(.A1(new_n10801), .A2(new_n10706), .B(new_n10820), .C(new_n11113), .D(new_n11115), .Y(new_n11118));
  NAND2xp33_ASAP7_75t_L     g10862(.A(\b[21] ), .B(new_n4916), .Y(new_n11119));
  OAI221xp5_ASAP7_75t_L     g10863(.A1(new_n4908), .A2(new_n2045), .B1(new_n1745), .B2(new_n5144), .C(new_n11119), .Y(new_n11120));
  A2O1A1Ixp33_ASAP7_75t_L   g10864(.A1(new_n2056), .A2(new_n4912), .B(new_n11120), .C(\a[38] ), .Y(new_n11121));
  AOI211xp5_ASAP7_75t_L     g10865(.A1(new_n2056), .A2(new_n4912), .B(new_n11120), .C(new_n4906), .Y(new_n11122));
  A2O1A1O1Ixp25_ASAP7_75t_L g10866(.A1(new_n4912), .A2(new_n2056), .B(new_n11120), .C(new_n11121), .D(new_n11122), .Y(new_n11123));
  A2O1A1Ixp33_ASAP7_75t_L   g10867(.A1(new_n11118), .A2(new_n11113), .B(new_n11117), .C(new_n11123), .Y(new_n11124));
  A2O1A1Ixp33_ASAP7_75t_L   g10868(.A1(new_n10799), .A2(new_n10800), .B(new_n10807), .C(new_n10809), .Y(new_n11125));
  XNOR2x2_ASAP7_75t_L       g10869(.A(\a[44] ), .B(new_n11025), .Y(new_n11126));
  A2O1A1Ixp33_ASAP7_75t_L   g10870(.A1(new_n11103), .A2(new_n11098), .B(new_n11101), .C(new_n11126), .Y(new_n11127));
  A2O1A1O1Ixp25_ASAP7_75t_L g10871(.A1(new_n11094), .A2(new_n11097), .B(new_n11028), .C(new_n11099), .D(new_n11126), .Y(new_n11128));
  AOI21xp33_ASAP7_75t_L     g10872(.A1(new_n11127), .A2(new_n11126), .B(new_n11128), .Y(new_n11129));
  NAND2xp33_ASAP7_75t_L     g10873(.A(new_n11108), .B(new_n11129), .Y(new_n11130));
  A2O1A1Ixp33_ASAP7_75t_L   g10874(.A1(new_n10792), .A2(new_n10714), .B(new_n10796), .C(new_n11105), .Y(new_n11131));
  XNOR2x2_ASAP7_75t_L       g10875(.A(\a[41] ), .B(new_n11111), .Y(new_n11132));
  AOI21xp33_ASAP7_75t_L     g10876(.A1(new_n11131), .A2(new_n11130), .B(new_n11132), .Y(new_n11133));
  OAI21xp33_ASAP7_75t_L     g10877(.A1(new_n11115), .A2(new_n11133), .B(new_n11125), .Y(new_n11134));
  NAND3xp33_ASAP7_75t_L     g10878(.A(new_n11114), .B(new_n11116), .C(new_n11113), .Y(new_n11135));
  INVx1_ASAP7_75t_L         g10879(.A(new_n11123), .Y(new_n11136));
  NAND3xp33_ASAP7_75t_L     g10880(.A(new_n11135), .B(new_n11134), .C(new_n11136), .Y(new_n11137));
  A2O1A1O1Ixp25_ASAP7_75t_L g10881(.A1(new_n10481), .A2(new_n10699), .B(new_n10700), .C(new_n10822), .D(new_n10805), .Y(new_n11138));
  NAND3xp33_ASAP7_75t_L     g10882(.A(new_n11138), .B(new_n11137), .C(new_n11124), .Y(new_n11139));
  O2A1O1Ixp33_ASAP7_75t_L   g10883(.A1(new_n10807), .A2(new_n10811), .B(new_n10809), .C(new_n11133), .Y(new_n11140));
  A2O1A1Ixp33_ASAP7_75t_L   g10884(.A1(new_n11116), .A2(new_n11140), .B(new_n11114), .C(new_n11135), .Y(new_n11141));
  A2O1A1Ixp33_ASAP7_75t_L   g10885(.A1(new_n11118), .A2(new_n11113), .B(new_n11117), .C(new_n11136), .Y(new_n11142));
  NOR3xp33_ASAP7_75t_L      g10886(.A(new_n11125), .B(new_n11115), .C(new_n11133), .Y(new_n11143));
  NOR3xp33_ASAP7_75t_L      g10887(.A(new_n11117), .B(new_n11143), .C(new_n11123), .Y(new_n11144));
  A2O1A1Ixp33_ASAP7_75t_L   g10888(.A1(new_n10818), .A2(new_n10492), .B(new_n10813), .C(new_n10819), .Y(new_n11145));
  A2O1A1Ixp33_ASAP7_75t_L   g10889(.A1(new_n11142), .A2(new_n11141), .B(new_n11144), .C(new_n11145), .Y(new_n11146));
  OAI22xp33_ASAP7_75t_L     g10890(.A1(new_n4397), .A2(new_n2188), .B1(new_n2205), .B2(new_n4142), .Y(new_n11147));
  AOI221xp5_ASAP7_75t_L     g10891(.A1(new_n4156), .A2(\b[25] ), .B1(new_n4151), .B2(new_n5001), .C(new_n11147), .Y(new_n11148));
  XNOR2x2_ASAP7_75t_L       g10892(.A(new_n4145), .B(new_n11148), .Y(new_n11149));
  NAND3xp33_ASAP7_75t_L     g10893(.A(new_n11139), .B(new_n11146), .C(new_n11149), .Y(new_n11150));
  A2O1A1O1Ixp25_ASAP7_75t_L g10894(.A1(new_n11116), .A2(new_n11140), .B(new_n11114), .C(new_n11135), .D(new_n11136), .Y(new_n11151));
  NOR3xp33_ASAP7_75t_L      g10895(.A(new_n11145), .B(new_n11151), .C(new_n11144), .Y(new_n11152));
  AOI21xp33_ASAP7_75t_L     g10896(.A1(new_n11137), .A2(new_n11124), .B(new_n11138), .Y(new_n11153));
  INVx1_ASAP7_75t_L         g10897(.A(new_n11149), .Y(new_n11154));
  OAI21xp33_ASAP7_75t_L     g10898(.A1(new_n11152), .A2(new_n11153), .B(new_n11154), .Y(new_n11155));
  NAND2xp33_ASAP7_75t_L     g10899(.A(new_n11150), .B(new_n11155), .Y(new_n11156));
  NOR2xp33_ASAP7_75t_L      g10900(.A(new_n10832), .B(new_n10830), .Y(new_n11157));
  NAND2xp33_ASAP7_75t_L     g10901(.A(new_n10833), .B(new_n11157), .Y(new_n11158));
  A2O1A1Ixp33_ASAP7_75t_L   g10902(.A1(new_n10827), .A2(new_n10828), .B(new_n10837), .C(new_n11158), .Y(new_n11159));
  NOR2xp33_ASAP7_75t_L      g10903(.A(new_n11159), .B(new_n11156), .Y(new_n11160));
  NAND3xp33_ASAP7_75t_L     g10904(.A(new_n11154), .B(new_n11139), .C(new_n11146), .Y(new_n11161));
  INVx1_ASAP7_75t_L         g10905(.A(new_n11161), .Y(new_n11162));
  MAJIxp5_ASAP7_75t_L       g10906(.A(new_n10841), .B(new_n10833), .C(new_n11157), .Y(new_n11163));
  O2A1O1Ixp33_ASAP7_75t_L   g10907(.A1(new_n11149), .A2(new_n11162), .B(new_n11150), .C(new_n11163), .Y(new_n11164));
  NOR2xp33_ASAP7_75t_L      g10908(.A(new_n3079), .B(new_n3510), .Y(new_n11165));
  AOI221xp5_ASAP7_75t_L     g10909(.A1(\b[26] ), .A2(new_n3708), .B1(\b[27] ), .B2(new_n3499), .C(new_n11165), .Y(new_n11166));
  O2A1O1Ixp33_ASAP7_75t_L   g10910(.A1(new_n3513), .A2(new_n3087), .B(new_n11166), .C(new_n3493), .Y(new_n11167));
  OAI21xp33_ASAP7_75t_L     g10911(.A1(new_n3513), .A2(new_n3087), .B(new_n11166), .Y(new_n11168));
  NAND2xp33_ASAP7_75t_L     g10912(.A(new_n3493), .B(new_n11168), .Y(new_n11169));
  OAI21xp33_ASAP7_75t_L     g10913(.A1(new_n3493), .A2(new_n11167), .B(new_n11169), .Y(new_n11170));
  NOR3xp33_ASAP7_75t_L      g10914(.A(new_n11164), .B(new_n11160), .C(new_n11170), .Y(new_n11171));
  NOR2xp33_ASAP7_75t_L      g10915(.A(new_n11152), .B(new_n11153), .Y(new_n11172));
  AOI21xp33_ASAP7_75t_L     g10916(.A1(new_n11139), .A2(new_n11146), .B(new_n11149), .Y(new_n11173));
  AOI21xp33_ASAP7_75t_L     g10917(.A1(new_n11161), .A2(new_n11172), .B(new_n11173), .Y(new_n11174));
  NAND2xp33_ASAP7_75t_L     g10918(.A(new_n11163), .B(new_n11174), .Y(new_n11175));
  NAND2xp33_ASAP7_75t_L     g10919(.A(new_n11159), .B(new_n11156), .Y(new_n11176));
  INVx1_ASAP7_75t_L         g10920(.A(new_n11170), .Y(new_n11177));
  AOI21xp33_ASAP7_75t_L     g10921(.A1(new_n11175), .A2(new_n11176), .B(new_n11177), .Y(new_n11178));
  NOR3xp33_ASAP7_75t_L      g10922(.A(new_n11023), .B(new_n11171), .C(new_n11178), .Y(new_n11179));
  A2O1A1Ixp33_ASAP7_75t_L   g10923(.A1(new_n10696), .A2(new_n10181), .B(new_n10509), .C(new_n10512), .Y(new_n11180));
  A2O1A1Ixp33_ASAP7_75t_L   g10924(.A1(new_n11180), .A2(new_n10511), .B(new_n10846), .C(new_n10853), .Y(new_n11181));
  NAND3xp33_ASAP7_75t_L     g10925(.A(new_n11175), .B(new_n11176), .C(new_n11177), .Y(new_n11182));
  OAI21xp33_ASAP7_75t_L     g10926(.A1(new_n11160), .A2(new_n11164), .B(new_n11170), .Y(new_n11183));
  AOI21xp33_ASAP7_75t_L     g10927(.A1(new_n11183), .A2(new_n11182), .B(new_n11181), .Y(new_n11184));
  OAI22xp33_ASAP7_75t_L     g10928(.A1(new_n3133), .A2(new_n3098), .B1(new_n3456), .B2(new_n2925), .Y(new_n11185));
  AOI221xp5_ASAP7_75t_L     g10929(.A1(new_n2938), .A2(\b[31] ), .B1(new_n2932), .B2(new_n4317), .C(new_n11185), .Y(new_n11186));
  XNOR2x2_ASAP7_75t_L       g10930(.A(\a[29] ), .B(new_n11186), .Y(new_n11187));
  OAI21xp33_ASAP7_75t_L     g10931(.A1(new_n11184), .A2(new_n11179), .B(new_n11187), .Y(new_n11188));
  NAND3xp33_ASAP7_75t_L     g10932(.A(new_n11181), .B(new_n11182), .C(new_n11183), .Y(new_n11189));
  NAND3xp33_ASAP7_75t_L     g10933(.A(new_n11175), .B(new_n11176), .C(new_n11170), .Y(new_n11190));
  A2O1A1Ixp33_ASAP7_75t_L   g10934(.A1(new_n11170), .A2(new_n11190), .B(new_n11171), .C(new_n11023), .Y(new_n11191));
  XNOR2x2_ASAP7_75t_L       g10935(.A(new_n2928), .B(new_n11186), .Y(new_n11192));
  NAND3xp33_ASAP7_75t_L     g10936(.A(new_n11192), .B(new_n11191), .C(new_n11189), .Y(new_n11193));
  AOI221xp5_ASAP7_75t_L     g10937(.A1(new_n10691), .A2(new_n10864), .B1(new_n11188), .B2(new_n11193), .C(new_n10855), .Y(new_n11194));
  A2O1A1O1Ixp25_ASAP7_75t_L g10938(.A1(new_n10517), .A2(new_n10365), .B(new_n10690), .C(new_n10864), .D(new_n10855), .Y(new_n11195));
  AOI21xp33_ASAP7_75t_L     g10939(.A1(new_n11189), .A2(new_n11191), .B(new_n11192), .Y(new_n11196));
  NOR3xp33_ASAP7_75t_L      g10940(.A(new_n11187), .B(new_n11184), .C(new_n11179), .Y(new_n11197));
  NOR3xp33_ASAP7_75t_L      g10941(.A(new_n11195), .B(new_n11197), .C(new_n11196), .Y(new_n11198));
  OAI22xp33_ASAP7_75t_L     g10942(.A1(new_n2572), .A2(new_n3891), .B1(new_n4101), .B2(new_n2410), .Y(new_n11199));
  AOI221xp5_ASAP7_75t_L     g10943(.A1(new_n2423), .A2(\b[34] ), .B1(new_n2417), .B2(new_n5599), .C(new_n11199), .Y(new_n11200));
  XNOR2x2_ASAP7_75t_L       g10944(.A(\a[26] ), .B(new_n11200), .Y(new_n11201));
  NOR3xp33_ASAP7_75t_L      g10945(.A(new_n11201), .B(new_n11194), .C(new_n11198), .Y(new_n11202));
  OA21x2_ASAP7_75t_L        g10946(.A1(new_n11198), .A2(new_n11194), .B(new_n11201), .Y(new_n11203));
  NOR2xp33_ASAP7_75t_L      g10947(.A(new_n11202), .B(new_n11203), .Y(new_n11204));
  NAND2xp33_ASAP7_75t_L     g10948(.A(new_n10866), .B(new_n10861), .Y(new_n11205));
  MAJx2_ASAP7_75t_L         g10949(.A(new_n10881), .B(new_n11205), .C(new_n10873), .Y(new_n11206));
  NAND2xp33_ASAP7_75t_L     g10950(.A(new_n11206), .B(new_n11204), .Y(new_n11207));
  NOR2xp33_ASAP7_75t_L      g10951(.A(new_n11198), .B(new_n11194), .Y(new_n11208));
  NAND2xp33_ASAP7_75t_L     g10952(.A(new_n11201), .B(new_n11208), .Y(new_n11209));
  MAJIxp5_ASAP7_75t_L       g10953(.A(new_n10881), .B(new_n10873), .C(new_n11205), .Y(new_n11210));
  A2O1A1Ixp33_ASAP7_75t_L   g10954(.A1(new_n11209), .A2(new_n11208), .B(new_n11203), .C(new_n11210), .Y(new_n11211));
  OAI22xp33_ASAP7_75t_L     g10955(.A1(new_n2089), .A2(new_n4581), .B1(new_n4613), .B2(new_n1962), .Y(new_n11212));
  AOI221xp5_ASAP7_75t_L     g10956(.A1(new_n1955), .A2(\b[37] ), .B1(new_n1964), .B2(new_n10229), .C(new_n11212), .Y(new_n11213));
  XNOR2x2_ASAP7_75t_L       g10957(.A(new_n1952), .B(new_n11213), .Y(new_n11214));
  NAND3xp33_ASAP7_75t_L     g10958(.A(new_n11207), .B(new_n11211), .C(new_n11214), .Y(new_n11215));
  AO21x2_ASAP7_75t_L        g10959(.A1(new_n11211), .A2(new_n11207), .B(new_n11214), .Y(new_n11216));
  A2O1A1O1Ixp25_ASAP7_75t_L g10960(.A1(new_n10540), .A2(new_n10542), .B(new_n10544), .C(new_n10904), .D(new_n10888), .Y(new_n11217));
  NAND3xp33_ASAP7_75t_L     g10961(.A(new_n11217), .B(new_n11216), .C(new_n11215), .Y(new_n11218));
  AO21x2_ASAP7_75t_L        g10962(.A1(new_n11215), .A2(new_n11216), .B(new_n11217), .Y(new_n11219));
  NOR2xp33_ASAP7_75t_L      g10963(.A(new_n5570), .B(new_n1517), .Y(new_n11220));
  AOI221xp5_ASAP7_75t_L     g10964(.A1(\b[38] ), .A2(new_n1659), .B1(\b[40] ), .B2(new_n1511), .C(new_n11220), .Y(new_n11221));
  O2A1O1Ixp33_ASAP7_75t_L   g10965(.A1(new_n1521), .A2(new_n5862), .B(new_n11221), .C(new_n1501), .Y(new_n11222));
  INVx1_ASAP7_75t_L         g10966(.A(new_n11221), .Y(new_n11223));
  A2O1A1Ixp33_ASAP7_75t_L   g10967(.A1(new_n6651), .A2(new_n1513), .B(new_n11223), .C(new_n1501), .Y(new_n11224));
  OAI21xp33_ASAP7_75t_L     g10968(.A1(new_n1501), .A2(new_n11222), .B(new_n11224), .Y(new_n11225));
  INVx1_ASAP7_75t_L         g10969(.A(new_n11225), .Y(new_n11226));
  NAND3xp33_ASAP7_75t_L     g10970(.A(new_n11219), .B(new_n11218), .C(new_n11226), .Y(new_n11227));
  AND3x1_ASAP7_75t_L        g10971(.A(new_n11217), .B(new_n11216), .C(new_n11215), .Y(new_n11228));
  AOI21xp33_ASAP7_75t_L     g10972(.A1(new_n11216), .A2(new_n11215), .B(new_n11217), .Y(new_n11229));
  OAI21xp33_ASAP7_75t_L     g10973(.A1(new_n11229), .A2(new_n11228), .B(new_n11225), .Y(new_n11230));
  NAND2xp33_ASAP7_75t_L     g10974(.A(new_n11227), .B(new_n11230), .Y(new_n11231));
  NOR2xp33_ASAP7_75t_L      g10975(.A(new_n10905), .B(new_n10907), .Y(new_n11232));
  A2O1A1Ixp33_ASAP7_75t_L   g10976(.A1(\a[20] ), .A2(new_n10899), .B(new_n10900), .C(new_n11232), .Y(new_n11233));
  A2O1A1Ixp33_ASAP7_75t_L   g10977(.A1(new_n10902), .A2(new_n10909), .B(new_n10911), .C(new_n11233), .Y(new_n11234));
  NOR2xp33_ASAP7_75t_L      g10978(.A(new_n11231), .B(new_n11234), .Y(new_n11235));
  NAND2xp33_ASAP7_75t_L     g10979(.A(new_n10893), .B(new_n10895), .Y(new_n11236));
  NAND3xp33_ASAP7_75t_L     g10980(.A(new_n11219), .B(new_n11218), .C(new_n11225), .Y(new_n11237));
  NOR3xp33_ASAP7_75t_L      g10981(.A(new_n11228), .B(new_n11229), .C(new_n11225), .Y(new_n11238));
  AOI21xp33_ASAP7_75t_L     g10982(.A1(new_n11237), .A2(new_n11225), .B(new_n11238), .Y(new_n11239));
  O2A1O1Ixp33_ASAP7_75t_L   g10983(.A1(new_n11236), .A2(new_n10901), .B(new_n10921), .C(new_n11239), .Y(new_n11240));
  OAI22xp33_ASAP7_75t_L     g10984(.A1(new_n1285), .A2(new_n6110), .B1(new_n6378), .B2(new_n2118), .Y(new_n11241));
  AOI221xp5_ASAP7_75t_L     g10985(.A1(new_n1209), .A2(\b[43] ), .B1(new_n1216), .B2(new_n6682), .C(new_n11241), .Y(new_n11242));
  XNOR2x2_ASAP7_75t_L       g10986(.A(new_n1206), .B(new_n11242), .Y(new_n11243));
  OAI21xp33_ASAP7_75t_L     g10987(.A1(new_n11235), .A2(new_n11240), .B(new_n11243), .Y(new_n11244));
  A2O1A1O1Ixp25_ASAP7_75t_L g10988(.A1(new_n10581), .A2(new_n10590), .B(new_n10593), .C(new_n10916), .D(new_n10931), .Y(new_n11245));
  INVx1_ASAP7_75t_L         g10989(.A(new_n10900), .Y(new_n11246));
  O2A1O1Ixp33_ASAP7_75t_L   g10990(.A1(new_n10898), .A2(new_n1501), .B(new_n11246), .C(new_n11236), .Y(new_n11247));
  A2O1A1O1Ixp25_ASAP7_75t_L g10991(.A1(new_n10919), .A2(new_n10558), .B(new_n10918), .C(new_n10920), .D(new_n11247), .Y(new_n11248));
  NAND2xp33_ASAP7_75t_L     g10992(.A(new_n11239), .B(new_n11248), .Y(new_n11249));
  NAND2xp33_ASAP7_75t_L     g10993(.A(new_n11231), .B(new_n11234), .Y(new_n11250));
  INVx1_ASAP7_75t_L         g10994(.A(new_n11243), .Y(new_n11251));
  NAND3xp33_ASAP7_75t_L     g10995(.A(new_n11251), .B(new_n11249), .C(new_n11250), .Y(new_n11252));
  AOI21xp33_ASAP7_75t_L     g10996(.A1(new_n11252), .A2(new_n11244), .B(new_n11245), .Y(new_n11253));
  NOR3xp33_ASAP7_75t_L      g10997(.A(new_n11240), .B(new_n11243), .C(new_n11235), .Y(new_n11254));
  A2O1A1O1Ixp25_ASAP7_75t_L g10998(.A1(new_n10932), .A2(new_n10929), .B(new_n10931), .C(new_n11244), .D(new_n11254), .Y(new_n11255));
  OAI22xp33_ASAP7_75t_L     g10999(.A1(new_n980), .A2(new_n6944), .B1(new_n7249), .B2(new_n864), .Y(new_n11256));
  AOI221xp5_ASAP7_75t_L     g11000(.A1(new_n886), .A2(\b[46] ), .B1(new_n873), .B2(new_n7278), .C(new_n11256), .Y(new_n11257));
  XNOR2x2_ASAP7_75t_L       g11001(.A(new_n867), .B(new_n11257), .Y(new_n11258));
  INVx1_ASAP7_75t_L         g11002(.A(new_n11258), .Y(new_n11259));
  AOI211xp5_ASAP7_75t_L     g11003(.A1(new_n11255), .A2(new_n11244), .B(new_n11259), .C(new_n11253), .Y(new_n11260));
  AOI21xp33_ASAP7_75t_L     g11004(.A1(new_n11249), .A2(new_n11250), .B(new_n11251), .Y(new_n11261));
  AO21x2_ASAP7_75t_L        g11005(.A1(new_n11244), .A2(new_n11252), .B(new_n11245), .Y(new_n11262));
  OAI21xp33_ASAP7_75t_L     g11006(.A1(new_n11261), .A2(new_n11245), .B(new_n11252), .Y(new_n11263));
  O2A1O1Ixp33_ASAP7_75t_L   g11007(.A1(new_n11261), .A2(new_n11263), .B(new_n11262), .C(new_n11258), .Y(new_n11264));
  AOI211xp5_ASAP7_75t_L     g11008(.A1(new_n10943), .A2(new_n11022), .B(new_n11260), .C(new_n11264), .Y(new_n11265));
  INVx1_ASAP7_75t_L         g11009(.A(new_n11022), .Y(new_n11266));
  OAI211xp5_ASAP7_75t_L     g11010(.A1(new_n11261), .A2(new_n11263), .B(new_n11262), .C(new_n11258), .Y(new_n11267));
  A2O1A1Ixp33_ASAP7_75t_L   g11011(.A1(new_n11255), .A2(new_n11244), .B(new_n11253), .C(new_n11259), .Y(new_n11268));
  AOI221xp5_ASAP7_75t_L     g11012(.A1(new_n10936), .A2(new_n10671), .B1(new_n11268), .B2(new_n11267), .C(new_n11266), .Y(new_n11269));
  OAI21xp33_ASAP7_75t_L     g11013(.A1(new_n11269), .A2(new_n11265), .B(new_n11021), .Y(new_n11270));
  INVx1_ASAP7_75t_L         g11014(.A(new_n11021), .Y(new_n11271));
  A2O1A1Ixp33_ASAP7_75t_L   g11015(.A1(new_n10927), .A2(new_n10935), .B(new_n10620), .C(new_n11022), .Y(new_n11272));
  NAND3xp33_ASAP7_75t_L     g11016(.A(new_n11272), .B(new_n11267), .C(new_n11268), .Y(new_n11273));
  O2A1O1Ixp33_ASAP7_75t_L   g11017(.A1(new_n10937), .A2(new_n10938), .B(new_n10671), .C(new_n11266), .Y(new_n11274));
  OAI21xp33_ASAP7_75t_L     g11018(.A1(new_n11260), .A2(new_n11264), .B(new_n11274), .Y(new_n11275));
  NAND3xp33_ASAP7_75t_L     g11019(.A(new_n11273), .B(new_n11271), .C(new_n11275), .Y(new_n11276));
  NAND3xp33_ASAP7_75t_L     g11020(.A(new_n11018), .B(new_n11270), .C(new_n11276), .Y(new_n11277));
  A2O1A1Ixp33_ASAP7_75t_L   g11021(.A1(new_n10683), .A2(new_n11022), .B(new_n10944), .C(new_n10943), .Y(new_n11278));
  O2A1O1Ixp33_ASAP7_75t_L   g11022(.A1(new_n637), .A2(new_n10674), .B(new_n10676), .C(new_n11278), .Y(new_n11279));
  O2A1O1Ixp33_ASAP7_75t_L   g11023(.A1(new_n10953), .A2(new_n10941), .B(new_n10952), .C(new_n11279), .Y(new_n11280));
  NAND2xp33_ASAP7_75t_L     g11024(.A(new_n11270), .B(new_n11276), .Y(new_n11281));
  NAND2xp33_ASAP7_75t_L     g11025(.A(new_n11280), .B(new_n11281), .Y(new_n11282));
  AOI21xp33_ASAP7_75t_L     g11026(.A1(new_n11277), .A2(new_n11282), .B(new_n11015), .Y(new_n11283));
  O2A1O1Ixp33_ASAP7_75t_L   g11027(.A1(new_n10942), .A2(new_n11278), .B(new_n10947), .C(new_n11281), .Y(new_n11284));
  AOI21xp33_ASAP7_75t_L     g11028(.A1(new_n11276), .A2(new_n11270), .B(new_n11018), .Y(new_n11285));
  NOR3xp33_ASAP7_75t_L      g11029(.A(new_n11284), .B(new_n11285), .C(new_n11014), .Y(new_n11286));
  NOR3xp33_ASAP7_75t_L      g11030(.A(new_n11011), .B(new_n11283), .C(new_n11286), .Y(new_n11287));
  OAI21xp33_ASAP7_75t_L     g11031(.A1(new_n11285), .A2(new_n11284), .B(new_n11014), .Y(new_n11288));
  NAND3xp33_ASAP7_75t_L     g11032(.A(new_n11277), .B(new_n11282), .C(new_n11015), .Y(new_n11289));
  AOI221xp5_ASAP7_75t_L     g11033(.A1(new_n10972), .A2(new_n10958), .B1(new_n11289), .B2(new_n11288), .C(new_n10971), .Y(new_n11290));
  OAI21xp33_ASAP7_75t_L     g11034(.A1(new_n11290), .A2(new_n11287), .B(new_n11010), .Y(new_n11291));
  INVx1_ASAP7_75t_L         g11035(.A(new_n11010), .Y(new_n11292));
  A2O1A1Ixp33_ASAP7_75t_L   g11036(.A1(new_n10637), .A2(new_n10629), .B(new_n10956), .C(new_n10961), .Y(new_n11293));
  NAND3xp33_ASAP7_75t_L     g11037(.A(new_n11293), .B(new_n11288), .C(new_n11289), .Y(new_n11294));
  OAI21xp33_ASAP7_75t_L     g11038(.A1(new_n11283), .A2(new_n11286), .B(new_n11011), .Y(new_n11295));
  NAND3xp33_ASAP7_75t_L     g11039(.A(new_n11294), .B(new_n11292), .C(new_n11295), .Y(new_n11296));
  NAND3xp33_ASAP7_75t_L     g11040(.A(new_n11007), .B(new_n11291), .C(new_n11296), .Y(new_n11297));
  NOR2xp33_ASAP7_75t_L      g11041(.A(new_n10970), .B(new_n10973), .Y(new_n11298));
  AOI21xp33_ASAP7_75t_L     g11042(.A1(new_n11294), .A2(new_n11295), .B(new_n11292), .Y(new_n11299));
  NOR3xp33_ASAP7_75t_L      g11043(.A(new_n11287), .B(new_n11290), .C(new_n11010), .Y(new_n11300));
  OAI221xp5_ASAP7_75t_L     g11044(.A1(new_n11298), .A2(new_n10969), .B1(new_n11300), .B2(new_n11299), .C(new_n10975), .Y(new_n11301));
  NAND2xp33_ASAP7_75t_L     g11045(.A(new_n11301), .B(new_n11297), .Y(new_n11302));
  INVx1_ASAP7_75t_L         g11046(.A(\b[58] ), .Y(new_n11303));
  NAND2xp33_ASAP7_75t_L     g11047(.A(\b[56] ), .B(new_n286), .Y(new_n11304));
  OAI221xp5_ASAP7_75t_L     g11048(.A1(new_n285), .A2(new_n10978), .B1(new_n11303), .B2(new_n269), .C(new_n11304), .Y(new_n11305));
  INVx1_ASAP7_75t_L         g11049(.A(new_n10983), .Y(new_n11306));
  NOR2xp33_ASAP7_75t_L      g11050(.A(\b[57] ), .B(\b[58] ), .Y(new_n11307));
  NOR2xp33_ASAP7_75t_L      g11051(.A(new_n10978), .B(new_n11303), .Y(new_n11308));
  NOR2xp33_ASAP7_75t_L      g11052(.A(new_n11307), .B(new_n11308), .Y(new_n11309));
  INVx1_ASAP7_75t_L         g11053(.A(new_n11309), .Y(new_n11310));
  A2O1A1O1Ixp25_ASAP7_75t_L g11054(.A1(new_n10988), .A2(new_n10335), .B(new_n10982), .C(new_n11306), .D(new_n11310), .Y(new_n11311));
  A2O1A1Ixp33_ASAP7_75t_L   g11055(.A1(new_n10335), .A2(new_n10988), .B(new_n10982), .C(new_n11306), .Y(new_n11312));
  NOR2xp33_ASAP7_75t_L      g11056(.A(new_n11309), .B(new_n11312), .Y(new_n11313));
  NOR2xp33_ASAP7_75t_L      g11057(.A(new_n11311), .B(new_n11313), .Y(new_n11314));
  A2O1A1Ixp33_ASAP7_75t_L   g11058(.A1(new_n11314), .A2(new_n273), .B(new_n11305), .C(\a[2] ), .Y(new_n11315));
  AOI211xp5_ASAP7_75t_L     g11059(.A1(new_n11314), .A2(new_n273), .B(new_n11305), .C(new_n257), .Y(new_n11316));
  A2O1A1O1Ixp25_ASAP7_75t_L g11060(.A1(new_n273), .A2(new_n11314), .B(new_n11305), .C(new_n11315), .D(new_n11316), .Y(new_n11317));
  XNOR2x2_ASAP7_75t_L       g11061(.A(new_n11317), .B(new_n11302), .Y(new_n11318));
  O2A1O1Ixp33_ASAP7_75t_L   g11062(.A1(new_n10997), .A2(new_n10994), .B(new_n11001), .C(new_n11318), .Y(new_n11319));
  MAJIxp5_ASAP7_75t_L       g11063(.A(new_n11003), .B(new_n10998), .C(new_n10996), .Y(new_n11320));
  AND2x2_ASAP7_75t_L        g11064(.A(new_n11320), .B(new_n11318), .Y(new_n11321));
  NOR2xp33_ASAP7_75t_L      g11065(.A(new_n11321), .B(new_n11319), .Y(\f[58] ));
  AOI21xp33_ASAP7_75t_L     g11066(.A1(new_n11007), .A2(new_n11291), .B(new_n11300), .Y(new_n11323));
  A2O1A1O1Ixp25_ASAP7_75t_L g11067(.A1(new_n10958), .A2(new_n10972), .B(new_n10971), .C(new_n11288), .D(new_n11286), .Y(new_n11324));
  OAI22xp33_ASAP7_75t_L     g11068(.A1(new_n513), .A2(new_n9355), .B1(new_n8779), .B2(new_n506), .Y(new_n11325));
  AOI221xp5_ASAP7_75t_L     g11069(.A1(new_n475), .A2(\b[53] ), .B1(new_n483), .B2(new_n9690), .C(new_n11325), .Y(new_n11326));
  XNOR2x2_ASAP7_75t_L       g11070(.A(new_n466), .B(new_n11326), .Y(new_n11327));
  NOR3xp33_ASAP7_75t_L      g11071(.A(new_n11265), .B(new_n11269), .C(new_n11021), .Y(new_n11328));
  A2O1A1O1Ixp25_ASAP7_75t_L g11072(.A1(new_n10946), .A2(new_n10952), .B(new_n11279), .C(new_n11270), .D(new_n11328), .Y(new_n11329));
  A2O1A1Ixp33_ASAP7_75t_L   g11073(.A1(new_n10943), .A2(new_n11022), .B(new_n11260), .C(new_n11268), .Y(new_n11330));
  OAI21xp33_ASAP7_75t_L     g11074(.A1(new_n11197), .A2(new_n11195), .B(new_n11188), .Y(new_n11331));
  A2O1A1Ixp33_ASAP7_75t_L   g11075(.A1(new_n11182), .A2(new_n11177), .B(new_n11023), .C(new_n11190), .Y(new_n11332));
  A2O1A1O1Ixp25_ASAP7_75t_L g11076(.A1(new_n11116), .A2(new_n11140), .B(new_n11114), .C(new_n11135), .D(new_n11123), .Y(new_n11333));
  O2A1O1Ixp33_ASAP7_75t_L   g11077(.A1(new_n11144), .A2(new_n11141), .B(new_n11145), .C(new_n11333), .Y(new_n11334));
  NOR2xp33_ASAP7_75t_L      g11078(.A(new_n1150), .B(new_n7304), .Y(new_n11335));
  AOI221xp5_ASAP7_75t_L     g11079(.A1(\b[15] ), .A2(new_n6742), .B1(\b[17] ), .B2(new_n6442), .C(new_n11335), .Y(new_n11336));
  INVx1_ASAP7_75t_L         g11080(.A(new_n11336), .Y(new_n11337));
  A2O1A1Ixp33_ASAP7_75t_L   g11081(.A1(new_n1633), .A2(new_n6450), .B(new_n11337), .C(\a[44] ), .Y(new_n11338));
  INVx1_ASAP7_75t_L         g11082(.A(new_n11338), .Y(new_n11339));
  O2A1O1Ixp33_ASAP7_75t_L   g11083(.A1(new_n6443), .A2(new_n1356), .B(new_n11336), .C(\a[44] ), .Y(new_n11340));
  INVx1_ASAP7_75t_L         g11084(.A(new_n11340), .Y(new_n11341));
  OAI21xp33_ASAP7_75t_L     g11085(.A1(new_n6439), .A2(new_n11339), .B(new_n11341), .Y(new_n11342));
  INVx1_ASAP7_75t_L         g11086(.A(new_n10785), .Y(new_n11343));
  A2O1A1Ixp33_ASAP7_75t_L   g11087(.A1(new_n11343), .A2(new_n11027), .B(new_n10782), .C(new_n11098), .Y(new_n11344));
  A2O1A1Ixp33_ASAP7_75t_L   g11088(.A1(new_n11081), .A2(new_n11082), .B(new_n11084), .C(new_n11087), .Y(new_n11345));
  OAI22xp33_ASAP7_75t_L     g11089(.A1(new_n8483), .A2(new_n590), .B1(new_n680), .B2(new_n10065), .Y(new_n11346));
  AOI221xp5_ASAP7_75t_L     g11090(.A1(new_n8175), .A2(\b[11] ), .B1(new_n8490), .B2(new_n976), .C(new_n11346), .Y(new_n11347));
  XNOR2x2_ASAP7_75t_L       g11091(.A(new_n8172), .B(new_n11347), .Y(new_n11348));
  AOI21xp33_ASAP7_75t_L     g11092(.A1(new_n11029), .A2(new_n11070), .B(new_n11077), .Y(new_n11349));
  OAI21xp33_ASAP7_75t_L     g11093(.A1(new_n11060), .A2(new_n11037), .B(new_n11061), .Y(new_n11350));
  INVx1_ASAP7_75t_L         g11094(.A(new_n11053), .Y(new_n11351));
  INVx1_ASAP7_75t_L         g11095(.A(new_n11045), .Y(new_n11352));
  NAND2xp33_ASAP7_75t_L     g11096(.A(\b[2] ), .B(new_n11051), .Y(new_n11353));
  NAND3xp33_ASAP7_75t_L     g11097(.A(new_n10732), .B(new_n11044), .C(new_n11050), .Y(new_n11354));
  OAI221xp5_ASAP7_75t_L     g11098(.A1(new_n11352), .A2(new_n262), .B1(new_n11354), .B2(new_n284), .C(new_n11353), .Y(new_n11355));
  A2O1A1Ixp33_ASAP7_75t_L   g11099(.A1(new_n294), .A2(new_n11351), .B(new_n11355), .C(\a[59] ), .Y(new_n11356));
  AOI21xp33_ASAP7_75t_L     g11100(.A1(new_n11351), .A2(new_n294), .B(new_n11355), .Y(new_n11357));
  NOR2xp33_ASAP7_75t_L      g11101(.A(\a[59] ), .B(new_n11357), .Y(new_n11358));
  A2O1A1O1Ixp25_ASAP7_75t_L g11102(.A1(new_n11055), .A2(new_n10734), .B(new_n11356), .C(\a[59] ), .D(new_n11358), .Y(new_n11359));
  AND4x1_ASAP7_75t_L        g11103(.A(new_n11357), .B(new_n11055), .C(new_n10734), .D(\a[59] ), .Y(new_n11360));
  INVx1_ASAP7_75t_L         g11104(.A(new_n10390), .Y(new_n11361));
  NOR2xp33_ASAP7_75t_L      g11105(.A(new_n332), .B(new_n10388), .Y(new_n11362));
  AOI221xp5_ASAP7_75t_L     g11106(.A1(new_n10086), .A2(\b[5] ), .B1(new_n11361), .B2(\b[3] ), .C(new_n11362), .Y(new_n11363));
  O2A1O1Ixp33_ASAP7_75t_L   g11107(.A1(new_n728), .A2(new_n10088), .B(new_n11363), .C(new_n10083), .Y(new_n11364));
  NOR2xp33_ASAP7_75t_L      g11108(.A(new_n10083), .B(new_n11364), .Y(new_n11365));
  O2A1O1Ixp33_ASAP7_75t_L   g11109(.A1(new_n728), .A2(new_n10088), .B(new_n11363), .C(\a[56] ), .Y(new_n11366));
  NOR2xp33_ASAP7_75t_L      g11110(.A(new_n11366), .B(new_n11365), .Y(new_n11367));
  NOR3xp33_ASAP7_75t_L      g11111(.A(new_n11359), .B(new_n11367), .C(new_n11360), .Y(new_n11368));
  OA21x2_ASAP7_75t_L        g11112(.A1(new_n11360), .A2(new_n11359), .B(new_n11367), .Y(new_n11369));
  OA21x2_ASAP7_75t_L        g11113(.A1(new_n11368), .A2(new_n11369), .B(new_n11350), .Y(new_n11370));
  NOR3xp33_ASAP7_75t_L      g11114(.A(new_n11350), .B(new_n11369), .C(new_n11368), .Y(new_n11371));
  OAI22xp33_ASAP7_75t_L     g11115(.A1(new_n9440), .A2(new_n427), .B1(new_n448), .B2(new_n10400), .Y(new_n11372));
  AOI221xp5_ASAP7_75t_L     g11116(.A1(new_n9102), .A2(\b[8] ), .B1(new_n9437), .B2(new_n1684), .C(new_n11372), .Y(new_n11373));
  XNOR2x2_ASAP7_75t_L       g11117(.A(\a[53] ), .B(new_n11373), .Y(new_n11374));
  NOR3xp33_ASAP7_75t_L      g11118(.A(new_n11370), .B(new_n11374), .C(new_n11371), .Y(new_n11375));
  OA21x2_ASAP7_75t_L        g11119(.A1(new_n11371), .A2(new_n11370), .B(new_n11374), .Y(new_n11376));
  NOR3xp33_ASAP7_75t_L      g11120(.A(new_n11349), .B(new_n11375), .C(new_n11376), .Y(new_n11377));
  AO21x2_ASAP7_75t_L        g11121(.A1(new_n11070), .A2(new_n11029), .B(new_n11077), .Y(new_n11378));
  NOR2xp33_ASAP7_75t_L      g11122(.A(new_n11375), .B(new_n11376), .Y(new_n11379));
  NOR2xp33_ASAP7_75t_L      g11123(.A(new_n11378), .B(new_n11379), .Y(new_n11380));
  OAI21xp33_ASAP7_75t_L     g11124(.A1(new_n11377), .A2(new_n11380), .B(new_n11348), .Y(new_n11381));
  INVx1_ASAP7_75t_L         g11125(.A(new_n11348), .Y(new_n11382));
  A2O1A1Ixp33_ASAP7_75t_L   g11126(.A1(new_n11070), .A2(new_n11029), .B(new_n11077), .C(new_n11379), .Y(new_n11383));
  OAI21xp33_ASAP7_75t_L     g11127(.A1(new_n11375), .A2(new_n11376), .B(new_n11349), .Y(new_n11384));
  NAND3xp33_ASAP7_75t_L     g11128(.A(new_n11382), .B(new_n11383), .C(new_n11384), .Y(new_n11385));
  NAND3xp33_ASAP7_75t_L     g11129(.A(new_n11385), .B(new_n11345), .C(new_n11381), .Y(new_n11386));
  AND3x1_ASAP7_75t_L        g11130(.A(new_n11074), .B(new_n11086), .C(new_n11078), .Y(new_n11387));
  O2A1O1Ixp33_ASAP7_75t_L   g11131(.A1(new_n11086), .A2(new_n11088), .B(new_n11089), .C(new_n11387), .Y(new_n11388));
  AOI21xp33_ASAP7_75t_L     g11132(.A1(new_n11383), .A2(new_n11384), .B(new_n11382), .Y(new_n11389));
  NOR3xp33_ASAP7_75t_L      g11133(.A(new_n11380), .B(new_n11377), .C(new_n11348), .Y(new_n11390));
  OAI21xp33_ASAP7_75t_L     g11134(.A1(new_n11390), .A2(new_n11389), .B(new_n11388), .Y(new_n11391));
  NOR2xp33_ASAP7_75t_L      g11135(.A(new_n936), .B(new_n7312), .Y(new_n11392));
  AOI221xp5_ASAP7_75t_L     g11136(.A1(\b[12] ), .A2(new_n7609), .B1(\b[14] ), .B2(new_n7334), .C(new_n11392), .Y(new_n11393));
  INVx1_ASAP7_75t_L         g11137(.A(new_n11393), .Y(new_n11394));
  A2O1A1Ixp33_ASAP7_75t_L   g11138(.A1(new_n971), .A2(new_n7322), .B(new_n11394), .C(\a[47] ), .Y(new_n11395));
  O2A1O1Ixp33_ASAP7_75t_L   g11139(.A1(new_n7321), .A2(new_n1268), .B(new_n11393), .C(\a[47] ), .Y(new_n11396));
  AOI21xp33_ASAP7_75t_L     g11140(.A1(new_n11395), .A2(\a[47] ), .B(new_n11396), .Y(new_n11397));
  NAND3xp33_ASAP7_75t_L     g11141(.A(new_n11391), .B(new_n11386), .C(new_n11397), .Y(new_n11398));
  AO21x2_ASAP7_75t_L        g11142(.A1(new_n11386), .A2(new_n11391), .B(new_n11397), .Y(new_n11399));
  AOI22xp33_ASAP7_75t_L     g11143(.A1(new_n11398), .A2(new_n11399), .B1(new_n11094), .B2(new_n11344), .Y(new_n11400));
  AND3x1_ASAP7_75t_L        g11144(.A(new_n11391), .B(new_n11386), .C(new_n11397), .Y(new_n11401));
  AOI21xp33_ASAP7_75t_L     g11145(.A1(new_n11391), .A2(new_n11386), .B(new_n11397), .Y(new_n11402));
  NOR4xp25_ASAP7_75t_L      g11146(.A(new_n11401), .B(new_n11097), .C(new_n11102), .D(new_n11402), .Y(new_n11403));
  OAI21xp33_ASAP7_75t_L     g11147(.A1(new_n11403), .A2(new_n11400), .B(new_n11342), .Y(new_n11404));
  AOI21xp33_ASAP7_75t_L     g11148(.A1(new_n11338), .A2(\a[44] ), .B(new_n11340), .Y(new_n11405));
  OAI22xp33_ASAP7_75t_L     g11149(.A1(new_n11401), .A2(new_n11402), .B1(new_n11102), .B2(new_n11097), .Y(new_n11406));
  NAND4xp25_ASAP7_75t_L     g11150(.A(new_n11344), .B(new_n11398), .C(new_n11399), .D(new_n11094), .Y(new_n11407));
  NAND3xp33_ASAP7_75t_L     g11151(.A(new_n11407), .B(new_n11406), .C(new_n11405), .Y(new_n11408));
  NAND2xp33_ASAP7_75t_L     g11152(.A(new_n11408), .B(new_n11404), .Y(new_n11409));
  O2A1O1Ixp33_ASAP7_75t_L   g11153(.A1(new_n11108), .A2(new_n11129), .B(new_n11127), .C(new_n11409), .Y(new_n11410));
  AOI221xp5_ASAP7_75t_L     g11154(.A1(new_n11408), .A2(new_n11404), .B1(new_n11105), .B2(new_n11106), .C(new_n11100), .Y(new_n11411));
  NOR2xp33_ASAP7_75t_L      g11155(.A(new_n1599), .B(new_n5640), .Y(new_n11412));
  AOI221xp5_ASAP7_75t_L     g11156(.A1(\b[18] ), .A2(new_n5920), .B1(\b[20] ), .B2(new_n5629), .C(new_n11412), .Y(new_n11413));
  INVx1_ASAP7_75t_L         g11157(.A(new_n11413), .Y(new_n11414));
  A2O1A1Ixp33_ASAP7_75t_L   g11158(.A1(new_n1752), .A2(new_n5637), .B(new_n11414), .C(\a[41] ), .Y(new_n11415));
  O2A1O1Ixp33_ASAP7_75t_L   g11159(.A1(new_n5630), .A2(new_n1754), .B(new_n11413), .C(\a[41] ), .Y(new_n11416));
  AOI21xp33_ASAP7_75t_L     g11160(.A1(new_n11415), .A2(\a[41] ), .B(new_n11416), .Y(new_n11417));
  OAI21xp33_ASAP7_75t_L     g11161(.A1(new_n11410), .A2(new_n11411), .B(new_n11417), .Y(new_n11418));
  AOI21xp33_ASAP7_75t_L     g11162(.A1(new_n11407), .A2(new_n11406), .B(new_n11405), .Y(new_n11419));
  NOR3xp33_ASAP7_75t_L      g11163(.A(new_n11400), .B(new_n11342), .C(new_n11403), .Y(new_n11420));
  NOR2xp33_ASAP7_75t_L      g11164(.A(new_n11419), .B(new_n11420), .Y(new_n11421));
  A2O1A1Ixp33_ASAP7_75t_L   g11165(.A1(new_n11105), .A2(new_n11106), .B(new_n11100), .C(new_n11421), .Y(new_n11422));
  OAI211xp5_ASAP7_75t_L     g11166(.A1(new_n11129), .A2(new_n11108), .B(new_n11409), .C(new_n11127), .Y(new_n11423));
  INVx1_ASAP7_75t_L         g11167(.A(new_n11417), .Y(new_n11424));
  NAND3xp33_ASAP7_75t_L     g11168(.A(new_n11422), .B(new_n11423), .C(new_n11424), .Y(new_n11425));
  NAND2xp33_ASAP7_75t_L     g11169(.A(new_n11418), .B(new_n11425), .Y(new_n11426));
  O2A1O1Ixp33_ASAP7_75t_L   g11170(.A1(new_n11114), .A2(new_n11133), .B(new_n11116), .C(new_n11426), .Y(new_n11427));
  AOI211xp5_ASAP7_75t_L     g11171(.A1(new_n11425), .A2(new_n11418), .B(new_n11115), .C(new_n11140), .Y(new_n11428));
  NOR2xp33_ASAP7_75t_L      g11172(.A(new_n2188), .B(new_n4908), .Y(new_n11429));
  AOI221xp5_ASAP7_75t_L     g11173(.A1(\b[21] ), .A2(new_n5139), .B1(\b[22] ), .B2(new_n4916), .C(new_n11429), .Y(new_n11430));
  O2A1O1Ixp33_ASAP7_75t_L   g11174(.A1(new_n4911), .A2(new_n2194), .B(new_n11430), .C(new_n4906), .Y(new_n11431));
  OAI21xp33_ASAP7_75t_L     g11175(.A1(new_n4911), .A2(new_n2194), .B(new_n11430), .Y(new_n11432));
  NAND2xp33_ASAP7_75t_L     g11176(.A(new_n4906), .B(new_n11432), .Y(new_n11433));
  OAI21xp33_ASAP7_75t_L     g11177(.A1(new_n4906), .A2(new_n11431), .B(new_n11433), .Y(new_n11434));
  OAI21xp33_ASAP7_75t_L     g11178(.A1(new_n11428), .A2(new_n11427), .B(new_n11434), .Y(new_n11435));
  AOI21xp33_ASAP7_75t_L     g11179(.A1(new_n11422), .A2(new_n11423), .B(new_n11424), .Y(new_n11436));
  NOR3xp33_ASAP7_75t_L      g11180(.A(new_n11411), .B(new_n11410), .C(new_n11417), .Y(new_n11437));
  NOR2xp33_ASAP7_75t_L      g11181(.A(new_n11437), .B(new_n11436), .Y(new_n11438));
  OAI21xp33_ASAP7_75t_L     g11182(.A1(new_n11115), .A2(new_n11140), .B(new_n11438), .Y(new_n11439));
  NAND2xp33_ASAP7_75t_L     g11183(.A(new_n11426), .B(new_n11118), .Y(new_n11440));
  OA21x2_ASAP7_75t_L        g11184(.A1(new_n4906), .A2(new_n11431), .B(new_n11433), .Y(new_n11441));
  NAND3xp33_ASAP7_75t_L     g11185(.A(new_n11440), .B(new_n11439), .C(new_n11441), .Y(new_n11442));
  NAND2xp33_ASAP7_75t_L     g11186(.A(new_n11442), .B(new_n11435), .Y(new_n11443));
  NAND2xp33_ASAP7_75t_L     g11187(.A(new_n11443), .B(new_n11334), .Y(new_n11444));
  NAND2xp33_ASAP7_75t_L     g11188(.A(new_n11137), .B(new_n11124), .Y(new_n11445));
  AOI21xp33_ASAP7_75t_L     g11189(.A1(new_n11440), .A2(new_n11439), .B(new_n11441), .Y(new_n11446));
  NOR3xp33_ASAP7_75t_L      g11190(.A(new_n11427), .B(new_n11428), .C(new_n11434), .Y(new_n11447));
  NOR2xp33_ASAP7_75t_L      g11191(.A(new_n11446), .B(new_n11447), .Y(new_n11448));
  A2O1A1Ixp33_ASAP7_75t_L   g11192(.A1(new_n11445), .A2(new_n11145), .B(new_n11333), .C(new_n11448), .Y(new_n11449));
  OAI22xp33_ASAP7_75t_L     g11193(.A1(new_n4397), .A2(new_n2205), .B1(new_n2377), .B2(new_n4142), .Y(new_n11450));
  AOI221xp5_ASAP7_75t_L     g11194(.A1(new_n4156), .A2(\b[26] ), .B1(new_n4151), .B2(new_n2709), .C(new_n11450), .Y(new_n11451));
  XNOR2x2_ASAP7_75t_L       g11195(.A(new_n4145), .B(new_n11451), .Y(new_n11452));
  NAND3xp33_ASAP7_75t_L     g11196(.A(new_n11449), .B(new_n11444), .C(new_n11452), .Y(new_n11453));
  AOI221xp5_ASAP7_75t_L     g11197(.A1(new_n11442), .A2(new_n11435), .B1(new_n11145), .B2(new_n11445), .C(new_n11333), .Y(new_n11454));
  NOR2xp33_ASAP7_75t_L      g11198(.A(new_n11443), .B(new_n11334), .Y(new_n11455));
  XNOR2x2_ASAP7_75t_L       g11199(.A(\a[35] ), .B(new_n11451), .Y(new_n11456));
  OAI21xp33_ASAP7_75t_L     g11200(.A1(new_n11454), .A2(new_n11455), .B(new_n11456), .Y(new_n11457));
  NAND2xp33_ASAP7_75t_L     g11201(.A(new_n11457), .B(new_n11453), .Y(new_n11458));
  A2O1A1Ixp33_ASAP7_75t_L   g11202(.A1(new_n11149), .A2(new_n11150), .B(new_n11163), .C(new_n11161), .Y(new_n11459));
  NOR2xp33_ASAP7_75t_L      g11203(.A(new_n11458), .B(new_n11459), .Y(new_n11460));
  AND2x2_ASAP7_75t_L        g11204(.A(new_n11457), .B(new_n11453), .Y(new_n11461));
  O2A1O1Ixp33_ASAP7_75t_L   g11205(.A1(new_n11174), .A2(new_n11163), .B(new_n11161), .C(new_n11461), .Y(new_n11462));
  NAND2xp33_ASAP7_75t_L     g11206(.A(\b[28] ), .B(new_n3499), .Y(new_n11463));
  OAI221xp5_ASAP7_75t_L     g11207(.A1(new_n3510), .A2(new_n3098), .B1(new_n2879), .B2(new_n3703), .C(new_n11463), .Y(new_n11464));
  A2O1A1Ixp33_ASAP7_75t_L   g11208(.A1(new_n3873), .A2(new_n3505), .B(new_n11464), .C(\a[32] ), .Y(new_n11465));
  NAND2xp33_ASAP7_75t_L     g11209(.A(\a[32] ), .B(new_n11465), .Y(new_n11466));
  A2O1A1Ixp33_ASAP7_75t_L   g11210(.A1(new_n3873), .A2(new_n3505), .B(new_n11464), .C(new_n3493), .Y(new_n11467));
  NAND2xp33_ASAP7_75t_L     g11211(.A(new_n11467), .B(new_n11466), .Y(new_n11468));
  INVx1_ASAP7_75t_L         g11212(.A(new_n11468), .Y(new_n11469));
  NOR3xp33_ASAP7_75t_L      g11213(.A(new_n11462), .B(new_n11469), .C(new_n11460), .Y(new_n11470));
  O2A1O1Ixp33_ASAP7_75t_L   g11214(.A1(new_n11173), .A2(new_n11172), .B(new_n11159), .C(new_n11162), .Y(new_n11471));
  NAND2xp33_ASAP7_75t_L     g11215(.A(new_n11461), .B(new_n11471), .Y(new_n11472));
  A2O1A1Ixp33_ASAP7_75t_L   g11216(.A1(new_n11156), .A2(new_n11159), .B(new_n11162), .C(new_n11458), .Y(new_n11473));
  AOI21xp33_ASAP7_75t_L     g11217(.A1(new_n11472), .A2(new_n11473), .B(new_n11468), .Y(new_n11474));
  OAI21xp33_ASAP7_75t_L     g11218(.A1(new_n11470), .A2(new_n11474), .B(new_n11332), .Y(new_n11475));
  OAI21xp33_ASAP7_75t_L     g11219(.A1(new_n11178), .A2(new_n11171), .B(new_n11181), .Y(new_n11476));
  NAND3xp33_ASAP7_75t_L     g11220(.A(new_n11472), .B(new_n11473), .C(new_n11468), .Y(new_n11477));
  OAI21xp33_ASAP7_75t_L     g11221(.A1(new_n11460), .A2(new_n11462), .B(new_n11469), .Y(new_n11478));
  NAND4xp25_ASAP7_75t_L     g11222(.A(new_n11476), .B(new_n11478), .C(new_n11190), .D(new_n11477), .Y(new_n11479));
  OAI22xp33_ASAP7_75t_L     g11223(.A1(new_n3133), .A2(new_n3456), .B1(new_n3674), .B2(new_n2925), .Y(new_n11480));
  AOI221xp5_ASAP7_75t_L     g11224(.A1(new_n2938), .A2(\b[32] ), .B1(new_n2932), .B2(new_n3900), .C(new_n11480), .Y(new_n11481));
  XNOR2x2_ASAP7_75t_L       g11225(.A(new_n2928), .B(new_n11481), .Y(new_n11482));
  NAND3xp33_ASAP7_75t_L     g11226(.A(new_n11475), .B(new_n11479), .C(new_n11482), .Y(new_n11483));
  AO21x2_ASAP7_75t_L        g11227(.A1(new_n11479), .A2(new_n11475), .B(new_n11482), .Y(new_n11484));
  NAND3xp33_ASAP7_75t_L     g11228(.A(new_n11331), .B(new_n11483), .C(new_n11484), .Y(new_n11485));
  A2O1A1O1Ixp25_ASAP7_75t_L g11229(.A1(new_n10864), .A2(new_n10691), .B(new_n10855), .C(new_n11193), .D(new_n11196), .Y(new_n11486));
  AND3x1_ASAP7_75t_L        g11230(.A(new_n11475), .B(new_n11482), .C(new_n11479), .Y(new_n11487));
  AOI21xp33_ASAP7_75t_L     g11231(.A1(new_n11475), .A2(new_n11479), .B(new_n11482), .Y(new_n11488));
  OAI21xp33_ASAP7_75t_L     g11232(.A1(new_n11487), .A2(new_n11488), .B(new_n11486), .Y(new_n11489));
  OAI22xp33_ASAP7_75t_L     g11233(.A1(new_n2572), .A2(new_n4101), .B1(new_n4344), .B2(new_n2410), .Y(new_n11490));
  AOI221xp5_ASAP7_75t_L     g11234(.A1(new_n2423), .A2(\b[35] ), .B1(new_n2417), .B2(new_n7773), .C(new_n11490), .Y(new_n11491));
  XNOR2x2_ASAP7_75t_L       g11235(.A(new_n2413), .B(new_n11491), .Y(new_n11492));
  NAND3xp33_ASAP7_75t_L     g11236(.A(new_n11485), .B(new_n11492), .C(new_n11489), .Y(new_n11493));
  AO21x2_ASAP7_75t_L        g11237(.A1(new_n11489), .A2(new_n11485), .B(new_n11492), .Y(new_n11494));
  NAND2xp33_ASAP7_75t_L     g11238(.A(new_n11493), .B(new_n11494), .Y(new_n11495));
  OAI21xp33_ASAP7_75t_L     g11239(.A1(new_n11206), .A2(new_n11204), .B(new_n11209), .Y(new_n11496));
  NOR2xp33_ASAP7_75t_L      g11240(.A(new_n11495), .B(new_n11496), .Y(new_n11497));
  NOR3xp33_ASAP7_75t_L      g11241(.A(new_n11486), .B(new_n11487), .C(new_n11488), .Y(new_n11498));
  AOI21xp33_ASAP7_75t_L     g11242(.A1(new_n11484), .A2(new_n11483), .B(new_n11331), .Y(new_n11499));
  NOR3xp33_ASAP7_75t_L      g11243(.A(new_n11498), .B(new_n11499), .C(new_n11492), .Y(new_n11500));
  MAJIxp5_ASAP7_75t_L       g11244(.A(new_n11210), .B(new_n11208), .C(new_n11201), .Y(new_n11501));
  O2A1O1Ixp33_ASAP7_75t_L   g11245(.A1(new_n11492), .A2(new_n11500), .B(new_n11493), .C(new_n11501), .Y(new_n11502));
  OAI22xp33_ASAP7_75t_L     g11246(.A1(new_n2089), .A2(new_n4613), .B1(new_n5074), .B2(new_n1962), .Y(new_n11503));
  AOI221xp5_ASAP7_75t_L     g11247(.A1(new_n1955), .A2(\b[38] ), .B1(new_n1964), .B2(new_n6083), .C(new_n11503), .Y(new_n11504));
  XNOR2x2_ASAP7_75t_L       g11248(.A(\a[23] ), .B(new_n11504), .Y(new_n11505));
  NOR3xp33_ASAP7_75t_L      g11249(.A(new_n11497), .B(new_n11502), .C(new_n11505), .Y(new_n11506));
  OA21x2_ASAP7_75t_L        g11250(.A1(new_n11502), .A2(new_n11497), .B(new_n11505), .Y(new_n11507));
  INVx1_ASAP7_75t_L         g11251(.A(new_n11214), .Y(new_n11508));
  NAND3xp33_ASAP7_75t_L     g11252(.A(new_n11508), .B(new_n11211), .C(new_n11207), .Y(new_n11509));
  A2O1A1Ixp33_ASAP7_75t_L   g11253(.A1(new_n11215), .A2(new_n11216), .B(new_n11217), .C(new_n11509), .Y(new_n11510));
  NOR3xp33_ASAP7_75t_L      g11254(.A(new_n11510), .B(new_n11507), .C(new_n11506), .Y(new_n11511));
  OA21x2_ASAP7_75t_L        g11255(.A1(new_n11506), .A2(new_n11507), .B(new_n11510), .Y(new_n11512));
  NOR2xp33_ASAP7_75t_L      g11256(.A(new_n6110), .B(new_n1518), .Y(new_n11513));
  AOI221xp5_ASAP7_75t_L     g11257(.A1(\b[39] ), .A2(new_n1659), .B1(\b[40] ), .B2(new_n1507), .C(new_n11513), .Y(new_n11514));
  O2A1O1Ixp33_ASAP7_75t_L   g11258(.A1(new_n1521), .A2(new_n6117), .B(new_n11514), .C(new_n1501), .Y(new_n11515));
  OAI21xp33_ASAP7_75t_L     g11259(.A1(new_n1521), .A2(new_n6117), .B(new_n11514), .Y(new_n11516));
  NAND2xp33_ASAP7_75t_L     g11260(.A(new_n1501), .B(new_n11516), .Y(new_n11517));
  OAI21xp33_ASAP7_75t_L     g11261(.A1(new_n1501), .A2(new_n11515), .B(new_n11517), .Y(new_n11518));
  INVx1_ASAP7_75t_L         g11262(.A(new_n11518), .Y(new_n11519));
  OAI21xp33_ASAP7_75t_L     g11263(.A1(new_n11511), .A2(new_n11512), .B(new_n11519), .Y(new_n11520));
  NOR3xp33_ASAP7_75t_L      g11264(.A(new_n11512), .B(new_n11519), .C(new_n11511), .Y(new_n11521));
  INVx1_ASAP7_75t_L         g11265(.A(new_n11521), .Y(new_n11522));
  AOI22xp33_ASAP7_75t_L     g11266(.A1(new_n11522), .A2(new_n11520), .B1(new_n11237), .B2(new_n11250), .Y(new_n11523));
  INVx1_ASAP7_75t_L         g11267(.A(new_n11237), .Y(new_n11524));
  A2O1A1O1Ixp25_ASAP7_75t_L g11268(.A1(new_n11231), .A2(new_n11234), .B(new_n11524), .C(new_n11520), .D(new_n11521), .Y(new_n11525));
  NOR2xp33_ASAP7_75t_L      g11269(.A(new_n6671), .B(new_n2118), .Y(new_n11526));
  AOI221xp5_ASAP7_75t_L     g11270(.A1(\b[42] ), .A2(new_n1290), .B1(\b[44] ), .B2(new_n1209), .C(new_n11526), .Y(new_n11527));
  INVx1_ASAP7_75t_L         g11271(.A(new_n11527), .Y(new_n11528));
  A2O1A1Ixp33_ASAP7_75t_L   g11272(.A1(new_n7824), .A2(new_n1216), .B(new_n11528), .C(\a[17] ), .Y(new_n11529));
  O2A1O1Ixp33_ASAP7_75t_L   g11273(.A1(new_n1210), .A2(new_n6951), .B(new_n11527), .C(new_n1206), .Y(new_n11530));
  NOR2xp33_ASAP7_75t_L      g11274(.A(new_n1206), .B(new_n11530), .Y(new_n11531));
  A2O1A1O1Ixp25_ASAP7_75t_L g11275(.A1(new_n7824), .A2(new_n1216), .B(new_n11528), .C(new_n11529), .D(new_n11531), .Y(new_n11532));
  A2O1A1Ixp33_ASAP7_75t_L   g11276(.A1(new_n11525), .A2(new_n11520), .B(new_n11523), .C(new_n11532), .Y(new_n11533));
  A2O1A1Ixp33_ASAP7_75t_L   g11277(.A1(new_n10921), .A2(new_n11233), .B(new_n11239), .C(new_n11237), .Y(new_n11534));
  OA21x2_ASAP7_75t_L        g11278(.A1(new_n11511), .A2(new_n11512), .B(new_n11519), .Y(new_n11535));
  OAI21xp33_ASAP7_75t_L     g11279(.A1(new_n11521), .A2(new_n11535), .B(new_n11534), .Y(new_n11536));
  NAND4xp25_ASAP7_75t_L     g11280(.A(new_n11250), .B(new_n11522), .C(new_n11520), .D(new_n11237), .Y(new_n11537));
  INVx1_ASAP7_75t_L         g11281(.A(new_n11532), .Y(new_n11538));
  NAND3xp33_ASAP7_75t_L     g11282(.A(new_n11536), .B(new_n11537), .C(new_n11538), .Y(new_n11539));
  NAND2xp33_ASAP7_75t_L     g11283(.A(new_n11539), .B(new_n11533), .Y(new_n11540));
  O2A1O1Ixp33_ASAP7_75t_L   g11284(.A1(new_n11245), .A2(new_n11261), .B(new_n11252), .C(new_n11540), .Y(new_n11541));
  NOR2xp33_ASAP7_75t_L      g11285(.A(new_n11511), .B(new_n11512), .Y(new_n11542));
  O2A1O1Ixp33_ASAP7_75t_L   g11286(.A1(new_n11518), .A2(new_n11542), .B(new_n11525), .C(new_n11523), .Y(new_n11543));
  A2O1A1Ixp33_ASAP7_75t_L   g11287(.A1(new_n11525), .A2(new_n11520), .B(new_n11523), .C(new_n11538), .Y(new_n11544));
  INVx1_ASAP7_75t_L         g11288(.A(new_n11544), .Y(new_n11545));
  O2A1O1Ixp33_ASAP7_75t_L   g11289(.A1(new_n11543), .A2(new_n11545), .B(new_n11539), .C(new_n11263), .Y(new_n11546));
  OAI22xp33_ASAP7_75t_L     g11290(.A1(new_n980), .A2(new_n7249), .B1(new_n7270), .B2(new_n864), .Y(new_n11547));
  AOI221xp5_ASAP7_75t_L     g11291(.A1(new_n886), .A2(\b[47] ), .B1(new_n873), .B2(new_n8726), .C(new_n11547), .Y(new_n11548));
  XNOR2x2_ASAP7_75t_L       g11292(.A(new_n867), .B(new_n11548), .Y(new_n11549));
  INVx1_ASAP7_75t_L         g11293(.A(new_n11549), .Y(new_n11550));
  OAI21xp33_ASAP7_75t_L     g11294(.A1(new_n11541), .A2(new_n11546), .B(new_n11550), .Y(new_n11551));
  O2A1O1Ixp33_ASAP7_75t_L   g11295(.A1(new_n11238), .A2(new_n11225), .B(new_n11234), .C(new_n11524), .Y(new_n11552));
  O2A1O1Ixp33_ASAP7_75t_L   g11296(.A1(new_n11239), .A2(new_n11248), .B(new_n11237), .C(new_n11535), .Y(new_n11553));
  A2O1A1O1Ixp25_ASAP7_75t_L g11297(.A1(new_n11522), .A2(new_n11553), .B(new_n11552), .C(new_n11537), .D(new_n11538), .Y(new_n11554));
  AOI211xp5_ASAP7_75t_L     g11298(.A1(new_n11525), .A2(new_n11520), .B(new_n11532), .C(new_n11523), .Y(new_n11555));
  NOR2xp33_ASAP7_75t_L      g11299(.A(new_n11554), .B(new_n11555), .Y(new_n11556));
  NAND2xp33_ASAP7_75t_L     g11300(.A(new_n11263), .B(new_n11556), .Y(new_n11557));
  A2O1A1Ixp33_ASAP7_75t_L   g11301(.A1(new_n11522), .A2(new_n11553), .B(new_n11552), .C(new_n11537), .Y(new_n11558));
  A2O1A1Ixp33_ASAP7_75t_L   g11302(.A1(new_n11558), .A2(new_n11544), .B(new_n11555), .C(new_n11255), .Y(new_n11559));
  NAND3xp33_ASAP7_75t_L     g11303(.A(new_n11557), .B(new_n11559), .C(new_n11549), .Y(new_n11560));
  NAND3xp33_ASAP7_75t_L     g11304(.A(new_n11330), .B(new_n11551), .C(new_n11560), .Y(new_n11561));
  A2O1A1O1Ixp25_ASAP7_75t_L g11305(.A1(new_n10671), .A2(new_n10936), .B(new_n11266), .C(new_n11267), .D(new_n11264), .Y(new_n11562));
  AOI21xp33_ASAP7_75t_L     g11306(.A1(new_n11557), .A2(new_n11559), .B(new_n11549), .Y(new_n11563));
  NOR3xp33_ASAP7_75t_L      g11307(.A(new_n11546), .B(new_n11541), .C(new_n11550), .Y(new_n11564));
  OAI21xp33_ASAP7_75t_L     g11308(.A1(new_n11563), .A2(new_n11564), .B(new_n11562), .Y(new_n11565));
  OAI22xp33_ASAP7_75t_L     g11309(.A1(new_n1550), .A2(new_n8427), .B1(new_n7860), .B2(new_n712), .Y(new_n11566));
  AOI221xp5_ASAP7_75t_L     g11310(.A1(new_n640), .A2(\b[50] ), .B1(new_n718), .B2(new_n8763), .C(new_n11566), .Y(new_n11567));
  XNOR2x2_ASAP7_75t_L       g11311(.A(new_n637), .B(new_n11567), .Y(new_n11568));
  NAND3xp33_ASAP7_75t_L     g11312(.A(new_n11561), .B(new_n11565), .C(new_n11568), .Y(new_n11569));
  AO21x2_ASAP7_75t_L        g11313(.A1(new_n11565), .A2(new_n11561), .B(new_n11568), .Y(new_n11570));
  AO21x2_ASAP7_75t_L        g11314(.A1(new_n11570), .A2(new_n11569), .B(new_n11329), .Y(new_n11571));
  NAND3xp33_ASAP7_75t_L     g11315(.A(new_n11329), .B(new_n11569), .C(new_n11570), .Y(new_n11572));
  AOI21xp33_ASAP7_75t_L     g11316(.A1(new_n11571), .A2(new_n11572), .B(new_n11327), .Y(new_n11573));
  NAND3xp33_ASAP7_75t_L     g11317(.A(new_n11571), .B(new_n11327), .C(new_n11572), .Y(new_n11574));
  INVx1_ASAP7_75t_L         g11318(.A(new_n11574), .Y(new_n11575));
  NOR3xp33_ASAP7_75t_L      g11319(.A(new_n11324), .B(new_n11575), .C(new_n11573), .Y(new_n11576));
  AO21x2_ASAP7_75t_L        g11320(.A1(new_n11572), .A2(new_n11571), .B(new_n11327), .Y(new_n11577));
  AOI221xp5_ASAP7_75t_L     g11321(.A1(new_n11577), .A2(new_n11574), .B1(new_n11288), .B2(new_n11293), .C(new_n11286), .Y(new_n11578));
  INVx1_ASAP7_75t_L         g11322(.A(new_n10339), .Y(new_n11579));
  OAI22xp33_ASAP7_75t_L     g11323(.A1(new_n350), .A2(new_n10309), .B1(new_n9709), .B2(new_n375), .Y(new_n11580));
  AOI221xp5_ASAP7_75t_L     g11324(.A1(new_n361), .A2(\b[56] ), .B1(new_n359), .B2(new_n11579), .C(new_n11580), .Y(new_n11581));
  XNOR2x2_ASAP7_75t_L       g11325(.A(new_n346), .B(new_n11581), .Y(new_n11582));
  OAI21xp33_ASAP7_75t_L     g11326(.A1(new_n11578), .A2(new_n11576), .B(new_n11582), .Y(new_n11583));
  AOI21xp33_ASAP7_75t_L     g11327(.A1(new_n11574), .A2(new_n11577), .B(new_n11324), .Y(new_n11584));
  OAI21xp33_ASAP7_75t_L     g11328(.A1(new_n11573), .A2(new_n11575), .B(new_n11324), .Y(new_n11585));
  INVx1_ASAP7_75t_L         g11329(.A(new_n11582), .Y(new_n11586));
  OAI211xp5_ASAP7_75t_L     g11330(.A1(new_n11324), .A2(new_n11584), .B(new_n11585), .C(new_n11586), .Y(new_n11587));
  NOR2xp33_ASAP7_75t_L      g11331(.A(new_n10978), .B(new_n287), .Y(new_n11588));
  AOI221xp5_ASAP7_75t_L     g11332(.A1(\b[58] ), .A2(new_n264), .B1(\b[59] ), .B2(new_n283), .C(new_n11588), .Y(new_n11589));
  NOR2xp33_ASAP7_75t_L      g11333(.A(\b[58] ), .B(\b[59] ), .Y(new_n11590));
  INVx1_ASAP7_75t_L         g11334(.A(\b[59] ), .Y(new_n11591));
  NOR2xp33_ASAP7_75t_L      g11335(.A(new_n11303), .B(new_n11591), .Y(new_n11592));
  NOR2xp33_ASAP7_75t_L      g11336(.A(new_n11590), .B(new_n11592), .Y(new_n11593));
  A2O1A1Ixp33_ASAP7_75t_L   g11337(.A1(new_n11312), .A2(new_n11309), .B(new_n11308), .C(new_n11593), .Y(new_n11594));
  A2O1A1O1Ixp25_ASAP7_75t_L g11338(.A1(new_n10984), .A2(new_n10989), .B(new_n10983), .C(new_n11309), .D(new_n11308), .Y(new_n11595));
  OAI21xp33_ASAP7_75t_L     g11339(.A1(new_n11590), .A2(new_n11592), .B(new_n11595), .Y(new_n11596));
  NAND2xp33_ASAP7_75t_L     g11340(.A(new_n11596), .B(new_n11594), .Y(new_n11597));
  O2A1O1Ixp33_ASAP7_75t_L   g11341(.A1(new_n279), .A2(new_n11597), .B(new_n11589), .C(new_n257), .Y(new_n11598));
  OAI21xp33_ASAP7_75t_L     g11342(.A1(new_n279), .A2(new_n11597), .B(new_n11589), .Y(new_n11599));
  NAND2xp33_ASAP7_75t_L     g11343(.A(new_n257), .B(new_n11599), .Y(new_n11600));
  OAI21xp33_ASAP7_75t_L     g11344(.A1(new_n257), .A2(new_n11598), .B(new_n11600), .Y(new_n11601));
  AOI21xp33_ASAP7_75t_L     g11345(.A1(new_n11587), .A2(new_n11583), .B(new_n11601), .Y(new_n11602));
  O2A1O1Ixp33_ASAP7_75t_L   g11346(.A1(new_n11324), .A2(new_n11584), .B(new_n11585), .C(new_n11586), .Y(new_n11603));
  NOR3xp33_ASAP7_75t_L      g11347(.A(new_n11576), .B(new_n11578), .C(new_n11582), .Y(new_n11604));
  INVx1_ASAP7_75t_L         g11348(.A(new_n11601), .Y(new_n11605));
  NOR3xp33_ASAP7_75t_L      g11349(.A(new_n11603), .B(new_n11604), .C(new_n11605), .Y(new_n11606));
  NOR2xp33_ASAP7_75t_L      g11350(.A(new_n11602), .B(new_n11606), .Y(new_n11607));
  A2O1A1O1Ixp25_ASAP7_75t_L g11351(.A1(new_n10976), .A2(new_n10975), .B(new_n11299), .C(new_n11296), .D(new_n11607), .Y(new_n11608));
  MAJIxp5_ASAP7_75t_L       g11352(.A(new_n11320), .B(new_n11317), .C(new_n11302), .Y(new_n11609));
  A2O1A1Ixp33_ASAP7_75t_L   g11353(.A1(new_n10976), .A2(new_n10975), .B(new_n11299), .C(new_n11296), .Y(new_n11610));
  INVx1_ASAP7_75t_L         g11354(.A(new_n11608), .Y(new_n11611));
  OAI21xp33_ASAP7_75t_L     g11355(.A1(new_n11602), .A2(new_n11606), .B(new_n11323), .Y(new_n11612));
  INVx1_ASAP7_75t_L         g11356(.A(new_n11612), .Y(new_n11613));
  A2O1A1Ixp33_ASAP7_75t_L   g11357(.A1(new_n11611), .A2(new_n11610), .B(new_n11613), .C(new_n11609), .Y(new_n11614));
  INVx1_ASAP7_75t_L         g11358(.A(new_n11614), .Y(new_n11615));
  O2A1O1Ixp33_ASAP7_75t_L   g11359(.A1(new_n11602), .A2(new_n11606), .B(new_n11323), .C(new_n11609), .Y(new_n11616));
  O2A1O1Ixp33_ASAP7_75t_L   g11360(.A1(new_n11608), .A2(new_n11323), .B(new_n11616), .C(new_n11615), .Y(\f[59] ));
  O2A1O1Ixp33_ASAP7_75t_L   g11361(.A1(new_n11613), .A2(new_n11610), .B(new_n11609), .C(new_n11608), .Y(new_n11618));
  A2O1A1Ixp33_ASAP7_75t_L   g11362(.A1(new_n11294), .A2(new_n11289), .B(new_n11584), .C(new_n11585), .Y(new_n11619));
  O2A1O1Ixp33_ASAP7_75t_L   g11363(.A1(new_n11324), .A2(new_n11584), .B(new_n11585), .C(new_n11582), .Y(new_n11620));
  O2A1O1Ixp33_ASAP7_75t_L   g11364(.A1(new_n11619), .A2(new_n11604), .B(new_n11601), .C(new_n11620), .Y(new_n11621));
  NOR2xp33_ASAP7_75t_L      g11365(.A(new_n11303), .B(new_n287), .Y(new_n11622));
  AOI221xp5_ASAP7_75t_L     g11366(.A1(\b[59] ), .A2(new_n264), .B1(\b[60] ), .B2(new_n283), .C(new_n11622), .Y(new_n11623));
  INVx1_ASAP7_75t_L         g11367(.A(new_n11592), .Y(new_n11624));
  NOR2xp33_ASAP7_75t_L      g11368(.A(\b[59] ), .B(\b[60] ), .Y(new_n11625));
  INVx1_ASAP7_75t_L         g11369(.A(\b[60] ), .Y(new_n11626));
  NOR2xp33_ASAP7_75t_L      g11370(.A(new_n11591), .B(new_n11626), .Y(new_n11627));
  NOR2xp33_ASAP7_75t_L      g11371(.A(new_n11625), .B(new_n11627), .Y(new_n11628));
  INVx1_ASAP7_75t_L         g11372(.A(new_n11628), .Y(new_n11629));
  O2A1O1Ixp33_ASAP7_75t_L   g11373(.A1(new_n11590), .A2(new_n11595), .B(new_n11624), .C(new_n11629), .Y(new_n11630));
  INVx1_ASAP7_75t_L         g11374(.A(new_n11630), .Y(new_n11631));
  A2O1A1O1Ixp25_ASAP7_75t_L g11375(.A1(new_n11309), .A2(new_n11312), .B(new_n11308), .C(new_n11593), .D(new_n11592), .Y(new_n11632));
  NAND2xp33_ASAP7_75t_L     g11376(.A(new_n11629), .B(new_n11632), .Y(new_n11633));
  NAND2xp33_ASAP7_75t_L     g11377(.A(new_n11631), .B(new_n11633), .Y(new_n11634));
  O2A1O1Ixp33_ASAP7_75t_L   g11378(.A1(new_n279), .A2(new_n11634), .B(new_n11623), .C(new_n257), .Y(new_n11635));
  OAI21xp33_ASAP7_75t_L     g11379(.A1(new_n279), .A2(new_n11634), .B(new_n11623), .Y(new_n11636));
  NAND2xp33_ASAP7_75t_L     g11380(.A(new_n257), .B(new_n11636), .Y(new_n11637));
  OAI21xp33_ASAP7_75t_L     g11381(.A1(new_n257), .A2(new_n11635), .B(new_n11637), .Y(new_n11638));
  INVx1_ASAP7_75t_L         g11382(.A(new_n11638), .Y(new_n11639));
  OAI22xp33_ASAP7_75t_L     g11383(.A1(new_n350), .A2(new_n10332), .B1(new_n10309), .B2(new_n375), .Y(new_n11640));
  AOI221xp5_ASAP7_75t_L     g11384(.A1(new_n361), .A2(\b[57] ), .B1(new_n359), .B2(new_n10991), .C(new_n11640), .Y(new_n11641));
  XNOR2x2_ASAP7_75t_L       g11385(.A(new_n346), .B(new_n11641), .Y(new_n11642));
  NAND2xp33_ASAP7_75t_L     g11386(.A(new_n11572), .B(new_n11571), .Y(new_n11643));
  MAJIxp5_ASAP7_75t_L       g11387(.A(new_n11324), .B(new_n11327), .C(new_n11643), .Y(new_n11644));
  OAI22xp33_ASAP7_75t_L     g11388(.A1(new_n513), .A2(new_n9683), .B1(new_n9355), .B2(new_n506), .Y(new_n11645));
  AOI221xp5_ASAP7_75t_L     g11389(.A1(new_n475), .A2(\b[54] ), .B1(new_n483), .B2(new_n9717), .C(new_n11645), .Y(new_n11646));
  XNOR2x2_ASAP7_75t_L       g11390(.A(new_n466), .B(new_n11646), .Y(new_n11647));
  INVx1_ASAP7_75t_L         g11391(.A(new_n11647), .Y(new_n11648));
  NOR2xp33_ASAP7_75t_L      g11392(.A(new_n8779), .B(new_n710), .Y(new_n11649));
  AOI221xp5_ASAP7_75t_L     g11393(.A1(\b[50] ), .A2(new_n635), .B1(\b[49] ), .B2(new_n713), .C(new_n11649), .Y(new_n11650));
  O2A1O1Ixp33_ASAP7_75t_L   g11394(.A1(new_n641), .A2(new_n8789), .B(new_n11650), .C(new_n637), .Y(new_n11651));
  NOR2xp33_ASAP7_75t_L      g11395(.A(new_n637), .B(new_n11651), .Y(new_n11652));
  O2A1O1Ixp33_ASAP7_75t_L   g11396(.A1(new_n641), .A2(new_n8789), .B(new_n11650), .C(\a[11] ), .Y(new_n11653));
  NOR2xp33_ASAP7_75t_L      g11397(.A(new_n11653), .B(new_n11652), .Y(new_n11654));
  INVx1_ASAP7_75t_L         g11398(.A(new_n11654), .Y(new_n11655));
  INVx1_ASAP7_75t_L         g11399(.A(new_n7868), .Y(new_n11656));
  NOR2xp33_ASAP7_75t_L      g11400(.A(new_n7552), .B(new_n864), .Y(new_n11657));
  AOI221xp5_ASAP7_75t_L     g11401(.A1(\b[46] ), .A2(new_n985), .B1(\b[48] ), .B2(new_n886), .C(new_n11657), .Y(new_n11658));
  INVx1_ASAP7_75t_L         g11402(.A(new_n11658), .Y(new_n11659));
  O2A1O1Ixp33_ASAP7_75t_L   g11403(.A1(new_n872), .A2(new_n7868), .B(new_n11658), .C(new_n867), .Y(new_n11660));
  INVx1_ASAP7_75t_L         g11404(.A(new_n11660), .Y(new_n11661));
  NOR2xp33_ASAP7_75t_L      g11405(.A(new_n867), .B(new_n11660), .Y(new_n11662));
  A2O1A1O1Ixp25_ASAP7_75t_L g11406(.A1(new_n11656), .A2(new_n873), .B(new_n11659), .C(new_n11661), .D(new_n11662), .Y(new_n11663));
  INVx1_ASAP7_75t_L         g11407(.A(new_n11663), .Y(new_n11664));
  MAJIxp5_ASAP7_75t_L       g11408(.A(new_n11255), .B(new_n11532), .C(new_n11543), .Y(new_n11665));
  NOR2xp33_ASAP7_75t_L      g11409(.A(new_n7249), .B(new_n1284), .Y(new_n11666));
  AOI221xp5_ASAP7_75t_L     g11410(.A1(\b[43] ), .A2(new_n1290), .B1(\b[44] ), .B2(new_n1204), .C(new_n11666), .Y(new_n11667));
  O2A1O1Ixp33_ASAP7_75t_L   g11411(.A1(new_n1210), .A2(new_n7255), .B(new_n11667), .C(new_n1206), .Y(new_n11668));
  OAI21xp33_ASAP7_75t_L     g11412(.A1(new_n1210), .A2(new_n7255), .B(new_n11667), .Y(new_n11669));
  NAND2xp33_ASAP7_75t_L     g11413(.A(new_n1206), .B(new_n11669), .Y(new_n11670));
  OAI21xp33_ASAP7_75t_L     g11414(.A1(new_n1206), .A2(new_n11668), .B(new_n11670), .Y(new_n11671));
  INVx1_ASAP7_75t_L         g11415(.A(new_n11500), .Y(new_n11672));
  INVx1_ASAP7_75t_L         g11416(.A(new_n11495), .Y(new_n11673));
  OAI21xp33_ASAP7_75t_L     g11417(.A1(new_n10859), .A2(new_n10862), .B(new_n10863), .Y(new_n11674));
  A2O1A1O1Ixp25_ASAP7_75t_L g11418(.A1(new_n11193), .A2(new_n11674), .B(new_n11196), .C(new_n11483), .D(new_n11488), .Y(new_n11675));
  NOR2xp33_ASAP7_75t_L      g11419(.A(new_n4101), .B(new_n2930), .Y(new_n11676));
  AOI221xp5_ASAP7_75t_L     g11420(.A1(\b[31] ), .A2(new_n3129), .B1(\b[32] ), .B2(new_n2936), .C(new_n11676), .Y(new_n11677));
  O2A1O1Ixp33_ASAP7_75t_L   g11421(.A1(new_n2940), .A2(new_n4108), .B(new_n11677), .C(new_n2928), .Y(new_n11678));
  OAI21xp33_ASAP7_75t_L     g11422(.A1(new_n2940), .A2(new_n4108), .B(new_n11677), .Y(new_n11679));
  NAND2xp33_ASAP7_75t_L     g11423(.A(new_n2928), .B(new_n11679), .Y(new_n11680));
  OAI21xp33_ASAP7_75t_L     g11424(.A1(new_n2928), .A2(new_n11678), .B(new_n11680), .Y(new_n11681));
  A2O1A1Ixp33_ASAP7_75t_L   g11425(.A1(new_n11476), .A2(new_n11190), .B(new_n11474), .C(new_n11477), .Y(new_n11682));
  A2O1A1Ixp33_ASAP7_75t_L   g11426(.A1(new_n10706), .A2(new_n10801), .B(new_n10820), .C(new_n11113), .Y(new_n11683));
  O2A1O1Ixp33_ASAP7_75t_L   g11427(.A1(new_n11128), .A2(new_n11126), .B(new_n11106), .C(new_n11100), .Y(new_n11684));
  O2A1O1Ixp33_ASAP7_75t_L   g11428(.A1(new_n11129), .A2(new_n11108), .B(new_n11127), .C(new_n11421), .Y(new_n11685));
  O2A1O1Ixp33_ASAP7_75t_L   g11429(.A1(new_n11684), .A2(new_n11685), .B(new_n11423), .C(new_n11417), .Y(new_n11686));
  INVx1_ASAP7_75t_L         g11430(.A(new_n11686), .Y(new_n11687));
  A2O1A1Ixp33_ASAP7_75t_L   g11431(.A1(new_n11116), .A2(new_n11683), .B(new_n11438), .C(new_n11687), .Y(new_n11688));
  NAND2xp33_ASAP7_75t_L     g11432(.A(\b[20] ), .B(new_n5623), .Y(new_n11689));
  OAI221xp5_ASAP7_75t_L     g11433(.A1(new_n5641), .A2(new_n1895), .B1(new_n1599), .B2(new_n5925), .C(new_n11689), .Y(new_n11690));
  A2O1A1Ixp33_ASAP7_75t_L   g11434(.A1(new_n2836), .A2(new_n5637), .B(new_n11690), .C(\a[41] ), .Y(new_n11691));
  AOI211xp5_ASAP7_75t_L     g11435(.A1(new_n2836), .A2(new_n5637), .B(new_n11690), .C(new_n5626), .Y(new_n11692));
  A2O1A1O1Ixp25_ASAP7_75t_L g11436(.A1(new_n5637), .A2(new_n2836), .B(new_n11690), .C(new_n11691), .D(new_n11692), .Y(new_n11693));
  NOR2xp33_ASAP7_75t_L      g11437(.A(new_n1150), .B(new_n6741), .Y(new_n11694));
  AOI221xp5_ASAP7_75t_L     g11438(.A1(\b[18] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[17] ), .C(new_n11694), .Y(new_n11695));
  O2A1O1Ixp33_ASAP7_75t_L   g11439(.A1(new_n6443), .A2(new_n1464), .B(new_n11695), .C(new_n6439), .Y(new_n11696));
  OAI21xp33_ASAP7_75t_L     g11440(.A1(new_n6443), .A2(new_n1464), .B(new_n11695), .Y(new_n11697));
  NAND2xp33_ASAP7_75t_L     g11441(.A(new_n6439), .B(new_n11697), .Y(new_n11698));
  OAI21xp33_ASAP7_75t_L     g11442(.A1(new_n6439), .A2(new_n11696), .B(new_n11698), .Y(new_n11699));
  INVx1_ASAP7_75t_L         g11443(.A(new_n11397), .Y(new_n11700));
  NAND3xp33_ASAP7_75t_L     g11444(.A(new_n11700), .B(new_n11391), .C(new_n11386), .Y(new_n11701));
  OAI22xp33_ASAP7_75t_L     g11445(.A1(new_n7614), .A2(new_n936), .B1(new_n960), .B2(new_n7312), .Y(new_n11702));
  AOI221xp5_ASAP7_75t_L     g11446(.A1(new_n7334), .A2(\b[15] ), .B1(new_n7322), .B2(new_n1052), .C(new_n11702), .Y(new_n11703));
  XNOR2x2_ASAP7_75t_L       g11447(.A(new_n7316), .B(new_n11703), .Y(new_n11704));
  NAND2xp33_ASAP7_75t_L     g11448(.A(new_n11082), .B(new_n11083), .Y(new_n11705));
  A2O1A1O1Ixp25_ASAP7_75t_L g11449(.A1(new_n11089), .A2(new_n11705), .B(new_n11387), .C(new_n11381), .D(new_n11390), .Y(new_n11706));
  NOR2xp33_ASAP7_75t_L      g11450(.A(new_n748), .B(new_n10065), .Y(new_n11707));
  AOI221xp5_ASAP7_75t_L     g11451(.A1(new_n8175), .A2(\b[12] ), .B1(new_n8484), .B2(\b[10] ), .C(new_n11707), .Y(new_n11708));
  O2A1O1Ixp33_ASAP7_75t_L   g11452(.A1(new_n8176), .A2(new_n841), .B(new_n11708), .C(new_n8172), .Y(new_n11709));
  NOR2xp33_ASAP7_75t_L      g11453(.A(new_n8172), .B(new_n11709), .Y(new_n11710));
  O2A1O1Ixp33_ASAP7_75t_L   g11454(.A1(new_n8176), .A2(new_n841), .B(new_n11708), .C(\a[50] ), .Y(new_n11711));
  NOR2xp33_ASAP7_75t_L      g11455(.A(new_n11711), .B(new_n11710), .Y(new_n11712));
  OR3x1_ASAP7_75t_L         g11456(.A(new_n11370), .B(new_n11374), .C(new_n11371), .Y(new_n11713));
  A2O1A1O1Ixp25_ASAP7_75t_L g11457(.A1(new_n11070), .A2(new_n11029), .B(new_n11077), .C(new_n11713), .D(new_n11376), .Y(new_n11714));
  O2A1O1Ixp33_ASAP7_75t_L   g11458(.A1(new_n11037), .A2(new_n11060), .B(new_n11061), .C(new_n11369), .Y(new_n11715));
  NAND4xp25_ASAP7_75t_L     g11459(.A(new_n11357), .B(\a[59] ), .C(new_n10734), .D(new_n11055), .Y(new_n11716));
  INVx1_ASAP7_75t_L         g11460(.A(\a[60] ), .Y(new_n11717));
  NAND2xp33_ASAP7_75t_L     g11461(.A(\a[59] ), .B(new_n11717), .Y(new_n11718));
  NAND2xp33_ASAP7_75t_L     g11462(.A(\a[60] ), .B(new_n11048), .Y(new_n11719));
  AND2x2_ASAP7_75t_L        g11463(.A(new_n11718), .B(new_n11719), .Y(new_n11720));
  NOR2xp33_ASAP7_75t_L      g11464(.A(new_n284), .B(new_n11720), .Y(new_n11721));
  NAND2xp33_ASAP7_75t_L     g11465(.A(new_n11721), .B(new_n11716), .Y(new_n11722));
  A2O1A1Ixp33_ASAP7_75t_L   g11466(.A1(new_n11718), .A2(new_n11719), .B(new_n284), .C(new_n11360), .Y(new_n11723));
  NAND2xp33_ASAP7_75t_L     g11467(.A(\b[3] ), .B(new_n11051), .Y(new_n11724));
  OAI221xp5_ASAP7_75t_L     g11468(.A1(new_n11352), .A2(new_n289), .B1(new_n262), .B2(new_n11354), .C(new_n11724), .Y(new_n11725));
  A2O1A1Ixp33_ASAP7_75t_L   g11469(.A1(new_n312), .A2(new_n11351), .B(new_n11725), .C(\a[59] ), .Y(new_n11726));
  AOI211xp5_ASAP7_75t_L     g11470(.A1(new_n312), .A2(new_n11351), .B(new_n11048), .C(new_n11725), .Y(new_n11727));
  A2O1A1O1Ixp25_ASAP7_75t_L g11471(.A1(new_n11351), .A2(new_n312), .B(new_n11725), .C(new_n11726), .D(new_n11727), .Y(new_n11728));
  AO21x2_ASAP7_75t_L        g11472(.A1(new_n11722), .A2(new_n11723), .B(new_n11728), .Y(new_n11729));
  NAND3xp33_ASAP7_75t_L     g11473(.A(new_n11723), .B(new_n11728), .C(new_n11722), .Y(new_n11730));
  NOR2xp33_ASAP7_75t_L      g11474(.A(new_n384), .B(new_n10388), .Y(new_n11731));
  AOI221xp5_ASAP7_75t_L     g11475(.A1(new_n10086), .A2(\b[6] ), .B1(new_n11361), .B2(\b[4] ), .C(new_n11731), .Y(new_n11732));
  O2A1O1Ixp33_ASAP7_75t_L   g11476(.A1(new_n10088), .A2(new_n434), .B(new_n11732), .C(new_n10083), .Y(new_n11733));
  OAI21xp33_ASAP7_75t_L     g11477(.A1(new_n10088), .A2(new_n434), .B(new_n11732), .Y(new_n11734));
  NAND2xp33_ASAP7_75t_L     g11478(.A(new_n10083), .B(new_n11734), .Y(new_n11735));
  OAI21xp33_ASAP7_75t_L     g11479(.A1(new_n10083), .A2(new_n11733), .B(new_n11735), .Y(new_n11736));
  INVx1_ASAP7_75t_L         g11480(.A(new_n11736), .Y(new_n11737));
  NAND3xp33_ASAP7_75t_L     g11481(.A(new_n11729), .B(new_n11730), .C(new_n11737), .Y(new_n11738));
  AO21x2_ASAP7_75t_L        g11482(.A1(new_n11730), .A2(new_n11729), .B(new_n11737), .Y(new_n11739));
  OAI211xp5_ASAP7_75t_L     g11483(.A1(new_n11368), .A2(new_n11715), .B(new_n11739), .C(new_n11738), .Y(new_n11740));
  OAI21xp33_ASAP7_75t_L     g11484(.A1(new_n11360), .A2(new_n11359), .B(new_n11367), .Y(new_n11741));
  A2O1A1O1Ixp25_ASAP7_75t_L g11485(.A1(new_n11068), .A2(new_n11064), .B(new_n11062), .C(new_n11741), .D(new_n11368), .Y(new_n11742));
  NAND3xp33_ASAP7_75t_L     g11486(.A(new_n11729), .B(new_n11730), .C(new_n11736), .Y(new_n11743));
  AND3x1_ASAP7_75t_L        g11487(.A(new_n11729), .B(new_n11737), .C(new_n11730), .Y(new_n11744));
  A2O1A1Ixp33_ASAP7_75t_L   g11488(.A1(new_n11736), .A2(new_n11743), .B(new_n11744), .C(new_n11742), .Y(new_n11745));
  NAND2xp33_ASAP7_75t_L     g11489(.A(\b[8] ), .B(new_n9096), .Y(new_n11746));
  OAI221xp5_ASAP7_75t_L     g11490(.A1(new_n9440), .A2(new_n448), .B1(new_n590), .B2(new_n9439), .C(new_n11746), .Y(new_n11747));
  A2O1A1Ixp33_ASAP7_75t_L   g11491(.A1(new_n602), .A2(new_n9437), .B(new_n11747), .C(\a[53] ), .Y(new_n11748));
  AOI211xp5_ASAP7_75t_L     g11492(.A1(new_n602), .A2(new_n9437), .B(new_n11747), .C(new_n9099), .Y(new_n11749));
  A2O1A1O1Ixp25_ASAP7_75t_L g11493(.A1(new_n9437), .A2(new_n602), .B(new_n11747), .C(new_n11748), .D(new_n11749), .Y(new_n11750));
  AOI21xp33_ASAP7_75t_L     g11494(.A1(new_n11745), .A2(new_n11740), .B(new_n11750), .Y(new_n11751));
  AND3x1_ASAP7_75t_L        g11495(.A(new_n11745), .B(new_n11740), .C(new_n11750), .Y(new_n11752));
  NOR3xp33_ASAP7_75t_L      g11496(.A(new_n11714), .B(new_n11751), .C(new_n11752), .Y(new_n11753));
  OA21x2_ASAP7_75t_L        g11497(.A1(new_n11751), .A2(new_n11752), .B(new_n11714), .Y(new_n11754));
  OAI21xp33_ASAP7_75t_L     g11498(.A1(new_n11753), .A2(new_n11754), .B(new_n11712), .Y(new_n11755));
  INVx1_ASAP7_75t_L         g11499(.A(new_n11755), .Y(new_n11756));
  NOR3xp33_ASAP7_75t_L      g11500(.A(new_n11754), .B(new_n11753), .C(new_n11712), .Y(new_n11757));
  NOR3xp33_ASAP7_75t_L      g11501(.A(new_n11756), .B(new_n11757), .C(new_n11706), .Y(new_n11758));
  A2O1A1Ixp33_ASAP7_75t_L   g11502(.A1(new_n11090), .A2(new_n11087), .B(new_n11389), .C(new_n11385), .Y(new_n11759));
  INVx1_ASAP7_75t_L         g11503(.A(new_n11757), .Y(new_n11760));
  AOI21xp33_ASAP7_75t_L     g11504(.A1(new_n11760), .A2(new_n11755), .B(new_n11759), .Y(new_n11761));
  NOR3xp33_ASAP7_75t_L      g11505(.A(new_n11761), .B(new_n11704), .C(new_n11758), .Y(new_n11762));
  XNOR2x2_ASAP7_75t_L       g11506(.A(\a[47] ), .B(new_n11703), .Y(new_n11763));
  NAND3xp33_ASAP7_75t_L     g11507(.A(new_n11760), .B(new_n11759), .C(new_n11755), .Y(new_n11764));
  OAI21xp33_ASAP7_75t_L     g11508(.A1(new_n11757), .A2(new_n11756), .B(new_n11706), .Y(new_n11765));
  AOI21xp33_ASAP7_75t_L     g11509(.A1(new_n11765), .A2(new_n11764), .B(new_n11763), .Y(new_n11766));
  AOI211xp5_ASAP7_75t_L     g11510(.A1(new_n11406), .A2(new_n11701), .B(new_n11766), .C(new_n11762), .Y(new_n11767));
  A2O1A1Ixp33_ASAP7_75t_L   g11511(.A1(new_n11398), .A2(new_n11397), .B(new_n11103), .C(new_n11701), .Y(new_n11768));
  NAND3xp33_ASAP7_75t_L     g11512(.A(new_n11763), .B(new_n11765), .C(new_n11764), .Y(new_n11769));
  OAI21xp33_ASAP7_75t_L     g11513(.A1(new_n11758), .A2(new_n11761), .B(new_n11704), .Y(new_n11770));
  AOI21xp33_ASAP7_75t_L     g11514(.A1(new_n11770), .A2(new_n11769), .B(new_n11768), .Y(new_n11771));
  OAI21xp33_ASAP7_75t_L     g11515(.A1(new_n11767), .A2(new_n11771), .B(new_n11699), .Y(new_n11772));
  NAND2xp33_ASAP7_75t_L     g11516(.A(new_n11406), .B(new_n11407), .Y(new_n11773));
  O2A1O1Ixp33_ASAP7_75t_L   g11517(.A1(new_n6439), .A2(new_n11339), .B(new_n11341), .C(new_n11773), .Y(new_n11774));
  A2O1A1O1Ixp25_ASAP7_75t_L g11518(.A1(new_n11105), .A2(new_n11106), .B(new_n11100), .C(new_n11409), .D(new_n11774), .Y(new_n11775));
  OA21x2_ASAP7_75t_L        g11519(.A1(new_n6439), .A2(new_n11696), .B(new_n11698), .Y(new_n11776));
  NAND3xp33_ASAP7_75t_L     g11520(.A(new_n11768), .B(new_n11769), .C(new_n11770), .Y(new_n11777));
  OAI211xp5_ASAP7_75t_L     g11521(.A1(new_n11766), .A2(new_n11762), .B(new_n11406), .C(new_n11701), .Y(new_n11778));
  NAND3xp33_ASAP7_75t_L     g11522(.A(new_n11777), .B(new_n11776), .C(new_n11778), .Y(new_n11779));
  AOI21xp33_ASAP7_75t_L     g11523(.A1(new_n11779), .A2(new_n11772), .B(new_n11775), .Y(new_n11780));
  A2O1A1Ixp33_ASAP7_75t_L   g11524(.A1(new_n11026), .A2(new_n11104), .B(new_n11108), .C(new_n11127), .Y(new_n11781));
  NOR2xp33_ASAP7_75t_L      g11525(.A(new_n11767), .B(new_n11771), .Y(new_n11782));
  AOI221xp5_ASAP7_75t_L     g11526(.A1(new_n11782), .A2(new_n11776), .B1(new_n11409), .B2(new_n11781), .C(new_n11774), .Y(new_n11783));
  AOI211xp5_ASAP7_75t_L     g11527(.A1(new_n11772), .A2(new_n11783), .B(new_n11693), .C(new_n11780), .Y(new_n11784));
  INVx1_ASAP7_75t_L         g11528(.A(new_n11693), .Y(new_n11785));
  NAND2xp33_ASAP7_75t_L     g11529(.A(new_n11779), .B(new_n11772), .Y(new_n11786));
  OAI21xp33_ASAP7_75t_L     g11530(.A1(new_n11774), .A2(new_n11685), .B(new_n11786), .Y(new_n11787));
  NAND3xp33_ASAP7_75t_L     g11531(.A(new_n11775), .B(new_n11772), .C(new_n11779), .Y(new_n11788));
  AOI21xp33_ASAP7_75t_L     g11532(.A1(new_n11787), .A2(new_n11788), .B(new_n11785), .Y(new_n11789));
  NOR2xp33_ASAP7_75t_L      g11533(.A(new_n11789), .B(new_n11784), .Y(new_n11790));
  NAND2xp33_ASAP7_75t_L     g11534(.A(new_n11688), .B(new_n11790), .Y(new_n11791));
  O2A1O1Ixp33_ASAP7_75t_L   g11535(.A1(new_n11115), .A2(new_n11140), .B(new_n11426), .C(new_n11686), .Y(new_n11792));
  OAI21xp33_ASAP7_75t_L     g11536(.A1(new_n11784), .A2(new_n11789), .B(new_n11792), .Y(new_n11793));
  OAI22xp33_ASAP7_75t_L     g11537(.A1(new_n5144), .A2(new_n2045), .B1(new_n2188), .B2(new_n4903), .Y(new_n11794));
  AOI221xp5_ASAP7_75t_L     g11538(.A1(new_n4917), .A2(\b[24] ), .B1(new_n4912), .B2(new_n2216), .C(new_n11794), .Y(new_n11795));
  XNOR2x2_ASAP7_75t_L       g11539(.A(new_n4906), .B(new_n11795), .Y(new_n11796));
  NAND3xp33_ASAP7_75t_L     g11540(.A(new_n11791), .B(new_n11793), .C(new_n11796), .Y(new_n11797));
  NOR3xp33_ASAP7_75t_L      g11541(.A(new_n11792), .B(new_n11784), .C(new_n11789), .Y(new_n11798));
  NAND3xp33_ASAP7_75t_L     g11542(.A(new_n11785), .B(new_n11787), .C(new_n11788), .Y(new_n11799));
  A2O1A1Ixp33_ASAP7_75t_L   g11543(.A1(new_n11783), .A2(new_n11772), .B(new_n11780), .C(new_n11693), .Y(new_n11800));
  AOI21xp33_ASAP7_75t_L     g11544(.A1(new_n11800), .A2(new_n11799), .B(new_n11688), .Y(new_n11801));
  XNOR2x2_ASAP7_75t_L       g11545(.A(\a[38] ), .B(new_n11795), .Y(new_n11802));
  OAI21xp33_ASAP7_75t_L     g11546(.A1(new_n11801), .A2(new_n11798), .B(new_n11802), .Y(new_n11803));
  A2O1A1O1Ixp25_ASAP7_75t_L g11547(.A1(new_n11145), .A2(new_n11445), .B(new_n11333), .C(new_n11442), .D(new_n11446), .Y(new_n11804));
  NAND3xp33_ASAP7_75t_L     g11548(.A(new_n11804), .B(new_n11803), .C(new_n11797), .Y(new_n11805));
  INVx1_ASAP7_75t_L         g11549(.A(new_n11334), .Y(new_n11806));
  NAND2xp33_ASAP7_75t_L     g11550(.A(new_n11797), .B(new_n11803), .Y(new_n11807));
  A2O1A1Ixp33_ASAP7_75t_L   g11551(.A1(new_n11442), .A2(new_n11806), .B(new_n11446), .C(new_n11807), .Y(new_n11808));
  OAI22xp33_ASAP7_75t_L     g11552(.A1(new_n4397), .A2(new_n2377), .B1(new_n2703), .B2(new_n4142), .Y(new_n11809));
  AOI221xp5_ASAP7_75t_L     g11553(.A1(new_n4156), .A2(\b[27] ), .B1(new_n4151), .B2(new_n2887), .C(new_n11809), .Y(new_n11810));
  XNOR2x2_ASAP7_75t_L       g11554(.A(new_n4145), .B(new_n11810), .Y(new_n11811));
  NAND3xp33_ASAP7_75t_L     g11555(.A(new_n11808), .B(new_n11805), .C(new_n11811), .Y(new_n11812));
  A2O1A1Ixp33_ASAP7_75t_L   g11556(.A1(new_n11146), .A2(new_n11142), .B(new_n11443), .C(new_n11435), .Y(new_n11813));
  NOR2xp33_ASAP7_75t_L      g11557(.A(new_n11807), .B(new_n11813), .Y(new_n11814));
  NAND3xp33_ASAP7_75t_L     g11558(.A(new_n11791), .B(new_n11793), .C(new_n11802), .Y(new_n11815));
  INVx1_ASAP7_75t_L         g11559(.A(new_n11815), .Y(new_n11816));
  O2A1O1Ixp33_ASAP7_75t_L   g11560(.A1(new_n11796), .A2(new_n11816), .B(new_n11797), .C(new_n11804), .Y(new_n11817));
  XNOR2x2_ASAP7_75t_L       g11561(.A(\a[35] ), .B(new_n11810), .Y(new_n11818));
  OAI21xp33_ASAP7_75t_L     g11562(.A1(new_n11814), .A2(new_n11817), .B(new_n11818), .Y(new_n11819));
  NAND2xp33_ASAP7_75t_L     g11563(.A(new_n11812), .B(new_n11819), .Y(new_n11820));
  NAND3xp33_ASAP7_75t_L     g11564(.A(new_n11449), .B(new_n11444), .C(new_n11456), .Y(new_n11821));
  A2O1A1Ixp33_ASAP7_75t_L   g11565(.A1(new_n11176), .A2(new_n11161), .B(new_n11461), .C(new_n11821), .Y(new_n11822));
  NOR2xp33_ASAP7_75t_L      g11566(.A(new_n11820), .B(new_n11822), .Y(new_n11823));
  NAND3xp33_ASAP7_75t_L     g11567(.A(new_n11808), .B(new_n11805), .C(new_n11818), .Y(new_n11824));
  NOR3xp33_ASAP7_75t_L      g11568(.A(new_n11817), .B(new_n11814), .C(new_n11818), .Y(new_n11825));
  AOI21xp33_ASAP7_75t_L     g11569(.A1(new_n11824), .A2(new_n11818), .B(new_n11825), .Y(new_n11826));
  INVx1_ASAP7_75t_L         g11570(.A(new_n11821), .Y(new_n11827));
  A2O1A1O1Ixp25_ASAP7_75t_L g11571(.A1(new_n11156), .A2(new_n11159), .B(new_n11162), .C(new_n11458), .D(new_n11827), .Y(new_n11828));
  NOR2xp33_ASAP7_75t_L      g11572(.A(new_n11828), .B(new_n11826), .Y(new_n11829));
  OAI22xp33_ASAP7_75t_L     g11573(.A1(new_n3703), .A2(new_n3079), .B1(new_n3098), .B2(new_n3509), .Y(new_n11830));
  AOI221xp5_ASAP7_75t_L     g11574(.A1(new_n3503), .A2(\b[30] ), .B1(new_n3505), .B2(new_n4813), .C(new_n11830), .Y(new_n11831));
  XNOR2x2_ASAP7_75t_L       g11575(.A(new_n3493), .B(new_n11831), .Y(new_n11832));
  OAI21xp33_ASAP7_75t_L     g11576(.A1(new_n11829), .A2(new_n11823), .B(new_n11832), .Y(new_n11833));
  NAND2xp33_ASAP7_75t_L     g11577(.A(new_n11828), .B(new_n11826), .Y(new_n11834));
  A2O1A1Ixp33_ASAP7_75t_L   g11578(.A1(new_n11458), .A2(new_n11459), .B(new_n11827), .C(new_n11820), .Y(new_n11835));
  INVx1_ASAP7_75t_L         g11579(.A(new_n11832), .Y(new_n11836));
  NAND3xp33_ASAP7_75t_L     g11580(.A(new_n11836), .B(new_n11834), .C(new_n11835), .Y(new_n11837));
  NAND3xp33_ASAP7_75t_L     g11581(.A(new_n11682), .B(new_n11833), .C(new_n11837), .Y(new_n11838));
  INVx1_ASAP7_75t_L         g11582(.A(new_n11190), .Y(new_n11839));
  NAND2xp33_ASAP7_75t_L     g11583(.A(new_n11182), .B(new_n11183), .Y(new_n11840));
  A2O1A1O1Ixp25_ASAP7_75t_L g11584(.A1(new_n11181), .A2(new_n11840), .B(new_n11839), .C(new_n11478), .D(new_n11470), .Y(new_n11841));
  AOI21xp33_ASAP7_75t_L     g11585(.A1(new_n11834), .A2(new_n11835), .B(new_n11836), .Y(new_n11842));
  NOR3xp33_ASAP7_75t_L      g11586(.A(new_n11823), .B(new_n11829), .C(new_n11832), .Y(new_n11843));
  OAI21xp33_ASAP7_75t_L     g11587(.A1(new_n11842), .A2(new_n11843), .B(new_n11841), .Y(new_n11844));
  NAND3xp33_ASAP7_75t_L     g11588(.A(new_n11838), .B(new_n11844), .C(new_n11681), .Y(new_n11845));
  NOR3xp33_ASAP7_75t_L      g11589(.A(new_n11841), .B(new_n11842), .C(new_n11843), .Y(new_n11846));
  AOI21xp33_ASAP7_75t_L     g11590(.A1(new_n11837), .A2(new_n11833), .B(new_n11682), .Y(new_n11847));
  NOR3xp33_ASAP7_75t_L      g11591(.A(new_n11846), .B(new_n11847), .C(new_n11681), .Y(new_n11848));
  AOI211xp5_ASAP7_75t_L     g11592(.A1(new_n11681), .A2(new_n11845), .B(new_n11675), .C(new_n11848), .Y(new_n11849));
  OAI21xp33_ASAP7_75t_L     g11593(.A1(new_n11487), .A2(new_n11486), .B(new_n11484), .Y(new_n11850));
  INVx1_ASAP7_75t_L         g11594(.A(new_n11681), .Y(new_n11851));
  NAND3xp33_ASAP7_75t_L     g11595(.A(new_n11838), .B(new_n11844), .C(new_n11851), .Y(new_n11852));
  OAI21xp33_ASAP7_75t_L     g11596(.A1(new_n11847), .A2(new_n11846), .B(new_n11681), .Y(new_n11853));
  AOI21xp33_ASAP7_75t_L     g11597(.A1(new_n11853), .A2(new_n11852), .B(new_n11850), .Y(new_n11854));
  OAI22xp33_ASAP7_75t_L     g11598(.A1(new_n2572), .A2(new_n4344), .B1(new_n4581), .B2(new_n2410), .Y(new_n11855));
  AOI221xp5_ASAP7_75t_L     g11599(.A1(new_n2423), .A2(\b[36] ), .B1(new_n2417), .B2(new_n4621), .C(new_n11855), .Y(new_n11856));
  XNOR2x2_ASAP7_75t_L       g11600(.A(new_n2413), .B(new_n11856), .Y(new_n11857));
  INVx1_ASAP7_75t_L         g11601(.A(new_n11857), .Y(new_n11858));
  OAI21xp33_ASAP7_75t_L     g11602(.A1(new_n11854), .A2(new_n11849), .B(new_n11858), .Y(new_n11859));
  NAND3xp33_ASAP7_75t_L     g11603(.A(new_n11850), .B(new_n11852), .C(new_n11853), .Y(new_n11860));
  A2O1A1Ixp33_ASAP7_75t_L   g11604(.A1(new_n11681), .A2(new_n11845), .B(new_n11848), .C(new_n11675), .Y(new_n11861));
  NAND3xp33_ASAP7_75t_L     g11605(.A(new_n11860), .B(new_n11861), .C(new_n11857), .Y(new_n11862));
  NAND2xp33_ASAP7_75t_L     g11606(.A(new_n11862), .B(new_n11859), .Y(new_n11863));
  OAI211xp5_ASAP7_75t_L     g11607(.A1(new_n11673), .A2(new_n11501), .B(new_n11863), .C(new_n11672), .Y(new_n11864));
  AOI21xp33_ASAP7_75t_L     g11608(.A1(new_n11860), .A2(new_n11861), .B(new_n11857), .Y(new_n11865));
  NOR3xp33_ASAP7_75t_L      g11609(.A(new_n11849), .B(new_n11858), .C(new_n11854), .Y(new_n11866));
  NOR2xp33_ASAP7_75t_L      g11610(.A(new_n11865), .B(new_n11866), .Y(new_n11867));
  A2O1A1Ixp33_ASAP7_75t_L   g11611(.A1(new_n11495), .A2(new_n11496), .B(new_n11500), .C(new_n11867), .Y(new_n11868));
  INVx1_ASAP7_75t_L         g11612(.A(new_n5578), .Y(new_n11869));
  NAND2xp33_ASAP7_75t_L     g11613(.A(\b[39] ), .B(new_n1955), .Y(new_n11870));
  OAI221xp5_ASAP7_75t_L     g11614(.A1(new_n1962), .A2(new_n5311), .B1(new_n5074), .B2(new_n2089), .C(new_n11870), .Y(new_n11871));
  A2O1A1Ixp33_ASAP7_75t_L   g11615(.A1(new_n11869), .A2(new_n1964), .B(new_n11871), .C(\a[23] ), .Y(new_n11872));
  AOI211xp5_ASAP7_75t_L     g11616(.A1(new_n11869), .A2(new_n1964), .B(new_n11871), .C(new_n1952), .Y(new_n11873));
  A2O1A1O1Ixp25_ASAP7_75t_L g11617(.A1(new_n11869), .A2(new_n1964), .B(new_n11871), .C(new_n11872), .D(new_n11873), .Y(new_n11874));
  NAND3xp33_ASAP7_75t_L     g11618(.A(new_n11868), .B(new_n11864), .C(new_n11874), .Y(new_n11875));
  A2O1A1Ixp33_ASAP7_75t_L   g11619(.A1(new_n11493), .A2(new_n11494), .B(new_n11501), .C(new_n11672), .Y(new_n11876));
  NOR2xp33_ASAP7_75t_L      g11620(.A(new_n11867), .B(new_n11876), .Y(new_n11877));
  O2A1O1Ixp33_ASAP7_75t_L   g11621(.A1(new_n11501), .A2(new_n11673), .B(new_n11672), .C(new_n11863), .Y(new_n11878));
  INVx1_ASAP7_75t_L         g11622(.A(new_n11874), .Y(new_n11879));
  OAI21xp33_ASAP7_75t_L     g11623(.A1(new_n11878), .A2(new_n11877), .B(new_n11879), .Y(new_n11880));
  INVx1_ASAP7_75t_L         g11624(.A(new_n11505), .Y(new_n11881));
  NOR3xp33_ASAP7_75t_L      g11625(.A(new_n11881), .B(new_n11497), .C(new_n11502), .Y(new_n11882));
  O2A1O1Ixp33_ASAP7_75t_L   g11626(.A1(new_n11506), .A2(new_n11505), .B(new_n11510), .C(new_n11882), .Y(new_n11883));
  NAND3xp33_ASAP7_75t_L     g11627(.A(new_n11883), .B(new_n11880), .C(new_n11875), .Y(new_n11884));
  NAND2xp33_ASAP7_75t_L     g11628(.A(new_n11880), .B(new_n11875), .Y(new_n11885));
  OAI21xp33_ASAP7_75t_L     g11629(.A1(new_n11882), .A2(new_n11512), .B(new_n11885), .Y(new_n11886));
  OAI22xp33_ASAP7_75t_L     g11630(.A1(new_n1654), .A2(new_n5855), .B1(new_n6110), .B2(new_n1517), .Y(new_n11887));
  AOI221xp5_ASAP7_75t_L     g11631(.A1(new_n1511), .A2(\b[42] ), .B1(new_n1513), .B2(new_n6389), .C(new_n11887), .Y(new_n11888));
  XNOR2x2_ASAP7_75t_L       g11632(.A(\a[20] ), .B(new_n11888), .Y(new_n11889));
  AOI21xp33_ASAP7_75t_L     g11633(.A1(new_n11886), .A2(new_n11884), .B(new_n11889), .Y(new_n11890));
  INVx1_ASAP7_75t_L         g11634(.A(new_n11882), .Y(new_n11891));
  OAI21xp33_ASAP7_75t_L     g11635(.A1(new_n11506), .A2(new_n11507), .B(new_n11510), .Y(new_n11892));
  AND4x1_ASAP7_75t_L        g11636(.A(new_n11892), .B(new_n11891), .C(new_n11880), .D(new_n11875), .Y(new_n11893));
  AOI21xp33_ASAP7_75t_L     g11637(.A1(new_n11880), .A2(new_n11875), .B(new_n11883), .Y(new_n11894));
  INVx1_ASAP7_75t_L         g11638(.A(new_n11889), .Y(new_n11895));
  NOR3xp33_ASAP7_75t_L      g11639(.A(new_n11895), .B(new_n11893), .C(new_n11894), .Y(new_n11896));
  NOR3xp33_ASAP7_75t_L      g11640(.A(new_n11525), .B(new_n11890), .C(new_n11896), .Y(new_n11897));
  OAI21xp33_ASAP7_75t_L     g11641(.A1(new_n11894), .A2(new_n11893), .B(new_n11895), .Y(new_n11898));
  NAND3xp33_ASAP7_75t_L     g11642(.A(new_n11886), .B(new_n11884), .C(new_n11889), .Y(new_n11899));
  AOI221xp5_ASAP7_75t_L     g11643(.A1(new_n11899), .A2(new_n11898), .B1(new_n11520), .B2(new_n11534), .C(new_n11521), .Y(new_n11900));
  OAI21xp33_ASAP7_75t_L     g11644(.A1(new_n11897), .A2(new_n11900), .B(new_n11671), .Y(new_n11901));
  INVx1_ASAP7_75t_L         g11645(.A(new_n11671), .Y(new_n11902));
  OAI211xp5_ASAP7_75t_L     g11646(.A1(new_n11521), .A2(new_n11553), .B(new_n11898), .C(new_n11899), .Y(new_n11903));
  OAI21xp33_ASAP7_75t_L     g11647(.A1(new_n11890), .A2(new_n11896), .B(new_n11525), .Y(new_n11904));
  NAND3xp33_ASAP7_75t_L     g11648(.A(new_n11903), .B(new_n11904), .C(new_n11902), .Y(new_n11905));
  NAND2xp33_ASAP7_75t_L     g11649(.A(new_n11901), .B(new_n11905), .Y(new_n11906));
  AOI21xp33_ASAP7_75t_L     g11650(.A1(new_n11903), .A2(new_n11904), .B(new_n11902), .Y(new_n11907));
  NOR3xp33_ASAP7_75t_L      g11651(.A(new_n11900), .B(new_n11897), .C(new_n11671), .Y(new_n11908));
  NOR3xp33_ASAP7_75t_L      g11652(.A(new_n11665), .B(new_n11907), .C(new_n11908), .Y(new_n11909));
  A2O1A1Ixp33_ASAP7_75t_L   g11653(.A1(new_n11665), .A2(new_n11906), .B(new_n11909), .C(new_n11664), .Y(new_n11910));
  A2O1A1O1Ixp25_ASAP7_75t_L g11654(.A1(new_n11267), .A2(new_n11272), .B(new_n11264), .C(new_n11560), .D(new_n11563), .Y(new_n11911));
  NAND2xp33_ASAP7_75t_L     g11655(.A(new_n11906), .B(new_n11665), .Y(new_n11912));
  OAI211xp5_ASAP7_75t_L     g11656(.A1(new_n11255), .A2(new_n11556), .B(new_n11544), .C(new_n11905), .Y(new_n11913));
  OAI211xp5_ASAP7_75t_L     g11657(.A1(new_n11907), .A2(new_n11913), .B(new_n11912), .C(new_n11663), .Y(new_n11914));
  AOI21xp33_ASAP7_75t_L     g11658(.A1(new_n11914), .A2(new_n11910), .B(new_n11911), .Y(new_n11915));
  AOI211xp5_ASAP7_75t_L     g11659(.A1(new_n11540), .A2(new_n11263), .B(new_n11908), .C(new_n11545), .Y(new_n11916));
  AOI221xp5_ASAP7_75t_L     g11660(.A1(new_n11665), .A2(new_n11906), .B1(new_n11901), .B2(new_n11916), .C(new_n11664), .Y(new_n11917));
  AOI211xp5_ASAP7_75t_L     g11661(.A1(new_n11560), .A2(new_n11330), .B(new_n11563), .C(new_n11917), .Y(new_n11918));
  A2O1A1Ixp33_ASAP7_75t_L   g11662(.A1(new_n11918), .A2(new_n11910), .B(new_n11915), .C(new_n11655), .Y(new_n11919));
  INVx1_ASAP7_75t_L         g11663(.A(new_n11919), .Y(new_n11920));
  NAND2xp33_ASAP7_75t_L     g11664(.A(new_n11565), .B(new_n11561), .Y(new_n11921));
  MAJIxp5_ASAP7_75t_L       g11665(.A(new_n11329), .B(new_n11568), .C(new_n11921), .Y(new_n11922));
  O2A1O1Ixp33_ASAP7_75t_L   g11666(.A1(new_n11907), .A2(new_n11913), .B(new_n11912), .C(new_n11663), .Y(new_n11923));
  NOR2xp33_ASAP7_75t_L      g11667(.A(new_n11917), .B(new_n11923), .Y(new_n11924));
  OAI211xp5_ASAP7_75t_L     g11668(.A1(new_n11562), .A2(new_n11564), .B(new_n11914), .C(new_n11551), .Y(new_n11925));
  OAI221xp5_ASAP7_75t_L     g11669(.A1(new_n11924), .A2(new_n11911), .B1(new_n11925), .B2(new_n11923), .C(new_n11655), .Y(new_n11926));
  OAI21xp33_ASAP7_75t_L     g11670(.A1(new_n11564), .A2(new_n11562), .B(new_n11551), .Y(new_n11927));
  NAND2xp33_ASAP7_75t_L     g11671(.A(new_n11914), .B(new_n11910), .Y(new_n11928));
  AOI221xp5_ASAP7_75t_L     g11672(.A1(new_n11928), .A2(new_n11927), .B1(new_n11910), .B2(new_n11918), .C(new_n11655), .Y(new_n11929));
  A2O1A1Ixp33_ASAP7_75t_L   g11673(.A1(new_n11655), .A2(new_n11926), .B(new_n11929), .C(new_n11922), .Y(new_n11930));
  OR2x4_ASAP7_75t_L         g11674(.A(new_n11568), .B(new_n11921), .Y(new_n11931));
  OAI221xp5_ASAP7_75t_L     g11675(.A1(new_n11924), .A2(new_n11911), .B1(new_n11925), .B2(new_n11923), .C(new_n11654), .Y(new_n11932));
  NAND3xp33_ASAP7_75t_L     g11676(.A(new_n11571), .B(new_n11931), .C(new_n11932), .Y(new_n11933));
  OAI211xp5_ASAP7_75t_L     g11677(.A1(new_n11920), .A2(new_n11933), .B(new_n11930), .C(new_n11648), .Y(new_n11934));
  INVx1_ASAP7_75t_L         g11678(.A(new_n11930), .Y(new_n11935));
  NOR2xp33_ASAP7_75t_L      g11679(.A(new_n11929), .B(new_n11922), .Y(new_n11936));
  A2O1A1Ixp33_ASAP7_75t_L   g11680(.A1(new_n11936), .A2(new_n11919), .B(new_n11935), .C(new_n11647), .Y(new_n11937));
  AND3x1_ASAP7_75t_L        g11681(.A(new_n11644), .B(new_n11937), .C(new_n11934), .Y(new_n11938));
  AOI21xp33_ASAP7_75t_L     g11682(.A1(new_n11937), .A2(new_n11934), .B(new_n11644), .Y(new_n11939));
  NOR3xp33_ASAP7_75t_L      g11683(.A(new_n11938), .B(new_n11939), .C(new_n11642), .Y(new_n11940));
  INVx1_ASAP7_75t_L         g11684(.A(new_n11642), .Y(new_n11941));
  NAND3xp33_ASAP7_75t_L     g11685(.A(new_n11644), .B(new_n11934), .C(new_n11937), .Y(new_n11942));
  AO21x2_ASAP7_75t_L        g11686(.A1(new_n11937), .A2(new_n11934), .B(new_n11644), .Y(new_n11943));
  AOI21xp33_ASAP7_75t_L     g11687(.A1(new_n11943), .A2(new_n11942), .B(new_n11941), .Y(new_n11944));
  NOR3xp33_ASAP7_75t_L      g11688(.A(new_n11940), .B(new_n11944), .C(new_n11639), .Y(new_n11945));
  NAND3xp33_ASAP7_75t_L     g11689(.A(new_n11943), .B(new_n11942), .C(new_n11941), .Y(new_n11946));
  OAI21xp33_ASAP7_75t_L     g11690(.A1(new_n11939), .A2(new_n11938), .B(new_n11642), .Y(new_n11947));
  AOI21xp33_ASAP7_75t_L     g11691(.A1(new_n11947), .A2(new_n11946), .B(new_n11638), .Y(new_n11948));
  NOR3xp33_ASAP7_75t_L      g11692(.A(new_n11945), .B(new_n11948), .C(new_n11621), .Y(new_n11949));
  OAI21xp33_ASAP7_75t_L     g11693(.A1(new_n11948), .A2(new_n11945), .B(new_n11621), .Y(new_n11950));
  INVx1_ASAP7_75t_L         g11694(.A(new_n11950), .Y(new_n11951));
  NOR2xp33_ASAP7_75t_L      g11695(.A(new_n11949), .B(new_n11951), .Y(new_n11952));
  XNOR2x2_ASAP7_75t_L       g11696(.A(new_n11618), .B(new_n11952), .Y(\f[60] ));
  INVx1_ASAP7_75t_L         g11697(.A(new_n11618), .Y(new_n11954));
  A2O1A1Ixp33_ASAP7_75t_L   g11698(.A1(new_n11656), .A2(new_n873), .B(new_n11659), .C(new_n867), .Y(new_n11955));
  NAND3xp33_ASAP7_75t_L     g11699(.A(new_n11903), .B(new_n11904), .C(new_n11671), .Y(new_n11956));
  A2O1A1Ixp33_ASAP7_75t_L   g11700(.A1(new_n11671), .A2(new_n11956), .B(new_n11913), .C(new_n11912), .Y(new_n11957));
  O2A1O1Ixp33_ASAP7_75t_L   g11701(.A1(new_n867), .A2(new_n11660), .B(new_n11955), .C(new_n11957), .Y(new_n11958));
  O2A1O1Ixp33_ASAP7_75t_L   g11702(.A1(new_n11958), .A2(new_n11663), .B(new_n11918), .C(new_n11915), .Y(new_n11959));
  OAI22xp33_ASAP7_75t_L     g11703(.A1(new_n1550), .A2(new_n8779), .B1(new_n8755), .B2(new_n712), .Y(new_n11960));
  AOI221xp5_ASAP7_75t_L     g11704(.A1(new_n640), .A2(\b[52] ), .B1(new_n718), .B2(new_n9367), .C(new_n11960), .Y(new_n11961));
  XNOR2x2_ASAP7_75t_L       g11705(.A(new_n637), .B(new_n11961), .Y(new_n11962));
  INVx1_ASAP7_75t_L         g11706(.A(new_n11962), .Y(new_n11963));
  OAI22xp33_ASAP7_75t_L     g11707(.A1(new_n980), .A2(new_n7552), .B1(new_n7860), .B2(new_n864), .Y(new_n11964));
  AOI221xp5_ASAP7_75t_L     g11708(.A1(new_n886), .A2(\b[49] ), .B1(new_n873), .B2(new_n8438), .C(new_n11964), .Y(new_n11965));
  XNOR2x2_ASAP7_75t_L       g11709(.A(new_n867), .B(new_n11965), .Y(new_n11966));
  A2O1A1Ixp33_ASAP7_75t_L   g11710(.A1(new_n11234), .A2(new_n11231), .B(new_n11524), .C(new_n11520), .Y(new_n11967));
  A2O1A1Ixp33_ASAP7_75t_L   g11711(.A1(new_n11967), .A2(new_n11522), .B(new_n11890), .C(new_n11899), .Y(new_n11968));
  A2O1A1Ixp33_ASAP7_75t_L   g11712(.A1(new_n11852), .A2(new_n11851), .B(new_n11675), .C(new_n11845), .Y(new_n11969));
  A2O1A1O1Ixp25_ASAP7_75t_L g11713(.A1(new_n11332), .A2(new_n11478), .B(new_n11470), .C(new_n11833), .D(new_n11843), .Y(new_n11970));
  NAND2xp33_ASAP7_75t_L     g11714(.A(new_n11699), .B(new_n11782), .Y(new_n11971));
  A2O1A1Ixp33_ASAP7_75t_L   g11715(.A1(new_n11738), .A2(new_n11737), .B(new_n11742), .C(new_n11743), .Y(new_n11972));
  NOR2xp33_ASAP7_75t_L      g11716(.A(new_n427), .B(new_n10388), .Y(new_n11973));
  AOI221xp5_ASAP7_75t_L     g11717(.A1(new_n10086), .A2(\b[7] ), .B1(new_n11361), .B2(\b[5] ), .C(new_n11973), .Y(new_n11974));
  O2A1O1Ixp33_ASAP7_75t_L   g11718(.A1(new_n10088), .A2(new_n456), .B(new_n11974), .C(new_n10083), .Y(new_n11975));
  OAI21xp33_ASAP7_75t_L     g11719(.A1(new_n10088), .A2(new_n456), .B(new_n11974), .Y(new_n11976));
  NAND2xp33_ASAP7_75t_L     g11720(.A(new_n10083), .B(new_n11976), .Y(new_n11977));
  OAI21xp33_ASAP7_75t_L     g11721(.A1(new_n10083), .A2(new_n11975), .B(new_n11977), .Y(new_n11978));
  INVx1_ASAP7_75t_L         g11722(.A(new_n11978), .Y(new_n11979));
  INVx1_ASAP7_75t_L         g11723(.A(new_n11721), .Y(new_n11980));
  MAJx2_ASAP7_75t_L         g11724(.A(new_n11728), .B(new_n11980), .C(new_n11716), .Y(new_n11981));
  NAND2xp33_ASAP7_75t_L     g11725(.A(\b[4] ), .B(new_n11051), .Y(new_n11982));
  OAI221xp5_ASAP7_75t_L     g11726(.A1(new_n11352), .A2(new_n301), .B1(new_n289), .B2(new_n11354), .C(new_n11982), .Y(new_n11983));
  A2O1A1Ixp33_ASAP7_75t_L   g11727(.A1(new_n342), .A2(new_n11351), .B(new_n11983), .C(\a[59] ), .Y(new_n11984));
  AOI21xp33_ASAP7_75t_L     g11728(.A1(new_n342), .A2(new_n11351), .B(new_n11983), .Y(new_n11985));
  NOR2xp33_ASAP7_75t_L      g11729(.A(\a[59] ), .B(new_n11985), .Y(new_n11986));
  INVx1_ASAP7_75t_L         g11730(.A(\a[62] ), .Y(new_n11987));
  NOR2xp33_ASAP7_75t_L      g11731(.A(new_n11987), .B(new_n11721), .Y(new_n11988));
  XNOR2x2_ASAP7_75t_L       g11732(.A(\a[61] ), .B(\a[60] ), .Y(new_n11989));
  INVx1_ASAP7_75t_L         g11733(.A(new_n11989), .Y(new_n11990));
  INVx1_ASAP7_75t_L         g11734(.A(\a[61] ), .Y(new_n11991));
  NAND2xp33_ASAP7_75t_L     g11735(.A(\a[62] ), .B(new_n11991), .Y(new_n11992));
  NAND2xp33_ASAP7_75t_L     g11736(.A(\a[61] ), .B(new_n11987), .Y(new_n11993));
  NAND2xp33_ASAP7_75t_L     g11737(.A(new_n11993), .B(new_n11992), .Y(new_n11994));
  NOR2xp33_ASAP7_75t_L      g11738(.A(new_n11994), .B(new_n11720), .Y(new_n11995));
  AOI32xp33_ASAP7_75t_L     g11739(.A1(new_n11990), .A2(new_n11720), .A3(\b[0] ), .B1(new_n11995), .B2(\b[1] ), .Y(new_n11996));
  AOI21xp33_ASAP7_75t_L     g11740(.A1(new_n11993), .A2(new_n11992), .B(new_n11720), .Y(new_n11997));
  INVx1_ASAP7_75t_L         g11741(.A(new_n11997), .Y(new_n11998));
  O2A1O1Ixp33_ASAP7_75t_L   g11742(.A1(new_n11998), .A2(new_n274), .B(new_n11996), .C(new_n11987), .Y(new_n11999));
  INVx1_ASAP7_75t_L         g11743(.A(new_n11999), .Y(new_n12000));
  O2A1O1Ixp33_ASAP7_75t_L   g11744(.A1(new_n11998), .A2(new_n274), .B(new_n11996), .C(\a[62] ), .Y(new_n12001));
  A2O1A1Ixp33_ASAP7_75t_L   g11745(.A1(new_n12000), .A2(\a[62] ), .B(new_n12001), .C(new_n11988), .Y(new_n12002));
  INVx1_ASAP7_75t_L         g11746(.A(new_n12001), .Y(new_n12003));
  A2O1A1Ixp33_ASAP7_75t_L   g11747(.A1(new_n11721), .A2(new_n11999), .B(new_n11987), .C(new_n12003), .Y(new_n12004));
  AOI221xp5_ASAP7_75t_L     g11748(.A1(\a[59] ), .A2(new_n11984), .B1(new_n12004), .B2(new_n12002), .C(new_n11986), .Y(new_n12005));
  NOR2xp33_ASAP7_75t_L      g11749(.A(new_n11048), .B(new_n11985), .Y(new_n12006));
  A2O1A1Ixp33_ASAP7_75t_L   g11750(.A1(new_n342), .A2(new_n11351), .B(new_n11983), .C(new_n11048), .Y(new_n12007));
  NAND2xp33_ASAP7_75t_L     g11751(.A(new_n12004), .B(new_n12002), .Y(new_n12008));
  O2A1O1Ixp33_ASAP7_75t_L   g11752(.A1(new_n11048), .A2(new_n12006), .B(new_n12007), .C(new_n12008), .Y(new_n12009));
  NOR3xp33_ASAP7_75t_L      g11753(.A(new_n12009), .B(new_n12005), .C(new_n11981), .Y(new_n12010));
  INVx1_ASAP7_75t_L         g11754(.A(new_n11981), .Y(new_n12011));
  INVx1_ASAP7_75t_L         g11755(.A(new_n12005), .Y(new_n12012));
  A2O1A1Ixp33_ASAP7_75t_L   g11756(.A1(new_n11718), .A2(new_n11719), .B(new_n284), .C(\a[62] ), .Y(new_n12013));
  O2A1O1Ixp33_ASAP7_75t_L   g11757(.A1(new_n11999), .A2(new_n11987), .B(new_n12003), .C(new_n12013), .Y(new_n12014));
  O2A1O1Ixp33_ASAP7_75t_L   g11758(.A1(new_n11980), .A2(new_n12000), .B(\a[62] ), .C(new_n12001), .Y(new_n12015));
  NOR2xp33_ASAP7_75t_L      g11759(.A(new_n12014), .B(new_n12015), .Y(new_n12016));
  A2O1A1Ixp33_ASAP7_75t_L   g11760(.A1(new_n11984), .A2(\a[59] ), .B(new_n11986), .C(new_n12016), .Y(new_n12017));
  AOI21xp33_ASAP7_75t_L     g11761(.A1(new_n12017), .A2(new_n12012), .B(new_n12011), .Y(new_n12018));
  OAI21xp33_ASAP7_75t_L     g11762(.A1(new_n12010), .A2(new_n12018), .B(new_n11979), .Y(new_n12019));
  NAND3xp33_ASAP7_75t_L     g11763(.A(new_n12011), .B(new_n12017), .C(new_n12012), .Y(new_n12020));
  OAI21xp33_ASAP7_75t_L     g11764(.A1(new_n12005), .A2(new_n12009), .B(new_n11981), .Y(new_n12021));
  NAND3xp33_ASAP7_75t_L     g11765(.A(new_n12020), .B(new_n11978), .C(new_n12021), .Y(new_n12022));
  NAND3xp33_ASAP7_75t_L     g11766(.A(new_n11972), .B(new_n12019), .C(new_n12022), .Y(new_n12023));
  AO21x2_ASAP7_75t_L        g11767(.A1(new_n12022), .A2(new_n12019), .B(new_n11972), .Y(new_n12024));
  OAI22xp33_ASAP7_75t_L     g11768(.A1(new_n9440), .A2(new_n534), .B1(new_n590), .B2(new_n10400), .Y(new_n12025));
  AOI221xp5_ASAP7_75t_L     g11769(.A1(new_n9102), .A2(\b[10] ), .B1(new_n9437), .B2(new_n690), .C(new_n12025), .Y(new_n12026));
  XNOR2x2_ASAP7_75t_L       g11770(.A(new_n9099), .B(new_n12026), .Y(new_n12027));
  AND3x1_ASAP7_75t_L        g11771(.A(new_n12024), .B(new_n12027), .C(new_n12023), .Y(new_n12028));
  AOI21xp33_ASAP7_75t_L     g11772(.A1(new_n12024), .A2(new_n12023), .B(new_n12027), .Y(new_n12029));
  INVx1_ASAP7_75t_L         g11773(.A(new_n11751), .Y(new_n12030));
  OAI21xp33_ASAP7_75t_L     g11774(.A1(new_n11752), .A2(new_n11714), .B(new_n12030), .Y(new_n12031));
  NOR3xp33_ASAP7_75t_L      g11775(.A(new_n12031), .B(new_n12029), .C(new_n12028), .Y(new_n12032));
  NAND3xp33_ASAP7_75t_L     g11776(.A(new_n12024), .B(new_n12023), .C(new_n12027), .Y(new_n12033));
  AO21x2_ASAP7_75t_L        g11777(.A1(new_n12023), .A2(new_n12024), .B(new_n12027), .Y(new_n12034));
  NAND3xp33_ASAP7_75t_L     g11778(.A(new_n11745), .B(new_n11740), .C(new_n11750), .Y(new_n12035));
  A2O1A1O1Ixp25_ASAP7_75t_L g11779(.A1(new_n11713), .A2(new_n11378), .B(new_n11376), .C(new_n12035), .D(new_n11751), .Y(new_n12036));
  AOI21xp33_ASAP7_75t_L     g11780(.A1(new_n12034), .A2(new_n12033), .B(new_n12036), .Y(new_n12037));
  OAI22xp33_ASAP7_75t_L     g11781(.A1(new_n8483), .A2(new_n748), .B1(new_n833), .B2(new_n10065), .Y(new_n12038));
  AOI221xp5_ASAP7_75t_L     g11782(.A1(new_n8175), .A2(\b[13] ), .B1(new_n8490), .B2(new_n1166), .C(new_n12038), .Y(new_n12039));
  XNOR2x2_ASAP7_75t_L       g11783(.A(new_n8172), .B(new_n12039), .Y(new_n12040));
  OAI21xp33_ASAP7_75t_L     g11784(.A1(new_n12037), .A2(new_n12032), .B(new_n12040), .Y(new_n12041));
  A2O1A1O1Ixp25_ASAP7_75t_L g11785(.A1(new_n11381), .A2(new_n11345), .B(new_n11390), .C(new_n11755), .D(new_n11757), .Y(new_n12042));
  NAND3xp33_ASAP7_75t_L     g11786(.A(new_n12034), .B(new_n12036), .C(new_n12033), .Y(new_n12043));
  INVx1_ASAP7_75t_L         g11787(.A(new_n12027), .Y(new_n12044));
  NAND3xp33_ASAP7_75t_L     g11788(.A(new_n12024), .B(new_n12023), .C(new_n12044), .Y(new_n12045));
  A2O1A1Ixp33_ASAP7_75t_L   g11789(.A1(new_n12045), .A2(new_n12044), .B(new_n12028), .C(new_n12031), .Y(new_n12046));
  INVx1_ASAP7_75t_L         g11790(.A(new_n12040), .Y(new_n12047));
  NAND3xp33_ASAP7_75t_L     g11791(.A(new_n12047), .B(new_n12046), .C(new_n12043), .Y(new_n12048));
  AOI21xp33_ASAP7_75t_L     g11792(.A1(new_n12048), .A2(new_n12041), .B(new_n12042), .Y(new_n12049));
  NOR3xp33_ASAP7_75t_L      g11793(.A(new_n12032), .B(new_n12037), .C(new_n12040), .Y(new_n12050));
  A2O1A1O1Ixp25_ASAP7_75t_L g11794(.A1(new_n11755), .A2(new_n11759), .B(new_n11757), .C(new_n12041), .D(new_n12050), .Y(new_n12051));
  OAI22xp33_ASAP7_75t_L     g11795(.A1(new_n7614), .A2(new_n960), .B1(new_n1043), .B2(new_n7312), .Y(new_n12052));
  AOI221xp5_ASAP7_75t_L     g11796(.A1(new_n7334), .A2(\b[16] ), .B1(new_n7322), .B2(new_n1156), .C(new_n12052), .Y(new_n12053));
  XNOR2x2_ASAP7_75t_L       g11797(.A(\a[47] ), .B(new_n12053), .Y(new_n12054));
  A2O1A1Ixp33_ASAP7_75t_L   g11798(.A1(new_n12051), .A2(new_n12041), .B(new_n12049), .C(new_n12054), .Y(new_n12055));
  XNOR2x2_ASAP7_75t_L       g11799(.A(new_n7316), .B(new_n12053), .Y(new_n12056));
  AOI211xp5_ASAP7_75t_L     g11800(.A1(new_n12051), .A2(new_n12041), .B(new_n12049), .C(new_n12056), .Y(new_n12057));
  A2O1A1O1Ixp25_ASAP7_75t_L g11801(.A1(new_n12041), .A2(new_n12051), .B(new_n12049), .C(new_n12055), .D(new_n12057), .Y(new_n12058));
  A2O1A1Ixp33_ASAP7_75t_L   g11802(.A1(new_n11406), .A2(new_n11701), .B(new_n11766), .C(new_n11769), .Y(new_n12059));
  INVx1_ASAP7_75t_L         g11803(.A(new_n12059), .Y(new_n12060));
  NAND2xp33_ASAP7_75t_L     g11804(.A(new_n12060), .B(new_n12058), .Y(new_n12061));
  AOI21xp33_ASAP7_75t_L     g11805(.A1(new_n12046), .A2(new_n12043), .B(new_n12047), .Y(new_n12062));
  O2A1O1Ixp33_ASAP7_75t_L   g11806(.A1(new_n11706), .A2(new_n11756), .B(new_n11760), .C(new_n12062), .Y(new_n12063));
  NAND3xp33_ASAP7_75t_L     g11807(.A(new_n12042), .B(new_n12048), .C(new_n12041), .Y(new_n12064));
  A2O1A1Ixp33_ASAP7_75t_L   g11808(.A1(new_n12063), .A2(new_n12048), .B(new_n12042), .C(new_n12064), .Y(new_n12065));
  A2O1A1Ixp33_ASAP7_75t_L   g11809(.A1(new_n12055), .A2(new_n12065), .B(new_n12057), .C(new_n12059), .Y(new_n12066));
  OAI22xp33_ASAP7_75t_L     g11810(.A1(new_n7304), .A2(new_n1458), .B1(new_n1349), .B2(new_n6741), .Y(new_n12067));
  AOI221xp5_ASAP7_75t_L     g11811(.A1(new_n6442), .A2(\b[19] ), .B1(new_n6450), .B2(new_n1607), .C(new_n12067), .Y(new_n12068));
  XNOR2x2_ASAP7_75t_L       g11812(.A(\a[44] ), .B(new_n12068), .Y(new_n12069));
  NAND3xp33_ASAP7_75t_L     g11813(.A(new_n12061), .B(new_n12066), .C(new_n12069), .Y(new_n12070));
  A2O1A1O1Ixp25_ASAP7_75t_L g11814(.A1(new_n12048), .A2(new_n12063), .B(new_n12042), .C(new_n12064), .D(new_n12056), .Y(new_n12071));
  A2O1A1Ixp33_ASAP7_75t_L   g11815(.A1(new_n12051), .A2(new_n12041), .B(new_n12049), .C(new_n12056), .Y(new_n12072));
  OAI21xp33_ASAP7_75t_L     g11816(.A1(new_n12056), .A2(new_n12071), .B(new_n12072), .Y(new_n12073));
  NOR2xp33_ASAP7_75t_L      g11817(.A(new_n12059), .B(new_n12073), .Y(new_n12074));
  INVx1_ASAP7_75t_L         g11818(.A(new_n12066), .Y(new_n12075));
  INVx1_ASAP7_75t_L         g11819(.A(new_n12069), .Y(new_n12076));
  OAI21xp33_ASAP7_75t_L     g11820(.A1(new_n12075), .A2(new_n12074), .B(new_n12076), .Y(new_n12077));
  AOI22xp33_ASAP7_75t_L     g11821(.A1(new_n12070), .A2(new_n12077), .B1(new_n11971), .B2(new_n11787), .Y(new_n12078));
  A2O1A1Ixp33_ASAP7_75t_L   g11822(.A1(new_n11772), .A2(new_n11779), .B(new_n11775), .C(new_n11971), .Y(new_n12079));
  NOR3xp33_ASAP7_75t_L      g11823(.A(new_n12076), .B(new_n12075), .C(new_n12074), .Y(new_n12080));
  AOI21xp33_ASAP7_75t_L     g11824(.A1(new_n12061), .A2(new_n12066), .B(new_n12069), .Y(new_n12081));
  NOR3xp33_ASAP7_75t_L      g11825(.A(new_n12079), .B(new_n12080), .C(new_n12081), .Y(new_n12082));
  OAI22xp33_ASAP7_75t_L     g11826(.A1(new_n5640), .A2(new_n1895), .B1(new_n1745), .B2(new_n5925), .Y(new_n12083));
  AOI221xp5_ASAP7_75t_L     g11827(.A1(new_n5629), .A2(\b[22] ), .B1(new_n5637), .B2(new_n2056), .C(new_n12083), .Y(new_n12084));
  XNOR2x2_ASAP7_75t_L       g11828(.A(new_n5626), .B(new_n12084), .Y(new_n12085));
  OAI21xp33_ASAP7_75t_L     g11829(.A1(new_n12078), .A2(new_n12082), .B(new_n12085), .Y(new_n12086));
  A2O1A1O1Ixp25_ASAP7_75t_L g11830(.A1(new_n11779), .A2(new_n11776), .B(new_n11775), .C(new_n11971), .D(new_n12081), .Y(new_n12087));
  OAI21xp33_ASAP7_75t_L     g11831(.A1(new_n12081), .A2(new_n12080), .B(new_n12079), .Y(new_n12088));
  XNOR2x2_ASAP7_75t_L       g11832(.A(\a[41] ), .B(new_n12084), .Y(new_n12089));
  OAI311xp33_ASAP7_75t_L    g11833(.A1(new_n12087), .A2(new_n12081), .A3(new_n12080), .B1(new_n12089), .C1(new_n12088), .Y(new_n12090));
  A2O1A1Ixp33_ASAP7_75t_L   g11834(.A1(new_n10463), .A2(new_n10370), .B(new_n10465), .C(new_n10801), .Y(new_n12091));
  A2O1A1Ixp33_ASAP7_75t_L   g11835(.A1(new_n12091), .A2(new_n10809), .B(new_n11133), .C(new_n11116), .Y(new_n12092));
  A2O1A1O1Ixp25_ASAP7_75t_L g11836(.A1(new_n11426), .A2(new_n12092), .B(new_n11686), .C(new_n11800), .D(new_n11784), .Y(new_n12093));
  NAND3xp33_ASAP7_75t_L     g11837(.A(new_n12093), .B(new_n12090), .C(new_n12086), .Y(new_n12094));
  NAND2xp33_ASAP7_75t_L     g11838(.A(new_n12090), .B(new_n12086), .Y(new_n12095));
  A2O1A1Ixp33_ASAP7_75t_L   g11839(.A1(new_n11113), .A2(new_n11125), .B(new_n11115), .C(new_n11426), .Y(new_n12096));
  A2O1A1Ixp33_ASAP7_75t_L   g11840(.A1(new_n12096), .A2(new_n11687), .B(new_n11789), .C(new_n11799), .Y(new_n12097));
  NAND2xp33_ASAP7_75t_L     g11841(.A(new_n12097), .B(new_n12095), .Y(new_n12098));
  OAI22xp33_ASAP7_75t_L     g11842(.A1(new_n5144), .A2(new_n2188), .B1(new_n2205), .B2(new_n4903), .Y(new_n12099));
  AOI221xp5_ASAP7_75t_L     g11843(.A1(new_n4917), .A2(\b[25] ), .B1(new_n4912), .B2(new_n5001), .C(new_n12099), .Y(new_n12100));
  XNOR2x2_ASAP7_75t_L       g11844(.A(new_n4906), .B(new_n12100), .Y(new_n12101));
  NAND3xp33_ASAP7_75t_L     g11845(.A(new_n12094), .B(new_n12098), .C(new_n12101), .Y(new_n12102));
  NOR2xp33_ASAP7_75t_L      g11846(.A(new_n12097), .B(new_n12095), .Y(new_n12103));
  A2O1A1O1Ixp25_ASAP7_75t_L g11847(.A1(new_n11782), .A2(new_n11699), .B(new_n11780), .C(new_n12077), .D(new_n12080), .Y(new_n12104));
  A2O1A1O1Ixp25_ASAP7_75t_L g11848(.A1(new_n12066), .A2(new_n12061), .B(new_n12069), .C(new_n12104), .D(new_n12078), .Y(new_n12105));
  A2O1A1Ixp33_ASAP7_75t_L   g11849(.A1(new_n11787), .A2(new_n11971), .B(new_n12081), .C(new_n12070), .Y(new_n12106));
  O2A1O1Ixp33_ASAP7_75t_L   g11850(.A1(new_n12081), .A2(new_n12106), .B(new_n12088), .C(new_n12085), .Y(new_n12107));
  O2A1O1Ixp33_ASAP7_75t_L   g11851(.A1(new_n12105), .A2(new_n12107), .B(new_n12090), .C(new_n12093), .Y(new_n12108));
  XNOR2x2_ASAP7_75t_L       g11852(.A(\a[38] ), .B(new_n12100), .Y(new_n12109));
  OAI21xp33_ASAP7_75t_L     g11853(.A1(new_n12103), .A2(new_n12108), .B(new_n12109), .Y(new_n12110));
  NAND2xp33_ASAP7_75t_L     g11854(.A(new_n12102), .B(new_n12110), .Y(new_n12111));
  A2O1A1Ixp33_ASAP7_75t_L   g11855(.A1(new_n11796), .A2(new_n11797), .B(new_n11804), .C(new_n11815), .Y(new_n12112));
  NOR2xp33_ASAP7_75t_L      g11856(.A(new_n12111), .B(new_n12112), .Y(new_n12113));
  NOR3xp33_ASAP7_75t_L      g11857(.A(new_n12108), .B(new_n12103), .C(new_n12109), .Y(new_n12114));
  AOI21xp33_ASAP7_75t_L     g11858(.A1(new_n12094), .A2(new_n12098), .B(new_n12101), .Y(new_n12115));
  NOR2xp33_ASAP7_75t_L      g11859(.A(new_n12115), .B(new_n12114), .Y(new_n12116));
  O2A1O1Ixp33_ASAP7_75t_L   g11860(.A1(new_n11446), .A2(new_n11455), .B(new_n11807), .C(new_n11816), .Y(new_n12117));
  NOR2xp33_ASAP7_75t_L      g11861(.A(new_n12117), .B(new_n12116), .Y(new_n12118));
  NOR2xp33_ASAP7_75t_L      g11862(.A(new_n12113), .B(new_n12118), .Y(new_n12119));
  NAND2xp33_ASAP7_75t_L     g11863(.A(new_n12117), .B(new_n12116), .Y(new_n12120));
  NAND2xp33_ASAP7_75t_L     g11864(.A(new_n12111), .B(new_n12112), .Y(new_n12121));
  NOR2xp33_ASAP7_75t_L      g11865(.A(new_n3079), .B(new_n4147), .Y(new_n12122));
  AOI221xp5_ASAP7_75t_L     g11866(.A1(\b[26] ), .A2(new_n4402), .B1(\b[27] ), .B2(new_n4155), .C(new_n12122), .Y(new_n12123));
  O2A1O1Ixp33_ASAP7_75t_L   g11867(.A1(new_n4150), .A2(new_n3087), .B(new_n12123), .C(new_n4145), .Y(new_n12124));
  OAI21xp33_ASAP7_75t_L     g11868(.A1(new_n4150), .A2(new_n3087), .B(new_n12123), .Y(new_n12125));
  NAND2xp33_ASAP7_75t_L     g11869(.A(new_n4145), .B(new_n12125), .Y(new_n12126));
  OAI21xp33_ASAP7_75t_L     g11870(.A1(new_n4145), .A2(new_n12124), .B(new_n12126), .Y(new_n12127));
  NAND3xp33_ASAP7_75t_L     g11871(.A(new_n12120), .B(new_n12121), .C(new_n12127), .Y(new_n12128));
  INVx1_ASAP7_75t_L         g11872(.A(new_n12127), .Y(new_n12129));
  AOI21xp33_ASAP7_75t_L     g11873(.A1(new_n12120), .A2(new_n12121), .B(new_n12129), .Y(new_n12130));
  AOI21xp33_ASAP7_75t_L     g11874(.A1(new_n12128), .A2(new_n12119), .B(new_n12130), .Y(new_n12131));
  NAND3xp33_ASAP7_75t_L     g11875(.A(new_n12131), .B(new_n11835), .C(new_n11824), .Y(new_n12132));
  NAND3xp33_ASAP7_75t_L     g11876(.A(new_n12120), .B(new_n12121), .C(new_n12129), .Y(new_n12133));
  OAI21xp33_ASAP7_75t_L     g11877(.A1(new_n12113), .A2(new_n12118), .B(new_n12127), .Y(new_n12134));
  NAND2xp33_ASAP7_75t_L     g11878(.A(new_n12133), .B(new_n12134), .Y(new_n12135));
  A2O1A1Ixp33_ASAP7_75t_L   g11879(.A1(new_n11811), .A2(new_n11812), .B(new_n11828), .C(new_n11824), .Y(new_n12136));
  NAND2xp33_ASAP7_75t_L     g11880(.A(new_n12135), .B(new_n12136), .Y(new_n12137));
  OAI22xp33_ASAP7_75t_L     g11881(.A1(new_n3703), .A2(new_n3098), .B1(new_n3456), .B2(new_n3509), .Y(new_n12138));
  AOI221xp5_ASAP7_75t_L     g11882(.A1(new_n3503), .A2(\b[31] ), .B1(new_n3505), .B2(new_n4317), .C(new_n12138), .Y(new_n12139));
  XNOR2x2_ASAP7_75t_L       g11883(.A(new_n3493), .B(new_n12139), .Y(new_n12140));
  NAND3xp33_ASAP7_75t_L     g11884(.A(new_n12132), .B(new_n12137), .C(new_n12140), .Y(new_n12141));
  INVx1_ASAP7_75t_L         g11885(.A(new_n12141), .Y(new_n12142));
  AOI21xp33_ASAP7_75t_L     g11886(.A1(new_n12132), .A2(new_n12137), .B(new_n12140), .Y(new_n12143));
  NOR3xp33_ASAP7_75t_L      g11887(.A(new_n12142), .B(new_n12143), .C(new_n11970), .Y(new_n12144));
  A2O1A1Ixp33_ASAP7_75t_L   g11888(.A1(new_n11840), .A2(new_n11181), .B(new_n11839), .C(new_n11478), .Y(new_n12145));
  A2O1A1Ixp33_ASAP7_75t_L   g11889(.A1(new_n12145), .A2(new_n11477), .B(new_n11842), .C(new_n11837), .Y(new_n12146));
  NOR2xp33_ASAP7_75t_L      g11890(.A(new_n12135), .B(new_n12136), .Y(new_n12147));
  O2A1O1Ixp33_ASAP7_75t_L   g11891(.A1(new_n11826), .A2(new_n11828), .B(new_n11824), .C(new_n12131), .Y(new_n12148));
  INVx1_ASAP7_75t_L         g11892(.A(new_n12140), .Y(new_n12149));
  OAI21xp33_ASAP7_75t_L     g11893(.A1(new_n12147), .A2(new_n12148), .B(new_n12149), .Y(new_n12150));
  AOI21xp33_ASAP7_75t_L     g11894(.A1(new_n12150), .A2(new_n12141), .B(new_n12146), .Y(new_n12151));
  OAI22xp33_ASAP7_75t_L     g11895(.A1(new_n3133), .A2(new_n3891), .B1(new_n4101), .B2(new_n2925), .Y(new_n12152));
  AOI221xp5_ASAP7_75t_L     g11896(.A1(new_n2938), .A2(\b[34] ), .B1(new_n2932), .B2(new_n5599), .C(new_n12152), .Y(new_n12153));
  XNOR2x2_ASAP7_75t_L       g11897(.A(new_n2928), .B(new_n12153), .Y(new_n12154));
  INVx1_ASAP7_75t_L         g11898(.A(new_n12154), .Y(new_n12155));
  OAI21xp33_ASAP7_75t_L     g11899(.A1(new_n12151), .A2(new_n12144), .B(new_n12155), .Y(new_n12156));
  NAND3xp33_ASAP7_75t_L     g11900(.A(new_n12146), .B(new_n12141), .C(new_n12150), .Y(new_n12157));
  OAI21xp33_ASAP7_75t_L     g11901(.A1(new_n12143), .A2(new_n12142), .B(new_n11970), .Y(new_n12158));
  NAND3xp33_ASAP7_75t_L     g11902(.A(new_n12158), .B(new_n12157), .C(new_n12154), .Y(new_n12159));
  AOI21xp33_ASAP7_75t_L     g11903(.A1(new_n12156), .A2(new_n12159), .B(new_n11969), .Y(new_n12160));
  INVx1_ASAP7_75t_L         g11904(.A(new_n12160), .Y(new_n12161));
  NAND3xp33_ASAP7_75t_L     g11905(.A(new_n12156), .B(new_n11969), .C(new_n12159), .Y(new_n12162));
  OAI22xp33_ASAP7_75t_L     g11906(.A1(new_n2572), .A2(new_n4581), .B1(new_n4613), .B2(new_n2410), .Y(new_n12163));
  AOI221xp5_ASAP7_75t_L     g11907(.A1(new_n2423), .A2(\b[37] ), .B1(new_n2417), .B2(new_n10229), .C(new_n12163), .Y(new_n12164));
  XNOR2x2_ASAP7_75t_L       g11908(.A(new_n2413), .B(new_n12164), .Y(new_n12165));
  NAND3xp33_ASAP7_75t_L     g11909(.A(new_n12161), .B(new_n12162), .C(new_n12165), .Y(new_n12166));
  INVx1_ASAP7_75t_L         g11910(.A(new_n12162), .Y(new_n12167));
  INVx1_ASAP7_75t_L         g11911(.A(new_n12165), .Y(new_n12168));
  OAI21xp33_ASAP7_75t_L     g11912(.A1(new_n12160), .A2(new_n12167), .B(new_n12168), .Y(new_n12169));
  A2O1A1O1Ixp25_ASAP7_75t_L g11913(.A1(new_n11495), .A2(new_n11496), .B(new_n11500), .C(new_n11862), .D(new_n11865), .Y(new_n12170));
  NAND3xp33_ASAP7_75t_L     g11914(.A(new_n12170), .B(new_n12169), .C(new_n12166), .Y(new_n12171));
  AO21x2_ASAP7_75t_L        g11915(.A1(new_n12166), .A2(new_n12169), .B(new_n12170), .Y(new_n12172));
  OAI22xp33_ASAP7_75t_L     g11916(.A1(new_n2089), .A2(new_n5311), .B1(new_n5570), .B2(new_n1962), .Y(new_n12173));
  AOI221xp5_ASAP7_75t_L     g11917(.A1(new_n1955), .A2(\b[40] ), .B1(new_n1964), .B2(new_n6651), .C(new_n12173), .Y(new_n12174));
  XNOR2x2_ASAP7_75t_L       g11918(.A(new_n1952), .B(new_n12174), .Y(new_n12175));
  NAND3xp33_ASAP7_75t_L     g11919(.A(new_n12172), .B(new_n12171), .C(new_n12175), .Y(new_n12176));
  AND3x1_ASAP7_75t_L        g11920(.A(new_n12170), .B(new_n12169), .C(new_n12166), .Y(new_n12177));
  AOI21xp33_ASAP7_75t_L     g11921(.A1(new_n12169), .A2(new_n12166), .B(new_n12170), .Y(new_n12178));
  XNOR2x2_ASAP7_75t_L       g11922(.A(\a[23] ), .B(new_n12174), .Y(new_n12179));
  OAI21xp33_ASAP7_75t_L     g11923(.A1(new_n12178), .A2(new_n12177), .B(new_n12179), .Y(new_n12180));
  NAND2xp33_ASAP7_75t_L     g11924(.A(new_n12176), .B(new_n12180), .Y(new_n12181));
  NAND3xp33_ASAP7_75t_L     g11925(.A(new_n11879), .B(new_n11868), .C(new_n11864), .Y(new_n12182));
  A2O1A1Ixp33_ASAP7_75t_L   g11926(.A1(new_n11875), .A2(new_n11880), .B(new_n11883), .C(new_n12182), .Y(new_n12183));
  NOR2xp33_ASAP7_75t_L      g11927(.A(new_n12183), .B(new_n12181), .Y(new_n12184));
  NAND2xp33_ASAP7_75t_L     g11928(.A(new_n11864), .B(new_n11868), .Y(new_n12185));
  NAND3xp33_ASAP7_75t_L     g11929(.A(new_n12172), .B(new_n12171), .C(new_n12179), .Y(new_n12186));
  NOR3xp33_ASAP7_75t_L      g11930(.A(new_n12177), .B(new_n12178), .C(new_n12179), .Y(new_n12187));
  AOI21xp33_ASAP7_75t_L     g11931(.A1(new_n12186), .A2(new_n12179), .B(new_n12187), .Y(new_n12188));
  O2A1O1Ixp33_ASAP7_75t_L   g11932(.A1(new_n12185), .A2(new_n11874), .B(new_n11886), .C(new_n12188), .Y(new_n12189));
  OAI22xp33_ASAP7_75t_L     g11933(.A1(new_n1654), .A2(new_n6110), .B1(new_n6378), .B2(new_n1517), .Y(new_n12190));
  AOI221xp5_ASAP7_75t_L     g11934(.A1(new_n1511), .A2(\b[43] ), .B1(new_n1513), .B2(new_n6682), .C(new_n12190), .Y(new_n12191));
  XNOR2x2_ASAP7_75t_L       g11935(.A(new_n1501), .B(new_n12191), .Y(new_n12192));
  NOR3xp33_ASAP7_75t_L      g11936(.A(new_n12189), .B(new_n12192), .C(new_n12184), .Y(new_n12193));
  NAND3xp33_ASAP7_75t_L     g11937(.A(new_n12188), .B(new_n11886), .C(new_n12182), .Y(new_n12194));
  A2O1A1Ixp33_ASAP7_75t_L   g11938(.A1(new_n12186), .A2(new_n12179), .B(new_n12187), .C(new_n12183), .Y(new_n12195));
  INVx1_ASAP7_75t_L         g11939(.A(new_n12192), .Y(new_n12196));
  AOI21xp33_ASAP7_75t_L     g11940(.A1(new_n12194), .A2(new_n12195), .B(new_n12196), .Y(new_n12197));
  OAI21xp33_ASAP7_75t_L     g11941(.A1(new_n12197), .A2(new_n12193), .B(new_n11968), .Y(new_n12198));
  A2O1A1O1Ixp25_ASAP7_75t_L g11942(.A1(new_n11520), .A2(new_n11534), .B(new_n11521), .C(new_n11898), .D(new_n11896), .Y(new_n12199));
  NAND3xp33_ASAP7_75t_L     g11943(.A(new_n12194), .B(new_n12195), .C(new_n12196), .Y(new_n12200));
  OAI21xp33_ASAP7_75t_L     g11944(.A1(new_n12184), .A2(new_n12189), .B(new_n12192), .Y(new_n12201));
  NAND3xp33_ASAP7_75t_L     g11945(.A(new_n12199), .B(new_n12200), .C(new_n12201), .Y(new_n12202));
  OAI22xp33_ASAP7_75t_L     g11946(.A1(new_n1285), .A2(new_n6944), .B1(new_n7249), .B2(new_n2118), .Y(new_n12203));
  AOI221xp5_ASAP7_75t_L     g11947(.A1(new_n1209), .A2(\b[46] ), .B1(new_n1216), .B2(new_n7278), .C(new_n12203), .Y(new_n12204));
  XNOR2x2_ASAP7_75t_L       g11948(.A(new_n1206), .B(new_n12204), .Y(new_n12205));
  NAND3xp33_ASAP7_75t_L     g11949(.A(new_n12202), .B(new_n12198), .C(new_n12205), .Y(new_n12206));
  AOI21xp33_ASAP7_75t_L     g11950(.A1(new_n12201), .A2(new_n12200), .B(new_n12199), .Y(new_n12207));
  NOR3xp33_ASAP7_75t_L      g11951(.A(new_n11968), .B(new_n12193), .C(new_n12197), .Y(new_n12208));
  INVx1_ASAP7_75t_L         g11952(.A(new_n12205), .Y(new_n12209));
  OAI21xp33_ASAP7_75t_L     g11953(.A1(new_n12208), .A2(new_n12207), .B(new_n12209), .Y(new_n12210));
  NAND2xp33_ASAP7_75t_L     g11954(.A(new_n12206), .B(new_n12210), .Y(new_n12211));
  AOI21xp33_ASAP7_75t_L     g11955(.A1(new_n11912), .A2(new_n11956), .B(new_n12211), .Y(new_n12212));
  INVx1_ASAP7_75t_L         g11956(.A(new_n11956), .Y(new_n12213));
  AOI221xp5_ASAP7_75t_L     g11957(.A1(new_n11665), .A2(new_n11906), .B1(new_n12206), .B2(new_n12210), .C(new_n12213), .Y(new_n12214));
  OAI21xp33_ASAP7_75t_L     g11958(.A1(new_n12214), .A2(new_n12212), .B(new_n11966), .Y(new_n12215));
  INVx1_ASAP7_75t_L         g11959(.A(new_n11966), .Y(new_n12216));
  MAJIxp5_ASAP7_75t_L       g11960(.A(new_n11263), .B(new_n11558), .C(new_n11538), .Y(new_n12217));
  NOR2xp33_ASAP7_75t_L      g11961(.A(new_n11908), .B(new_n11907), .Y(new_n12218));
  OAI21xp33_ASAP7_75t_L     g11962(.A1(new_n12218), .A2(new_n12217), .B(new_n11956), .Y(new_n12219));
  NOR3xp33_ASAP7_75t_L      g11963(.A(new_n12207), .B(new_n12208), .C(new_n12209), .Y(new_n12220));
  AOI21xp33_ASAP7_75t_L     g11964(.A1(new_n12202), .A2(new_n12198), .B(new_n12205), .Y(new_n12221));
  NOR2xp33_ASAP7_75t_L      g11965(.A(new_n12221), .B(new_n12220), .Y(new_n12222));
  NAND2xp33_ASAP7_75t_L     g11966(.A(new_n12222), .B(new_n12219), .Y(new_n12223));
  OAI221xp5_ASAP7_75t_L     g11967(.A1(new_n12217), .A2(new_n12218), .B1(new_n12220), .B2(new_n12221), .C(new_n11956), .Y(new_n12224));
  NAND3xp33_ASAP7_75t_L     g11968(.A(new_n12223), .B(new_n12216), .C(new_n12224), .Y(new_n12225));
  OAI211xp5_ASAP7_75t_L     g11969(.A1(new_n11958), .A2(new_n11915), .B(new_n12215), .C(new_n12225), .Y(new_n12226));
  AOI221xp5_ASAP7_75t_L     g11970(.A1(new_n12225), .A2(new_n12215), .B1(new_n11928), .B2(new_n11927), .C(new_n11958), .Y(new_n12227));
  INVx1_ASAP7_75t_L         g11971(.A(new_n12227), .Y(new_n12228));
  AOI21xp33_ASAP7_75t_L     g11972(.A1(new_n12228), .A2(new_n12226), .B(new_n11963), .Y(new_n12229));
  O2A1O1Ixp33_ASAP7_75t_L   g11973(.A1(new_n11543), .A2(new_n11545), .B(new_n11539), .C(new_n11255), .Y(new_n12230));
  O2A1O1Ixp33_ASAP7_75t_L   g11974(.A1(new_n11545), .A2(new_n12230), .B(new_n11906), .C(new_n11909), .Y(new_n12231));
  MAJIxp5_ASAP7_75t_L       g11975(.A(new_n11927), .B(new_n11664), .C(new_n12231), .Y(new_n12232));
  NAND2xp33_ASAP7_75t_L     g11976(.A(new_n12215), .B(new_n12225), .Y(new_n12233));
  NOR2xp33_ASAP7_75t_L      g11977(.A(new_n12232), .B(new_n12233), .Y(new_n12234));
  NOR3xp33_ASAP7_75t_L      g11978(.A(new_n12234), .B(new_n12227), .C(new_n11962), .Y(new_n12235));
  NOR2xp33_ASAP7_75t_L      g11979(.A(new_n12235), .B(new_n12229), .Y(new_n12236));
  A2O1A1Ixp33_ASAP7_75t_L   g11980(.A1(new_n11959), .A2(new_n11655), .B(new_n11935), .C(new_n12236), .Y(new_n12237));
  INVx1_ASAP7_75t_L         g11981(.A(new_n11926), .Y(new_n12238));
  O2A1O1Ixp33_ASAP7_75t_L   g11982(.A1(new_n11929), .A2(new_n11655), .B(new_n11922), .C(new_n12238), .Y(new_n12239));
  OAI21xp33_ASAP7_75t_L     g11983(.A1(new_n12229), .A2(new_n12235), .B(new_n12239), .Y(new_n12240));
  OAI22xp33_ASAP7_75t_L     g11984(.A1(new_n513), .A2(new_n9709), .B1(new_n9683), .B2(new_n506), .Y(new_n12241));
  AOI221xp5_ASAP7_75t_L     g11985(.A1(new_n475), .A2(\b[55] ), .B1(new_n483), .B2(new_n10320), .C(new_n12241), .Y(new_n12242));
  XNOR2x2_ASAP7_75t_L       g11986(.A(new_n466), .B(new_n12242), .Y(new_n12243));
  NAND3xp33_ASAP7_75t_L     g11987(.A(new_n12237), .B(new_n12240), .C(new_n12243), .Y(new_n12244));
  AO21x2_ASAP7_75t_L        g11988(.A1(new_n12240), .A2(new_n12237), .B(new_n12243), .Y(new_n12245));
  INVx1_ASAP7_75t_L         g11989(.A(new_n11934), .Y(new_n12246));
  AOI21xp33_ASAP7_75t_L     g11990(.A1(new_n11644), .A2(new_n11937), .B(new_n12246), .Y(new_n12247));
  NAND3xp33_ASAP7_75t_L     g11991(.A(new_n12245), .B(new_n12247), .C(new_n12244), .Y(new_n12248));
  AO21x2_ASAP7_75t_L        g11992(.A1(new_n12244), .A2(new_n12245), .B(new_n12247), .Y(new_n12249));
  OAI22xp33_ASAP7_75t_L     g11993(.A1(new_n350), .A2(new_n10978), .B1(new_n10332), .B2(new_n375), .Y(new_n12250));
  AOI221xp5_ASAP7_75t_L     g11994(.A1(new_n361), .A2(\b[58] ), .B1(new_n359), .B2(new_n11314), .C(new_n12250), .Y(new_n12251));
  XNOR2x2_ASAP7_75t_L       g11995(.A(new_n346), .B(new_n12251), .Y(new_n12252));
  INVx1_ASAP7_75t_L         g11996(.A(new_n12252), .Y(new_n12253));
  AOI21xp33_ASAP7_75t_L     g11997(.A1(new_n12249), .A2(new_n12248), .B(new_n12253), .Y(new_n12254));
  AND3x1_ASAP7_75t_L        g11998(.A(new_n12245), .B(new_n12247), .C(new_n12244), .Y(new_n12255));
  AOI21xp33_ASAP7_75t_L     g11999(.A1(new_n12245), .A2(new_n12244), .B(new_n12247), .Y(new_n12256));
  NOR3xp33_ASAP7_75t_L      g12000(.A(new_n12255), .B(new_n12256), .C(new_n12252), .Y(new_n12257));
  INVx1_ASAP7_75t_L         g12001(.A(\b[61] ), .Y(new_n12258));
  NAND2xp33_ASAP7_75t_L     g12002(.A(\b[59] ), .B(new_n286), .Y(new_n12259));
  OAI221xp5_ASAP7_75t_L     g12003(.A1(new_n285), .A2(new_n11626), .B1(new_n12258), .B2(new_n269), .C(new_n12259), .Y(new_n12260));
  NOR2xp33_ASAP7_75t_L      g12004(.A(\b[60] ), .B(\b[61] ), .Y(new_n12261));
  NOR2xp33_ASAP7_75t_L      g12005(.A(new_n11626), .B(new_n12258), .Y(new_n12262));
  NOR2xp33_ASAP7_75t_L      g12006(.A(new_n12261), .B(new_n12262), .Y(new_n12263));
  A2O1A1Ixp33_ASAP7_75t_L   g12007(.A1(\b[60] ), .A2(\b[59] ), .B(new_n11630), .C(new_n12263), .Y(new_n12264));
  INVx1_ASAP7_75t_L         g12008(.A(new_n12264), .Y(new_n12265));
  INVx1_ASAP7_75t_L         g12009(.A(new_n11627), .Y(new_n12266));
  A2O1A1Ixp33_ASAP7_75t_L   g12010(.A1(new_n11594), .A2(new_n11624), .B(new_n11625), .C(new_n12266), .Y(new_n12267));
  NOR2xp33_ASAP7_75t_L      g12011(.A(new_n12263), .B(new_n12267), .Y(new_n12268));
  NOR2xp33_ASAP7_75t_L      g12012(.A(new_n12265), .B(new_n12268), .Y(new_n12269));
  AOI21xp33_ASAP7_75t_L     g12013(.A1(new_n12269), .A2(new_n273), .B(new_n12260), .Y(new_n12270));
  NAND2xp33_ASAP7_75t_L     g12014(.A(\a[2] ), .B(new_n12270), .Y(new_n12271));
  A2O1A1Ixp33_ASAP7_75t_L   g12015(.A1(new_n12269), .A2(new_n273), .B(new_n12260), .C(new_n257), .Y(new_n12272));
  NAND2xp33_ASAP7_75t_L     g12016(.A(new_n12272), .B(new_n12271), .Y(new_n12273));
  NOR3xp33_ASAP7_75t_L      g12017(.A(new_n12257), .B(new_n12254), .C(new_n12273), .Y(new_n12274));
  OAI21xp33_ASAP7_75t_L     g12018(.A1(new_n12256), .A2(new_n12255), .B(new_n12252), .Y(new_n12275));
  NAND3xp33_ASAP7_75t_L     g12019(.A(new_n12249), .B(new_n12248), .C(new_n12253), .Y(new_n12276));
  AOI22xp33_ASAP7_75t_L     g12020(.A1(new_n12271), .A2(new_n12272), .B1(new_n12276), .B2(new_n12275), .Y(new_n12277));
  OAI21xp33_ASAP7_75t_L     g12021(.A1(new_n11639), .A2(new_n11944), .B(new_n11946), .Y(new_n12278));
  NOR3xp33_ASAP7_75t_L      g12022(.A(new_n12274), .B(new_n12277), .C(new_n12278), .Y(new_n12279));
  OAI21xp33_ASAP7_75t_L     g12023(.A1(new_n12277), .A2(new_n12274), .B(new_n12278), .Y(new_n12280));
  INVx1_ASAP7_75t_L         g12024(.A(new_n12280), .Y(new_n12281));
  NOR2xp33_ASAP7_75t_L      g12025(.A(new_n12279), .B(new_n12281), .Y(new_n12282));
  A2O1A1Ixp33_ASAP7_75t_L   g12026(.A1(new_n11954), .A2(new_n11952), .B(new_n11949), .C(new_n12282), .Y(new_n12283));
  INVx1_ASAP7_75t_L         g12027(.A(new_n12283), .Y(new_n12284));
  OAI21xp33_ASAP7_75t_L     g12028(.A1(new_n11604), .A2(new_n11603), .B(new_n11605), .Y(new_n12285));
  NAND3xp33_ASAP7_75t_L     g12029(.A(new_n11587), .B(new_n11583), .C(new_n11601), .Y(new_n12286));
  NAND3xp33_ASAP7_75t_L     g12030(.A(new_n12285), .B(new_n12286), .C(new_n11610), .Y(new_n12287));
  NAND2xp33_ASAP7_75t_L     g12031(.A(new_n12287), .B(new_n11612), .Y(new_n12288));
  A2O1A1O1Ixp25_ASAP7_75t_L g12032(.A1(new_n12288), .A2(new_n11609), .B(new_n11608), .C(new_n11950), .D(new_n11949), .Y(new_n12289));
  INVx1_ASAP7_75t_L         g12033(.A(new_n12289), .Y(new_n12290));
  NOR2xp33_ASAP7_75t_L      g12034(.A(new_n12290), .B(new_n12282), .Y(new_n12291));
  NOR2xp33_ASAP7_75t_L      g12035(.A(new_n12291), .B(new_n12284), .Y(\f[61] ));
  A2O1A1Ixp33_ASAP7_75t_L   g12036(.A1(new_n12269), .A2(new_n273), .B(new_n12260), .C(\a[2] ), .Y(new_n12293));
  INVx1_ASAP7_75t_L         g12037(.A(new_n12272), .Y(new_n12294));
  A2O1A1O1Ixp25_ASAP7_75t_L g12038(.A1(new_n12293), .A2(\a[2] ), .B(new_n12294), .C(new_n12275), .D(new_n12257), .Y(new_n12295));
  NAND2xp33_ASAP7_75t_L     g12039(.A(new_n11932), .B(new_n11919), .Y(new_n12296));
  OAI21xp33_ASAP7_75t_L     g12040(.A1(new_n12227), .A2(new_n12234), .B(new_n11962), .Y(new_n12297));
  A2O1A1O1Ixp25_ASAP7_75t_L g12041(.A1(new_n11922), .A2(new_n12296), .B(new_n12238), .C(new_n12297), .D(new_n12235), .Y(new_n12298));
  INVx1_ASAP7_75t_L         g12042(.A(new_n12232), .Y(new_n12299));
  NOR3xp33_ASAP7_75t_L      g12043(.A(new_n12212), .B(new_n12214), .C(new_n11966), .Y(new_n12300));
  A2O1A1O1Ixp25_ASAP7_75t_L g12044(.A1(new_n11906), .A2(new_n11665), .B(new_n12213), .C(new_n12206), .D(new_n12221), .Y(new_n12301));
  O2A1O1Ixp33_ASAP7_75t_L   g12045(.A1(new_n11525), .A2(new_n11890), .B(new_n11899), .C(new_n12197), .Y(new_n12302));
  OAI22xp33_ASAP7_75t_L     g12046(.A1(new_n2572), .A2(new_n4613), .B1(new_n5074), .B2(new_n2410), .Y(new_n12303));
  AOI221xp5_ASAP7_75t_L     g12047(.A1(new_n2423), .A2(\b[38] ), .B1(new_n2417), .B2(new_n6083), .C(new_n12303), .Y(new_n12304));
  XNOR2x2_ASAP7_75t_L       g12048(.A(new_n2413), .B(new_n12304), .Y(new_n12305));
  INVx1_ASAP7_75t_L         g12049(.A(new_n12079), .Y(new_n12306));
  OAI22xp33_ASAP7_75t_L     g12050(.A1(new_n7614), .A2(new_n1043), .B1(new_n1150), .B2(new_n7312), .Y(new_n12307));
  AOI221xp5_ASAP7_75t_L     g12051(.A1(new_n7334), .A2(\b[17] ), .B1(new_n7322), .B2(new_n1633), .C(new_n12307), .Y(new_n12308));
  XNOR2x2_ASAP7_75t_L       g12052(.A(\a[47] ), .B(new_n12308), .Y(new_n12309));
  A2O1A1Ixp33_ASAP7_75t_L   g12053(.A1(new_n12027), .A2(new_n12033), .B(new_n12036), .C(new_n12045), .Y(new_n12310));
  OAI22xp33_ASAP7_75t_L     g12054(.A1(new_n9440), .A2(new_n590), .B1(new_n680), .B2(new_n10400), .Y(new_n12311));
  AOI221xp5_ASAP7_75t_L     g12055(.A1(new_n9102), .A2(\b[11] ), .B1(new_n9437), .B2(new_n976), .C(new_n12311), .Y(new_n12312));
  XNOR2x2_ASAP7_75t_L       g12056(.A(new_n9099), .B(new_n12312), .Y(new_n12313));
  INVx1_ASAP7_75t_L         g12057(.A(new_n12022), .Y(new_n12314));
  AOI21xp33_ASAP7_75t_L     g12058(.A1(new_n11972), .A2(new_n12019), .B(new_n12314), .Y(new_n12315));
  OAI21xp33_ASAP7_75t_L     g12059(.A1(new_n11998), .A2(new_n274), .B(new_n11996), .Y(new_n12316));
  INVx1_ASAP7_75t_L         g12060(.A(new_n12316), .Y(new_n12317));
  NAND2xp33_ASAP7_75t_L     g12061(.A(new_n11990), .B(new_n11720), .Y(new_n12318));
  NAND2xp33_ASAP7_75t_L     g12062(.A(\b[2] ), .B(new_n11995), .Y(new_n12319));
  NAND3xp33_ASAP7_75t_L     g12063(.A(new_n11720), .B(new_n11989), .C(new_n11994), .Y(new_n12320));
  OAI221xp5_ASAP7_75t_L     g12064(.A1(new_n12318), .A2(new_n262), .B1(new_n12320), .B2(new_n284), .C(new_n12319), .Y(new_n12321));
  A2O1A1Ixp33_ASAP7_75t_L   g12065(.A1(new_n294), .A2(new_n11997), .B(new_n12321), .C(\a[62] ), .Y(new_n12322));
  A2O1A1Ixp33_ASAP7_75t_L   g12066(.A1(new_n294), .A2(new_n11997), .B(new_n12321), .C(new_n11987), .Y(new_n12323));
  INVx1_ASAP7_75t_L         g12067(.A(new_n12323), .Y(new_n12324));
  A2O1A1O1Ixp25_ASAP7_75t_L g12068(.A1(new_n12317), .A2(new_n11980), .B(new_n12322), .C(\a[62] ), .D(new_n12324), .Y(new_n12325));
  AOI21xp33_ASAP7_75t_L     g12069(.A1(new_n11997), .A2(new_n294), .B(new_n12321), .Y(new_n12326));
  NAND4xp25_ASAP7_75t_L     g12070(.A(new_n12326), .B(new_n12317), .C(\a[62] ), .D(new_n11980), .Y(new_n12327));
  INVx1_ASAP7_75t_L         g12071(.A(new_n12327), .Y(new_n12328));
  NOR2xp33_ASAP7_75t_L      g12072(.A(new_n301), .B(new_n11354), .Y(new_n12329));
  AOI221xp5_ASAP7_75t_L     g12073(.A1(\b[5] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[4] ), .C(new_n12329), .Y(new_n12330));
  O2A1O1Ixp33_ASAP7_75t_L   g12074(.A1(new_n728), .A2(new_n11053), .B(new_n12330), .C(new_n11048), .Y(new_n12331));
  NOR2xp33_ASAP7_75t_L      g12075(.A(new_n11048), .B(new_n12331), .Y(new_n12332));
  O2A1O1Ixp33_ASAP7_75t_L   g12076(.A1(new_n728), .A2(new_n11053), .B(new_n12330), .C(\a[59] ), .Y(new_n12333));
  NOR2xp33_ASAP7_75t_L      g12077(.A(new_n12333), .B(new_n12332), .Y(new_n12334));
  OAI21xp33_ASAP7_75t_L     g12078(.A1(new_n12328), .A2(new_n12325), .B(new_n12334), .Y(new_n12335));
  NAND2xp33_ASAP7_75t_L     g12079(.A(new_n11721), .B(new_n11360), .Y(new_n12336));
  A2O1A1Ixp33_ASAP7_75t_L   g12080(.A1(new_n11729), .A2(new_n12336), .B(new_n12005), .C(new_n12017), .Y(new_n12337));
  NOR3xp33_ASAP7_75t_L      g12081(.A(new_n12334), .B(new_n12328), .C(new_n12325), .Y(new_n12338));
  INVx1_ASAP7_75t_L         g12082(.A(new_n12335), .Y(new_n12339));
  OA21x2_ASAP7_75t_L        g12083(.A1(new_n12338), .A2(new_n12339), .B(new_n12337), .Y(new_n12340));
  A2O1A1O1Ixp25_ASAP7_75t_L g12084(.A1(new_n12012), .A2(new_n12011), .B(new_n12009), .C(new_n12335), .D(new_n12338), .Y(new_n12341));
  OAI22xp33_ASAP7_75t_L     g12085(.A1(new_n10390), .A2(new_n427), .B1(new_n448), .B2(new_n10388), .Y(new_n12342));
  AOI221xp5_ASAP7_75t_L     g12086(.A1(new_n10086), .A2(\b[8] ), .B1(new_n10386), .B2(new_n1684), .C(new_n12342), .Y(new_n12343));
  XNOR2x2_ASAP7_75t_L       g12087(.A(new_n10083), .B(new_n12343), .Y(new_n12344));
  INVx1_ASAP7_75t_L         g12088(.A(new_n12344), .Y(new_n12345));
  AOI211xp5_ASAP7_75t_L     g12089(.A1(new_n12341), .A2(new_n12335), .B(new_n12345), .C(new_n12340), .Y(new_n12346));
  INVx1_ASAP7_75t_L         g12090(.A(new_n12337), .Y(new_n12347));
  A2O1A1Ixp33_ASAP7_75t_L   g12091(.A1(new_n12011), .A2(new_n12012), .B(new_n12009), .C(new_n12335), .Y(new_n12348));
  NOR2xp33_ASAP7_75t_L      g12092(.A(new_n12338), .B(new_n12348), .Y(new_n12349));
  NAND2xp33_ASAP7_75t_L     g12093(.A(new_n12335), .B(new_n12341), .Y(new_n12350));
  O2A1O1Ixp33_ASAP7_75t_L   g12094(.A1(new_n12347), .A2(new_n12349), .B(new_n12350), .C(new_n12344), .Y(new_n12351));
  NOR3xp33_ASAP7_75t_L      g12095(.A(new_n12315), .B(new_n12346), .C(new_n12351), .Y(new_n12352));
  AO21x2_ASAP7_75t_L        g12096(.A1(new_n12019), .A2(new_n11972), .B(new_n12314), .Y(new_n12353));
  OAI211xp5_ASAP7_75t_L     g12097(.A1(new_n12349), .A2(new_n12347), .B(new_n12350), .C(new_n12344), .Y(new_n12354));
  A2O1A1Ixp33_ASAP7_75t_L   g12098(.A1(new_n12341), .A2(new_n12335), .B(new_n12340), .C(new_n12345), .Y(new_n12355));
  AOI21xp33_ASAP7_75t_L     g12099(.A1(new_n12355), .A2(new_n12354), .B(new_n12353), .Y(new_n12356));
  OAI21xp33_ASAP7_75t_L     g12100(.A1(new_n12352), .A2(new_n12356), .B(new_n12313), .Y(new_n12357));
  INVx1_ASAP7_75t_L         g12101(.A(new_n12313), .Y(new_n12358));
  NAND3xp33_ASAP7_75t_L     g12102(.A(new_n12353), .B(new_n12354), .C(new_n12355), .Y(new_n12359));
  OAI21xp33_ASAP7_75t_L     g12103(.A1(new_n12351), .A2(new_n12346), .B(new_n12315), .Y(new_n12360));
  NAND3xp33_ASAP7_75t_L     g12104(.A(new_n12359), .B(new_n12358), .C(new_n12360), .Y(new_n12361));
  NAND3xp33_ASAP7_75t_L     g12105(.A(new_n12357), .B(new_n12361), .C(new_n12310), .Y(new_n12362));
  AND3x1_ASAP7_75t_L        g12106(.A(new_n12024), .B(new_n12044), .C(new_n12023), .Y(new_n12363));
  O2A1O1Ixp33_ASAP7_75t_L   g12107(.A1(new_n12044), .A2(new_n12028), .B(new_n12031), .C(new_n12363), .Y(new_n12364));
  AOI21xp33_ASAP7_75t_L     g12108(.A1(new_n12359), .A2(new_n12360), .B(new_n12358), .Y(new_n12365));
  NOR3xp33_ASAP7_75t_L      g12109(.A(new_n12356), .B(new_n12352), .C(new_n12313), .Y(new_n12366));
  OAI21xp33_ASAP7_75t_L     g12110(.A1(new_n12366), .A2(new_n12365), .B(new_n12364), .Y(new_n12367));
  OAI22xp33_ASAP7_75t_L     g12111(.A1(new_n8483), .A2(new_n833), .B1(new_n936), .B2(new_n10065), .Y(new_n12368));
  AOI221xp5_ASAP7_75t_L     g12112(.A1(new_n8175), .A2(\b[14] ), .B1(new_n8490), .B2(new_n971), .C(new_n12368), .Y(new_n12369));
  XNOR2x2_ASAP7_75t_L       g12113(.A(new_n8172), .B(new_n12369), .Y(new_n12370));
  NAND3xp33_ASAP7_75t_L     g12114(.A(new_n12367), .B(new_n12362), .C(new_n12370), .Y(new_n12371));
  NOR3xp33_ASAP7_75t_L      g12115(.A(new_n12364), .B(new_n12365), .C(new_n12366), .Y(new_n12372));
  AOI21xp33_ASAP7_75t_L     g12116(.A1(new_n12357), .A2(new_n12361), .B(new_n12310), .Y(new_n12373));
  XNOR2x2_ASAP7_75t_L       g12117(.A(\a[50] ), .B(new_n12369), .Y(new_n12374));
  OAI21xp33_ASAP7_75t_L     g12118(.A1(new_n12373), .A2(new_n12372), .B(new_n12374), .Y(new_n12375));
  AOI21xp33_ASAP7_75t_L     g12119(.A1(new_n12375), .A2(new_n12371), .B(new_n12051), .Y(new_n12376));
  NOR3xp33_ASAP7_75t_L      g12120(.A(new_n12372), .B(new_n12373), .C(new_n12374), .Y(new_n12377));
  AOI21xp33_ASAP7_75t_L     g12121(.A1(new_n12367), .A2(new_n12362), .B(new_n12370), .Y(new_n12378));
  NOR4xp25_ASAP7_75t_L      g12122(.A(new_n12063), .B(new_n12377), .C(new_n12378), .D(new_n12050), .Y(new_n12379));
  OAI21xp33_ASAP7_75t_L     g12123(.A1(new_n12376), .A2(new_n12379), .B(new_n12309), .Y(new_n12380));
  XNOR2x2_ASAP7_75t_L       g12124(.A(new_n7316), .B(new_n12308), .Y(new_n12381));
  OAI22xp33_ASAP7_75t_L     g12125(.A1(new_n12063), .A2(new_n12050), .B1(new_n12378), .B2(new_n12377), .Y(new_n12382));
  NAND3xp33_ASAP7_75t_L     g12126(.A(new_n12051), .B(new_n12371), .C(new_n12375), .Y(new_n12383));
  NAND3xp33_ASAP7_75t_L     g12127(.A(new_n12382), .B(new_n12381), .C(new_n12383), .Y(new_n12384));
  NAND2xp33_ASAP7_75t_L     g12128(.A(new_n12384), .B(new_n12380), .Y(new_n12385));
  O2A1O1Ixp33_ASAP7_75t_L   g12129(.A1(new_n12058), .A2(new_n12060), .B(new_n12055), .C(new_n12385), .Y(new_n12386));
  AOI221xp5_ASAP7_75t_L     g12130(.A1(new_n12384), .A2(new_n12380), .B1(new_n12059), .B2(new_n12073), .C(new_n12071), .Y(new_n12387));
  NOR2xp33_ASAP7_75t_L      g12131(.A(new_n1458), .B(new_n6741), .Y(new_n12388));
  AOI221xp5_ASAP7_75t_L     g12132(.A1(\b[20] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[19] ), .C(new_n12388), .Y(new_n12389));
  O2A1O1Ixp33_ASAP7_75t_L   g12133(.A1(new_n6443), .A2(new_n1754), .B(new_n12389), .C(new_n6439), .Y(new_n12390));
  OAI21xp33_ASAP7_75t_L     g12134(.A1(new_n6443), .A2(new_n1754), .B(new_n12389), .Y(new_n12391));
  NAND2xp33_ASAP7_75t_L     g12135(.A(new_n6439), .B(new_n12391), .Y(new_n12392));
  OAI21xp33_ASAP7_75t_L     g12136(.A1(new_n6439), .A2(new_n12390), .B(new_n12392), .Y(new_n12393));
  INVx1_ASAP7_75t_L         g12137(.A(new_n12393), .Y(new_n12394));
  OAI21xp33_ASAP7_75t_L     g12138(.A1(new_n12387), .A2(new_n12386), .B(new_n12394), .Y(new_n12395));
  NAND3xp33_ASAP7_75t_L     g12139(.A(new_n12382), .B(new_n12309), .C(new_n12383), .Y(new_n12396));
  NOR3xp33_ASAP7_75t_L      g12140(.A(new_n12379), .B(new_n12309), .C(new_n12376), .Y(new_n12397));
  AOI21xp33_ASAP7_75t_L     g12141(.A1(new_n12396), .A2(new_n12309), .B(new_n12397), .Y(new_n12398));
  A2O1A1Ixp33_ASAP7_75t_L   g12142(.A1(new_n12073), .A2(new_n12059), .B(new_n12071), .C(new_n12398), .Y(new_n12399));
  A2O1A1O1Ixp25_ASAP7_75t_L g12143(.A1(new_n12048), .A2(new_n12063), .B(new_n12042), .C(new_n12064), .D(new_n12054), .Y(new_n12400));
  O2A1O1Ixp33_ASAP7_75t_L   g12144(.A1(new_n12400), .A2(new_n12054), .B(new_n12059), .C(new_n12071), .Y(new_n12401));
  A2O1A1Ixp33_ASAP7_75t_L   g12145(.A1(new_n12309), .A2(new_n12396), .B(new_n12397), .C(new_n12401), .Y(new_n12402));
  NAND3xp33_ASAP7_75t_L     g12146(.A(new_n12399), .B(new_n12402), .C(new_n12393), .Y(new_n12403));
  NAND2xp33_ASAP7_75t_L     g12147(.A(new_n12395), .B(new_n12403), .Y(new_n12404));
  O2A1O1Ixp33_ASAP7_75t_L   g12148(.A1(new_n12306), .A2(new_n12081), .B(new_n12070), .C(new_n12404), .Y(new_n12405));
  AOI21xp33_ASAP7_75t_L     g12149(.A1(new_n12403), .A2(new_n12395), .B(new_n12106), .Y(new_n12406));
  NAND2xp33_ASAP7_75t_L     g12150(.A(\b[22] ), .B(new_n5623), .Y(new_n12407));
  OAI221xp5_ASAP7_75t_L     g12151(.A1(new_n5641), .A2(new_n2188), .B1(new_n1895), .B2(new_n5925), .C(new_n12407), .Y(new_n12408));
  A2O1A1Ixp33_ASAP7_75t_L   g12152(.A1(new_n2679), .A2(new_n5637), .B(new_n12408), .C(\a[41] ), .Y(new_n12409));
  AOI211xp5_ASAP7_75t_L     g12153(.A1(new_n2679), .A2(new_n5637), .B(new_n12408), .C(new_n5626), .Y(new_n12410));
  A2O1A1O1Ixp25_ASAP7_75t_L g12154(.A1(new_n5637), .A2(new_n2679), .B(new_n12408), .C(new_n12409), .D(new_n12410), .Y(new_n12411));
  INVx1_ASAP7_75t_L         g12155(.A(new_n12411), .Y(new_n12412));
  OAI21xp33_ASAP7_75t_L     g12156(.A1(new_n12406), .A2(new_n12405), .B(new_n12412), .Y(new_n12413));
  NAND3xp33_ASAP7_75t_L     g12157(.A(new_n12106), .B(new_n12395), .C(new_n12403), .Y(new_n12414));
  NAND2xp33_ASAP7_75t_L     g12158(.A(new_n12404), .B(new_n12104), .Y(new_n12415));
  NAND3xp33_ASAP7_75t_L     g12159(.A(new_n12414), .B(new_n12415), .C(new_n12411), .Y(new_n12416));
  AOI221xp5_ASAP7_75t_L     g12160(.A1(new_n12095), .A2(new_n12097), .B1(new_n12416), .B2(new_n12413), .C(new_n12107), .Y(new_n12417));
  NAND2xp33_ASAP7_75t_L     g12161(.A(new_n12416), .B(new_n12413), .Y(new_n12418));
  O2A1O1Ixp33_ASAP7_75t_L   g12162(.A1(new_n12105), .A2(new_n12085), .B(new_n12098), .C(new_n12418), .Y(new_n12419));
  OAI22xp33_ASAP7_75t_L     g12163(.A1(new_n5144), .A2(new_n2205), .B1(new_n2377), .B2(new_n4903), .Y(new_n12420));
  AOI221xp5_ASAP7_75t_L     g12164(.A1(new_n4917), .A2(\b[26] ), .B1(new_n4912), .B2(new_n2709), .C(new_n12420), .Y(new_n12421));
  XNOR2x2_ASAP7_75t_L       g12165(.A(\a[38] ), .B(new_n12421), .Y(new_n12422));
  NOR3xp33_ASAP7_75t_L      g12166(.A(new_n12419), .B(new_n12422), .C(new_n12417), .Y(new_n12423));
  INVx1_ASAP7_75t_L         g12167(.A(new_n12417), .Y(new_n12424));
  AOI21xp33_ASAP7_75t_L     g12168(.A1(new_n12414), .A2(new_n12415), .B(new_n12411), .Y(new_n12425));
  NOR3xp33_ASAP7_75t_L      g12169(.A(new_n12405), .B(new_n12406), .C(new_n12412), .Y(new_n12426));
  NOR2xp33_ASAP7_75t_L      g12170(.A(new_n12425), .B(new_n12426), .Y(new_n12427));
  A2O1A1Ixp33_ASAP7_75t_L   g12171(.A1(new_n12095), .A2(new_n12097), .B(new_n12107), .C(new_n12427), .Y(new_n12428));
  XNOR2x2_ASAP7_75t_L       g12172(.A(new_n4906), .B(new_n12421), .Y(new_n12429));
  AOI21xp33_ASAP7_75t_L     g12173(.A1(new_n12424), .A2(new_n12428), .B(new_n12429), .Y(new_n12430));
  NOR2xp33_ASAP7_75t_L      g12174(.A(new_n12423), .B(new_n12430), .Y(new_n12431));
  NOR3xp33_ASAP7_75t_L      g12175(.A(new_n12108), .B(new_n12103), .C(new_n12101), .Y(new_n12432));
  O2A1O1Ixp33_ASAP7_75t_L   g12176(.A1(new_n12114), .A2(new_n12109), .B(new_n12112), .C(new_n12432), .Y(new_n12433));
  NAND2xp33_ASAP7_75t_L     g12177(.A(new_n12433), .B(new_n12431), .Y(new_n12434));
  NOR3xp33_ASAP7_75t_L      g12178(.A(new_n12419), .B(new_n12429), .C(new_n12417), .Y(new_n12435));
  INVx1_ASAP7_75t_L         g12179(.A(new_n12435), .Y(new_n12436));
  INVx1_ASAP7_75t_L         g12180(.A(new_n12432), .Y(new_n12437));
  A2O1A1Ixp33_ASAP7_75t_L   g12181(.A1(new_n12101), .A2(new_n12102), .B(new_n12117), .C(new_n12437), .Y(new_n12438));
  A2O1A1Ixp33_ASAP7_75t_L   g12182(.A1(new_n12436), .A2(new_n12422), .B(new_n12423), .C(new_n12438), .Y(new_n12439));
  OAI22xp33_ASAP7_75t_L     g12183(.A1(new_n4397), .A2(new_n2879), .B1(new_n3079), .B2(new_n4142), .Y(new_n12440));
  AOI221xp5_ASAP7_75t_L     g12184(.A1(new_n4156), .A2(\b[29] ), .B1(new_n4151), .B2(new_n3873), .C(new_n12440), .Y(new_n12441));
  XNOR2x2_ASAP7_75t_L       g12185(.A(new_n4145), .B(new_n12441), .Y(new_n12442));
  NAND3xp33_ASAP7_75t_L     g12186(.A(new_n12439), .B(new_n12434), .C(new_n12442), .Y(new_n12443));
  AO21x2_ASAP7_75t_L        g12187(.A1(new_n12434), .A2(new_n12439), .B(new_n12442), .Y(new_n12444));
  NAND2xp33_ASAP7_75t_L     g12188(.A(new_n12443), .B(new_n12444), .Y(new_n12445));
  A2O1A1Ixp33_ASAP7_75t_L   g12189(.A1(new_n11835), .A2(new_n11824), .B(new_n12131), .C(new_n12128), .Y(new_n12446));
  NOR2xp33_ASAP7_75t_L      g12190(.A(new_n12446), .B(new_n12445), .Y(new_n12447));
  INVx1_ASAP7_75t_L         g12191(.A(new_n12442), .Y(new_n12448));
  NAND3xp33_ASAP7_75t_L     g12192(.A(new_n12439), .B(new_n12434), .C(new_n12448), .Y(new_n12449));
  INVx1_ASAP7_75t_L         g12193(.A(new_n12449), .Y(new_n12450));
  INVx1_ASAP7_75t_L         g12194(.A(new_n12128), .Y(new_n12451));
  O2A1O1Ixp33_ASAP7_75t_L   g12195(.A1(new_n12130), .A2(new_n12119), .B(new_n12136), .C(new_n12451), .Y(new_n12452));
  O2A1O1Ixp33_ASAP7_75t_L   g12196(.A1(new_n12442), .A2(new_n12450), .B(new_n12443), .C(new_n12452), .Y(new_n12453));
  OAI22xp33_ASAP7_75t_L     g12197(.A1(new_n3703), .A2(new_n3456), .B1(new_n3674), .B2(new_n3509), .Y(new_n12454));
  AOI221xp5_ASAP7_75t_L     g12198(.A1(new_n3503), .A2(\b[32] ), .B1(new_n3505), .B2(new_n3900), .C(new_n12454), .Y(new_n12455));
  XNOR2x2_ASAP7_75t_L       g12199(.A(new_n3493), .B(new_n12455), .Y(new_n12456));
  OAI21xp33_ASAP7_75t_L     g12200(.A1(new_n12453), .A2(new_n12447), .B(new_n12456), .Y(new_n12457));
  NOR2xp33_ASAP7_75t_L      g12201(.A(new_n12147), .B(new_n12148), .Y(new_n12458));
  MAJIxp5_ASAP7_75t_L       g12202(.A(new_n12146), .B(new_n12149), .C(new_n12458), .Y(new_n12459));
  AND3x1_ASAP7_75t_L        g12203(.A(new_n12439), .B(new_n12434), .C(new_n12442), .Y(new_n12460));
  AOI21xp33_ASAP7_75t_L     g12204(.A1(new_n12449), .A2(new_n12448), .B(new_n12460), .Y(new_n12461));
  NAND2xp33_ASAP7_75t_L     g12205(.A(new_n12452), .B(new_n12461), .Y(new_n12462));
  A2O1A1Ixp33_ASAP7_75t_L   g12206(.A1(new_n12449), .A2(new_n12448), .B(new_n12460), .C(new_n12446), .Y(new_n12463));
  INVx1_ASAP7_75t_L         g12207(.A(new_n12456), .Y(new_n12464));
  NAND3xp33_ASAP7_75t_L     g12208(.A(new_n12462), .B(new_n12463), .C(new_n12464), .Y(new_n12465));
  AOI21xp33_ASAP7_75t_L     g12209(.A1(new_n12457), .A2(new_n12465), .B(new_n12459), .Y(new_n12466));
  NAND2xp33_ASAP7_75t_L     g12210(.A(new_n12137), .B(new_n12132), .Y(new_n12467));
  MAJIxp5_ASAP7_75t_L       g12211(.A(new_n11970), .B(new_n12140), .C(new_n12467), .Y(new_n12468));
  NOR3xp33_ASAP7_75t_L      g12212(.A(new_n12447), .B(new_n12453), .C(new_n12456), .Y(new_n12469));
  AOI21xp33_ASAP7_75t_L     g12213(.A1(new_n12468), .A2(new_n12457), .B(new_n12469), .Y(new_n12470));
  OAI22xp33_ASAP7_75t_L     g12214(.A1(new_n3133), .A2(new_n4101), .B1(new_n4344), .B2(new_n2925), .Y(new_n12471));
  AOI221xp5_ASAP7_75t_L     g12215(.A1(new_n2938), .A2(\b[35] ), .B1(new_n2932), .B2(new_n7773), .C(new_n12471), .Y(new_n12472));
  AND2x2_ASAP7_75t_L        g12216(.A(\a[29] ), .B(new_n12472), .Y(new_n12473));
  NOR2xp33_ASAP7_75t_L      g12217(.A(\a[29] ), .B(new_n12472), .Y(new_n12474));
  NOR2xp33_ASAP7_75t_L      g12218(.A(new_n12474), .B(new_n12473), .Y(new_n12475));
  A2O1A1Ixp33_ASAP7_75t_L   g12219(.A1(new_n12470), .A2(new_n12457), .B(new_n12466), .C(new_n12475), .Y(new_n12476));
  AOI21xp33_ASAP7_75t_L     g12220(.A1(new_n12462), .A2(new_n12463), .B(new_n12464), .Y(new_n12477));
  OAI21xp33_ASAP7_75t_L     g12221(.A1(new_n12469), .A2(new_n12477), .B(new_n12468), .Y(new_n12478));
  NAND3xp33_ASAP7_75t_L     g12222(.A(new_n12459), .B(new_n12465), .C(new_n12457), .Y(new_n12479));
  INVx1_ASAP7_75t_L         g12223(.A(new_n12475), .Y(new_n12480));
  NAND3xp33_ASAP7_75t_L     g12224(.A(new_n12480), .B(new_n12479), .C(new_n12478), .Y(new_n12481));
  AOI21xp33_ASAP7_75t_L     g12225(.A1(new_n12158), .A2(new_n12157), .B(new_n12154), .Y(new_n12482));
  AOI21xp33_ASAP7_75t_L     g12226(.A1(new_n11969), .A2(new_n12159), .B(new_n12482), .Y(new_n12483));
  AND3x1_ASAP7_75t_L        g12227(.A(new_n12483), .B(new_n12481), .C(new_n12476), .Y(new_n12484));
  AOI21xp33_ASAP7_75t_L     g12228(.A1(new_n12476), .A2(new_n12481), .B(new_n12483), .Y(new_n12485));
  NOR3xp33_ASAP7_75t_L      g12229(.A(new_n12484), .B(new_n12485), .C(new_n12305), .Y(new_n12486));
  NAND3xp33_ASAP7_75t_L     g12230(.A(new_n12483), .B(new_n12476), .C(new_n12481), .Y(new_n12487));
  AO21x2_ASAP7_75t_L        g12231(.A1(new_n12476), .A2(new_n12481), .B(new_n12483), .Y(new_n12488));
  NAND3xp33_ASAP7_75t_L     g12232(.A(new_n12488), .B(new_n12487), .C(new_n12305), .Y(new_n12489));
  OAI21xp33_ASAP7_75t_L     g12233(.A1(new_n12305), .A2(new_n12486), .B(new_n12489), .Y(new_n12490));
  NAND3xp33_ASAP7_75t_L     g12234(.A(new_n12161), .B(new_n12168), .C(new_n12162), .Y(new_n12491));
  A2O1A1Ixp33_ASAP7_75t_L   g12235(.A1(new_n12165), .A2(new_n12166), .B(new_n12170), .C(new_n12491), .Y(new_n12492));
  NOR2xp33_ASAP7_75t_L      g12236(.A(new_n12492), .B(new_n12490), .Y(new_n12493));
  AND2x2_ASAP7_75t_L        g12237(.A(new_n12492), .B(new_n12490), .Y(new_n12494));
  NOR2xp33_ASAP7_75t_L      g12238(.A(new_n5855), .B(new_n1962), .Y(new_n12495));
  AOI221xp5_ASAP7_75t_L     g12239(.A1(new_n1955), .A2(\b[41] ), .B1(new_n2093), .B2(\b[39] ), .C(new_n12495), .Y(new_n12496));
  O2A1O1Ixp33_ASAP7_75t_L   g12240(.A1(new_n1956), .A2(new_n6117), .B(new_n12496), .C(new_n1952), .Y(new_n12497));
  NOR2xp33_ASAP7_75t_L      g12241(.A(new_n1952), .B(new_n12497), .Y(new_n12498));
  O2A1O1Ixp33_ASAP7_75t_L   g12242(.A1(new_n1956), .A2(new_n6117), .B(new_n12496), .C(\a[23] ), .Y(new_n12499));
  NOR2xp33_ASAP7_75t_L      g12243(.A(new_n12499), .B(new_n12498), .Y(new_n12500));
  OAI21xp33_ASAP7_75t_L     g12244(.A1(new_n12493), .A2(new_n12494), .B(new_n12500), .Y(new_n12501));
  INVx1_ASAP7_75t_L         g12245(.A(new_n12186), .Y(new_n12502));
  O2A1O1Ixp33_ASAP7_75t_L   g12246(.A1(new_n12187), .A2(new_n12179), .B(new_n12183), .C(new_n12502), .Y(new_n12503));
  OR3x1_ASAP7_75t_L         g12247(.A(new_n12494), .B(new_n12493), .C(new_n12500), .Y(new_n12504));
  AOI21xp33_ASAP7_75t_L     g12248(.A1(new_n12504), .A2(new_n12501), .B(new_n12503), .Y(new_n12505));
  NOR3xp33_ASAP7_75t_L      g12249(.A(new_n12494), .B(new_n12500), .C(new_n12493), .Y(new_n12506));
  A2O1A1O1Ixp25_ASAP7_75t_L g12250(.A1(new_n12181), .A2(new_n12183), .B(new_n12502), .C(new_n12501), .D(new_n12506), .Y(new_n12507));
  NOR2xp33_ASAP7_75t_L      g12251(.A(new_n6944), .B(new_n1518), .Y(new_n12508));
  AOI221xp5_ASAP7_75t_L     g12252(.A1(\b[42] ), .A2(new_n1659), .B1(\b[43] ), .B2(new_n1507), .C(new_n12508), .Y(new_n12509));
  O2A1O1Ixp33_ASAP7_75t_L   g12253(.A1(new_n1521), .A2(new_n6951), .B(new_n12509), .C(new_n1501), .Y(new_n12510));
  OAI21xp33_ASAP7_75t_L     g12254(.A1(new_n1521), .A2(new_n6951), .B(new_n12509), .Y(new_n12511));
  NAND2xp33_ASAP7_75t_L     g12255(.A(new_n1501), .B(new_n12511), .Y(new_n12512));
  OAI21xp33_ASAP7_75t_L     g12256(.A1(new_n1501), .A2(new_n12510), .B(new_n12512), .Y(new_n12513));
  INVx1_ASAP7_75t_L         g12257(.A(new_n12513), .Y(new_n12514));
  A2O1A1Ixp33_ASAP7_75t_L   g12258(.A1(new_n12507), .A2(new_n12501), .B(new_n12505), .C(new_n12514), .Y(new_n12515));
  AO21x2_ASAP7_75t_L        g12259(.A1(new_n12501), .A2(new_n12504), .B(new_n12503), .Y(new_n12516));
  NAND3xp33_ASAP7_75t_L     g12260(.A(new_n12503), .B(new_n12504), .C(new_n12501), .Y(new_n12517));
  NAND3xp33_ASAP7_75t_L     g12261(.A(new_n12516), .B(new_n12517), .C(new_n12513), .Y(new_n12518));
  OAI211xp5_ASAP7_75t_L     g12262(.A1(new_n12193), .A2(new_n12302), .B(new_n12518), .C(new_n12515), .Y(new_n12519));
  INVx1_ASAP7_75t_L         g12263(.A(new_n11525), .Y(new_n12520));
  A2O1A1O1Ixp25_ASAP7_75t_L g12264(.A1(new_n11898), .A2(new_n12520), .B(new_n11896), .C(new_n12201), .D(new_n12193), .Y(new_n12521));
  A2O1A1Ixp33_ASAP7_75t_L   g12265(.A1(new_n12507), .A2(new_n12501), .B(new_n12505), .C(new_n12513), .Y(new_n12522));
  AOI21xp33_ASAP7_75t_L     g12266(.A1(new_n12516), .A2(new_n12517), .B(new_n12513), .Y(new_n12523));
  A2O1A1Ixp33_ASAP7_75t_L   g12267(.A1(new_n12513), .A2(new_n12522), .B(new_n12523), .C(new_n12521), .Y(new_n12524));
  OAI22xp33_ASAP7_75t_L     g12268(.A1(new_n1285), .A2(new_n7249), .B1(new_n7270), .B2(new_n2118), .Y(new_n12525));
  AOI221xp5_ASAP7_75t_L     g12269(.A1(new_n1209), .A2(\b[47] ), .B1(new_n1216), .B2(new_n8726), .C(new_n12525), .Y(new_n12526));
  XNOR2x2_ASAP7_75t_L       g12270(.A(new_n1206), .B(new_n12526), .Y(new_n12527));
  AOI21xp33_ASAP7_75t_L     g12271(.A1(new_n12524), .A2(new_n12519), .B(new_n12527), .Y(new_n12528));
  AOI211xp5_ASAP7_75t_L     g12272(.A1(new_n12507), .A2(new_n12501), .B(new_n12514), .C(new_n12505), .Y(new_n12529));
  NOR3xp33_ASAP7_75t_L      g12273(.A(new_n12521), .B(new_n12523), .C(new_n12529), .Y(new_n12530));
  AOI211xp5_ASAP7_75t_L     g12274(.A1(new_n12518), .A2(new_n12515), .B(new_n12193), .C(new_n12302), .Y(new_n12531));
  INVx1_ASAP7_75t_L         g12275(.A(new_n12527), .Y(new_n12532));
  NOR3xp33_ASAP7_75t_L      g12276(.A(new_n12531), .B(new_n12530), .C(new_n12532), .Y(new_n12533));
  NOR3xp33_ASAP7_75t_L      g12277(.A(new_n12301), .B(new_n12528), .C(new_n12533), .Y(new_n12534));
  OAI21xp33_ASAP7_75t_L     g12278(.A1(new_n12530), .A2(new_n12531), .B(new_n12532), .Y(new_n12535));
  NAND3xp33_ASAP7_75t_L     g12279(.A(new_n12524), .B(new_n12519), .C(new_n12527), .Y(new_n12536));
  AOI221xp5_ASAP7_75t_L     g12280(.A1(new_n12219), .A2(new_n12222), .B1(new_n12535), .B2(new_n12536), .C(new_n12221), .Y(new_n12537));
  OAI22xp33_ASAP7_75t_L     g12281(.A1(new_n980), .A2(new_n7860), .B1(new_n8427), .B2(new_n864), .Y(new_n12538));
  AOI221xp5_ASAP7_75t_L     g12282(.A1(new_n886), .A2(\b[50] ), .B1(new_n873), .B2(new_n8763), .C(new_n12538), .Y(new_n12539));
  XNOR2x2_ASAP7_75t_L       g12283(.A(new_n867), .B(new_n12539), .Y(new_n12540));
  INVx1_ASAP7_75t_L         g12284(.A(new_n12540), .Y(new_n12541));
  NOR3xp33_ASAP7_75t_L      g12285(.A(new_n12537), .B(new_n12534), .C(new_n12541), .Y(new_n12542));
  OA21x2_ASAP7_75t_L        g12286(.A1(new_n12534), .A2(new_n12537), .B(new_n12541), .Y(new_n12543));
  NOR2xp33_ASAP7_75t_L      g12287(.A(new_n12542), .B(new_n12543), .Y(new_n12544));
  A2O1A1Ixp33_ASAP7_75t_L   g12288(.A1(new_n12215), .A2(new_n12299), .B(new_n12300), .C(new_n12544), .Y(new_n12545));
  A2O1A1O1Ixp25_ASAP7_75t_L g12289(.A1(new_n11927), .A2(new_n11928), .B(new_n11958), .C(new_n12215), .D(new_n12300), .Y(new_n12546));
  NOR3xp33_ASAP7_75t_L      g12290(.A(new_n12537), .B(new_n12534), .C(new_n12540), .Y(new_n12547));
  INVx1_ASAP7_75t_L         g12291(.A(new_n12547), .Y(new_n12548));
  A2O1A1Ixp33_ASAP7_75t_L   g12292(.A1(new_n12548), .A2(new_n12541), .B(new_n12542), .C(new_n12546), .Y(new_n12549));
  OAI22xp33_ASAP7_75t_L     g12293(.A1(new_n1550), .A2(new_n9355), .B1(new_n8779), .B2(new_n712), .Y(new_n12550));
  AOI221xp5_ASAP7_75t_L     g12294(.A1(new_n640), .A2(\b[53] ), .B1(new_n718), .B2(new_n9690), .C(new_n12550), .Y(new_n12551));
  XNOR2x2_ASAP7_75t_L       g12295(.A(new_n637), .B(new_n12551), .Y(new_n12552));
  AOI21xp33_ASAP7_75t_L     g12296(.A1(new_n12545), .A2(new_n12549), .B(new_n12552), .Y(new_n12553));
  NAND2xp33_ASAP7_75t_L     g12297(.A(new_n12536), .B(new_n12535), .Y(new_n12554));
  XNOR2x2_ASAP7_75t_L       g12298(.A(new_n12301), .B(new_n12554), .Y(new_n12555));
  OAI21xp33_ASAP7_75t_L     g12299(.A1(new_n12534), .A2(new_n12537), .B(new_n12541), .Y(new_n12556));
  OAI21xp33_ASAP7_75t_L     g12300(.A1(new_n12547), .A2(new_n12555), .B(new_n12556), .Y(new_n12557));
  NOR2xp33_ASAP7_75t_L      g12301(.A(new_n12546), .B(new_n12557), .Y(new_n12558));
  OAI21xp33_ASAP7_75t_L     g12302(.A1(new_n12232), .A2(new_n12233), .B(new_n12225), .Y(new_n12559));
  NOR2xp33_ASAP7_75t_L      g12303(.A(new_n12544), .B(new_n12559), .Y(new_n12560));
  INVx1_ASAP7_75t_L         g12304(.A(new_n12552), .Y(new_n12561));
  NOR3xp33_ASAP7_75t_L      g12305(.A(new_n12558), .B(new_n12560), .C(new_n12561), .Y(new_n12562));
  NOR3xp33_ASAP7_75t_L      g12306(.A(new_n12298), .B(new_n12562), .C(new_n12553), .Y(new_n12563));
  NAND3xp33_ASAP7_75t_L     g12307(.A(new_n12228), .B(new_n12226), .C(new_n11963), .Y(new_n12564));
  A2O1A1Ixp33_ASAP7_75t_L   g12308(.A1(new_n11930), .A2(new_n11926), .B(new_n12229), .C(new_n12564), .Y(new_n12565));
  OAI21xp33_ASAP7_75t_L     g12309(.A1(new_n12560), .A2(new_n12558), .B(new_n12561), .Y(new_n12566));
  NAND3xp33_ASAP7_75t_L     g12310(.A(new_n12545), .B(new_n12549), .C(new_n12552), .Y(new_n12567));
  AOI21xp33_ASAP7_75t_L     g12311(.A1(new_n12567), .A2(new_n12566), .B(new_n12565), .Y(new_n12568));
  OAI22xp33_ASAP7_75t_L     g12312(.A1(new_n513), .A2(new_n10309), .B1(new_n9709), .B2(new_n506), .Y(new_n12569));
  AOI221xp5_ASAP7_75t_L     g12313(.A1(new_n475), .A2(\b[56] ), .B1(new_n483), .B2(new_n11579), .C(new_n12569), .Y(new_n12570));
  XNOR2x2_ASAP7_75t_L       g12314(.A(new_n466), .B(new_n12570), .Y(new_n12571));
  OAI21xp33_ASAP7_75t_L     g12315(.A1(new_n12563), .A2(new_n12568), .B(new_n12571), .Y(new_n12572));
  NAND3xp33_ASAP7_75t_L     g12316(.A(new_n12565), .B(new_n12566), .C(new_n12567), .Y(new_n12573));
  OAI21xp33_ASAP7_75t_L     g12317(.A1(new_n12553), .A2(new_n12562), .B(new_n12298), .Y(new_n12574));
  INVx1_ASAP7_75t_L         g12318(.A(new_n12571), .Y(new_n12575));
  NAND3xp33_ASAP7_75t_L     g12319(.A(new_n12573), .B(new_n12574), .C(new_n12575), .Y(new_n12576));
  INVx1_ASAP7_75t_L         g12320(.A(new_n11597), .Y(new_n12577));
  NOR2xp33_ASAP7_75t_L      g12321(.A(new_n10978), .B(new_n375), .Y(new_n12578));
  AOI221xp5_ASAP7_75t_L     g12322(.A1(\b[59] ), .A2(new_n361), .B1(new_n349), .B2(\b[58] ), .C(new_n12578), .Y(new_n12579));
  INVx1_ASAP7_75t_L         g12323(.A(new_n12579), .Y(new_n12580));
  A2O1A1Ixp33_ASAP7_75t_L   g12324(.A1(new_n12577), .A2(new_n359), .B(new_n12580), .C(\a[5] ), .Y(new_n12581));
  O2A1O1Ixp33_ASAP7_75t_L   g12325(.A1(new_n356), .A2(new_n11597), .B(new_n12579), .C(new_n346), .Y(new_n12582));
  NOR2xp33_ASAP7_75t_L      g12326(.A(new_n346), .B(new_n12582), .Y(new_n12583));
  A2O1A1O1Ixp25_ASAP7_75t_L g12327(.A1(new_n12577), .A2(new_n359), .B(new_n12580), .C(new_n12581), .D(new_n12583), .Y(new_n12584));
  NAND3xp33_ASAP7_75t_L     g12328(.A(new_n12572), .B(new_n12576), .C(new_n12584), .Y(new_n12585));
  AOI21xp33_ASAP7_75t_L     g12329(.A1(new_n12573), .A2(new_n12574), .B(new_n12575), .Y(new_n12586));
  NOR3xp33_ASAP7_75t_L      g12330(.A(new_n12568), .B(new_n12571), .C(new_n12563), .Y(new_n12587));
  NAND2xp33_ASAP7_75t_L     g12331(.A(\a[5] ), .B(new_n12581), .Y(new_n12588));
  O2A1O1Ixp33_ASAP7_75t_L   g12332(.A1(new_n356), .A2(new_n11597), .B(new_n12579), .C(\a[5] ), .Y(new_n12589));
  INVx1_ASAP7_75t_L         g12333(.A(new_n12589), .Y(new_n12590));
  NAND2xp33_ASAP7_75t_L     g12334(.A(new_n12590), .B(new_n12588), .Y(new_n12591));
  OAI21xp33_ASAP7_75t_L     g12335(.A1(new_n12587), .A2(new_n12586), .B(new_n12591), .Y(new_n12592));
  NAND2xp33_ASAP7_75t_L     g12336(.A(new_n12240), .B(new_n12237), .Y(new_n12593));
  MAJx2_ASAP7_75t_L         g12337(.A(new_n12247), .B(new_n12243), .C(new_n12593), .Y(new_n12594));
  NAND3xp33_ASAP7_75t_L     g12338(.A(new_n12594), .B(new_n12592), .C(new_n12585), .Y(new_n12595));
  NOR3xp33_ASAP7_75t_L      g12339(.A(new_n12586), .B(new_n12587), .C(new_n12591), .Y(new_n12596));
  AOI21xp33_ASAP7_75t_L     g12340(.A1(new_n12572), .A2(new_n12576), .B(new_n12584), .Y(new_n12597));
  MAJIxp5_ASAP7_75t_L       g12341(.A(new_n12247), .B(new_n12243), .C(new_n12593), .Y(new_n12598));
  OAI21xp33_ASAP7_75t_L     g12342(.A1(new_n12597), .A2(new_n12596), .B(new_n12598), .Y(new_n12599));
  NOR2xp33_ASAP7_75t_L      g12343(.A(new_n11626), .B(new_n287), .Y(new_n12600));
  AOI221xp5_ASAP7_75t_L     g12344(.A1(\b[61] ), .A2(new_n264), .B1(\b[62] ), .B2(new_n283), .C(new_n12600), .Y(new_n12601));
  NOR2xp33_ASAP7_75t_L      g12345(.A(\b[61] ), .B(\b[62] ), .Y(new_n12602));
  INVx1_ASAP7_75t_L         g12346(.A(\b[62] ), .Y(new_n12603));
  NOR2xp33_ASAP7_75t_L      g12347(.A(new_n12258), .B(new_n12603), .Y(new_n12604));
  NOR2xp33_ASAP7_75t_L      g12348(.A(new_n12602), .B(new_n12604), .Y(new_n12605));
  A2O1A1Ixp33_ASAP7_75t_L   g12349(.A1(new_n12267), .A2(new_n12263), .B(new_n12262), .C(new_n12605), .Y(new_n12606));
  O2A1O1Ixp33_ASAP7_75t_L   g12350(.A1(new_n11627), .A2(new_n11630), .B(new_n12263), .C(new_n12262), .Y(new_n12607));
  INVx1_ASAP7_75t_L         g12351(.A(new_n12605), .Y(new_n12608));
  NAND2xp33_ASAP7_75t_L     g12352(.A(new_n12608), .B(new_n12607), .Y(new_n12609));
  NAND2xp33_ASAP7_75t_L     g12353(.A(new_n12609), .B(new_n12606), .Y(new_n12610));
  O2A1O1Ixp33_ASAP7_75t_L   g12354(.A1(new_n279), .A2(new_n12610), .B(new_n12601), .C(new_n257), .Y(new_n12611));
  NOR2xp33_ASAP7_75t_L      g12355(.A(new_n257), .B(new_n12611), .Y(new_n12612));
  O2A1O1Ixp33_ASAP7_75t_L   g12356(.A1(new_n279), .A2(new_n12610), .B(new_n12601), .C(\a[2] ), .Y(new_n12613));
  NOR2xp33_ASAP7_75t_L      g12357(.A(new_n12613), .B(new_n12612), .Y(new_n12614));
  INVx1_ASAP7_75t_L         g12358(.A(new_n12614), .Y(new_n12615));
  AOI21xp33_ASAP7_75t_L     g12359(.A1(new_n12595), .A2(new_n12599), .B(new_n12615), .Y(new_n12616));
  NOR3xp33_ASAP7_75t_L      g12360(.A(new_n12596), .B(new_n12597), .C(new_n12598), .Y(new_n12617));
  AOI21xp33_ASAP7_75t_L     g12361(.A1(new_n12592), .A2(new_n12585), .B(new_n12594), .Y(new_n12618));
  NOR3xp33_ASAP7_75t_L      g12362(.A(new_n12618), .B(new_n12617), .C(new_n12614), .Y(new_n12619));
  NOR3xp33_ASAP7_75t_L      g12363(.A(new_n12619), .B(new_n12295), .C(new_n12616), .Y(new_n12620));
  A2O1A1Ixp33_ASAP7_75t_L   g12364(.A1(new_n12271), .A2(new_n12272), .B(new_n12254), .C(new_n12276), .Y(new_n12621));
  OAI21xp33_ASAP7_75t_L     g12365(.A1(new_n12617), .A2(new_n12618), .B(new_n12614), .Y(new_n12622));
  NAND3xp33_ASAP7_75t_L     g12366(.A(new_n12595), .B(new_n12615), .C(new_n12599), .Y(new_n12623));
  AOI21xp33_ASAP7_75t_L     g12367(.A1(new_n12622), .A2(new_n12623), .B(new_n12621), .Y(new_n12624));
  NOR2xp33_ASAP7_75t_L      g12368(.A(new_n12624), .B(new_n12620), .Y(new_n12625));
  INVx1_ASAP7_75t_L         g12369(.A(new_n12625), .Y(new_n12626));
  O2A1O1Ixp33_ASAP7_75t_L   g12370(.A1(new_n12279), .A2(new_n12289), .B(new_n12280), .C(new_n12626), .Y(new_n12627));
  OAI21xp33_ASAP7_75t_L     g12371(.A1(new_n12279), .A2(new_n12289), .B(new_n12280), .Y(new_n12628));
  NOR2xp33_ASAP7_75t_L      g12372(.A(new_n12625), .B(new_n12628), .Y(new_n12629));
  NOR2xp33_ASAP7_75t_L      g12373(.A(new_n12629), .B(new_n12627), .Y(\f[62] ));
  OAI21xp33_ASAP7_75t_L     g12374(.A1(new_n12614), .A2(new_n12617), .B(new_n12599), .Y(new_n12631));
  INVx1_ASAP7_75t_L         g12375(.A(new_n12631), .Y(new_n12632));
  NOR2xp33_ASAP7_75t_L      g12376(.A(new_n8779), .B(new_n869), .Y(new_n12633));
  AOI221xp5_ASAP7_75t_L     g12377(.A1(\b[49] ), .A2(new_n985), .B1(\b[50] ), .B2(new_n885), .C(new_n12633), .Y(new_n12634));
  NAND2xp33_ASAP7_75t_L     g12378(.A(new_n873), .B(new_n8790), .Y(new_n12635));
  O2A1O1Ixp33_ASAP7_75t_L   g12379(.A1(new_n872), .A2(new_n8789), .B(new_n12634), .C(new_n867), .Y(new_n12636));
  OA21x2_ASAP7_75t_L        g12380(.A1(new_n872), .A2(new_n8789), .B(new_n12634), .Y(new_n12637));
  NAND2xp33_ASAP7_75t_L     g12381(.A(\a[14] ), .B(new_n12637), .Y(new_n12638));
  A2O1A1Ixp33_ASAP7_75t_L   g12382(.A1(new_n12635), .A2(new_n12634), .B(new_n12636), .C(new_n12638), .Y(new_n12639));
  OAI22xp33_ASAP7_75t_L     g12383(.A1(new_n1285), .A2(new_n7270), .B1(new_n7552), .B2(new_n2118), .Y(new_n12640));
  AOI221xp5_ASAP7_75t_L     g12384(.A1(new_n1209), .A2(\b[48] ), .B1(new_n1216), .B2(new_n11656), .C(new_n12640), .Y(new_n12641));
  XNOR2x2_ASAP7_75t_L       g12385(.A(new_n1206), .B(new_n12641), .Y(new_n12642));
  A2O1A1Ixp33_ASAP7_75t_L   g12386(.A1(new_n12515), .A2(new_n12514), .B(new_n12521), .C(new_n12522), .Y(new_n12643));
  INVx1_ASAP7_75t_L         g12387(.A(new_n12643), .Y(new_n12644));
  OAI22xp33_ASAP7_75t_L     g12388(.A1(new_n1654), .A2(new_n6671), .B1(new_n6944), .B2(new_n1517), .Y(new_n12645));
  AOI221xp5_ASAP7_75t_L     g12389(.A1(new_n1511), .A2(\b[45] ), .B1(new_n1513), .B2(new_n7256), .C(new_n12645), .Y(new_n12646));
  XNOR2x2_ASAP7_75t_L       g12390(.A(new_n1501), .B(new_n12646), .Y(new_n12647));
  INVx1_ASAP7_75t_L         g12391(.A(new_n12647), .Y(new_n12648));
  OAI22xp33_ASAP7_75t_L     g12392(.A1(new_n2089), .A2(new_n5855), .B1(new_n6110), .B2(new_n1962), .Y(new_n12649));
  AOI221xp5_ASAP7_75t_L     g12393(.A1(new_n1955), .A2(\b[42] ), .B1(new_n1964), .B2(new_n6389), .C(new_n12649), .Y(new_n12650));
  XNOR2x2_ASAP7_75t_L       g12394(.A(new_n1952), .B(new_n12650), .Y(new_n12651));
  A2O1A1Ixp33_ASAP7_75t_L   g12395(.A1(new_n12470), .A2(new_n12457), .B(new_n12466), .C(new_n12480), .Y(new_n12652));
  A2O1A1Ixp33_ASAP7_75t_L   g12396(.A1(new_n12476), .A2(new_n12475), .B(new_n12483), .C(new_n12652), .Y(new_n12653));
  INVx1_ASAP7_75t_L         g12397(.A(new_n12401), .Y(new_n12654));
  A2O1A1Ixp33_ASAP7_75t_L   g12398(.A1(new_n12073), .A2(new_n12059), .B(new_n12071), .C(new_n12385), .Y(new_n12655));
  A2O1A1Ixp33_ASAP7_75t_L   g12399(.A1(new_n12655), .A2(new_n12654), .B(new_n12387), .C(new_n12393), .Y(new_n12656));
  INVx1_ASAP7_75t_L         g12400(.A(new_n12656), .Y(new_n12657));
  OAI22xp33_ASAP7_75t_L     g12401(.A1(new_n7304), .A2(new_n1745), .B1(new_n1599), .B2(new_n6741), .Y(new_n12658));
  AOI221xp5_ASAP7_75t_L     g12402(.A1(new_n6442), .A2(\b[21] ), .B1(new_n6450), .B2(new_n2836), .C(new_n12658), .Y(new_n12659));
  XNOR2x2_ASAP7_75t_L       g12403(.A(new_n6439), .B(new_n12659), .Y(new_n12660));
  INVx1_ASAP7_75t_L         g12404(.A(new_n12396), .Y(new_n12661));
  A2O1A1O1Ixp25_ASAP7_75t_L g12405(.A1(new_n12073), .A2(new_n12059), .B(new_n12071), .C(new_n12385), .D(new_n12661), .Y(new_n12662));
  NAND2xp33_ASAP7_75t_L     g12406(.A(new_n12362), .B(new_n12367), .Y(new_n12663));
  NOR2xp33_ASAP7_75t_L      g12407(.A(new_n12370), .B(new_n12663), .Y(new_n12664));
  INVx1_ASAP7_75t_L         g12408(.A(new_n12664), .Y(new_n12665));
  A2O1A1Ixp33_ASAP7_75t_L   g12409(.A1(new_n12046), .A2(new_n12045), .B(new_n12365), .C(new_n12361), .Y(new_n12666));
  A2O1A1Ixp33_ASAP7_75t_L   g12410(.A1(new_n12023), .A2(new_n12022), .B(new_n12346), .C(new_n12355), .Y(new_n12667));
  O2A1O1Ixp33_ASAP7_75t_L   g12411(.A1(new_n11981), .A2(new_n12005), .B(new_n12017), .C(new_n12339), .Y(new_n12668));
  NOR2xp33_ASAP7_75t_L      g12412(.A(\a[63] ), .B(new_n11987), .Y(new_n12669));
  INVx1_ASAP7_75t_L         g12413(.A(\a[63] ), .Y(new_n12670));
  NOR2xp33_ASAP7_75t_L      g12414(.A(\a[62] ), .B(new_n12670), .Y(new_n12671));
  NOR2xp33_ASAP7_75t_L      g12415(.A(new_n12669), .B(new_n12671), .Y(new_n12672));
  NOR2xp33_ASAP7_75t_L      g12416(.A(new_n284), .B(new_n12672), .Y(new_n12673));
  NOR3xp33_ASAP7_75t_L      g12417(.A(new_n12327), .B(new_n12672), .C(new_n284), .Y(new_n12674));
  INVx1_ASAP7_75t_L         g12418(.A(new_n12674), .Y(new_n12675));
  O2A1O1Ixp33_ASAP7_75t_L   g12419(.A1(new_n12669), .A2(new_n12671), .B(\b[0] ), .C(new_n12327), .Y(new_n12676));
  NAND2xp33_ASAP7_75t_L     g12420(.A(\b[3] ), .B(new_n11995), .Y(new_n12677));
  OAI221xp5_ASAP7_75t_L     g12421(.A1(new_n12318), .A2(new_n289), .B1(new_n262), .B2(new_n12320), .C(new_n12677), .Y(new_n12678));
  A2O1A1Ixp33_ASAP7_75t_L   g12422(.A1(new_n312), .A2(new_n11997), .B(new_n12678), .C(\a[62] ), .Y(new_n12679));
  NAND2xp33_ASAP7_75t_L     g12423(.A(\a[62] ), .B(new_n12679), .Y(new_n12680));
  A2O1A1Ixp33_ASAP7_75t_L   g12424(.A1(new_n312), .A2(new_n11997), .B(new_n12678), .C(new_n11987), .Y(new_n12681));
  NAND2xp33_ASAP7_75t_L     g12425(.A(new_n12681), .B(new_n12680), .Y(new_n12682));
  INVx1_ASAP7_75t_L         g12426(.A(new_n12682), .Y(new_n12683));
  A2O1A1Ixp33_ASAP7_75t_L   g12427(.A1(new_n12675), .A2(new_n12673), .B(new_n12676), .C(new_n12683), .Y(new_n12684));
  INVx1_ASAP7_75t_L         g12428(.A(new_n12669), .Y(new_n12685));
  INVx1_ASAP7_75t_L         g12429(.A(new_n12671), .Y(new_n12686));
  A2O1A1Ixp33_ASAP7_75t_L   g12430(.A1(new_n12685), .A2(new_n12686), .B(new_n284), .C(new_n12328), .Y(new_n12687));
  NAND2xp33_ASAP7_75t_L     g12431(.A(new_n12673), .B(new_n12327), .Y(new_n12688));
  NAND3xp33_ASAP7_75t_L     g12432(.A(new_n12687), .B(new_n12688), .C(new_n12682), .Y(new_n12689));
  NOR2xp33_ASAP7_75t_L      g12433(.A(new_n332), .B(new_n11354), .Y(new_n12690));
  AOI221xp5_ASAP7_75t_L     g12434(.A1(\b[6] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[5] ), .C(new_n12690), .Y(new_n12691));
  O2A1O1Ixp33_ASAP7_75t_L   g12435(.A1(new_n11053), .A2(new_n434), .B(new_n12691), .C(new_n11048), .Y(new_n12692));
  OAI21xp33_ASAP7_75t_L     g12436(.A1(new_n11053), .A2(new_n434), .B(new_n12691), .Y(new_n12693));
  NAND2xp33_ASAP7_75t_L     g12437(.A(new_n11048), .B(new_n12693), .Y(new_n12694));
  OAI21xp33_ASAP7_75t_L     g12438(.A1(new_n11048), .A2(new_n12692), .B(new_n12694), .Y(new_n12695));
  INVx1_ASAP7_75t_L         g12439(.A(new_n12695), .Y(new_n12696));
  NAND3xp33_ASAP7_75t_L     g12440(.A(new_n12684), .B(new_n12689), .C(new_n12696), .Y(new_n12697));
  O2A1O1Ixp33_ASAP7_75t_L   g12441(.A1(new_n12327), .A2(new_n12674), .B(new_n12688), .C(new_n12682), .Y(new_n12698));
  AND3x1_ASAP7_75t_L        g12442(.A(new_n12687), .B(new_n12682), .C(new_n12688), .Y(new_n12699));
  OAI21xp33_ASAP7_75t_L     g12443(.A1(new_n12698), .A2(new_n12699), .B(new_n12695), .Y(new_n12700));
  OAI211xp5_ASAP7_75t_L     g12444(.A1(new_n12338), .A2(new_n12668), .B(new_n12700), .C(new_n12697), .Y(new_n12701));
  NOR3xp33_ASAP7_75t_L      g12445(.A(new_n12699), .B(new_n12695), .C(new_n12698), .Y(new_n12702));
  O2A1O1Ixp33_ASAP7_75t_L   g12446(.A1(new_n12327), .A2(new_n12674), .B(new_n12688), .C(new_n12683), .Y(new_n12703));
  A2O1A1O1Ixp25_ASAP7_75t_L g12447(.A1(new_n12688), .A2(new_n12687), .B(new_n12703), .C(new_n12689), .D(new_n12696), .Y(new_n12704));
  OAI21xp33_ASAP7_75t_L     g12448(.A1(new_n12704), .A2(new_n12702), .B(new_n12341), .Y(new_n12705));
  AND2x2_ASAP7_75t_L        g12449(.A(new_n12705), .B(new_n12701), .Y(new_n12706));
  NAND2xp33_ASAP7_75t_L     g12450(.A(\b[9] ), .B(new_n10086), .Y(new_n12707));
  OAI221xp5_ASAP7_75t_L     g12451(.A1(new_n10388), .A2(new_n534), .B1(new_n448), .B2(new_n10390), .C(new_n12707), .Y(new_n12708));
  A2O1A1Ixp33_ASAP7_75t_L   g12452(.A1(new_n602), .A2(new_n10386), .B(new_n12708), .C(\a[56] ), .Y(new_n12709));
  NAND2xp33_ASAP7_75t_L     g12453(.A(\a[56] ), .B(new_n12709), .Y(new_n12710));
  A2O1A1Ixp33_ASAP7_75t_L   g12454(.A1(new_n602), .A2(new_n10386), .B(new_n12708), .C(new_n10083), .Y(new_n12711));
  NAND2xp33_ASAP7_75t_L     g12455(.A(new_n12711), .B(new_n12710), .Y(new_n12712));
  NAND3xp33_ASAP7_75t_L     g12456(.A(new_n12701), .B(new_n12705), .C(new_n12712), .Y(new_n12713));
  NAND2xp33_ASAP7_75t_L     g12457(.A(new_n12713), .B(new_n12706), .Y(new_n12714));
  INVx1_ASAP7_75t_L         g12458(.A(new_n12712), .Y(new_n12715));
  AOI21xp33_ASAP7_75t_L     g12459(.A1(new_n12701), .A2(new_n12705), .B(new_n12715), .Y(new_n12716));
  INVx1_ASAP7_75t_L         g12460(.A(new_n12716), .Y(new_n12717));
  NAND3xp33_ASAP7_75t_L     g12461(.A(new_n12667), .B(new_n12714), .C(new_n12717), .Y(new_n12718));
  A2O1A1O1Ixp25_ASAP7_75t_L g12462(.A1(new_n12019), .A2(new_n11972), .B(new_n12314), .C(new_n12354), .D(new_n12351), .Y(new_n12719));
  NAND2xp33_ASAP7_75t_L     g12463(.A(new_n12705), .B(new_n12701), .Y(new_n12720));
  NOR2xp33_ASAP7_75t_L      g12464(.A(new_n12712), .B(new_n12720), .Y(new_n12721));
  A2O1A1Ixp33_ASAP7_75t_L   g12465(.A1(new_n12712), .A2(new_n12713), .B(new_n12721), .C(new_n12719), .Y(new_n12722));
  NOR2xp33_ASAP7_75t_L      g12466(.A(new_n748), .B(new_n10400), .Y(new_n12723));
  AOI221xp5_ASAP7_75t_L     g12467(.A1(new_n9102), .A2(\b[12] ), .B1(new_n10398), .B2(\b[10] ), .C(new_n12723), .Y(new_n12724));
  O2A1O1Ixp33_ASAP7_75t_L   g12468(.A1(new_n9104), .A2(new_n841), .B(new_n12724), .C(new_n9099), .Y(new_n12725));
  OAI21xp33_ASAP7_75t_L     g12469(.A1(new_n9104), .A2(new_n841), .B(new_n12724), .Y(new_n12726));
  NAND2xp33_ASAP7_75t_L     g12470(.A(new_n9099), .B(new_n12726), .Y(new_n12727));
  OAI21xp33_ASAP7_75t_L     g12471(.A1(new_n9099), .A2(new_n12725), .B(new_n12727), .Y(new_n12728));
  INVx1_ASAP7_75t_L         g12472(.A(new_n12728), .Y(new_n12729));
  NAND3xp33_ASAP7_75t_L     g12473(.A(new_n12722), .B(new_n12718), .C(new_n12729), .Y(new_n12730));
  NOR3xp33_ASAP7_75t_L      g12474(.A(new_n12719), .B(new_n12721), .C(new_n12716), .Y(new_n12731));
  INVx1_ASAP7_75t_L         g12475(.A(new_n12713), .Y(new_n12732));
  O2A1O1Ixp33_ASAP7_75t_L   g12476(.A1(new_n12715), .A2(new_n12732), .B(new_n12714), .C(new_n12667), .Y(new_n12733));
  OAI21xp33_ASAP7_75t_L     g12477(.A1(new_n12733), .A2(new_n12731), .B(new_n12728), .Y(new_n12734));
  NAND3xp33_ASAP7_75t_L     g12478(.A(new_n12666), .B(new_n12730), .C(new_n12734), .Y(new_n12735));
  O2A1O1Ixp33_ASAP7_75t_L   g12479(.A1(new_n12363), .A2(new_n12037), .B(new_n12357), .C(new_n12366), .Y(new_n12736));
  NAND2xp33_ASAP7_75t_L     g12480(.A(new_n12730), .B(new_n12734), .Y(new_n12737));
  NAND2xp33_ASAP7_75t_L     g12481(.A(new_n12736), .B(new_n12737), .Y(new_n12738));
  OAI22xp33_ASAP7_75t_L     g12482(.A1(new_n8483), .A2(new_n936), .B1(new_n960), .B2(new_n10065), .Y(new_n12739));
  AOI221xp5_ASAP7_75t_L     g12483(.A1(new_n8175), .A2(\b[15] ), .B1(new_n8490), .B2(new_n1052), .C(new_n12739), .Y(new_n12740));
  XNOR2x2_ASAP7_75t_L       g12484(.A(new_n8172), .B(new_n12740), .Y(new_n12741));
  NAND3xp33_ASAP7_75t_L     g12485(.A(new_n12738), .B(new_n12735), .C(new_n12741), .Y(new_n12742));
  AO21x2_ASAP7_75t_L        g12486(.A1(new_n12735), .A2(new_n12738), .B(new_n12741), .Y(new_n12743));
  NAND4xp25_ASAP7_75t_L     g12487(.A(new_n12743), .B(new_n12665), .C(new_n12382), .D(new_n12742), .Y(new_n12744));
  INVx1_ASAP7_75t_L         g12488(.A(new_n12741), .Y(new_n12745));
  NAND3xp33_ASAP7_75t_L     g12489(.A(new_n12738), .B(new_n12745), .C(new_n12735), .Y(new_n12746));
  AND3x1_ASAP7_75t_L        g12490(.A(new_n12738), .B(new_n12741), .C(new_n12735), .Y(new_n12747));
  MAJIxp5_ASAP7_75t_L       g12491(.A(new_n12051), .B(new_n12370), .C(new_n12663), .Y(new_n12748));
  A2O1A1Ixp33_ASAP7_75t_L   g12492(.A1(new_n12746), .A2(new_n12745), .B(new_n12747), .C(new_n12748), .Y(new_n12749));
  NOR2xp33_ASAP7_75t_L      g12493(.A(new_n1458), .B(new_n7318), .Y(new_n12750));
  AOI221xp5_ASAP7_75t_L     g12494(.A1(new_n7333), .A2(\b[17] ), .B1(new_n7609), .B2(\b[16] ), .C(new_n12750), .Y(new_n12751));
  O2A1O1Ixp33_ASAP7_75t_L   g12495(.A1(new_n7321), .A2(new_n1464), .B(new_n12751), .C(new_n7316), .Y(new_n12752));
  OAI21xp33_ASAP7_75t_L     g12496(.A1(new_n7321), .A2(new_n1464), .B(new_n12751), .Y(new_n12753));
  NAND2xp33_ASAP7_75t_L     g12497(.A(new_n7316), .B(new_n12753), .Y(new_n12754));
  OAI21xp33_ASAP7_75t_L     g12498(.A1(new_n7316), .A2(new_n12752), .B(new_n12754), .Y(new_n12755));
  AOI21xp33_ASAP7_75t_L     g12499(.A1(new_n12749), .A2(new_n12744), .B(new_n12755), .Y(new_n12756));
  AOI211xp5_ASAP7_75t_L     g12500(.A1(new_n12746), .A2(new_n12745), .B(new_n12748), .C(new_n12747), .Y(new_n12757));
  AOI22xp33_ASAP7_75t_L     g12501(.A1(new_n12665), .A2(new_n12382), .B1(new_n12742), .B2(new_n12743), .Y(new_n12758));
  INVx1_ASAP7_75t_L         g12502(.A(new_n12755), .Y(new_n12759));
  NOR3xp33_ASAP7_75t_L      g12503(.A(new_n12757), .B(new_n12758), .C(new_n12759), .Y(new_n12760));
  NOR3xp33_ASAP7_75t_L      g12504(.A(new_n12662), .B(new_n12756), .C(new_n12760), .Y(new_n12761));
  A2O1A1Ixp33_ASAP7_75t_L   g12505(.A1(new_n12380), .A2(new_n12384), .B(new_n12401), .C(new_n12396), .Y(new_n12762));
  OAI21xp33_ASAP7_75t_L     g12506(.A1(new_n12758), .A2(new_n12757), .B(new_n12759), .Y(new_n12763));
  NAND3xp33_ASAP7_75t_L     g12507(.A(new_n12749), .B(new_n12744), .C(new_n12755), .Y(new_n12764));
  AOI21xp33_ASAP7_75t_L     g12508(.A1(new_n12764), .A2(new_n12763), .B(new_n12762), .Y(new_n12765));
  NOR3xp33_ASAP7_75t_L      g12509(.A(new_n12761), .B(new_n12765), .C(new_n12660), .Y(new_n12766));
  XNOR2x2_ASAP7_75t_L       g12510(.A(\a[44] ), .B(new_n12659), .Y(new_n12767));
  NAND3xp33_ASAP7_75t_L     g12511(.A(new_n12762), .B(new_n12763), .C(new_n12764), .Y(new_n12768));
  OAI21xp33_ASAP7_75t_L     g12512(.A1(new_n12756), .A2(new_n12760), .B(new_n12662), .Y(new_n12769));
  AOI21xp33_ASAP7_75t_L     g12513(.A1(new_n12769), .A2(new_n12768), .B(new_n12767), .Y(new_n12770));
  NOR2xp33_ASAP7_75t_L      g12514(.A(new_n12770), .B(new_n12766), .Y(new_n12771));
  A2O1A1Ixp33_ASAP7_75t_L   g12515(.A1(new_n12404), .A2(new_n12106), .B(new_n12657), .C(new_n12771), .Y(new_n12772));
  O2A1O1Ixp33_ASAP7_75t_L   g12516(.A1(new_n12087), .A2(new_n12080), .B(new_n12404), .C(new_n12657), .Y(new_n12773));
  NAND3xp33_ASAP7_75t_L     g12517(.A(new_n12769), .B(new_n12768), .C(new_n12767), .Y(new_n12774));
  OAI21xp33_ASAP7_75t_L     g12518(.A1(new_n12765), .A2(new_n12761), .B(new_n12660), .Y(new_n12775));
  NAND2xp33_ASAP7_75t_L     g12519(.A(new_n12774), .B(new_n12775), .Y(new_n12776));
  NAND2xp33_ASAP7_75t_L     g12520(.A(new_n12773), .B(new_n12776), .Y(new_n12777));
  OAI22xp33_ASAP7_75t_L     g12521(.A1(new_n5640), .A2(new_n2188), .B1(new_n2045), .B2(new_n5925), .Y(new_n12778));
  AOI221xp5_ASAP7_75t_L     g12522(.A1(new_n5629), .A2(\b[24] ), .B1(new_n5637), .B2(new_n2216), .C(new_n12778), .Y(new_n12779));
  XNOR2x2_ASAP7_75t_L       g12523(.A(new_n5626), .B(new_n12779), .Y(new_n12780));
  NAND3xp33_ASAP7_75t_L     g12524(.A(new_n12772), .B(new_n12777), .C(new_n12780), .Y(new_n12781));
  O2A1O1Ixp33_ASAP7_75t_L   g12525(.A1(new_n12071), .A2(new_n12075), .B(new_n12655), .C(new_n12387), .Y(new_n12782));
  A2O1A1Ixp33_ASAP7_75t_L   g12526(.A1(new_n12077), .A2(new_n12079), .B(new_n12080), .C(new_n12404), .Y(new_n12783));
  O2A1O1Ixp33_ASAP7_75t_L   g12527(.A1(new_n12782), .A2(new_n12394), .B(new_n12783), .C(new_n12776), .Y(new_n12784));
  A2O1A1Ixp33_ASAP7_75t_L   g12528(.A1(new_n12395), .A2(new_n12403), .B(new_n12104), .C(new_n12656), .Y(new_n12785));
  NOR2xp33_ASAP7_75t_L      g12529(.A(new_n12771), .B(new_n12785), .Y(new_n12786));
  INVx1_ASAP7_75t_L         g12530(.A(new_n12780), .Y(new_n12787));
  OAI21xp33_ASAP7_75t_L     g12531(.A1(new_n12786), .A2(new_n12784), .B(new_n12787), .Y(new_n12788));
  A2O1A1O1Ixp25_ASAP7_75t_L g12532(.A1(new_n12097), .A2(new_n12095), .B(new_n12107), .C(new_n12416), .D(new_n12425), .Y(new_n12789));
  NAND3xp33_ASAP7_75t_L     g12533(.A(new_n12789), .B(new_n12788), .C(new_n12781), .Y(new_n12790));
  O2A1O1Ixp33_ASAP7_75t_L   g12534(.A1(new_n11784), .A2(new_n11798), .B(new_n12095), .C(new_n12107), .Y(new_n12791));
  INVx1_ASAP7_75t_L         g12535(.A(new_n12791), .Y(new_n12792));
  NAND2xp33_ASAP7_75t_L     g12536(.A(new_n12781), .B(new_n12788), .Y(new_n12793));
  A2O1A1Ixp33_ASAP7_75t_L   g12537(.A1(new_n12416), .A2(new_n12792), .B(new_n12425), .C(new_n12793), .Y(new_n12794));
  OAI22xp33_ASAP7_75t_L     g12538(.A1(new_n5144), .A2(new_n2377), .B1(new_n2703), .B2(new_n4903), .Y(new_n12795));
  AOI221xp5_ASAP7_75t_L     g12539(.A1(new_n4917), .A2(\b[27] ), .B1(new_n4912), .B2(new_n2887), .C(new_n12795), .Y(new_n12796));
  XNOR2x2_ASAP7_75t_L       g12540(.A(\a[38] ), .B(new_n12796), .Y(new_n12797));
  INVx1_ASAP7_75t_L         g12541(.A(new_n12797), .Y(new_n12798));
  NAND3xp33_ASAP7_75t_L     g12542(.A(new_n12794), .B(new_n12798), .C(new_n12790), .Y(new_n12799));
  INVx1_ASAP7_75t_L         g12543(.A(new_n12790), .Y(new_n12800));
  NAND2xp33_ASAP7_75t_L     g12544(.A(new_n12777), .B(new_n12772), .Y(new_n12801));
  NOR2xp33_ASAP7_75t_L      g12545(.A(new_n12780), .B(new_n12801), .Y(new_n12802));
  O2A1O1Ixp33_ASAP7_75t_L   g12546(.A1(new_n12780), .A2(new_n12802), .B(new_n12781), .C(new_n12789), .Y(new_n12803));
  OAI21xp33_ASAP7_75t_L     g12547(.A1(new_n12800), .A2(new_n12803), .B(new_n12797), .Y(new_n12804));
  NAND2xp33_ASAP7_75t_L     g12548(.A(new_n12799), .B(new_n12804), .Y(new_n12805));
  NAND3xp33_ASAP7_75t_L     g12549(.A(new_n12424), .B(new_n12428), .C(new_n12429), .Y(new_n12806));
  A2O1A1Ixp33_ASAP7_75t_L   g12550(.A1(new_n12429), .A2(new_n12806), .B(new_n12433), .C(new_n12436), .Y(new_n12807));
  NOR2xp33_ASAP7_75t_L      g12551(.A(new_n12807), .B(new_n12805), .Y(new_n12808));
  NAND3xp33_ASAP7_75t_L     g12552(.A(new_n12794), .B(new_n12790), .C(new_n12797), .Y(new_n12809));
  NOR3xp33_ASAP7_75t_L      g12553(.A(new_n12803), .B(new_n12797), .C(new_n12800), .Y(new_n12810));
  AOI21xp33_ASAP7_75t_L     g12554(.A1(new_n12809), .A2(new_n12797), .B(new_n12810), .Y(new_n12811));
  O2A1O1Ixp33_ASAP7_75t_L   g12555(.A1(new_n12423), .A2(new_n12430), .B(new_n12438), .C(new_n12435), .Y(new_n12812));
  NOR2xp33_ASAP7_75t_L      g12556(.A(new_n12812), .B(new_n12811), .Y(new_n12813));
  OAI22xp33_ASAP7_75t_L     g12557(.A1(new_n4397), .A2(new_n3079), .B1(new_n3098), .B2(new_n4142), .Y(new_n12814));
  AOI221xp5_ASAP7_75t_L     g12558(.A1(new_n4156), .A2(\b[30] ), .B1(new_n4151), .B2(new_n4813), .C(new_n12814), .Y(new_n12815));
  XNOR2x2_ASAP7_75t_L       g12559(.A(new_n4145), .B(new_n12815), .Y(new_n12816));
  OAI21xp33_ASAP7_75t_L     g12560(.A1(new_n12808), .A2(new_n12813), .B(new_n12816), .Y(new_n12817));
  NAND2xp33_ASAP7_75t_L     g12561(.A(new_n12812), .B(new_n12811), .Y(new_n12818));
  A2O1A1Ixp33_ASAP7_75t_L   g12562(.A1(new_n12809), .A2(new_n12797), .B(new_n12810), .C(new_n12807), .Y(new_n12819));
  INVx1_ASAP7_75t_L         g12563(.A(new_n12816), .Y(new_n12820));
  NAND3xp33_ASAP7_75t_L     g12564(.A(new_n12818), .B(new_n12819), .C(new_n12820), .Y(new_n12821));
  NAND2xp33_ASAP7_75t_L     g12565(.A(new_n12821), .B(new_n12817), .Y(new_n12822));
  O2A1O1Ixp33_ASAP7_75t_L   g12566(.A1(new_n12461), .A2(new_n12452), .B(new_n12449), .C(new_n12822), .Y(new_n12823));
  AOI21xp33_ASAP7_75t_L     g12567(.A1(new_n12818), .A2(new_n12819), .B(new_n12820), .Y(new_n12824));
  NOR3xp33_ASAP7_75t_L      g12568(.A(new_n12813), .B(new_n12808), .C(new_n12816), .Y(new_n12825));
  NOR2xp33_ASAP7_75t_L      g12569(.A(new_n12824), .B(new_n12825), .Y(new_n12826));
  A2O1A1Ixp33_ASAP7_75t_L   g12570(.A1(new_n12442), .A2(new_n12443), .B(new_n12452), .C(new_n12449), .Y(new_n12827));
  NOR2xp33_ASAP7_75t_L      g12571(.A(new_n12827), .B(new_n12826), .Y(new_n12828));
  NOR2xp33_ASAP7_75t_L      g12572(.A(new_n4101), .B(new_n3510), .Y(new_n12829));
  AOI221xp5_ASAP7_75t_L     g12573(.A1(\b[31] ), .A2(new_n3708), .B1(\b[32] ), .B2(new_n3499), .C(new_n12829), .Y(new_n12830));
  O2A1O1Ixp33_ASAP7_75t_L   g12574(.A1(new_n3513), .A2(new_n4108), .B(new_n12830), .C(new_n3493), .Y(new_n12831));
  OAI21xp33_ASAP7_75t_L     g12575(.A1(new_n3513), .A2(new_n4108), .B(new_n12830), .Y(new_n12832));
  NAND2xp33_ASAP7_75t_L     g12576(.A(new_n3493), .B(new_n12832), .Y(new_n12833));
  OAI21xp33_ASAP7_75t_L     g12577(.A1(new_n3493), .A2(new_n12831), .B(new_n12833), .Y(new_n12834));
  NOR3xp33_ASAP7_75t_L      g12578(.A(new_n12823), .B(new_n12828), .C(new_n12834), .Y(new_n12835));
  A2O1A1Ixp33_ASAP7_75t_L   g12579(.A1(new_n12445), .A2(new_n12446), .B(new_n12450), .C(new_n12826), .Y(new_n12836));
  O2A1O1Ixp33_ASAP7_75t_L   g12580(.A1(new_n12460), .A2(new_n12448), .B(new_n12446), .C(new_n12450), .Y(new_n12837));
  NAND2xp33_ASAP7_75t_L     g12581(.A(new_n12837), .B(new_n12822), .Y(new_n12838));
  INVx1_ASAP7_75t_L         g12582(.A(new_n12834), .Y(new_n12839));
  AOI21xp33_ASAP7_75t_L     g12583(.A1(new_n12836), .A2(new_n12838), .B(new_n12839), .Y(new_n12840));
  NOR3xp33_ASAP7_75t_L      g12584(.A(new_n12840), .B(new_n12835), .C(new_n12470), .Y(new_n12841));
  O2A1O1Ixp33_ASAP7_75t_L   g12585(.A1(new_n12447), .A2(new_n12453), .B(new_n12456), .C(new_n12459), .Y(new_n12842));
  NAND3xp33_ASAP7_75t_L     g12586(.A(new_n12836), .B(new_n12838), .C(new_n12839), .Y(new_n12843));
  OAI21xp33_ASAP7_75t_L     g12587(.A1(new_n12828), .A2(new_n12823), .B(new_n12834), .Y(new_n12844));
  AOI211xp5_ASAP7_75t_L     g12588(.A1(new_n12844), .A2(new_n12843), .B(new_n12469), .C(new_n12842), .Y(new_n12845));
  NOR2xp33_ASAP7_75t_L      g12589(.A(new_n4613), .B(new_n2930), .Y(new_n12846));
  AOI221xp5_ASAP7_75t_L     g12590(.A1(\b[34] ), .A2(new_n3129), .B1(\b[35] ), .B2(new_n2936), .C(new_n12846), .Y(new_n12847));
  O2A1O1Ixp33_ASAP7_75t_L   g12591(.A1(new_n2940), .A2(new_n4622), .B(new_n12847), .C(new_n2928), .Y(new_n12848));
  OAI21xp33_ASAP7_75t_L     g12592(.A1(new_n2940), .A2(new_n4622), .B(new_n12847), .Y(new_n12849));
  NAND2xp33_ASAP7_75t_L     g12593(.A(new_n2928), .B(new_n12849), .Y(new_n12850));
  OAI21xp33_ASAP7_75t_L     g12594(.A1(new_n2928), .A2(new_n12848), .B(new_n12850), .Y(new_n12851));
  OAI21xp33_ASAP7_75t_L     g12595(.A1(new_n12841), .A2(new_n12845), .B(new_n12851), .Y(new_n12852));
  OAI211xp5_ASAP7_75t_L     g12596(.A1(new_n12469), .A2(new_n12842), .B(new_n12843), .C(new_n12844), .Y(new_n12853));
  NAND3xp33_ASAP7_75t_L     g12597(.A(new_n12836), .B(new_n12838), .C(new_n12834), .Y(new_n12854));
  A2O1A1Ixp33_ASAP7_75t_L   g12598(.A1(new_n12854), .A2(new_n12834), .B(new_n12835), .C(new_n12470), .Y(new_n12855));
  INVx1_ASAP7_75t_L         g12599(.A(new_n12851), .Y(new_n12856));
  NAND3xp33_ASAP7_75t_L     g12600(.A(new_n12853), .B(new_n12855), .C(new_n12856), .Y(new_n12857));
  AO21x2_ASAP7_75t_L        g12601(.A1(new_n12857), .A2(new_n12852), .B(new_n12653), .Y(new_n12858));
  NAND3xp33_ASAP7_75t_L     g12602(.A(new_n12653), .B(new_n12857), .C(new_n12852), .Y(new_n12859));
  OAI22xp33_ASAP7_75t_L     g12603(.A1(new_n2572), .A2(new_n5074), .B1(new_n5311), .B2(new_n2410), .Y(new_n12860));
  AOI221xp5_ASAP7_75t_L     g12604(.A1(new_n2423), .A2(\b[39] ), .B1(new_n2417), .B2(new_n11869), .C(new_n12860), .Y(new_n12861));
  XNOR2x2_ASAP7_75t_L       g12605(.A(\a[26] ), .B(new_n12861), .Y(new_n12862));
  AOI21xp33_ASAP7_75t_L     g12606(.A1(new_n12858), .A2(new_n12859), .B(new_n12862), .Y(new_n12863));
  AND3x1_ASAP7_75t_L        g12607(.A(new_n12858), .B(new_n12862), .C(new_n12859), .Y(new_n12864));
  NOR2xp33_ASAP7_75t_L      g12608(.A(new_n12863), .B(new_n12864), .Y(new_n12865));
  A2O1A1Ixp33_ASAP7_75t_L   g12609(.A1(new_n12490), .A2(new_n12492), .B(new_n12486), .C(new_n12865), .Y(new_n12866));
  NOR2xp33_ASAP7_75t_L      g12610(.A(new_n12160), .B(new_n12167), .Y(new_n12867));
  A2O1A1O1Ixp25_ASAP7_75t_L g12611(.A1(new_n12168), .A2(new_n12867), .B(new_n12178), .C(new_n12490), .D(new_n12486), .Y(new_n12868));
  OAI21xp33_ASAP7_75t_L     g12612(.A1(new_n12863), .A2(new_n12864), .B(new_n12868), .Y(new_n12869));
  AO21x2_ASAP7_75t_L        g12613(.A1(new_n12869), .A2(new_n12866), .B(new_n12651), .Y(new_n12870));
  NAND3xp33_ASAP7_75t_L     g12614(.A(new_n12866), .B(new_n12869), .C(new_n12651), .Y(new_n12871));
  AOI21xp33_ASAP7_75t_L     g12615(.A1(new_n12870), .A2(new_n12871), .B(new_n12507), .Y(new_n12872));
  AND3x1_ASAP7_75t_L        g12616(.A(new_n12870), .B(new_n12507), .C(new_n12871), .Y(new_n12873));
  OAI21xp33_ASAP7_75t_L     g12617(.A1(new_n12872), .A2(new_n12873), .B(new_n12648), .Y(new_n12874));
  AO21x2_ASAP7_75t_L        g12618(.A1(new_n12871), .A2(new_n12870), .B(new_n12507), .Y(new_n12875));
  NAND3xp33_ASAP7_75t_L     g12619(.A(new_n12870), .B(new_n12507), .C(new_n12871), .Y(new_n12876));
  NAND3xp33_ASAP7_75t_L     g12620(.A(new_n12875), .B(new_n12647), .C(new_n12876), .Y(new_n12877));
  NAND2xp33_ASAP7_75t_L     g12621(.A(new_n12877), .B(new_n12874), .Y(new_n12878));
  INVx1_ASAP7_75t_L         g12622(.A(new_n12878), .Y(new_n12879));
  A2O1A1Ixp33_ASAP7_75t_L   g12623(.A1(new_n11903), .A2(new_n11899), .B(new_n12197), .C(new_n12200), .Y(new_n12880));
  OAI21xp33_ASAP7_75t_L     g12624(.A1(new_n12523), .A2(new_n12529), .B(new_n12880), .Y(new_n12881));
  NAND4xp25_ASAP7_75t_L     g12625(.A(new_n12881), .B(new_n12874), .C(new_n12877), .D(new_n12522), .Y(new_n12882));
  O2A1O1Ixp33_ASAP7_75t_L   g12626(.A1(new_n12644), .A2(new_n12879), .B(new_n12882), .C(new_n12642), .Y(new_n12883));
  OAI21xp33_ASAP7_75t_L     g12627(.A1(new_n12533), .A2(new_n12301), .B(new_n12535), .Y(new_n12884));
  INVx1_ASAP7_75t_L         g12628(.A(new_n12642), .Y(new_n12885));
  OAI211xp5_ASAP7_75t_L     g12629(.A1(new_n12644), .A2(new_n12879), .B(new_n12882), .C(new_n12885), .Y(new_n12886));
  AOI22xp33_ASAP7_75t_L     g12630(.A1(new_n12874), .A2(new_n12877), .B1(new_n12522), .B2(new_n12881), .Y(new_n12887));
  INVx1_ASAP7_75t_L         g12631(.A(new_n12877), .Y(new_n12888));
  NOR2xp33_ASAP7_75t_L      g12632(.A(new_n12643), .B(new_n12888), .Y(new_n12889));
  AOI211xp5_ASAP7_75t_L     g12633(.A1(new_n12874), .A2(new_n12889), .B(new_n12885), .C(new_n12887), .Y(new_n12890));
  A2O1A1Ixp33_ASAP7_75t_L   g12634(.A1(new_n12886), .A2(new_n12885), .B(new_n12890), .C(new_n12884), .Y(new_n12891));
  A2O1A1O1Ixp25_ASAP7_75t_L g12635(.A1(new_n12206), .A2(new_n12219), .B(new_n12221), .C(new_n12536), .D(new_n12528), .Y(new_n12892));
  OAI211xp5_ASAP7_75t_L     g12636(.A1(new_n12644), .A2(new_n12879), .B(new_n12882), .C(new_n12642), .Y(new_n12893));
  NAND2xp33_ASAP7_75t_L     g12637(.A(new_n12893), .B(new_n12892), .Y(new_n12894));
  OAI211xp5_ASAP7_75t_L     g12638(.A1(new_n12883), .A2(new_n12894), .B(new_n12891), .C(new_n12639), .Y(new_n12895));
  INVx1_ASAP7_75t_L         g12639(.A(new_n12639), .Y(new_n12896));
  A2O1A1Ixp33_ASAP7_75t_L   g12640(.A1(new_n12889), .A2(new_n12874), .B(new_n12887), .C(new_n12885), .Y(new_n12897));
  NAND2xp33_ASAP7_75t_L     g12641(.A(new_n12897), .B(new_n12893), .Y(new_n12898));
  NOR3xp33_ASAP7_75t_L      g12642(.A(new_n12884), .B(new_n12890), .C(new_n12883), .Y(new_n12899));
  A2O1A1Ixp33_ASAP7_75t_L   g12643(.A1(new_n12884), .A2(new_n12898), .B(new_n12899), .C(new_n12896), .Y(new_n12900));
  NAND2xp33_ASAP7_75t_L     g12644(.A(new_n12895), .B(new_n12900), .Y(new_n12901));
  O2A1O1Ixp33_ASAP7_75t_L   g12645(.A1(new_n12546), .A2(new_n12544), .B(new_n12548), .C(new_n12901), .Y(new_n12902));
  A2O1A1Ixp33_ASAP7_75t_L   g12646(.A1(new_n12556), .A2(new_n12555), .B(new_n12546), .C(new_n12548), .Y(new_n12903));
  AOI211xp5_ASAP7_75t_L     g12647(.A1(new_n12884), .A2(new_n12898), .B(new_n12896), .C(new_n12899), .Y(new_n12904));
  O2A1O1Ixp33_ASAP7_75t_L   g12648(.A1(new_n12883), .A2(new_n12894), .B(new_n12891), .C(new_n12639), .Y(new_n12905));
  NOR2xp33_ASAP7_75t_L      g12649(.A(new_n12905), .B(new_n12904), .Y(new_n12906));
  NOR2xp33_ASAP7_75t_L      g12650(.A(new_n12903), .B(new_n12906), .Y(new_n12907));
  OAI22xp33_ASAP7_75t_L     g12651(.A1(new_n1550), .A2(new_n9683), .B1(new_n9355), .B2(new_n712), .Y(new_n12908));
  AOI221xp5_ASAP7_75t_L     g12652(.A1(new_n640), .A2(\b[54] ), .B1(new_n718), .B2(new_n9717), .C(new_n12908), .Y(new_n12909));
  XNOR2x2_ASAP7_75t_L       g12653(.A(new_n637), .B(new_n12909), .Y(new_n12910));
  INVx1_ASAP7_75t_L         g12654(.A(new_n12910), .Y(new_n12911));
  NOR3xp33_ASAP7_75t_L      g12655(.A(new_n12902), .B(new_n12907), .C(new_n12911), .Y(new_n12912));
  A2O1A1Ixp33_ASAP7_75t_L   g12656(.A1(new_n12557), .A2(new_n12559), .B(new_n12547), .C(new_n12906), .Y(new_n12913));
  O2A1O1Ixp33_ASAP7_75t_L   g12657(.A1(new_n12542), .A2(new_n12543), .B(new_n12559), .C(new_n12547), .Y(new_n12914));
  NAND2xp33_ASAP7_75t_L     g12658(.A(new_n12901), .B(new_n12914), .Y(new_n12915));
  AOI21xp33_ASAP7_75t_L     g12659(.A1(new_n12915), .A2(new_n12913), .B(new_n12910), .Y(new_n12916));
  OAI21xp33_ASAP7_75t_L     g12660(.A1(new_n12562), .A2(new_n12298), .B(new_n12566), .Y(new_n12917));
  NOR3xp33_ASAP7_75t_L      g12661(.A(new_n12917), .B(new_n12916), .C(new_n12912), .Y(new_n12918));
  NAND3xp33_ASAP7_75t_L     g12662(.A(new_n12915), .B(new_n12913), .C(new_n12910), .Y(new_n12919));
  OAI21xp33_ASAP7_75t_L     g12663(.A1(new_n12907), .A2(new_n12902), .B(new_n12911), .Y(new_n12920));
  AOI21xp33_ASAP7_75t_L     g12664(.A1(new_n11926), .A2(new_n11655), .B(new_n11929), .Y(new_n12921));
  A2O1A1Ixp33_ASAP7_75t_L   g12665(.A1(new_n11571), .A2(new_n11931), .B(new_n12921), .C(new_n11926), .Y(new_n12922));
  A2O1A1O1Ixp25_ASAP7_75t_L g12666(.A1(new_n12297), .A2(new_n12922), .B(new_n12235), .C(new_n12567), .D(new_n12553), .Y(new_n12923));
  AOI21xp33_ASAP7_75t_L     g12667(.A1(new_n12920), .A2(new_n12919), .B(new_n12923), .Y(new_n12924));
  OAI22xp33_ASAP7_75t_L     g12668(.A1(new_n513), .A2(new_n10332), .B1(new_n10309), .B2(new_n506), .Y(new_n12925));
  AOI221xp5_ASAP7_75t_L     g12669(.A1(new_n475), .A2(\b[57] ), .B1(new_n483), .B2(new_n10991), .C(new_n12925), .Y(new_n12926));
  XNOR2x2_ASAP7_75t_L       g12670(.A(new_n466), .B(new_n12926), .Y(new_n12927));
  INVx1_ASAP7_75t_L         g12671(.A(new_n12927), .Y(new_n12928));
  NOR3xp33_ASAP7_75t_L      g12672(.A(new_n12924), .B(new_n12918), .C(new_n12928), .Y(new_n12929));
  NAND3xp33_ASAP7_75t_L     g12673(.A(new_n12923), .B(new_n12920), .C(new_n12919), .Y(new_n12930));
  NAND3xp33_ASAP7_75t_L     g12674(.A(new_n12915), .B(new_n12913), .C(new_n12911), .Y(new_n12931));
  A2O1A1Ixp33_ASAP7_75t_L   g12675(.A1(new_n12931), .A2(new_n12911), .B(new_n12912), .C(new_n12917), .Y(new_n12932));
  AOI21xp33_ASAP7_75t_L     g12676(.A1(new_n12930), .A2(new_n12932), .B(new_n12927), .Y(new_n12933));
  NOR2xp33_ASAP7_75t_L      g12677(.A(new_n11303), .B(new_n375), .Y(new_n12934));
  AOI221xp5_ASAP7_75t_L     g12678(.A1(\b[60] ), .A2(new_n361), .B1(new_n349), .B2(\b[59] ), .C(new_n12934), .Y(new_n12935));
  O2A1O1Ixp33_ASAP7_75t_L   g12679(.A1(new_n356), .A2(new_n11634), .B(new_n12935), .C(new_n346), .Y(new_n12936));
  OAI21xp33_ASAP7_75t_L     g12680(.A1(new_n356), .A2(new_n11634), .B(new_n12935), .Y(new_n12937));
  NAND2xp33_ASAP7_75t_L     g12681(.A(new_n346), .B(new_n12937), .Y(new_n12938));
  OAI21xp33_ASAP7_75t_L     g12682(.A1(new_n346), .A2(new_n12936), .B(new_n12938), .Y(new_n12939));
  INVx1_ASAP7_75t_L         g12683(.A(new_n12939), .Y(new_n12940));
  OAI21xp33_ASAP7_75t_L     g12684(.A1(new_n12933), .A2(new_n12929), .B(new_n12940), .Y(new_n12941));
  NAND3xp33_ASAP7_75t_L     g12685(.A(new_n12930), .B(new_n12932), .C(new_n12927), .Y(new_n12942));
  OAI21xp33_ASAP7_75t_L     g12686(.A1(new_n12918), .A2(new_n12924), .B(new_n12928), .Y(new_n12943));
  NAND3xp33_ASAP7_75t_L     g12687(.A(new_n12943), .B(new_n12942), .C(new_n12939), .Y(new_n12944));
  O2A1O1Ixp33_ASAP7_75t_L   g12688(.A1(new_n12583), .A2(new_n12589), .B(new_n12572), .C(new_n12587), .Y(new_n12945));
  NAND3xp33_ASAP7_75t_L     g12689(.A(new_n12941), .B(new_n12944), .C(new_n12945), .Y(new_n12946));
  AOI21xp33_ASAP7_75t_L     g12690(.A1(new_n12943), .A2(new_n12942), .B(new_n12939), .Y(new_n12947));
  NOR3xp33_ASAP7_75t_L      g12691(.A(new_n12929), .B(new_n12933), .C(new_n12940), .Y(new_n12948));
  A2O1A1Ixp33_ASAP7_75t_L   g12692(.A1(new_n12588), .A2(new_n12590), .B(new_n12586), .C(new_n12576), .Y(new_n12949));
  OAI21xp33_ASAP7_75t_L     g12693(.A1(new_n12947), .A2(new_n12948), .B(new_n12949), .Y(new_n12950));
  NOR2xp33_ASAP7_75t_L      g12694(.A(new_n12258), .B(new_n287), .Y(new_n12951));
  AOI221xp5_ASAP7_75t_L     g12695(.A1(\b[62] ), .A2(new_n264), .B1(\b[63] ), .B2(new_n283), .C(new_n12951), .Y(new_n12952));
  INVx1_ASAP7_75t_L         g12696(.A(new_n12952), .Y(new_n12953));
  INVx1_ASAP7_75t_L         g12697(.A(new_n12604), .Y(new_n12954));
  NOR2xp33_ASAP7_75t_L      g12698(.A(\b[63] ), .B(new_n12603), .Y(new_n12955));
  INVx1_ASAP7_75t_L         g12699(.A(\b[63] ), .Y(new_n12956));
  NOR2xp33_ASAP7_75t_L      g12700(.A(\b[62] ), .B(new_n12956), .Y(new_n12957));
  NOR2xp33_ASAP7_75t_L      g12701(.A(new_n12955), .B(new_n12957), .Y(new_n12958));
  O2A1O1Ixp33_ASAP7_75t_L   g12702(.A1(new_n12608), .A2(new_n12607), .B(new_n12954), .C(new_n12958), .Y(new_n12959));
  AND3x1_ASAP7_75t_L        g12703(.A(new_n12606), .B(new_n12958), .C(new_n12954), .Y(new_n12960));
  NOR2xp33_ASAP7_75t_L      g12704(.A(new_n12959), .B(new_n12960), .Y(new_n12961));
  A2O1A1Ixp33_ASAP7_75t_L   g12705(.A1(new_n12961), .A2(new_n273), .B(new_n12953), .C(\a[2] ), .Y(new_n12962));
  A2O1A1Ixp33_ASAP7_75t_L   g12706(.A1(new_n12961), .A2(new_n273), .B(new_n12953), .C(new_n257), .Y(new_n12963));
  INVx1_ASAP7_75t_L         g12707(.A(new_n12963), .Y(new_n12964));
  AOI21xp33_ASAP7_75t_L     g12708(.A1(new_n12962), .A2(\a[2] ), .B(new_n12964), .Y(new_n12965));
  NAND3xp33_ASAP7_75t_L     g12709(.A(new_n12950), .B(new_n12946), .C(new_n12965), .Y(new_n12966));
  NOR3xp33_ASAP7_75t_L      g12710(.A(new_n12948), .B(new_n12949), .C(new_n12947), .Y(new_n12967));
  AOI21xp33_ASAP7_75t_L     g12711(.A1(new_n12941), .A2(new_n12944), .B(new_n12945), .Y(new_n12968));
  NAND2xp33_ASAP7_75t_L     g12712(.A(\a[2] ), .B(new_n12962), .Y(new_n12969));
  NAND2xp33_ASAP7_75t_L     g12713(.A(new_n12963), .B(new_n12969), .Y(new_n12970));
  OAI21xp33_ASAP7_75t_L     g12714(.A1(new_n12968), .A2(new_n12967), .B(new_n12970), .Y(new_n12971));
  AOI21xp33_ASAP7_75t_L     g12715(.A1(new_n12971), .A2(new_n12966), .B(new_n12632), .Y(new_n12972));
  NOR3xp33_ASAP7_75t_L      g12716(.A(new_n12967), .B(new_n12968), .C(new_n12970), .Y(new_n12973));
  AOI21xp33_ASAP7_75t_L     g12717(.A1(new_n12950), .A2(new_n12946), .B(new_n12965), .Y(new_n12974));
  OAI21xp33_ASAP7_75t_L     g12718(.A1(new_n12974), .A2(new_n12973), .B(new_n12632), .Y(new_n12975));
  A2O1A1O1Ixp25_ASAP7_75t_L g12719(.A1(new_n12290), .A2(new_n12282), .B(new_n12281), .C(new_n12625), .D(new_n12620), .Y(new_n12976));
  O2A1O1Ixp33_ASAP7_75t_L   g12720(.A1(new_n12632), .A2(new_n12972), .B(new_n12975), .C(new_n12976), .Y(new_n12977));
  NAND3xp33_ASAP7_75t_L     g12721(.A(new_n12971), .B(new_n12966), .C(new_n12631), .Y(new_n12978));
  NAND2xp33_ASAP7_75t_L     g12722(.A(new_n12978), .B(new_n12975), .Y(new_n12979));
  NOR3xp33_ASAP7_75t_L      g12723(.A(new_n12627), .B(new_n12979), .C(new_n12620), .Y(new_n12980));
  NOR2xp33_ASAP7_75t_L      g12724(.A(new_n12980), .B(new_n12977), .Y(\f[63] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g12725(.A1(new_n12625), .A2(new_n12628), .B(new_n12620), .C(new_n12979), .D(new_n12972), .Y(new_n12982));
  A2O1A1O1Ixp25_ASAP7_75t_L g12726(.A1(new_n12962), .A2(\a[2] ), .B(new_n12964), .C(new_n12946), .D(new_n12968), .Y(new_n12983));
  INVx1_ASAP7_75t_L         g12727(.A(new_n12983), .Y(new_n12984));
  AOI22xp33_ASAP7_75t_L     g12728(.A1(new_n264), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n286), .Y(new_n12985));
  O2A1O1Ixp33_ASAP7_75t_L   g12729(.A1(new_n12258), .A2(new_n12607), .B(new_n12603), .C(new_n12956), .Y(new_n12986));
  NOR2xp33_ASAP7_75t_L      g12730(.A(new_n12956), .B(new_n12986), .Y(new_n12987));
  INVx1_ASAP7_75t_L         g12731(.A(new_n12987), .Y(new_n12988));
  INVx1_ASAP7_75t_L         g12732(.A(new_n12606), .Y(new_n12989));
  A2O1A1Ixp33_ASAP7_75t_L   g12733(.A1(\b[62] ), .A2(\b[61] ), .B(new_n12989), .C(new_n12955), .Y(new_n12990));
  A2O1A1Ixp33_ASAP7_75t_L   g12734(.A1(new_n12990), .A2(new_n12988), .B(new_n279), .C(new_n12985), .Y(new_n12991));
  NOR2xp33_ASAP7_75t_L      g12735(.A(new_n257), .B(new_n12991), .Y(new_n12992));
  O2A1O1Ixp33_ASAP7_75t_L   g12736(.A1(new_n12604), .A2(new_n12989), .B(new_n12955), .C(new_n12987), .Y(new_n12993));
  O2A1O1Ixp33_ASAP7_75t_L   g12737(.A1(new_n279), .A2(new_n12993), .B(new_n12985), .C(\a[2] ), .Y(new_n12994));
  NOR2xp33_ASAP7_75t_L      g12738(.A(new_n12994), .B(new_n12992), .Y(new_n12995));
  INVx1_ASAP7_75t_L         g12739(.A(new_n12995), .Y(new_n12996));
  NOR2xp33_ASAP7_75t_L      g12740(.A(new_n12918), .B(new_n12924), .Y(new_n12997));
  NOR3xp33_ASAP7_75t_L      g12741(.A(new_n12924), .B(new_n12918), .C(new_n12927), .Y(new_n12998));
  O2A1O1Ixp33_ASAP7_75t_L   g12742(.A1(new_n12997), .A2(new_n12933), .B(new_n12939), .C(new_n12998), .Y(new_n12999));
  INVx1_ASAP7_75t_L         g12743(.A(new_n12999), .Y(new_n13000));
  A2O1A1Ixp33_ASAP7_75t_L   g12744(.A1(new_n12910), .A2(new_n12919), .B(new_n12923), .C(new_n12931), .Y(new_n13001));
  OAI22xp33_ASAP7_75t_L     g12745(.A1(new_n1550), .A2(new_n9709), .B1(new_n9683), .B2(new_n712), .Y(new_n13002));
  AOI221xp5_ASAP7_75t_L     g12746(.A1(new_n640), .A2(\b[55] ), .B1(new_n718), .B2(new_n10320), .C(new_n13002), .Y(new_n13003));
  XNOR2x2_ASAP7_75t_L       g12747(.A(new_n637), .B(new_n13003), .Y(new_n13004));
  INVx1_ASAP7_75t_L         g12748(.A(new_n13004), .Y(new_n13005));
  A2O1A1O1Ixp25_ASAP7_75t_L g12749(.A1(new_n12559), .A2(new_n12557), .B(new_n12547), .C(new_n12900), .D(new_n12904), .Y(new_n13006));
  OAI22xp33_ASAP7_75t_L     g12750(.A1(new_n980), .A2(new_n8755), .B1(new_n8779), .B2(new_n864), .Y(new_n13007));
  AOI221xp5_ASAP7_75t_L     g12751(.A1(new_n886), .A2(\b[52] ), .B1(new_n873), .B2(new_n9367), .C(new_n13007), .Y(new_n13008));
  XNOR2x2_ASAP7_75t_L       g12752(.A(new_n867), .B(new_n13008), .Y(new_n13009));
  A2O1A1Ixp33_ASAP7_75t_L   g12753(.A1(new_n12893), .A2(new_n12642), .B(new_n12892), .C(new_n12886), .Y(new_n13010));
  OAI22xp33_ASAP7_75t_L     g12754(.A1(new_n1285), .A2(new_n7552), .B1(new_n7860), .B2(new_n2118), .Y(new_n13011));
  AOI221xp5_ASAP7_75t_L     g12755(.A1(new_n1209), .A2(\b[49] ), .B1(new_n1216), .B2(new_n8438), .C(new_n13011), .Y(new_n13012));
  XNOR2x2_ASAP7_75t_L       g12756(.A(new_n1206), .B(new_n13012), .Y(new_n13013));
  INVx1_ASAP7_75t_L         g12757(.A(new_n13013), .Y(new_n13014));
  OAI22xp33_ASAP7_75t_L     g12758(.A1(new_n1654), .A2(new_n6944), .B1(new_n7249), .B2(new_n1517), .Y(new_n13015));
  AOI221xp5_ASAP7_75t_L     g12759(.A1(new_n1511), .A2(\b[46] ), .B1(new_n1513), .B2(new_n7278), .C(new_n13015), .Y(new_n13016));
  XNOR2x2_ASAP7_75t_L       g12760(.A(new_n1501), .B(new_n13016), .Y(new_n13017));
  INVx1_ASAP7_75t_L         g12761(.A(new_n13017), .Y(new_n13018));
  NAND2xp33_ASAP7_75t_L     g12762(.A(new_n12869), .B(new_n12866), .Y(new_n13019));
  AO21x2_ASAP7_75t_L        g12763(.A1(new_n12859), .A2(new_n12858), .B(new_n12862), .Y(new_n13020));
  A2O1A1O1Ixp25_ASAP7_75t_L g12764(.A1(new_n12492), .A2(new_n12490), .B(new_n12486), .C(new_n13020), .D(new_n12864), .Y(new_n13021));
  NOR2xp33_ASAP7_75t_L      g12765(.A(new_n3079), .B(new_n4908), .Y(new_n13022));
  AOI221xp5_ASAP7_75t_L     g12766(.A1(\b[26] ), .A2(new_n5139), .B1(\b[27] ), .B2(new_n4916), .C(new_n13022), .Y(new_n13023));
  OAI21xp33_ASAP7_75t_L     g12767(.A1(new_n4911), .A2(new_n3087), .B(new_n13023), .Y(new_n13024));
  NOR2xp33_ASAP7_75t_L      g12768(.A(new_n4906), .B(new_n13024), .Y(new_n13025));
  O2A1O1Ixp33_ASAP7_75t_L   g12769(.A1(new_n4911), .A2(new_n3087), .B(new_n13023), .C(\a[38] ), .Y(new_n13026));
  O2A1O1Ixp33_ASAP7_75t_L   g12770(.A1(new_n12338), .A2(new_n12668), .B(new_n12697), .C(new_n12704), .Y(new_n13027));
  INVx1_ASAP7_75t_L         g12771(.A(new_n12672), .Y(new_n13028));
  NOR2xp33_ASAP7_75t_L      g12772(.A(new_n11987), .B(new_n12670), .Y(new_n13029));
  INVx1_ASAP7_75t_L         g12773(.A(new_n13029), .Y(new_n13030));
  NOR2xp33_ASAP7_75t_L      g12774(.A(new_n284), .B(new_n13030), .Y(new_n13031));
  O2A1O1Ixp33_ASAP7_75t_L   g12775(.A1(new_n12669), .A2(new_n12671), .B(\b[1] ), .C(new_n13031), .Y(new_n13032));
  INVx1_ASAP7_75t_L         g12776(.A(new_n13032), .Y(new_n13033));
  NAND2xp33_ASAP7_75t_L     g12777(.A(\b[4] ), .B(new_n11995), .Y(new_n13034));
  OAI221xp5_ASAP7_75t_L     g12778(.A1(new_n12318), .A2(new_n301), .B1(new_n289), .B2(new_n12320), .C(new_n13034), .Y(new_n13035));
  A2O1A1Ixp33_ASAP7_75t_L   g12779(.A1(new_n342), .A2(new_n11997), .B(new_n13035), .C(\a[62] ), .Y(new_n13036));
  A2O1A1Ixp33_ASAP7_75t_L   g12780(.A1(new_n342), .A2(new_n11997), .B(new_n13035), .C(new_n11987), .Y(new_n13037));
  INVx1_ASAP7_75t_L         g12781(.A(new_n13037), .Y(new_n13038));
  A2O1A1Ixp33_ASAP7_75t_L   g12782(.A1(\a[62] ), .A2(new_n13036), .B(new_n13038), .C(new_n13033), .Y(new_n13039));
  A2O1A1Ixp33_ASAP7_75t_L   g12783(.A1(\a[62] ), .A2(new_n13036), .B(new_n13038), .C(new_n13032), .Y(new_n13040));
  INVx1_ASAP7_75t_L         g12784(.A(new_n13040), .Y(new_n13041));
  A2O1A1O1Ixp25_ASAP7_75t_L g12785(.A1(new_n13028), .A2(\b[1] ), .B(new_n13031), .C(new_n13039), .D(new_n13041), .Y(new_n13042));
  O2A1O1Ixp33_ASAP7_75t_L   g12786(.A1(new_n12673), .A2(new_n12676), .B(new_n12682), .C(new_n12674), .Y(new_n13043));
  NAND2xp33_ASAP7_75t_L     g12787(.A(new_n13043), .B(new_n13042), .Y(new_n13044));
  INVx1_ASAP7_75t_L         g12788(.A(new_n13043), .Y(new_n13045));
  A2O1A1Ixp33_ASAP7_75t_L   g12789(.A1(new_n13039), .A2(new_n13033), .B(new_n13041), .C(new_n13045), .Y(new_n13046));
  NOR2xp33_ASAP7_75t_L      g12790(.A(new_n384), .B(new_n11354), .Y(new_n13047));
  AOI221xp5_ASAP7_75t_L     g12791(.A1(\b[7] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[6] ), .C(new_n13047), .Y(new_n13048));
  O2A1O1Ixp33_ASAP7_75t_L   g12792(.A1(new_n11053), .A2(new_n456), .B(new_n13048), .C(new_n11048), .Y(new_n13049));
  OAI21xp33_ASAP7_75t_L     g12793(.A1(new_n11053), .A2(new_n456), .B(new_n13048), .Y(new_n13050));
  NAND2xp33_ASAP7_75t_L     g12794(.A(new_n11048), .B(new_n13050), .Y(new_n13051));
  OAI21xp33_ASAP7_75t_L     g12795(.A1(new_n11048), .A2(new_n13049), .B(new_n13051), .Y(new_n13052));
  AOI21xp33_ASAP7_75t_L     g12796(.A1(new_n13046), .A2(new_n13044), .B(new_n13052), .Y(new_n13053));
  NAND3xp33_ASAP7_75t_L     g12797(.A(new_n13046), .B(new_n13044), .C(new_n13052), .Y(new_n13054));
  INVx1_ASAP7_75t_L         g12798(.A(new_n13054), .Y(new_n13055));
  NOR3xp33_ASAP7_75t_L      g12799(.A(new_n13055), .B(new_n13053), .C(new_n13027), .Y(new_n13056));
  INVx1_ASAP7_75t_L         g12800(.A(new_n13027), .Y(new_n13057));
  INVx1_ASAP7_75t_L         g12801(.A(new_n13053), .Y(new_n13058));
  AOI21xp33_ASAP7_75t_L     g12802(.A1(new_n13058), .A2(new_n13054), .B(new_n13057), .Y(new_n13059));
  OAI22xp33_ASAP7_75t_L     g12803(.A1(new_n10390), .A2(new_n534), .B1(new_n590), .B2(new_n10388), .Y(new_n13060));
  AOI221xp5_ASAP7_75t_L     g12804(.A1(new_n10086), .A2(\b[10] ), .B1(new_n10386), .B2(new_n690), .C(new_n13060), .Y(new_n13061));
  XNOR2x2_ASAP7_75t_L       g12805(.A(new_n10083), .B(new_n13061), .Y(new_n13062));
  INVx1_ASAP7_75t_L         g12806(.A(new_n13062), .Y(new_n13063));
  OR3x1_ASAP7_75t_L         g12807(.A(new_n13059), .B(new_n13056), .C(new_n13063), .Y(new_n13064));
  OAI21xp33_ASAP7_75t_L     g12808(.A1(new_n13056), .A2(new_n13059), .B(new_n13063), .Y(new_n13065));
  O2A1O1Ixp33_ASAP7_75t_L   g12809(.A1(new_n12716), .A2(new_n12706), .B(new_n12667), .C(new_n12732), .Y(new_n13066));
  NAND3xp33_ASAP7_75t_L     g12810(.A(new_n13066), .B(new_n13064), .C(new_n13065), .Y(new_n13067));
  NOR3xp33_ASAP7_75t_L      g12811(.A(new_n13059), .B(new_n13056), .C(new_n13062), .Y(new_n13068));
  O2A1O1Ixp33_ASAP7_75t_L   g12812(.A1(new_n13062), .A2(new_n13068), .B(new_n13064), .C(new_n13066), .Y(new_n13069));
  INVx1_ASAP7_75t_L         g12813(.A(new_n13069), .Y(new_n13070));
  OAI22xp33_ASAP7_75t_L     g12814(.A1(new_n9440), .A2(new_n748), .B1(new_n833), .B2(new_n10400), .Y(new_n13071));
  AOI221xp5_ASAP7_75t_L     g12815(.A1(new_n9102), .A2(\b[13] ), .B1(new_n9437), .B2(new_n1166), .C(new_n13071), .Y(new_n13072));
  XNOR2x2_ASAP7_75t_L       g12816(.A(new_n9099), .B(new_n13072), .Y(new_n13073));
  INVx1_ASAP7_75t_L         g12817(.A(new_n13073), .Y(new_n13074));
  AOI21xp33_ASAP7_75t_L     g12818(.A1(new_n13070), .A2(new_n13067), .B(new_n13074), .Y(new_n13075));
  INVx1_ASAP7_75t_L         g12819(.A(new_n13067), .Y(new_n13076));
  NOR3xp33_ASAP7_75t_L      g12820(.A(new_n13076), .B(new_n13069), .C(new_n13073), .Y(new_n13077));
  INVx1_ASAP7_75t_L         g12821(.A(new_n12734), .Y(new_n13078));
  O2A1O1Ixp33_ASAP7_75t_L   g12822(.A1(new_n12366), .A2(new_n12372), .B(new_n12730), .C(new_n13078), .Y(new_n13079));
  NOR3xp33_ASAP7_75t_L      g12823(.A(new_n13075), .B(new_n13079), .C(new_n13077), .Y(new_n13080));
  OAI21xp33_ASAP7_75t_L     g12824(.A1(new_n13069), .A2(new_n13076), .B(new_n13073), .Y(new_n13081));
  NAND3xp33_ASAP7_75t_L     g12825(.A(new_n13070), .B(new_n13067), .C(new_n13074), .Y(new_n13082));
  A2O1A1Ixp33_ASAP7_75t_L   g12826(.A1(new_n12361), .A2(new_n12362), .B(new_n12737), .C(new_n12734), .Y(new_n13083));
  AOI21xp33_ASAP7_75t_L     g12827(.A1(new_n13082), .A2(new_n13081), .B(new_n13083), .Y(new_n13084));
  OAI22xp33_ASAP7_75t_L     g12828(.A1(new_n8483), .A2(new_n960), .B1(new_n1043), .B2(new_n10065), .Y(new_n13085));
  AOI221xp5_ASAP7_75t_L     g12829(.A1(new_n8175), .A2(\b[16] ), .B1(new_n8490), .B2(new_n1156), .C(new_n13085), .Y(new_n13086));
  XNOR2x2_ASAP7_75t_L       g12830(.A(\a[50] ), .B(new_n13086), .Y(new_n13087));
  OR3x1_ASAP7_75t_L         g12831(.A(new_n13084), .B(new_n13080), .C(new_n13087), .Y(new_n13088));
  OAI21xp33_ASAP7_75t_L     g12832(.A1(new_n13080), .A2(new_n13084), .B(new_n13087), .Y(new_n13089));
  NAND4xp25_ASAP7_75t_L     g12833(.A(new_n13088), .B(new_n12746), .C(new_n12749), .D(new_n13089), .Y(new_n13090));
  NOR3xp33_ASAP7_75t_L      g12834(.A(new_n13084), .B(new_n13080), .C(new_n13087), .Y(new_n13091));
  OA21x2_ASAP7_75t_L        g12835(.A1(new_n13080), .A2(new_n13084), .B(new_n13087), .Y(new_n13092));
  INVx1_ASAP7_75t_L         g12836(.A(new_n12748), .Y(new_n13093));
  A2O1A1Ixp33_ASAP7_75t_L   g12837(.A1(new_n12742), .A2(new_n12743), .B(new_n13093), .C(new_n12746), .Y(new_n13094));
  OAI21xp33_ASAP7_75t_L     g12838(.A1(new_n13091), .A2(new_n13092), .B(new_n13094), .Y(new_n13095));
  OAI22xp33_ASAP7_75t_L     g12839(.A1(new_n7614), .A2(new_n1349), .B1(new_n1458), .B2(new_n7312), .Y(new_n13096));
  AOI221xp5_ASAP7_75t_L     g12840(.A1(new_n7334), .A2(\b[19] ), .B1(new_n7322), .B2(new_n1607), .C(new_n13096), .Y(new_n13097));
  XNOR2x2_ASAP7_75t_L       g12841(.A(\a[47] ), .B(new_n13097), .Y(new_n13098));
  AOI21xp33_ASAP7_75t_L     g12842(.A1(new_n13090), .A2(new_n13095), .B(new_n13098), .Y(new_n13099));
  AND3x1_ASAP7_75t_L        g12843(.A(new_n13090), .B(new_n13095), .C(new_n13098), .Y(new_n13100));
  A2O1A1O1Ixp25_ASAP7_75t_L g12844(.A1(new_n12385), .A2(new_n12654), .B(new_n12661), .C(new_n12763), .D(new_n12760), .Y(new_n13101));
  NOR3xp33_ASAP7_75t_L      g12845(.A(new_n13100), .B(new_n13101), .C(new_n13099), .Y(new_n13102));
  AO21x2_ASAP7_75t_L        g12846(.A1(new_n13095), .A2(new_n13090), .B(new_n13098), .Y(new_n13103));
  NAND3xp33_ASAP7_75t_L     g12847(.A(new_n13090), .B(new_n13095), .C(new_n13098), .Y(new_n13104));
  A2O1A1Ixp33_ASAP7_75t_L   g12848(.A1(new_n12655), .A2(new_n12396), .B(new_n12756), .C(new_n12764), .Y(new_n13105));
  AOI21xp33_ASAP7_75t_L     g12849(.A1(new_n13104), .A2(new_n13103), .B(new_n13105), .Y(new_n13106));
  OAI22xp33_ASAP7_75t_L     g12850(.A1(new_n7304), .A2(new_n1895), .B1(new_n1745), .B2(new_n6741), .Y(new_n13107));
  AOI221xp5_ASAP7_75t_L     g12851(.A1(new_n6442), .A2(\b[22] ), .B1(new_n6450), .B2(new_n2056), .C(new_n13107), .Y(new_n13108));
  XNOR2x2_ASAP7_75t_L       g12852(.A(\a[44] ), .B(new_n13108), .Y(new_n13109));
  NOR3xp33_ASAP7_75t_L      g12853(.A(new_n13106), .B(new_n13102), .C(new_n13109), .Y(new_n13110));
  OA21x2_ASAP7_75t_L        g12854(.A1(new_n13102), .A2(new_n13106), .B(new_n13109), .Y(new_n13111));
  A2O1A1O1Ixp25_ASAP7_75t_L g12855(.A1(new_n12404), .A2(new_n12106), .B(new_n12657), .C(new_n12775), .D(new_n12766), .Y(new_n13112));
  INVx1_ASAP7_75t_L         g12856(.A(new_n13112), .Y(new_n13113));
  NOR3xp33_ASAP7_75t_L      g12857(.A(new_n13113), .B(new_n13111), .C(new_n13110), .Y(new_n13114));
  NOR2xp33_ASAP7_75t_L      g12858(.A(new_n13110), .B(new_n13111), .Y(new_n13115));
  O2A1O1Ixp33_ASAP7_75t_L   g12859(.A1(new_n12773), .A2(new_n12776), .B(new_n12774), .C(new_n13115), .Y(new_n13116));
  NOR2xp33_ASAP7_75t_L      g12860(.A(new_n13114), .B(new_n13116), .Y(new_n13117));
  NAND2xp33_ASAP7_75t_L     g12861(.A(new_n13112), .B(new_n13115), .Y(new_n13118));
  NOR2xp33_ASAP7_75t_L      g12862(.A(new_n13102), .B(new_n13106), .Y(new_n13119));
  INVx1_ASAP7_75t_L         g12863(.A(new_n13109), .Y(new_n13120));
  NOR3xp33_ASAP7_75t_L      g12864(.A(new_n13120), .B(new_n13106), .C(new_n13102), .Y(new_n13121));
  INVx1_ASAP7_75t_L         g12865(.A(new_n13121), .Y(new_n13122));
  A2O1A1Ixp33_ASAP7_75t_L   g12866(.A1(new_n13122), .A2(new_n13119), .B(new_n13111), .C(new_n13113), .Y(new_n13123));
  OAI22xp33_ASAP7_75t_L     g12867(.A1(new_n5640), .A2(new_n2205), .B1(new_n2188), .B2(new_n5925), .Y(new_n13124));
  AOI221xp5_ASAP7_75t_L     g12868(.A1(new_n5629), .A2(\b[25] ), .B1(new_n5637), .B2(new_n5001), .C(new_n13124), .Y(new_n13125));
  XNOR2x2_ASAP7_75t_L       g12869(.A(new_n5626), .B(new_n13125), .Y(new_n13126));
  INVx1_ASAP7_75t_L         g12870(.A(new_n13126), .Y(new_n13127));
  NAND3xp33_ASAP7_75t_L     g12871(.A(new_n13123), .B(new_n13118), .C(new_n13127), .Y(new_n13128));
  AOI21xp33_ASAP7_75t_L     g12872(.A1(new_n13123), .A2(new_n13118), .B(new_n13126), .Y(new_n13129));
  AOI21xp33_ASAP7_75t_L     g12873(.A1(new_n13128), .A2(new_n13117), .B(new_n13129), .Y(new_n13130));
  O2A1O1Ixp33_ASAP7_75t_L   g12874(.A1(new_n12425), .A2(new_n12419), .B(new_n12793), .C(new_n12802), .Y(new_n13131));
  NAND2xp33_ASAP7_75t_L     g12875(.A(new_n13131), .B(new_n13130), .Y(new_n13132));
  INVx1_ASAP7_75t_L         g12876(.A(new_n12802), .Y(new_n13133));
  A2O1A1Ixp33_ASAP7_75t_L   g12877(.A1(new_n12801), .A2(new_n12788), .B(new_n12789), .C(new_n13133), .Y(new_n13134));
  A2O1A1Ixp33_ASAP7_75t_L   g12878(.A1(new_n13117), .A2(new_n13128), .B(new_n13129), .C(new_n13134), .Y(new_n13135));
  O2A1O1Ixp33_ASAP7_75t_L   g12879(.A1(new_n4911), .A2(new_n3087), .B(new_n13023), .C(new_n4906), .Y(new_n13136));
  NAND2xp33_ASAP7_75t_L     g12880(.A(new_n4906), .B(new_n13024), .Y(new_n13137));
  OAI21xp33_ASAP7_75t_L     g12881(.A1(new_n4906), .A2(new_n13136), .B(new_n13137), .Y(new_n13138));
  NAND3xp33_ASAP7_75t_L     g12882(.A(new_n13135), .B(new_n13132), .C(new_n13138), .Y(new_n13139));
  NAND3xp33_ASAP7_75t_L     g12883(.A(new_n13123), .B(new_n13118), .C(new_n13126), .Y(new_n13140));
  OAI21xp33_ASAP7_75t_L     g12884(.A1(new_n13114), .A2(new_n13116), .B(new_n13127), .Y(new_n13141));
  AND3x1_ASAP7_75t_L        g12885(.A(new_n13131), .B(new_n13141), .C(new_n13140), .Y(new_n13142));
  O2A1O1Ixp33_ASAP7_75t_L   g12886(.A1(new_n12801), .A2(new_n12780), .B(new_n12794), .C(new_n13130), .Y(new_n13143));
  NOR3xp33_ASAP7_75t_L      g12887(.A(new_n13142), .B(new_n13143), .C(new_n13138), .Y(new_n13144));
  O2A1O1Ixp33_ASAP7_75t_L   g12888(.A1(new_n13025), .A2(new_n13026), .B(new_n13139), .C(new_n13144), .Y(new_n13145));
  NAND3xp33_ASAP7_75t_L     g12889(.A(new_n13145), .B(new_n12819), .C(new_n12809), .Y(new_n13146));
  A2O1A1Ixp33_ASAP7_75t_L   g12890(.A1(new_n12798), .A2(new_n12799), .B(new_n12812), .C(new_n12809), .Y(new_n13147));
  A2O1A1Ixp33_ASAP7_75t_L   g12891(.A1(new_n13139), .A2(new_n13138), .B(new_n13144), .C(new_n13147), .Y(new_n13148));
  OAI22xp33_ASAP7_75t_L     g12892(.A1(new_n4397), .A2(new_n3098), .B1(new_n3456), .B2(new_n4142), .Y(new_n13149));
  AOI221xp5_ASAP7_75t_L     g12893(.A1(new_n4156), .A2(\b[31] ), .B1(new_n4151), .B2(new_n4317), .C(new_n13149), .Y(new_n13150));
  XNOR2x2_ASAP7_75t_L       g12894(.A(new_n4145), .B(new_n13150), .Y(new_n13151));
  INVx1_ASAP7_75t_L         g12895(.A(new_n13151), .Y(new_n13152));
  AOI21xp33_ASAP7_75t_L     g12896(.A1(new_n13146), .A2(new_n13148), .B(new_n13152), .Y(new_n13153));
  AO21x2_ASAP7_75t_L        g12897(.A1(new_n13138), .A2(new_n13139), .B(new_n13144), .Y(new_n13154));
  NOR2xp33_ASAP7_75t_L      g12898(.A(new_n13147), .B(new_n13154), .Y(new_n13155));
  INVx1_ASAP7_75t_L         g12899(.A(new_n13148), .Y(new_n13156));
  NOR3xp33_ASAP7_75t_L      g12900(.A(new_n13155), .B(new_n13156), .C(new_n13151), .Y(new_n13157));
  NOR2xp33_ASAP7_75t_L      g12901(.A(new_n13153), .B(new_n13157), .Y(new_n13158));
  A2O1A1O1Ixp25_ASAP7_75t_L g12902(.A1(new_n12446), .A2(new_n12445), .B(new_n12450), .C(new_n12817), .D(new_n12825), .Y(new_n13159));
  INVx1_ASAP7_75t_L         g12903(.A(new_n13159), .Y(new_n13160));
  NAND2xp33_ASAP7_75t_L     g12904(.A(new_n13160), .B(new_n13158), .Y(new_n13161));
  OAI21xp33_ASAP7_75t_L     g12905(.A1(new_n13156), .A2(new_n13155), .B(new_n13151), .Y(new_n13162));
  NAND3xp33_ASAP7_75t_L     g12906(.A(new_n13146), .B(new_n13148), .C(new_n13152), .Y(new_n13163));
  NAND2xp33_ASAP7_75t_L     g12907(.A(new_n13163), .B(new_n13162), .Y(new_n13164));
  NAND2xp33_ASAP7_75t_L     g12908(.A(new_n13159), .B(new_n13164), .Y(new_n13165));
  OAI22xp33_ASAP7_75t_L     g12909(.A1(new_n3703), .A2(new_n3891), .B1(new_n4101), .B2(new_n3509), .Y(new_n13166));
  AOI221xp5_ASAP7_75t_L     g12910(.A1(new_n3503), .A2(\b[34] ), .B1(new_n3505), .B2(new_n5599), .C(new_n13166), .Y(new_n13167));
  XNOR2x2_ASAP7_75t_L       g12911(.A(new_n3493), .B(new_n13167), .Y(new_n13168));
  NAND3xp33_ASAP7_75t_L     g12912(.A(new_n13161), .B(new_n13165), .C(new_n13168), .Y(new_n13169));
  NOR2xp33_ASAP7_75t_L      g12913(.A(new_n13159), .B(new_n13164), .Y(new_n13170));
  NOR2xp33_ASAP7_75t_L      g12914(.A(new_n13160), .B(new_n13158), .Y(new_n13171));
  INVx1_ASAP7_75t_L         g12915(.A(new_n13168), .Y(new_n13172));
  OAI21xp33_ASAP7_75t_L     g12916(.A1(new_n13170), .A2(new_n13171), .B(new_n13172), .Y(new_n13173));
  OAI22xp33_ASAP7_75t_L     g12917(.A1(new_n12842), .A2(new_n12469), .B1(new_n12840), .B2(new_n12835), .Y(new_n13174));
  NAND4xp25_ASAP7_75t_L     g12918(.A(new_n13173), .B(new_n13169), .C(new_n12854), .D(new_n13174), .Y(new_n13175));
  NOR3xp33_ASAP7_75t_L      g12919(.A(new_n13171), .B(new_n13170), .C(new_n13172), .Y(new_n13176));
  AOI21xp33_ASAP7_75t_L     g12920(.A1(new_n13161), .A2(new_n13165), .B(new_n13168), .Y(new_n13177));
  A2O1A1Ixp33_ASAP7_75t_L   g12921(.A1(new_n12843), .A2(new_n12839), .B(new_n12470), .C(new_n12854), .Y(new_n13178));
  OAI21xp33_ASAP7_75t_L     g12922(.A1(new_n13177), .A2(new_n13176), .B(new_n13178), .Y(new_n13179));
  OAI22xp33_ASAP7_75t_L     g12923(.A1(new_n3133), .A2(new_n4581), .B1(new_n4613), .B2(new_n2925), .Y(new_n13180));
  AOI221xp5_ASAP7_75t_L     g12924(.A1(new_n2938), .A2(\b[37] ), .B1(new_n2932), .B2(new_n10229), .C(new_n13180), .Y(new_n13181));
  XNOR2x2_ASAP7_75t_L       g12925(.A(new_n2928), .B(new_n13181), .Y(new_n13182));
  NAND3xp33_ASAP7_75t_L     g12926(.A(new_n13179), .B(new_n13175), .C(new_n13182), .Y(new_n13183));
  NOR3xp33_ASAP7_75t_L      g12927(.A(new_n13176), .B(new_n13177), .C(new_n13178), .Y(new_n13184));
  INVx1_ASAP7_75t_L         g12928(.A(new_n13178), .Y(new_n13185));
  AOI21xp33_ASAP7_75t_L     g12929(.A1(new_n13173), .A2(new_n13169), .B(new_n13185), .Y(new_n13186));
  INVx1_ASAP7_75t_L         g12930(.A(new_n13182), .Y(new_n13187));
  OAI21xp33_ASAP7_75t_L     g12931(.A1(new_n13184), .A2(new_n13186), .B(new_n13187), .Y(new_n13188));
  A2O1A1Ixp33_ASAP7_75t_L   g12932(.A1(new_n12842), .A2(new_n12465), .B(new_n12459), .C(new_n12479), .Y(new_n13189));
  AOI21xp33_ASAP7_75t_L     g12933(.A1(new_n12853), .A2(new_n12855), .B(new_n12856), .Y(new_n13190));
  A2O1A1O1Ixp25_ASAP7_75t_L g12934(.A1(new_n12480), .A2(new_n13189), .B(new_n12485), .C(new_n12857), .D(new_n13190), .Y(new_n13191));
  NAND3xp33_ASAP7_75t_L     g12935(.A(new_n13188), .B(new_n13191), .C(new_n13183), .Y(new_n13192));
  AO21x2_ASAP7_75t_L        g12936(.A1(new_n13183), .A2(new_n13188), .B(new_n13191), .Y(new_n13193));
  OAI22xp33_ASAP7_75t_L     g12937(.A1(new_n2572), .A2(new_n5311), .B1(new_n5570), .B2(new_n2410), .Y(new_n13194));
  AOI221xp5_ASAP7_75t_L     g12938(.A1(new_n2423), .A2(\b[40] ), .B1(new_n2417), .B2(new_n6651), .C(new_n13194), .Y(new_n13195));
  XNOR2x2_ASAP7_75t_L       g12939(.A(new_n2413), .B(new_n13195), .Y(new_n13196));
  NAND3xp33_ASAP7_75t_L     g12940(.A(new_n13193), .B(new_n13192), .C(new_n13196), .Y(new_n13197));
  AND3x1_ASAP7_75t_L        g12941(.A(new_n13188), .B(new_n13191), .C(new_n13183), .Y(new_n13198));
  AOI21xp33_ASAP7_75t_L     g12942(.A1(new_n13188), .A2(new_n13183), .B(new_n13191), .Y(new_n13199));
  INVx1_ASAP7_75t_L         g12943(.A(new_n13196), .Y(new_n13200));
  OAI21xp33_ASAP7_75t_L     g12944(.A1(new_n13199), .A2(new_n13198), .B(new_n13200), .Y(new_n13201));
  AOI21xp33_ASAP7_75t_L     g12945(.A1(new_n13201), .A2(new_n13197), .B(new_n13021), .Y(new_n13202));
  NOR3xp33_ASAP7_75t_L      g12946(.A(new_n13198), .B(new_n13199), .C(new_n13200), .Y(new_n13203));
  AOI21xp33_ASAP7_75t_L     g12947(.A1(new_n13193), .A2(new_n13192), .B(new_n13196), .Y(new_n13204));
  OAI21xp33_ASAP7_75t_L     g12948(.A1(new_n13204), .A2(new_n13203), .B(new_n13021), .Y(new_n13205));
  OAI22xp33_ASAP7_75t_L     g12949(.A1(new_n2089), .A2(new_n6110), .B1(new_n6378), .B2(new_n1962), .Y(new_n13206));
  AOI221xp5_ASAP7_75t_L     g12950(.A1(new_n1955), .A2(\b[43] ), .B1(new_n1964), .B2(new_n6682), .C(new_n13206), .Y(new_n13207));
  XNOR2x2_ASAP7_75t_L       g12951(.A(new_n1952), .B(new_n13207), .Y(new_n13208));
  INVx1_ASAP7_75t_L         g12952(.A(new_n13208), .Y(new_n13209));
  O2A1O1Ixp33_ASAP7_75t_L   g12953(.A1(new_n13021), .A2(new_n13202), .B(new_n13205), .C(new_n13209), .Y(new_n13210));
  OA21x2_ASAP7_75t_L        g12954(.A1(new_n13204), .A2(new_n13203), .B(new_n13021), .Y(new_n13211));
  NOR3xp33_ASAP7_75t_L      g12955(.A(new_n13021), .B(new_n13203), .C(new_n13204), .Y(new_n13212));
  NOR3xp33_ASAP7_75t_L      g12956(.A(new_n13211), .B(new_n13212), .C(new_n13208), .Y(new_n13213));
  NOR2xp33_ASAP7_75t_L      g12957(.A(new_n13210), .B(new_n13213), .Y(new_n13214));
  O2A1O1Ixp33_ASAP7_75t_L   g12958(.A1(new_n12651), .A2(new_n13019), .B(new_n12875), .C(new_n13214), .Y(new_n13215));
  MAJIxp5_ASAP7_75t_L       g12959(.A(new_n12507), .B(new_n12651), .C(new_n13019), .Y(new_n13216));
  OAI21xp33_ASAP7_75t_L     g12960(.A1(new_n13212), .A2(new_n13211), .B(new_n13208), .Y(new_n13217));
  OAI211xp5_ASAP7_75t_L     g12961(.A1(new_n13021), .A2(new_n13202), .B(new_n13205), .C(new_n13209), .Y(new_n13218));
  NAND2xp33_ASAP7_75t_L     g12962(.A(new_n13218), .B(new_n13217), .Y(new_n13219));
  NOR2xp33_ASAP7_75t_L      g12963(.A(new_n13216), .B(new_n13219), .Y(new_n13220));
  OAI21xp33_ASAP7_75t_L     g12964(.A1(new_n13220), .A2(new_n13215), .B(new_n13018), .Y(new_n13221));
  NAND2xp33_ASAP7_75t_L     g12965(.A(new_n12876), .B(new_n12875), .Y(new_n13222));
  NOR2xp33_ASAP7_75t_L      g12966(.A(new_n12647), .B(new_n13222), .Y(new_n13223));
  O2A1O1Ixp33_ASAP7_75t_L   g12967(.A1(new_n12648), .A2(new_n12888), .B(new_n12643), .C(new_n13223), .Y(new_n13224));
  NOR3xp33_ASAP7_75t_L      g12968(.A(new_n13215), .B(new_n13220), .C(new_n13017), .Y(new_n13225));
  NAND2xp33_ASAP7_75t_L     g12969(.A(new_n13216), .B(new_n13219), .Y(new_n13226));
  OR2x4_ASAP7_75t_L         g12970(.A(new_n12651), .B(new_n13019), .Y(new_n13227));
  NAND3xp33_ASAP7_75t_L     g12971(.A(new_n13214), .B(new_n12875), .C(new_n13227), .Y(new_n13228));
  NAND3xp33_ASAP7_75t_L     g12972(.A(new_n13228), .B(new_n13226), .C(new_n13017), .Y(new_n13229));
  O2A1O1Ixp33_ASAP7_75t_L   g12973(.A1(new_n13017), .A2(new_n13225), .B(new_n13229), .C(new_n13224), .Y(new_n13230));
  NOR2xp33_ASAP7_75t_L      g12974(.A(new_n13220), .B(new_n13215), .Y(new_n13231));
  AOI221xp5_ASAP7_75t_L     g12975(.A1(new_n12878), .A2(new_n12643), .B1(new_n13231), .B2(new_n13017), .C(new_n13223), .Y(new_n13232));
  A2O1A1Ixp33_ASAP7_75t_L   g12976(.A1(new_n13232), .A2(new_n13221), .B(new_n13230), .C(new_n13014), .Y(new_n13233));
  INVx1_ASAP7_75t_L         g12977(.A(new_n13221), .Y(new_n13234));
  NAND2xp33_ASAP7_75t_L     g12978(.A(new_n13229), .B(new_n13221), .Y(new_n13235));
  A2O1A1Ixp33_ASAP7_75t_L   g12979(.A1(new_n12878), .A2(new_n12643), .B(new_n13223), .C(new_n13235), .Y(new_n13236));
  NAND2xp33_ASAP7_75t_L     g12980(.A(new_n13229), .B(new_n13224), .Y(new_n13237));
  OAI211xp5_ASAP7_75t_L     g12981(.A1(new_n13234), .A2(new_n13237), .B(new_n13236), .C(new_n13013), .Y(new_n13238));
  NAND2xp33_ASAP7_75t_L     g12982(.A(new_n13233), .B(new_n13238), .Y(new_n13239));
  AOI211xp5_ASAP7_75t_L     g12983(.A1(new_n13221), .A2(new_n13232), .B(new_n13014), .C(new_n13230), .Y(new_n13240));
  NOR2xp33_ASAP7_75t_L      g12984(.A(new_n13010), .B(new_n13240), .Y(new_n13241));
  AOI221xp5_ASAP7_75t_L     g12985(.A1(new_n13239), .A2(new_n13010), .B1(new_n13233), .B2(new_n13241), .C(new_n13009), .Y(new_n13242));
  INVx1_ASAP7_75t_L         g12986(.A(new_n13009), .Y(new_n13243));
  INVx1_ASAP7_75t_L         g12987(.A(new_n13010), .Y(new_n13244));
  INVx1_ASAP7_75t_L         g12988(.A(new_n13225), .Y(new_n13245));
  A2O1A1O1Ixp25_ASAP7_75t_L g12989(.A1(new_n13245), .A2(new_n13018), .B(new_n13237), .C(new_n13236), .D(new_n13013), .Y(new_n13246));
  NOR2xp33_ASAP7_75t_L      g12990(.A(new_n13240), .B(new_n13246), .Y(new_n13247));
  NAND4xp25_ASAP7_75t_L     g12991(.A(new_n13233), .B(new_n13238), .C(new_n12891), .D(new_n12886), .Y(new_n13248));
  O2A1O1Ixp33_ASAP7_75t_L   g12992(.A1(new_n13244), .A2(new_n13247), .B(new_n13248), .C(new_n13243), .Y(new_n13249));
  OR3x1_ASAP7_75t_L         g12993(.A(new_n13006), .B(new_n13242), .C(new_n13249), .Y(new_n13250));
  OAI21xp33_ASAP7_75t_L     g12994(.A1(new_n13242), .A2(new_n13249), .B(new_n13006), .Y(new_n13251));
  NAND3xp33_ASAP7_75t_L     g12995(.A(new_n13250), .B(new_n13005), .C(new_n13251), .Y(new_n13252));
  NOR3xp33_ASAP7_75t_L      g12996(.A(new_n13006), .B(new_n13242), .C(new_n13249), .Y(new_n13253));
  INVx1_ASAP7_75t_L         g12997(.A(new_n13251), .Y(new_n13254));
  OAI21xp33_ASAP7_75t_L     g12998(.A1(new_n13253), .A2(new_n13254), .B(new_n13004), .Y(new_n13255));
  NAND3xp33_ASAP7_75t_L     g12999(.A(new_n13001), .B(new_n13252), .C(new_n13255), .Y(new_n13256));
  NOR2xp33_ASAP7_75t_L      g13000(.A(new_n12907), .B(new_n12902), .Y(new_n13257));
  MAJIxp5_ASAP7_75t_L       g13001(.A(new_n12917), .B(new_n12911), .C(new_n13257), .Y(new_n13258));
  NOR3xp33_ASAP7_75t_L      g13002(.A(new_n13254), .B(new_n13253), .C(new_n13004), .Y(new_n13259));
  AOI21xp33_ASAP7_75t_L     g13003(.A1(new_n13250), .A2(new_n13251), .B(new_n13005), .Y(new_n13260));
  OAI21xp33_ASAP7_75t_L     g13004(.A1(new_n13260), .A2(new_n13259), .B(new_n13258), .Y(new_n13261));
  OAI22xp33_ASAP7_75t_L     g13005(.A1(new_n513), .A2(new_n10978), .B1(new_n10332), .B2(new_n506), .Y(new_n13262));
  AOI221xp5_ASAP7_75t_L     g13006(.A1(new_n475), .A2(\b[58] ), .B1(new_n483), .B2(new_n11314), .C(new_n13262), .Y(new_n13263));
  XNOR2x2_ASAP7_75t_L       g13007(.A(new_n466), .B(new_n13263), .Y(new_n13264));
  NAND3xp33_ASAP7_75t_L     g13008(.A(new_n13256), .B(new_n13261), .C(new_n13264), .Y(new_n13265));
  NOR3xp33_ASAP7_75t_L      g13009(.A(new_n13258), .B(new_n13259), .C(new_n13260), .Y(new_n13266));
  AOI21xp33_ASAP7_75t_L     g13010(.A1(new_n13255), .A2(new_n13252), .B(new_n13001), .Y(new_n13267));
  INVx1_ASAP7_75t_L         g13011(.A(new_n13264), .Y(new_n13268));
  OAI21xp33_ASAP7_75t_L     g13012(.A1(new_n13266), .A2(new_n13267), .B(new_n13268), .Y(new_n13269));
  OAI22xp33_ASAP7_75t_L     g13013(.A1(new_n350), .A2(new_n11626), .B1(new_n11591), .B2(new_n375), .Y(new_n13270));
  AOI221xp5_ASAP7_75t_L     g13014(.A1(new_n361), .A2(\b[61] ), .B1(new_n359), .B2(new_n12269), .C(new_n13270), .Y(new_n13271));
  XNOR2x2_ASAP7_75t_L       g13015(.A(\a[5] ), .B(new_n13271), .Y(new_n13272));
  AOI21xp33_ASAP7_75t_L     g13016(.A1(new_n13269), .A2(new_n13265), .B(new_n13272), .Y(new_n13273));
  NOR3xp33_ASAP7_75t_L      g13017(.A(new_n13267), .B(new_n13266), .C(new_n13268), .Y(new_n13274));
  AOI21xp33_ASAP7_75t_L     g13018(.A1(new_n13256), .A2(new_n13261), .B(new_n13264), .Y(new_n13275));
  XNOR2x2_ASAP7_75t_L       g13019(.A(new_n346), .B(new_n13271), .Y(new_n13276));
  NOR3xp33_ASAP7_75t_L      g13020(.A(new_n13274), .B(new_n13275), .C(new_n13276), .Y(new_n13277));
  OAI21xp33_ASAP7_75t_L     g13021(.A1(new_n13273), .A2(new_n13277), .B(new_n13000), .Y(new_n13278));
  OAI21xp33_ASAP7_75t_L     g13022(.A1(new_n13275), .A2(new_n13274), .B(new_n13276), .Y(new_n13279));
  NAND3xp33_ASAP7_75t_L     g13023(.A(new_n13269), .B(new_n13265), .C(new_n13272), .Y(new_n13280));
  NAND3xp33_ASAP7_75t_L     g13024(.A(new_n13279), .B(new_n13280), .C(new_n12999), .Y(new_n13281));
  NAND3xp33_ASAP7_75t_L     g13025(.A(new_n13278), .B(new_n12996), .C(new_n13281), .Y(new_n13282));
  AOI21xp33_ASAP7_75t_L     g13026(.A1(new_n13279), .A2(new_n13280), .B(new_n12999), .Y(new_n13283));
  NOR3xp33_ASAP7_75t_L      g13027(.A(new_n13277), .B(new_n13273), .C(new_n13000), .Y(new_n13284));
  OAI21xp33_ASAP7_75t_L     g13028(.A1(new_n13283), .A2(new_n13284), .B(new_n12995), .Y(new_n13285));
  NAND3xp33_ASAP7_75t_L     g13029(.A(new_n13285), .B(new_n13282), .C(new_n12984), .Y(new_n13286));
  NOR3xp33_ASAP7_75t_L      g13030(.A(new_n13284), .B(new_n13283), .C(new_n12995), .Y(new_n13287));
  AOI21xp33_ASAP7_75t_L     g13031(.A1(new_n13278), .A2(new_n13281), .B(new_n12996), .Y(new_n13288));
  OAI21xp33_ASAP7_75t_L     g13032(.A1(new_n13288), .A2(new_n13287), .B(new_n12983), .Y(new_n13289));
  NAND2xp33_ASAP7_75t_L     g13033(.A(new_n13286), .B(new_n13289), .Y(new_n13290));
  XOR2x2_ASAP7_75t_L        g13034(.A(new_n13290), .B(new_n12982), .Y(\f[64] ));
  O2A1O1Ixp33_ASAP7_75t_L   g13035(.A1(new_n13231), .A2(new_n13017), .B(new_n13232), .C(new_n13230), .Y(new_n13292));
  NAND2xp33_ASAP7_75t_L     g13036(.A(new_n13014), .B(new_n13292), .Y(new_n13293));
  A2O1A1Ixp33_ASAP7_75t_L   g13037(.A1(new_n13233), .A2(new_n13238), .B(new_n13244), .C(new_n13293), .Y(new_n13294));
  O2A1O1Ixp33_ASAP7_75t_L   g13038(.A1(new_n13223), .A2(new_n12887), .B(new_n13235), .C(new_n13225), .Y(new_n13295));
  OAI22xp33_ASAP7_75t_L     g13039(.A1(new_n1654), .A2(new_n7249), .B1(new_n7270), .B2(new_n1517), .Y(new_n13296));
  AOI221xp5_ASAP7_75t_L     g13040(.A1(new_n1511), .A2(\b[47] ), .B1(new_n1513), .B2(new_n8726), .C(new_n13296), .Y(new_n13297));
  XNOR2x2_ASAP7_75t_L       g13041(.A(new_n1501), .B(new_n13297), .Y(new_n13298));
  NAND2xp33_ASAP7_75t_L     g13042(.A(new_n13192), .B(new_n13193), .Y(new_n13299));
  INVx1_ASAP7_75t_L         g13043(.A(new_n13299), .Y(new_n13300));
  NAND2xp33_ASAP7_75t_L     g13044(.A(new_n13200), .B(new_n13300), .Y(new_n13301));
  A2O1A1Ixp33_ASAP7_75t_L   g13045(.A1(new_n13299), .A2(new_n13201), .B(new_n13021), .C(new_n13301), .Y(new_n13302));
  O2A1O1Ixp33_ASAP7_75t_L   g13046(.A1(new_n13111), .A2(new_n13119), .B(new_n13113), .C(new_n13121), .Y(new_n13303));
  A2O1A1O1Ixp25_ASAP7_75t_L g13047(.A1(new_n12763), .A2(new_n12762), .B(new_n12760), .C(new_n13103), .D(new_n13100), .Y(new_n13304));
  NOR2xp33_ASAP7_75t_L      g13048(.A(new_n13080), .B(new_n13084), .Y(new_n13305));
  AND2x2_ASAP7_75t_L        g13049(.A(new_n13087), .B(new_n13305), .Y(new_n13306));
  INVx1_ASAP7_75t_L         g13050(.A(new_n13095), .Y(new_n13307));
  A2O1A1O1Ixp25_ASAP7_75t_L g13051(.A1(new_n12730), .A2(new_n12666), .B(new_n13078), .C(new_n13081), .D(new_n13077), .Y(new_n13308));
  NAND2xp33_ASAP7_75t_L     g13052(.A(new_n13065), .B(new_n13064), .Y(new_n13309));
  O2A1O1Ixp33_ASAP7_75t_L   g13053(.A1(new_n12715), .A2(new_n12732), .B(new_n12714), .C(new_n12719), .Y(new_n13310));
  O2A1O1Ixp33_ASAP7_75t_L   g13054(.A1(new_n12732), .A2(new_n13310), .B(new_n13309), .C(new_n13068), .Y(new_n13311));
  NOR2xp33_ASAP7_75t_L      g13055(.A(new_n262), .B(new_n13030), .Y(new_n13312));
  O2A1O1Ixp33_ASAP7_75t_L   g13056(.A1(new_n12669), .A2(new_n12671), .B(\b[2] ), .C(new_n13312), .Y(new_n13313));
  INVx1_ASAP7_75t_L         g13057(.A(new_n12320), .Y(new_n13314));
  NOR2xp33_ASAP7_75t_L      g13058(.A(new_n332), .B(new_n12318), .Y(new_n13315));
  AOI221xp5_ASAP7_75t_L     g13059(.A1(new_n11995), .A2(\b[5] ), .B1(new_n13314), .B2(\b[3] ), .C(new_n13315), .Y(new_n13316));
  O2A1O1Ixp33_ASAP7_75t_L   g13060(.A1(new_n728), .A2(new_n11998), .B(new_n13316), .C(new_n11987), .Y(new_n13317));
  O2A1O1Ixp33_ASAP7_75t_L   g13061(.A1(new_n728), .A2(new_n11998), .B(new_n13316), .C(\a[62] ), .Y(new_n13318));
  INVx1_ASAP7_75t_L         g13062(.A(new_n13318), .Y(new_n13319));
  O2A1O1Ixp33_ASAP7_75t_L   g13063(.A1(new_n13317), .A2(new_n11987), .B(new_n13319), .C(new_n13313), .Y(new_n13320));
  INVx1_ASAP7_75t_L         g13064(.A(new_n13320), .Y(new_n13321));
  INVx1_ASAP7_75t_L         g13065(.A(new_n13313), .Y(new_n13322));
  O2A1O1Ixp33_ASAP7_75t_L   g13066(.A1(new_n13317), .A2(new_n11987), .B(new_n13319), .C(new_n13322), .Y(new_n13323));
  A2O1A1O1Ixp25_ASAP7_75t_L g13067(.A1(new_n13028), .A2(\b[2] ), .B(new_n13312), .C(new_n13321), .D(new_n13323), .Y(new_n13324));
  A2O1A1Ixp33_ASAP7_75t_L   g13068(.A1(new_n13028), .A2(\b[1] ), .B(new_n13031), .C(new_n13039), .Y(new_n13325));
  A2O1A1Ixp33_ASAP7_75t_L   g13069(.A1(new_n13325), .A2(new_n13040), .B(new_n13043), .C(new_n13039), .Y(new_n13326));
  INVx1_ASAP7_75t_L         g13070(.A(new_n13326), .Y(new_n13327));
  NAND2xp33_ASAP7_75t_L     g13071(.A(new_n13324), .B(new_n13327), .Y(new_n13328));
  A2O1A1Ixp33_ASAP7_75t_L   g13072(.A1(new_n13321), .A2(new_n13322), .B(new_n13323), .C(new_n13326), .Y(new_n13329));
  NAND2xp33_ASAP7_75t_L     g13073(.A(new_n13329), .B(new_n13328), .Y(new_n13330));
  NOR2xp33_ASAP7_75t_L      g13074(.A(new_n427), .B(new_n11354), .Y(new_n13331));
  AOI221xp5_ASAP7_75t_L     g13075(.A1(\b[8] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[7] ), .C(new_n13331), .Y(new_n13332));
  O2A1O1Ixp33_ASAP7_75t_L   g13076(.A1(new_n11053), .A2(new_n540), .B(new_n13332), .C(new_n11048), .Y(new_n13333));
  INVx1_ASAP7_75t_L         g13077(.A(new_n13333), .Y(new_n13334));
  O2A1O1Ixp33_ASAP7_75t_L   g13078(.A1(new_n11053), .A2(new_n540), .B(new_n13332), .C(\a[59] ), .Y(new_n13335));
  AOI21xp33_ASAP7_75t_L     g13079(.A1(new_n13334), .A2(\a[59] ), .B(new_n13335), .Y(new_n13336));
  A2O1A1Ixp33_ASAP7_75t_L   g13080(.A1(new_n12701), .A2(new_n12700), .B(new_n13053), .C(new_n13054), .Y(new_n13337));
  INVx1_ASAP7_75t_L         g13081(.A(new_n13335), .Y(new_n13338));
  O2A1O1Ixp33_ASAP7_75t_L   g13082(.A1(new_n13333), .A2(new_n11048), .B(new_n13338), .C(new_n13330), .Y(new_n13339));
  NAND2xp33_ASAP7_75t_L     g13083(.A(new_n13336), .B(new_n13330), .Y(new_n13340));
  INVx1_ASAP7_75t_L         g13084(.A(new_n13340), .Y(new_n13341));
  OAI21xp33_ASAP7_75t_L     g13085(.A1(new_n13339), .A2(new_n13341), .B(new_n13337), .Y(new_n13342));
  A2O1A1Ixp33_ASAP7_75t_L   g13086(.A1(new_n13058), .A2(new_n13057), .B(new_n13055), .C(new_n13340), .Y(new_n13343));
  OAI21xp33_ASAP7_75t_L     g13087(.A1(new_n13330), .A2(new_n13336), .B(new_n13343), .Y(new_n13344));
  A2O1A1Ixp33_ASAP7_75t_L   g13088(.A1(new_n13330), .A2(new_n13336), .B(new_n13344), .C(new_n13342), .Y(new_n13345));
  OAI22xp33_ASAP7_75t_L     g13089(.A1(new_n10390), .A2(new_n590), .B1(new_n680), .B2(new_n10388), .Y(new_n13346));
  AOI221xp5_ASAP7_75t_L     g13090(.A1(new_n10086), .A2(\b[11] ), .B1(new_n10386), .B2(new_n976), .C(new_n13346), .Y(new_n13347));
  XNOR2x2_ASAP7_75t_L       g13091(.A(new_n10083), .B(new_n13347), .Y(new_n13348));
  INVx1_ASAP7_75t_L         g13092(.A(new_n13348), .Y(new_n13349));
  NOR2xp33_ASAP7_75t_L      g13093(.A(new_n13349), .B(new_n13345), .Y(new_n13350));
  O2A1O1Ixp33_ASAP7_75t_L   g13094(.A1(new_n13341), .A2(new_n13344), .B(new_n13342), .C(new_n13348), .Y(new_n13351));
  OR2x4_ASAP7_75t_L         g13095(.A(new_n13351), .B(new_n13350), .Y(new_n13352));
  NOR2xp33_ASAP7_75t_L      g13096(.A(new_n13311), .B(new_n13352), .Y(new_n13353));
  NOR2xp33_ASAP7_75t_L      g13097(.A(new_n13351), .B(new_n13350), .Y(new_n13354));
  NOR3xp33_ASAP7_75t_L      g13098(.A(new_n13354), .B(new_n13069), .C(new_n13068), .Y(new_n13355));
  OAI22xp33_ASAP7_75t_L     g13099(.A1(new_n9440), .A2(new_n833), .B1(new_n936), .B2(new_n10400), .Y(new_n13356));
  AOI221xp5_ASAP7_75t_L     g13100(.A1(new_n9102), .A2(\b[14] ), .B1(new_n9437), .B2(new_n971), .C(new_n13356), .Y(new_n13357));
  XNOR2x2_ASAP7_75t_L       g13101(.A(new_n9099), .B(new_n13357), .Y(new_n13358));
  INVx1_ASAP7_75t_L         g13102(.A(new_n13358), .Y(new_n13359));
  NOR3xp33_ASAP7_75t_L      g13103(.A(new_n13353), .B(new_n13355), .C(new_n13359), .Y(new_n13360));
  INVx1_ASAP7_75t_L         g13104(.A(new_n13066), .Y(new_n13361));
  A2O1A1Ixp33_ASAP7_75t_L   g13105(.A1(new_n13309), .A2(new_n13361), .B(new_n13068), .C(new_n13354), .Y(new_n13362));
  NAND2xp33_ASAP7_75t_L     g13106(.A(new_n13311), .B(new_n13352), .Y(new_n13363));
  AOI21xp33_ASAP7_75t_L     g13107(.A1(new_n13363), .A2(new_n13362), .B(new_n13358), .Y(new_n13364));
  NOR3xp33_ASAP7_75t_L      g13108(.A(new_n13360), .B(new_n13364), .C(new_n13308), .Y(new_n13365));
  INVx1_ASAP7_75t_L         g13109(.A(new_n13308), .Y(new_n13366));
  NAND3xp33_ASAP7_75t_L     g13110(.A(new_n13363), .B(new_n13362), .C(new_n13358), .Y(new_n13367));
  OAI21xp33_ASAP7_75t_L     g13111(.A1(new_n13355), .A2(new_n13353), .B(new_n13359), .Y(new_n13368));
  AOI21xp33_ASAP7_75t_L     g13112(.A1(new_n13368), .A2(new_n13367), .B(new_n13366), .Y(new_n13369));
  OAI22xp33_ASAP7_75t_L     g13113(.A1(new_n8483), .A2(new_n1043), .B1(new_n1150), .B2(new_n10065), .Y(new_n13370));
  AOI221xp5_ASAP7_75t_L     g13114(.A1(new_n8175), .A2(\b[17] ), .B1(new_n8490), .B2(new_n1633), .C(new_n13370), .Y(new_n13371));
  XNOR2x2_ASAP7_75t_L       g13115(.A(new_n8172), .B(new_n13371), .Y(new_n13372));
  INVx1_ASAP7_75t_L         g13116(.A(new_n13372), .Y(new_n13373));
  OAI21xp33_ASAP7_75t_L     g13117(.A1(new_n13369), .A2(new_n13365), .B(new_n13373), .Y(new_n13374));
  NAND3xp33_ASAP7_75t_L     g13118(.A(new_n13368), .B(new_n13367), .C(new_n13366), .Y(new_n13375));
  OAI21xp33_ASAP7_75t_L     g13119(.A1(new_n13364), .A2(new_n13360), .B(new_n13308), .Y(new_n13376));
  NAND3xp33_ASAP7_75t_L     g13120(.A(new_n13376), .B(new_n13375), .C(new_n13372), .Y(new_n13377));
  AOI211xp5_ASAP7_75t_L     g13121(.A1(new_n13374), .A2(new_n13377), .B(new_n13307), .C(new_n13306), .Y(new_n13378));
  OAI211xp5_ASAP7_75t_L     g13122(.A1(new_n13307), .A2(new_n13306), .B(new_n13374), .C(new_n13377), .Y(new_n13379));
  INVx1_ASAP7_75t_L         g13123(.A(new_n13379), .Y(new_n13380));
  NOR2xp33_ASAP7_75t_L      g13124(.A(new_n1745), .B(new_n7318), .Y(new_n13381));
  AOI221xp5_ASAP7_75t_L     g13125(.A1(new_n7333), .A2(\b[19] ), .B1(new_n7609), .B2(\b[18] ), .C(new_n13381), .Y(new_n13382));
  O2A1O1Ixp33_ASAP7_75t_L   g13126(.A1(new_n7321), .A2(new_n1754), .B(new_n13382), .C(new_n7316), .Y(new_n13383));
  OAI21xp33_ASAP7_75t_L     g13127(.A1(new_n7321), .A2(new_n1754), .B(new_n13382), .Y(new_n13384));
  NAND2xp33_ASAP7_75t_L     g13128(.A(new_n7316), .B(new_n13384), .Y(new_n13385));
  OA21x2_ASAP7_75t_L        g13129(.A1(new_n7316), .A2(new_n13383), .B(new_n13385), .Y(new_n13386));
  INVx1_ASAP7_75t_L         g13130(.A(new_n13386), .Y(new_n13387));
  NOR3xp33_ASAP7_75t_L      g13131(.A(new_n13380), .B(new_n13387), .C(new_n13378), .Y(new_n13388));
  O2A1O1Ixp33_ASAP7_75t_L   g13132(.A1(new_n13091), .A2(new_n13087), .B(new_n13094), .C(new_n13306), .Y(new_n13389));
  NAND2xp33_ASAP7_75t_L     g13133(.A(new_n13377), .B(new_n13374), .Y(new_n13390));
  NAND2xp33_ASAP7_75t_L     g13134(.A(new_n13389), .B(new_n13390), .Y(new_n13391));
  AOI21xp33_ASAP7_75t_L     g13135(.A1(new_n13391), .A2(new_n13379), .B(new_n13386), .Y(new_n13392));
  NOR3xp33_ASAP7_75t_L      g13136(.A(new_n13388), .B(new_n13392), .C(new_n13304), .Y(new_n13393));
  INVx1_ASAP7_75t_L         g13137(.A(new_n13304), .Y(new_n13394));
  NAND3xp33_ASAP7_75t_L     g13138(.A(new_n13391), .B(new_n13379), .C(new_n13386), .Y(new_n13395));
  OAI21xp33_ASAP7_75t_L     g13139(.A1(new_n13378), .A2(new_n13380), .B(new_n13387), .Y(new_n13396));
  AOI21xp33_ASAP7_75t_L     g13140(.A1(new_n13396), .A2(new_n13395), .B(new_n13394), .Y(new_n13397));
  OAI22xp33_ASAP7_75t_L     g13141(.A1(new_n7304), .A2(new_n2045), .B1(new_n1895), .B2(new_n6741), .Y(new_n13398));
  AOI221xp5_ASAP7_75t_L     g13142(.A1(new_n6442), .A2(\b[23] ), .B1(new_n6450), .B2(new_n2679), .C(new_n13398), .Y(new_n13399));
  XNOR2x2_ASAP7_75t_L       g13143(.A(new_n6439), .B(new_n13399), .Y(new_n13400));
  INVx1_ASAP7_75t_L         g13144(.A(new_n13400), .Y(new_n13401));
  OAI21xp33_ASAP7_75t_L     g13145(.A1(new_n13397), .A2(new_n13393), .B(new_n13401), .Y(new_n13402));
  NAND3xp33_ASAP7_75t_L     g13146(.A(new_n13396), .B(new_n13395), .C(new_n13394), .Y(new_n13403));
  NAND3xp33_ASAP7_75t_L     g13147(.A(new_n13379), .B(new_n13391), .C(new_n13387), .Y(new_n13404));
  A2O1A1Ixp33_ASAP7_75t_L   g13148(.A1(new_n13404), .A2(new_n13387), .B(new_n13388), .C(new_n13304), .Y(new_n13405));
  NAND3xp33_ASAP7_75t_L     g13149(.A(new_n13405), .B(new_n13403), .C(new_n13400), .Y(new_n13406));
  NAND2xp33_ASAP7_75t_L     g13150(.A(new_n13402), .B(new_n13406), .Y(new_n13407));
  NAND2xp33_ASAP7_75t_L     g13151(.A(new_n13303), .B(new_n13407), .Y(new_n13408));
  AOI21xp33_ASAP7_75t_L     g13152(.A1(new_n13405), .A2(new_n13403), .B(new_n13400), .Y(new_n13409));
  NOR3xp33_ASAP7_75t_L      g13153(.A(new_n13393), .B(new_n13397), .C(new_n13401), .Y(new_n13410));
  NOR2xp33_ASAP7_75t_L      g13154(.A(new_n13410), .B(new_n13409), .Y(new_n13411));
  A2O1A1Ixp33_ASAP7_75t_L   g13155(.A1(new_n13109), .A2(new_n13119), .B(new_n13116), .C(new_n13411), .Y(new_n13412));
  OAI22xp33_ASAP7_75t_L     g13156(.A1(new_n5640), .A2(new_n2377), .B1(new_n2205), .B2(new_n5925), .Y(new_n13413));
  AOI221xp5_ASAP7_75t_L     g13157(.A1(new_n5629), .A2(\b[26] ), .B1(new_n5637), .B2(new_n2709), .C(new_n13413), .Y(new_n13414));
  XNOR2x2_ASAP7_75t_L       g13158(.A(new_n5626), .B(new_n13414), .Y(new_n13415));
  NAND3xp33_ASAP7_75t_L     g13159(.A(new_n13412), .B(new_n13408), .C(new_n13415), .Y(new_n13416));
  INVx1_ASAP7_75t_L         g13160(.A(new_n13303), .Y(new_n13417));
  NOR2xp33_ASAP7_75t_L      g13161(.A(new_n13417), .B(new_n13411), .Y(new_n13418));
  O2A1O1Ixp33_ASAP7_75t_L   g13162(.A1(new_n13115), .A2(new_n13112), .B(new_n13122), .C(new_n13407), .Y(new_n13419));
  INVx1_ASAP7_75t_L         g13163(.A(new_n13415), .Y(new_n13420));
  OAI21xp33_ASAP7_75t_L     g13164(.A1(new_n13418), .A2(new_n13419), .B(new_n13420), .Y(new_n13421));
  NAND4xp25_ASAP7_75t_L     g13165(.A(new_n13416), .B(new_n13421), .C(new_n13128), .D(new_n13135), .Y(new_n13422));
  AOI22xp33_ASAP7_75t_L     g13166(.A1(new_n13135), .A2(new_n13128), .B1(new_n13421), .B2(new_n13416), .Y(new_n13423));
  INVx1_ASAP7_75t_L         g13167(.A(new_n13423), .Y(new_n13424));
  OAI22xp33_ASAP7_75t_L     g13168(.A1(new_n5144), .A2(new_n2879), .B1(new_n3079), .B2(new_n4903), .Y(new_n13425));
  AOI221xp5_ASAP7_75t_L     g13169(.A1(new_n4917), .A2(\b[29] ), .B1(new_n4912), .B2(new_n3873), .C(new_n13425), .Y(new_n13426));
  XNOR2x2_ASAP7_75t_L       g13170(.A(new_n4906), .B(new_n13426), .Y(new_n13427));
  NAND3xp33_ASAP7_75t_L     g13171(.A(new_n13424), .B(new_n13422), .C(new_n13427), .Y(new_n13428));
  INVx1_ASAP7_75t_L         g13172(.A(new_n13422), .Y(new_n13429));
  INVx1_ASAP7_75t_L         g13173(.A(new_n13427), .Y(new_n13430));
  OAI21xp33_ASAP7_75t_L     g13174(.A1(new_n13423), .A2(new_n13429), .B(new_n13430), .Y(new_n13431));
  INVx1_ASAP7_75t_L         g13175(.A(new_n13139), .Y(new_n13432));
  O2A1O1Ixp33_ASAP7_75t_L   g13176(.A1(new_n13144), .A2(new_n13138), .B(new_n13147), .C(new_n13432), .Y(new_n13433));
  NAND3xp33_ASAP7_75t_L     g13177(.A(new_n13428), .B(new_n13431), .C(new_n13433), .Y(new_n13434));
  INVx1_ASAP7_75t_L         g13178(.A(new_n13434), .Y(new_n13435));
  AOI21xp33_ASAP7_75t_L     g13179(.A1(new_n13428), .A2(new_n13431), .B(new_n13433), .Y(new_n13436));
  OAI22xp33_ASAP7_75t_L     g13180(.A1(new_n4397), .A2(new_n3456), .B1(new_n3674), .B2(new_n4142), .Y(new_n13437));
  AOI221xp5_ASAP7_75t_L     g13181(.A1(new_n4156), .A2(\b[32] ), .B1(new_n4151), .B2(new_n3900), .C(new_n13437), .Y(new_n13438));
  XNOR2x2_ASAP7_75t_L       g13182(.A(new_n4145), .B(new_n13438), .Y(new_n13439));
  OAI21xp33_ASAP7_75t_L     g13183(.A1(new_n13436), .A2(new_n13435), .B(new_n13439), .Y(new_n13440));
  A2O1A1O1Ixp25_ASAP7_75t_L g13184(.A1(new_n12817), .A2(new_n12827), .B(new_n12825), .C(new_n13162), .D(new_n13157), .Y(new_n13441));
  INVx1_ASAP7_75t_L         g13185(.A(new_n13436), .Y(new_n13442));
  INVx1_ASAP7_75t_L         g13186(.A(new_n13439), .Y(new_n13443));
  NAND3xp33_ASAP7_75t_L     g13187(.A(new_n13442), .B(new_n13434), .C(new_n13443), .Y(new_n13444));
  AOI21xp33_ASAP7_75t_L     g13188(.A1(new_n13440), .A2(new_n13444), .B(new_n13441), .Y(new_n13445));
  NOR3xp33_ASAP7_75t_L      g13189(.A(new_n13435), .B(new_n13436), .C(new_n13439), .Y(new_n13446));
  A2O1A1O1Ixp25_ASAP7_75t_L g13190(.A1(new_n13158), .A2(new_n13160), .B(new_n13157), .C(new_n13440), .D(new_n13446), .Y(new_n13447));
  OAI22xp33_ASAP7_75t_L     g13191(.A1(new_n3703), .A2(new_n4101), .B1(new_n4344), .B2(new_n3509), .Y(new_n13448));
  AOI221xp5_ASAP7_75t_L     g13192(.A1(new_n3503), .A2(\b[35] ), .B1(new_n3505), .B2(new_n7773), .C(new_n13448), .Y(new_n13449));
  XNOR2x2_ASAP7_75t_L       g13193(.A(new_n3493), .B(new_n13449), .Y(new_n13450));
  A2O1A1Ixp33_ASAP7_75t_L   g13194(.A1(new_n13447), .A2(new_n13440), .B(new_n13445), .C(new_n13450), .Y(new_n13451));
  A2O1A1O1Ixp25_ASAP7_75t_L g13195(.A1(new_n13442), .A2(new_n13434), .B(new_n13443), .C(new_n13447), .D(new_n13445), .Y(new_n13452));
  INVx1_ASAP7_75t_L         g13196(.A(new_n13450), .Y(new_n13453));
  NAND2xp33_ASAP7_75t_L     g13197(.A(new_n13453), .B(new_n13452), .Y(new_n13454));
  NOR3xp33_ASAP7_75t_L      g13198(.A(new_n13171), .B(new_n13170), .C(new_n13168), .Y(new_n13455));
  O2A1O1Ixp33_ASAP7_75t_L   g13199(.A1(new_n13172), .A2(new_n13176), .B(new_n13178), .C(new_n13455), .Y(new_n13456));
  NAND3xp33_ASAP7_75t_L     g13200(.A(new_n13454), .B(new_n13451), .C(new_n13456), .Y(new_n13457));
  A2O1A1Ixp33_ASAP7_75t_L   g13201(.A1(new_n13447), .A2(new_n13440), .B(new_n13445), .C(new_n13453), .Y(new_n13458));
  INVx1_ASAP7_75t_L         g13202(.A(new_n13451), .Y(new_n13459));
  INVx1_ASAP7_75t_L         g13203(.A(new_n13456), .Y(new_n13460));
  A2O1A1Ixp33_ASAP7_75t_L   g13204(.A1(new_n13458), .A2(new_n13453), .B(new_n13459), .C(new_n13460), .Y(new_n13461));
  OAI22xp33_ASAP7_75t_L     g13205(.A1(new_n3133), .A2(new_n4613), .B1(new_n5074), .B2(new_n2925), .Y(new_n13462));
  AOI221xp5_ASAP7_75t_L     g13206(.A1(new_n2938), .A2(\b[38] ), .B1(new_n2932), .B2(new_n6083), .C(new_n13462), .Y(new_n13463));
  XNOR2x2_ASAP7_75t_L       g13207(.A(new_n2928), .B(new_n13463), .Y(new_n13464));
  NAND3xp33_ASAP7_75t_L     g13208(.A(new_n13457), .B(new_n13461), .C(new_n13464), .Y(new_n13465));
  AOI211xp5_ASAP7_75t_L     g13209(.A1(new_n13453), .A2(new_n13458), .B(new_n13459), .C(new_n13460), .Y(new_n13466));
  INVx1_ASAP7_75t_L         g13210(.A(new_n13458), .Y(new_n13467));
  O2A1O1Ixp33_ASAP7_75t_L   g13211(.A1(new_n13450), .A2(new_n13467), .B(new_n13451), .C(new_n13456), .Y(new_n13468));
  INVx1_ASAP7_75t_L         g13212(.A(new_n13464), .Y(new_n13469));
  OAI21xp33_ASAP7_75t_L     g13213(.A1(new_n13466), .A2(new_n13468), .B(new_n13469), .Y(new_n13470));
  NAND3xp33_ASAP7_75t_L     g13214(.A(new_n13179), .B(new_n13175), .C(new_n13187), .Y(new_n13471));
  A2O1A1Ixp33_ASAP7_75t_L   g13215(.A1(new_n13183), .A2(new_n13182), .B(new_n13191), .C(new_n13471), .Y(new_n13472));
  INVx1_ASAP7_75t_L         g13216(.A(new_n13472), .Y(new_n13473));
  NAND3xp33_ASAP7_75t_L     g13217(.A(new_n13470), .B(new_n13465), .C(new_n13473), .Y(new_n13474));
  INVx1_ASAP7_75t_L         g13218(.A(new_n13465), .Y(new_n13475));
  AOI21xp33_ASAP7_75t_L     g13219(.A1(new_n13457), .A2(new_n13461), .B(new_n13464), .Y(new_n13476));
  OAI21xp33_ASAP7_75t_L     g13220(.A1(new_n13476), .A2(new_n13475), .B(new_n13472), .Y(new_n13477));
  NOR2xp33_ASAP7_75t_L      g13221(.A(new_n6110), .B(new_n2415), .Y(new_n13478));
  AOI221xp5_ASAP7_75t_L     g13222(.A1(\b[39] ), .A2(new_n2577), .B1(\b[40] ), .B2(new_n2421), .C(new_n13478), .Y(new_n13479));
  O2A1O1Ixp33_ASAP7_75t_L   g13223(.A1(new_n2425), .A2(new_n6117), .B(new_n13479), .C(new_n2413), .Y(new_n13480));
  OAI21xp33_ASAP7_75t_L     g13224(.A1(new_n2425), .A2(new_n6117), .B(new_n13479), .Y(new_n13481));
  NAND2xp33_ASAP7_75t_L     g13225(.A(new_n2413), .B(new_n13481), .Y(new_n13482));
  OA21x2_ASAP7_75t_L        g13226(.A1(new_n2413), .A2(new_n13480), .B(new_n13482), .Y(new_n13483));
  INVx1_ASAP7_75t_L         g13227(.A(new_n13483), .Y(new_n13484));
  NAND3xp33_ASAP7_75t_L     g13228(.A(new_n13477), .B(new_n13474), .C(new_n13484), .Y(new_n13485));
  NOR3xp33_ASAP7_75t_L      g13229(.A(new_n13475), .B(new_n13476), .C(new_n13472), .Y(new_n13486));
  NOR3xp33_ASAP7_75t_L      g13230(.A(new_n13468), .B(new_n13466), .C(new_n13464), .Y(new_n13487));
  O2A1O1Ixp33_ASAP7_75t_L   g13231(.A1(new_n13464), .A2(new_n13487), .B(new_n13465), .C(new_n13473), .Y(new_n13488));
  OAI21xp33_ASAP7_75t_L     g13232(.A1(new_n13488), .A2(new_n13486), .B(new_n13483), .Y(new_n13489));
  NAND3xp33_ASAP7_75t_L     g13233(.A(new_n13302), .B(new_n13489), .C(new_n13485), .Y(new_n13490));
  NOR3xp33_ASAP7_75t_L      g13234(.A(new_n13486), .B(new_n13488), .C(new_n13483), .Y(new_n13491));
  AOI21xp33_ASAP7_75t_L     g13235(.A1(new_n13477), .A2(new_n13474), .B(new_n13484), .Y(new_n13492));
  NOR3xp33_ASAP7_75t_L      g13236(.A(new_n13491), .B(new_n13302), .C(new_n13492), .Y(new_n13493));
  NOR2xp33_ASAP7_75t_L      g13237(.A(new_n6671), .B(new_n1962), .Y(new_n13494));
  AOI221xp5_ASAP7_75t_L     g13238(.A1(new_n1955), .A2(\b[44] ), .B1(new_n2093), .B2(\b[42] ), .C(new_n13494), .Y(new_n13495));
  O2A1O1Ixp33_ASAP7_75t_L   g13239(.A1(new_n1956), .A2(new_n6951), .B(new_n13495), .C(new_n1952), .Y(new_n13496));
  OAI21xp33_ASAP7_75t_L     g13240(.A1(new_n1956), .A2(new_n6951), .B(new_n13495), .Y(new_n13497));
  NAND2xp33_ASAP7_75t_L     g13241(.A(new_n1952), .B(new_n13497), .Y(new_n13498));
  OA21x2_ASAP7_75t_L        g13242(.A1(new_n1952), .A2(new_n13496), .B(new_n13498), .Y(new_n13499));
  A2O1A1Ixp33_ASAP7_75t_L   g13243(.A1(new_n13490), .A2(new_n13302), .B(new_n13493), .C(new_n13499), .Y(new_n13500));
  A2O1A1O1Ixp25_ASAP7_75t_L g13244(.A1(new_n13197), .A2(new_n13196), .B(new_n13021), .C(new_n13301), .D(new_n13492), .Y(new_n13501));
  OAI21xp33_ASAP7_75t_L     g13245(.A1(new_n13492), .A2(new_n13491), .B(new_n13302), .Y(new_n13502));
  INVx1_ASAP7_75t_L         g13246(.A(new_n13499), .Y(new_n13503));
  OAI311xp33_ASAP7_75t_L    g13247(.A1(new_n13501), .A2(new_n13492), .A3(new_n13491), .B1(new_n13503), .C1(new_n13502), .Y(new_n13504));
  OAI21xp33_ASAP7_75t_L     g13248(.A1(new_n13212), .A2(new_n13211), .B(new_n13209), .Y(new_n13505));
  A2O1A1Ixp33_ASAP7_75t_L   g13249(.A1(new_n12875), .A2(new_n13227), .B(new_n13214), .C(new_n13505), .Y(new_n13506));
  INVx1_ASAP7_75t_L         g13250(.A(new_n13506), .Y(new_n13507));
  AOI21xp33_ASAP7_75t_L     g13251(.A1(new_n13504), .A2(new_n13500), .B(new_n13507), .Y(new_n13508));
  AND3x1_ASAP7_75t_L        g13252(.A(new_n13507), .B(new_n13504), .C(new_n13500), .Y(new_n13509));
  NOR3xp33_ASAP7_75t_L      g13253(.A(new_n13509), .B(new_n13508), .C(new_n13298), .Y(new_n13510));
  A2O1A1Ixp33_ASAP7_75t_L   g13254(.A1(new_n13490), .A2(new_n13302), .B(new_n13493), .C(new_n13503), .Y(new_n13511));
  INVx1_ASAP7_75t_L         g13255(.A(new_n13500), .Y(new_n13512));
  A2O1A1Ixp33_ASAP7_75t_L   g13256(.A1(new_n13511), .A2(new_n13503), .B(new_n13512), .C(new_n13506), .Y(new_n13513));
  NAND3xp33_ASAP7_75t_L     g13257(.A(new_n13507), .B(new_n13504), .C(new_n13500), .Y(new_n13514));
  NAND3xp33_ASAP7_75t_L     g13258(.A(new_n13513), .B(new_n13298), .C(new_n13514), .Y(new_n13515));
  O2A1O1Ixp33_ASAP7_75t_L   g13259(.A1(new_n13298), .A2(new_n13510), .B(new_n13515), .C(new_n13295), .Y(new_n13516));
  OAI21xp33_ASAP7_75t_L     g13260(.A1(new_n13298), .A2(new_n13510), .B(new_n13515), .Y(new_n13517));
  NAND2xp33_ASAP7_75t_L     g13261(.A(new_n13295), .B(new_n13517), .Y(new_n13518));
  OAI22xp33_ASAP7_75t_L     g13262(.A1(new_n1285), .A2(new_n7860), .B1(new_n8427), .B2(new_n2118), .Y(new_n13519));
  AOI221xp5_ASAP7_75t_L     g13263(.A1(new_n1209), .A2(\b[50] ), .B1(new_n1216), .B2(new_n8763), .C(new_n13519), .Y(new_n13520));
  XNOR2x2_ASAP7_75t_L       g13264(.A(new_n1206), .B(new_n13520), .Y(new_n13521));
  OAI211xp5_ASAP7_75t_L     g13265(.A1(new_n13516), .A2(new_n13295), .B(new_n13518), .C(new_n13521), .Y(new_n13522));
  NOR2xp33_ASAP7_75t_L      g13266(.A(new_n13295), .B(new_n13517), .Y(new_n13523));
  INVx1_ASAP7_75t_L         g13267(.A(new_n13295), .Y(new_n13524));
  O2A1O1Ixp33_ASAP7_75t_L   g13268(.A1(new_n13298), .A2(new_n13510), .B(new_n13515), .C(new_n13524), .Y(new_n13525));
  INVx1_ASAP7_75t_L         g13269(.A(new_n13521), .Y(new_n13526));
  OAI21xp33_ASAP7_75t_L     g13270(.A1(new_n13525), .A2(new_n13523), .B(new_n13526), .Y(new_n13527));
  NAND3xp33_ASAP7_75t_L     g13271(.A(new_n13522), .B(new_n13527), .C(new_n13294), .Y(new_n13528));
  AO21x2_ASAP7_75t_L        g13272(.A1(new_n13527), .A2(new_n13522), .B(new_n13294), .Y(new_n13529));
  OAI22xp33_ASAP7_75t_L     g13273(.A1(new_n980), .A2(new_n8779), .B1(new_n9355), .B2(new_n864), .Y(new_n13530));
  AOI221xp5_ASAP7_75t_L     g13274(.A1(new_n886), .A2(\b[53] ), .B1(new_n873), .B2(new_n9690), .C(new_n13530), .Y(new_n13531));
  XNOR2x2_ASAP7_75t_L       g13275(.A(new_n867), .B(new_n13531), .Y(new_n13532));
  NAND3xp33_ASAP7_75t_L     g13276(.A(new_n13529), .B(new_n13528), .C(new_n13532), .Y(new_n13533));
  AO21x2_ASAP7_75t_L        g13277(.A1(new_n13528), .A2(new_n13529), .B(new_n13532), .Y(new_n13534));
  INVx1_ASAP7_75t_L         g13278(.A(new_n13249), .Y(new_n13535));
  A2O1A1O1Ixp25_ASAP7_75t_L g13279(.A1(new_n12903), .A2(new_n12906), .B(new_n12904), .C(new_n13535), .D(new_n13242), .Y(new_n13536));
  AND3x1_ASAP7_75t_L        g13280(.A(new_n13534), .B(new_n13536), .C(new_n13533), .Y(new_n13537));
  AOI21xp33_ASAP7_75t_L     g13281(.A1(new_n13534), .A2(new_n13533), .B(new_n13536), .Y(new_n13538));
  OAI22xp33_ASAP7_75t_L     g13282(.A1(new_n1550), .A2(new_n10309), .B1(new_n9709), .B2(new_n712), .Y(new_n13539));
  AOI221xp5_ASAP7_75t_L     g13283(.A1(new_n640), .A2(\b[56] ), .B1(new_n718), .B2(new_n11579), .C(new_n13539), .Y(new_n13540));
  XNOR2x2_ASAP7_75t_L       g13284(.A(new_n637), .B(new_n13540), .Y(new_n13541));
  OAI21xp33_ASAP7_75t_L     g13285(.A1(new_n13538), .A2(new_n13537), .B(new_n13541), .Y(new_n13542));
  NAND3xp33_ASAP7_75t_L     g13286(.A(new_n13534), .B(new_n13536), .C(new_n13533), .Y(new_n13543));
  AO21x2_ASAP7_75t_L        g13287(.A1(new_n13533), .A2(new_n13534), .B(new_n13536), .Y(new_n13544));
  INVx1_ASAP7_75t_L         g13288(.A(new_n13541), .Y(new_n13545));
  NAND3xp33_ASAP7_75t_L     g13289(.A(new_n13544), .B(new_n13543), .C(new_n13545), .Y(new_n13546));
  OAI22xp33_ASAP7_75t_L     g13290(.A1(new_n513), .A2(new_n11303), .B1(new_n10978), .B2(new_n506), .Y(new_n13547));
  AOI221xp5_ASAP7_75t_L     g13291(.A1(new_n475), .A2(\b[59] ), .B1(new_n483), .B2(new_n12577), .C(new_n13547), .Y(new_n13548));
  XNOR2x2_ASAP7_75t_L       g13292(.A(new_n466), .B(new_n13548), .Y(new_n13549));
  NAND3xp33_ASAP7_75t_L     g13293(.A(new_n13542), .B(new_n13546), .C(new_n13549), .Y(new_n13550));
  AOI21xp33_ASAP7_75t_L     g13294(.A1(new_n13544), .A2(new_n13543), .B(new_n13545), .Y(new_n13551));
  NOR3xp33_ASAP7_75t_L      g13295(.A(new_n13537), .B(new_n13538), .C(new_n13541), .Y(new_n13552));
  INVx1_ASAP7_75t_L         g13296(.A(new_n13549), .Y(new_n13553));
  OAI21xp33_ASAP7_75t_L     g13297(.A1(new_n13551), .A2(new_n13552), .B(new_n13553), .Y(new_n13554));
  A2O1A1O1Ixp25_ASAP7_75t_L g13298(.A1(new_n12911), .A2(new_n13257), .B(new_n12924), .C(new_n13255), .D(new_n13259), .Y(new_n13555));
  NAND3xp33_ASAP7_75t_L     g13299(.A(new_n13554), .B(new_n13550), .C(new_n13555), .Y(new_n13556));
  AOI21xp33_ASAP7_75t_L     g13300(.A1(new_n13554), .A2(new_n13550), .B(new_n13555), .Y(new_n13557));
  INVx1_ASAP7_75t_L         g13301(.A(new_n13557), .Y(new_n13558));
  INVx1_ASAP7_75t_L         g13302(.A(new_n12610), .Y(new_n13559));
  OAI22xp33_ASAP7_75t_L     g13303(.A1(new_n350), .A2(new_n12258), .B1(new_n11626), .B2(new_n375), .Y(new_n13560));
  AOI221xp5_ASAP7_75t_L     g13304(.A1(new_n361), .A2(\b[62] ), .B1(new_n359), .B2(new_n13559), .C(new_n13560), .Y(new_n13561));
  XNOR2x2_ASAP7_75t_L       g13305(.A(new_n346), .B(new_n13561), .Y(new_n13562));
  NAND3xp33_ASAP7_75t_L     g13306(.A(new_n13558), .B(new_n13556), .C(new_n13562), .Y(new_n13563));
  INVx1_ASAP7_75t_L         g13307(.A(new_n13556), .Y(new_n13564));
  INVx1_ASAP7_75t_L         g13308(.A(new_n13562), .Y(new_n13565));
  OAI21xp33_ASAP7_75t_L     g13309(.A1(new_n13557), .A2(new_n13564), .B(new_n13565), .Y(new_n13566));
  NAND3xp33_ASAP7_75t_L     g13310(.A(new_n13256), .B(new_n13261), .C(new_n13268), .Y(new_n13567));
  NOR2xp33_ASAP7_75t_L      g13311(.A(new_n12956), .B(new_n287), .Y(new_n13568));
  A2O1A1Ixp33_ASAP7_75t_L   g13312(.A1(new_n12986), .A2(new_n273), .B(new_n13568), .C(\a[2] ), .Y(new_n13569));
  A2O1A1Ixp33_ASAP7_75t_L   g13313(.A1(new_n273), .A2(new_n12986), .B(\a[2] ), .C(new_n13569), .Y(new_n13570));
  A2O1A1O1Ixp25_ASAP7_75t_L g13314(.A1(new_n13264), .A2(new_n13265), .B(new_n13276), .C(new_n13567), .D(new_n13570), .Y(new_n13571));
  A2O1A1Ixp33_ASAP7_75t_L   g13315(.A1(new_n13265), .A2(new_n13264), .B(new_n13276), .C(new_n13567), .Y(new_n13572));
  INVx1_ASAP7_75t_L         g13316(.A(new_n12986), .Y(new_n13573));
  NOR2xp33_ASAP7_75t_L      g13317(.A(new_n279), .B(new_n13573), .Y(new_n13574));
  O2A1O1Ixp33_ASAP7_75t_L   g13318(.A1(new_n13574), .A2(\a[2] ), .B(new_n13569), .C(new_n13572), .Y(new_n13575));
  NOR2xp33_ASAP7_75t_L      g13319(.A(new_n13571), .B(new_n13575), .Y(new_n13576));
  AOI21xp33_ASAP7_75t_L     g13320(.A1(new_n13563), .A2(new_n13566), .B(new_n13576), .Y(new_n13577));
  NOR3xp33_ASAP7_75t_L      g13321(.A(new_n13564), .B(new_n13557), .C(new_n13565), .Y(new_n13578));
  AOI21xp33_ASAP7_75t_L     g13322(.A1(new_n13558), .A2(new_n13556), .B(new_n13562), .Y(new_n13579));
  XOR2x2_ASAP7_75t_L        g13323(.A(new_n13570), .B(new_n13572), .Y(new_n13580));
  NOR3xp33_ASAP7_75t_L      g13324(.A(new_n13579), .B(new_n13578), .C(new_n13580), .Y(new_n13581));
  O2A1O1Ixp33_ASAP7_75t_L   g13325(.A1(new_n12994), .A2(new_n12992), .B(new_n13281), .C(new_n13283), .Y(new_n13582));
  INVx1_ASAP7_75t_L         g13326(.A(new_n13582), .Y(new_n13583));
  NOR3xp33_ASAP7_75t_L      g13327(.A(new_n13581), .B(new_n13577), .C(new_n13583), .Y(new_n13584));
  OAI21xp33_ASAP7_75t_L     g13328(.A1(new_n13578), .A2(new_n13579), .B(new_n13580), .Y(new_n13585));
  NAND3xp33_ASAP7_75t_L     g13329(.A(new_n13576), .B(new_n13563), .C(new_n13566), .Y(new_n13586));
  AOI21xp33_ASAP7_75t_L     g13330(.A1(new_n13585), .A2(new_n13586), .B(new_n13582), .Y(new_n13587));
  NOR2xp33_ASAP7_75t_L      g13331(.A(new_n13587), .B(new_n13584), .Y(new_n13588));
  INVx1_ASAP7_75t_L         g13332(.A(new_n13588), .Y(new_n13589));
  O2A1O1Ixp33_ASAP7_75t_L   g13333(.A1(new_n12982), .A2(new_n13290), .B(new_n13286), .C(new_n13589), .Y(new_n13590));
  OAI21xp33_ASAP7_75t_L     g13334(.A1(new_n13290), .A2(new_n12982), .B(new_n13286), .Y(new_n13591));
  NOR2xp33_ASAP7_75t_L      g13335(.A(new_n13588), .B(new_n13591), .Y(new_n13592));
  NOR2xp33_ASAP7_75t_L      g13336(.A(new_n13592), .B(new_n13590), .Y(\f[65] ));
  OAI22xp33_ASAP7_75t_L     g13337(.A1(new_n350), .A2(new_n12603), .B1(new_n12258), .B2(new_n375), .Y(new_n13594));
  AOI221xp5_ASAP7_75t_L     g13338(.A1(new_n361), .A2(\b[63] ), .B1(new_n359), .B2(new_n12961), .C(new_n13594), .Y(new_n13595));
  XNOR2x2_ASAP7_75t_L       g13339(.A(new_n346), .B(new_n13595), .Y(new_n13596));
  A2O1A1Ixp33_ASAP7_75t_L   g13340(.A1(new_n13556), .A2(new_n13565), .B(new_n13557), .C(new_n13596), .Y(new_n13597));
  AOI21xp33_ASAP7_75t_L     g13341(.A1(new_n13556), .A2(new_n13565), .B(new_n13557), .Y(new_n13598));
  INVx1_ASAP7_75t_L         g13342(.A(new_n13596), .Y(new_n13599));
  NAND2xp33_ASAP7_75t_L     g13343(.A(new_n13599), .B(new_n13598), .Y(new_n13600));
  OAI22xp33_ASAP7_75t_L     g13344(.A1(new_n1550), .A2(new_n10332), .B1(new_n10309), .B2(new_n712), .Y(new_n13601));
  AOI221xp5_ASAP7_75t_L     g13345(.A1(new_n640), .A2(\b[57] ), .B1(new_n718), .B2(new_n10991), .C(new_n13601), .Y(new_n13602));
  XNOR2x2_ASAP7_75t_L       g13346(.A(new_n637), .B(new_n13602), .Y(new_n13603));
  INVx1_ASAP7_75t_L         g13347(.A(new_n13603), .Y(new_n13604));
  INVx1_ASAP7_75t_L         g13348(.A(new_n13532), .Y(new_n13605));
  NAND3xp33_ASAP7_75t_L     g13349(.A(new_n13529), .B(new_n13528), .C(new_n13605), .Y(new_n13606));
  A2O1A1Ixp33_ASAP7_75t_L   g13350(.A1(new_n13533), .A2(new_n13532), .B(new_n13536), .C(new_n13606), .Y(new_n13607));
  NOR2xp33_ASAP7_75t_L      g13351(.A(new_n13604), .B(new_n13607), .Y(new_n13608));
  A2O1A1O1Ixp25_ASAP7_75t_L g13352(.A1(new_n13532), .A2(new_n13533), .B(new_n13536), .C(new_n13606), .D(new_n13603), .Y(new_n13609));
  OAI22xp33_ASAP7_75t_L     g13353(.A1(new_n1285), .A2(new_n8427), .B1(new_n8755), .B2(new_n2118), .Y(new_n13610));
  AOI221xp5_ASAP7_75t_L     g13354(.A1(new_n1209), .A2(\b[51] ), .B1(new_n1216), .B2(new_n8790), .C(new_n13610), .Y(new_n13611));
  XNOR2x2_ASAP7_75t_L       g13355(.A(new_n1206), .B(new_n13611), .Y(new_n13612));
  O2A1O1Ixp33_ASAP7_75t_L   g13356(.A1(new_n13230), .A2(new_n13225), .B(new_n13517), .C(new_n13510), .Y(new_n13613));
  NAND2xp33_ASAP7_75t_L     g13357(.A(new_n13612), .B(new_n13613), .Y(new_n13614));
  INVx1_ASAP7_75t_L         g13358(.A(new_n13614), .Y(new_n13615));
  INVx1_ASAP7_75t_L         g13359(.A(new_n13510), .Y(new_n13616));
  A2O1A1O1Ixp25_ASAP7_75t_L g13360(.A1(new_n13515), .A2(new_n13298), .B(new_n13295), .C(new_n13616), .D(new_n13612), .Y(new_n13617));
  NOR2xp33_ASAP7_75t_L      g13361(.A(new_n13617), .B(new_n13615), .Y(new_n13618));
  OAI22xp33_ASAP7_75t_L     g13362(.A1(new_n1654), .A2(new_n7270), .B1(new_n7552), .B2(new_n1517), .Y(new_n13619));
  AOI221xp5_ASAP7_75t_L     g13363(.A1(new_n1511), .A2(\b[48] ), .B1(new_n1513), .B2(new_n11656), .C(new_n13619), .Y(new_n13620));
  XNOR2x2_ASAP7_75t_L       g13364(.A(new_n1501), .B(new_n13620), .Y(new_n13621));
  INVx1_ASAP7_75t_L         g13365(.A(new_n13621), .Y(new_n13622));
  A2O1A1O1Ixp25_ASAP7_75t_L g13366(.A1(new_n13490), .A2(new_n13302), .B(new_n13493), .C(new_n13503), .D(new_n13508), .Y(new_n13623));
  INVx1_ASAP7_75t_L         g13367(.A(new_n13623), .Y(new_n13624));
  NOR2xp33_ASAP7_75t_L      g13368(.A(new_n13622), .B(new_n13624), .Y(new_n13625));
  A2O1A1O1Ixp25_ASAP7_75t_L g13369(.A1(new_n13200), .A2(new_n13300), .B(new_n13202), .C(new_n13490), .D(new_n13493), .Y(new_n13626));
  A2O1A1O1Ixp25_ASAP7_75t_L g13370(.A1(new_n13504), .A2(new_n13626), .B(new_n13507), .C(new_n13511), .D(new_n13621), .Y(new_n13627));
  OAI22xp33_ASAP7_75t_L     g13371(.A1(new_n2089), .A2(new_n6671), .B1(new_n6944), .B2(new_n1962), .Y(new_n13628));
  AOI221xp5_ASAP7_75t_L     g13372(.A1(new_n1955), .A2(\b[45] ), .B1(new_n1964), .B2(new_n7256), .C(new_n13628), .Y(new_n13629));
  XNOR2x2_ASAP7_75t_L       g13373(.A(new_n1952), .B(new_n13629), .Y(new_n13630));
  A2O1A1Ixp33_ASAP7_75t_L   g13374(.A1(new_n13302), .A2(new_n13489), .B(new_n13491), .C(new_n13630), .Y(new_n13631));
  A2O1A1O1Ixp25_ASAP7_75t_L g13375(.A1(new_n13200), .A2(new_n13300), .B(new_n13202), .C(new_n13489), .D(new_n13491), .Y(new_n13632));
  INVx1_ASAP7_75t_L         g13376(.A(new_n13630), .Y(new_n13633));
  NAND2xp33_ASAP7_75t_L     g13377(.A(new_n13633), .B(new_n13632), .Y(new_n13634));
  NAND2xp33_ASAP7_75t_L     g13378(.A(new_n13631), .B(new_n13634), .Y(new_n13635));
  OAI22xp33_ASAP7_75t_L     g13379(.A1(new_n2572), .A2(new_n5855), .B1(new_n6110), .B2(new_n2410), .Y(new_n13636));
  AOI221xp5_ASAP7_75t_L     g13380(.A1(new_n2423), .A2(\b[42] ), .B1(new_n2417), .B2(new_n6389), .C(new_n13636), .Y(new_n13637));
  XNOR2x2_ASAP7_75t_L       g13381(.A(new_n2413), .B(new_n13637), .Y(new_n13638));
  INVx1_ASAP7_75t_L         g13382(.A(new_n13638), .Y(new_n13639));
  A2O1A1O1Ixp25_ASAP7_75t_L g13383(.A1(new_n13457), .A2(new_n13461), .B(new_n13476), .C(new_n13472), .D(new_n13487), .Y(new_n13640));
  INVx1_ASAP7_75t_L         g13384(.A(new_n13640), .Y(new_n13641));
  NOR2xp33_ASAP7_75t_L      g13385(.A(new_n13639), .B(new_n13641), .Y(new_n13642));
  NOR2xp33_ASAP7_75t_L      g13386(.A(new_n13466), .B(new_n13468), .Y(new_n13643));
  A2O1A1Ixp33_ASAP7_75t_L   g13387(.A1(new_n13469), .A2(new_n13643), .B(new_n13488), .C(new_n13639), .Y(new_n13644));
  INVx1_ASAP7_75t_L         g13388(.A(new_n13644), .Y(new_n13645));
  NOR2xp33_ASAP7_75t_L      g13389(.A(new_n13642), .B(new_n13645), .Y(new_n13646));
  INVx1_ASAP7_75t_L         g13390(.A(new_n13646), .Y(new_n13647));
  NOR2xp33_ASAP7_75t_L      g13391(.A(new_n5570), .B(new_n2930), .Y(new_n13648));
  AOI221xp5_ASAP7_75t_L     g13392(.A1(\b[37] ), .A2(new_n3129), .B1(\b[38] ), .B2(new_n2936), .C(new_n13648), .Y(new_n13649));
  OA211x2_ASAP7_75t_L       g13393(.A1(new_n2940), .A2(new_n5578), .B(new_n13649), .C(\a[29] ), .Y(new_n13650));
  O2A1O1Ixp33_ASAP7_75t_L   g13394(.A1(new_n2940), .A2(new_n5578), .B(new_n13649), .C(\a[29] ), .Y(new_n13651));
  NOR2xp33_ASAP7_75t_L      g13395(.A(new_n13651), .B(new_n13650), .Y(new_n13652));
  A2O1A1O1Ixp25_ASAP7_75t_L g13396(.A1(new_n13450), .A2(new_n13451), .B(new_n13456), .C(new_n13458), .D(new_n13652), .Y(new_n13653));
  AND3x1_ASAP7_75t_L        g13397(.A(new_n13461), .B(new_n13652), .C(new_n13458), .Y(new_n13654));
  NOR2xp33_ASAP7_75t_L      g13398(.A(new_n13653), .B(new_n13654), .Y(new_n13655));
  NOR2xp33_ASAP7_75t_L      g13399(.A(new_n4101), .B(new_n4147), .Y(new_n13656));
  AOI221xp5_ASAP7_75t_L     g13400(.A1(\b[31] ), .A2(new_n4402), .B1(\b[32] ), .B2(new_n4155), .C(new_n13656), .Y(new_n13657));
  OAI21xp33_ASAP7_75t_L     g13401(.A1(new_n4150), .A2(new_n4108), .B(new_n13657), .Y(new_n13658));
  NOR2xp33_ASAP7_75t_L      g13402(.A(new_n4145), .B(new_n13658), .Y(new_n13659));
  O2A1O1Ixp33_ASAP7_75t_L   g13403(.A1(new_n4150), .A2(new_n4108), .B(new_n13657), .C(\a[35] ), .Y(new_n13660));
  NOR2xp33_ASAP7_75t_L      g13404(.A(new_n13660), .B(new_n13659), .Y(new_n13661));
  INVx1_ASAP7_75t_L         g13405(.A(new_n13661), .Y(new_n13662));
  NAND3xp33_ASAP7_75t_L     g13406(.A(new_n13412), .B(new_n13408), .C(new_n13420), .Y(new_n13663));
  O2A1O1Ixp33_ASAP7_75t_L   g13407(.A1(new_n13069), .A2(new_n13068), .B(new_n13354), .C(new_n13351), .Y(new_n13664));
  NOR2xp33_ASAP7_75t_L      g13408(.A(new_n289), .B(new_n13030), .Y(new_n13665));
  A2O1A1Ixp33_ASAP7_75t_L   g13409(.A1(new_n13028), .A2(\b[3] ), .B(new_n13665), .C(\a[2] ), .Y(new_n13666));
  O2A1O1Ixp33_ASAP7_75t_L   g13410(.A1(new_n12669), .A2(new_n12671), .B(\b[3] ), .C(new_n13665), .Y(new_n13667));
  NAND2xp33_ASAP7_75t_L     g13411(.A(new_n257), .B(new_n13667), .Y(new_n13668));
  NAND2xp33_ASAP7_75t_L     g13412(.A(new_n13666), .B(new_n13668), .Y(new_n13669));
  NOR2xp33_ASAP7_75t_L      g13413(.A(new_n384), .B(new_n12318), .Y(new_n13670));
  AOI221xp5_ASAP7_75t_L     g13414(.A1(new_n11995), .A2(\b[6] ), .B1(new_n13314), .B2(\b[4] ), .C(new_n13670), .Y(new_n13671));
  INVx1_ASAP7_75t_L         g13415(.A(new_n13671), .Y(new_n13672));
  A2O1A1Ixp33_ASAP7_75t_L   g13416(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n13671), .Y(new_n13673));
  O2A1O1Ixp33_ASAP7_75t_L   g13417(.A1(new_n5363), .A2(new_n13672), .B(new_n13673), .C(new_n11987), .Y(new_n13674));
  O2A1O1Ixp33_ASAP7_75t_L   g13418(.A1(new_n11998), .A2(new_n434), .B(new_n13671), .C(\a[62] ), .Y(new_n13675));
  NOR2xp33_ASAP7_75t_L      g13419(.A(new_n13675), .B(new_n13674), .Y(new_n13676));
  NOR2xp33_ASAP7_75t_L      g13420(.A(new_n13669), .B(new_n13676), .Y(new_n13677));
  AOI211xp5_ASAP7_75t_L     g13421(.A1(new_n13668), .A2(new_n13666), .B(new_n13675), .C(new_n13674), .Y(new_n13678));
  NOR2xp33_ASAP7_75t_L      g13422(.A(new_n13678), .B(new_n13677), .Y(new_n13679));
  INVx1_ASAP7_75t_L         g13423(.A(new_n13679), .Y(new_n13680));
  O2A1O1Ixp33_ASAP7_75t_L   g13424(.A1(new_n13324), .A2(new_n13327), .B(new_n13321), .C(new_n13680), .Y(new_n13681));
  A2O1A1Ixp33_ASAP7_75t_L   g13425(.A1(new_n13046), .A2(new_n13039), .B(new_n13324), .C(new_n13321), .Y(new_n13682));
  NOR2xp33_ASAP7_75t_L      g13426(.A(new_n13679), .B(new_n13682), .Y(new_n13683));
  NOR2xp33_ASAP7_75t_L      g13427(.A(new_n13681), .B(new_n13683), .Y(new_n13684));
  NOR2xp33_ASAP7_75t_L      g13428(.A(new_n448), .B(new_n11354), .Y(new_n13685));
  AOI221xp5_ASAP7_75t_L     g13429(.A1(\b[9] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[8] ), .C(new_n13685), .Y(new_n13686));
  O2A1O1Ixp33_ASAP7_75t_L   g13430(.A1(new_n11053), .A2(new_n1066), .B(new_n13686), .C(new_n11048), .Y(new_n13687));
  INVx1_ASAP7_75t_L         g13431(.A(new_n13687), .Y(new_n13688));
  O2A1O1Ixp33_ASAP7_75t_L   g13432(.A1(new_n11053), .A2(new_n1066), .B(new_n13686), .C(\a[59] ), .Y(new_n13689));
  A2O1A1Ixp33_ASAP7_75t_L   g13433(.A1(\a[59] ), .A2(new_n13688), .B(new_n13689), .C(new_n13684), .Y(new_n13690));
  INVx1_ASAP7_75t_L         g13434(.A(new_n13689), .Y(new_n13691));
  O2A1O1Ixp33_ASAP7_75t_L   g13435(.A1(new_n13687), .A2(new_n11048), .B(new_n13691), .C(new_n13684), .Y(new_n13692));
  AOI21xp33_ASAP7_75t_L     g13436(.A1(new_n13690), .A2(new_n13684), .B(new_n13692), .Y(new_n13693));
  A2O1A1Ixp33_ASAP7_75t_L   g13437(.A1(new_n13340), .A2(new_n13337), .B(new_n13339), .C(new_n13693), .Y(new_n13694));
  INVx1_ASAP7_75t_L         g13438(.A(new_n13344), .Y(new_n13695));
  A2O1A1Ixp33_ASAP7_75t_L   g13439(.A1(new_n13690), .A2(new_n13684), .B(new_n13692), .C(new_n13695), .Y(new_n13696));
  NOR2xp33_ASAP7_75t_L      g13440(.A(new_n748), .B(new_n10388), .Y(new_n13697));
  AOI221xp5_ASAP7_75t_L     g13441(.A1(new_n10086), .A2(\b[12] ), .B1(new_n11361), .B2(\b[10] ), .C(new_n13697), .Y(new_n13698));
  INVx1_ASAP7_75t_L         g13442(.A(new_n13698), .Y(new_n13699));
  O2A1O1Ixp33_ASAP7_75t_L   g13443(.A1(new_n10088), .A2(new_n841), .B(new_n13698), .C(new_n10083), .Y(new_n13700));
  INVx1_ASAP7_75t_L         g13444(.A(new_n13700), .Y(new_n13701));
  NOR2xp33_ASAP7_75t_L      g13445(.A(new_n10083), .B(new_n13700), .Y(new_n13702));
  A2O1A1O1Ixp25_ASAP7_75t_L g13446(.A1(new_n10386), .A2(new_n1057), .B(new_n13699), .C(new_n13701), .D(new_n13702), .Y(new_n13703));
  NAND3xp33_ASAP7_75t_L     g13447(.A(new_n13696), .B(new_n13694), .C(new_n13703), .Y(new_n13704));
  NAND2xp33_ASAP7_75t_L     g13448(.A(new_n13694), .B(new_n13696), .Y(new_n13705));
  O2A1O1Ixp33_ASAP7_75t_L   g13449(.A1(new_n10088), .A2(new_n841), .B(new_n13698), .C(\a[56] ), .Y(new_n13706));
  A2O1A1Ixp33_ASAP7_75t_L   g13450(.A1(\a[56] ), .A2(new_n13701), .B(new_n13706), .C(new_n13705), .Y(new_n13707));
  NAND2xp33_ASAP7_75t_L     g13451(.A(new_n13704), .B(new_n13707), .Y(new_n13708));
  XNOR2x2_ASAP7_75t_L       g13452(.A(new_n13664), .B(new_n13708), .Y(new_n13709));
  OAI22xp33_ASAP7_75t_L     g13453(.A1(new_n9440), .A2(new_n936), .B1(new_n960), .B2(new_n10400), .Y(new_n13710));
  AOI221xp5_ASAP7_75t_L     g13454(.A1(new_n9102), .A2(\b[15] ), .B1(new_n9437), .B2(new_n1052), .C(new_n13710), .Y(new_n13711));
  XNOR2x2_ASAP7_75t_L       g13455(.A(new_n9099), .B(new_n13711), .Y(new_n13712));
  XOR2x2_ASAP7_75t_L        g13456(.A(new_n13712), .B(new_n13709), .Y(new_n13713));
  NAND3xp33_ASAP7_75t_L     g13457(.A(new_n13363), .B(new_n13362), .C(new_n13359), .Y(new_n13714));
  A2O1A1Ixp33_ASAP7_75t_L   g13458(.A1(new_n13367), .A2(new_n13358), .B(new_n13308), .C(new_n13714), .Y(new_n13715));
  XOR2x2_ASAP7_75t_L        g13459(.A(new_n13715), .B(new_n13713), .Y(new_n13716));
  NOR2xp33_ASAP7_75t_L      g13460(.A(new_n1349), .B(new_n10065), .Y(new_n13717));
  AOI221xp5_ASAP7_75t_L     g13461(.A1(new_n8175), .A2(\b[18] ), .B1(new_n8484), .B2(\b[16] ), .C(new_n13717), .Y(new_n13718));
  O2A1O1Ixp33_ASAP7_75t_L   g13462(.A1(new_n8176), .A2(new_n1464), .B(new_n13718), .C(new_n8172), .Y(new_n13719));
  OAI21xp33_ASAP7_75t_L     g13463(.A1(new_n8176), .A2(new_n1464), .B(new_n13718), .Y(new_n13720));
  NAND2xp33_ASAP7_75t_L     g13464(.A(new_n8172), .B(new_n13720), .Y(new_n13721));
  OA21x2_ASAP7_75t_L        g13465(.A1(new_n8172), .A2(new_n13719), .B(new_n13721), .Y(new_n13722));
  NAND2xp33_ASAP7_75t_L     g13466(.A(new_n13722), .B(new_n13716), .Y(new_n13723));
  O2A1O1Ixp33_ASAP7_75t_L   g13467(.A1(new_n13719), .A2(new_n8172), .B(new_n13721), .C(new_n13716), .Y(new_n13724));
  INVx1_ASAP7_75t_L         g13468(.A(new_n13724), .Y(new_n13725));
  NAND2xp33_ASAP7_75t_L     g13469(.A(new_n13723), .B(new_n13725), .Y(new_n13726));
  AOI21xp33_ASAP7_75t_L     g13470(.A1(new_n13376), .A2(new_n13375), .B(new_n13372), .Y(new_n13727));
  O2A1O1Ixp33_ASAP7_75t_L   g13471(.A1(new_n13306), .A2(new_n13307), .B(new_n13377), .C(new_n13727), .Y(new_n13728));
  INVx1_ASAP7_75t_L         g13472(.A(new_n13728), .Y(new_n13729));
  NOR2xp33_ASAP7_75t_L      g13473(.A(new_n13729), .B(new_n13726), .Y(new_n13730));
  INVx1_ASAP7_75t_L         g13474(.A(new_n13722), .Y(new_n13731));
  NAND2xp33_ASAP7_75t_L     g13475(.A(new_n13731), .B(new_n13716), .Y(new_n13732));
  A2O1A1Ixp33_ASAP7_75t_L   g13476(.A1(new_n13732), .A2(new_n13716), .B(new_n13724), .C(new_n13729), .Y(new_n13733));
  INVx1_ASAP7_75t_L         g13477(.A(new_n13733), .Y(new_n13734));
  NOR2xp33_ASAP7_75t_L      g13478(.A(new_n13734), .B(new_n13730), .Y(new_n13735));
  OAI22xp33_ASAP7_75t_L     g13479(.A1(new_n7614), .A2(new_n1599), .B1(new_n1745), .B2(new_n7312), .Y(new_n13736));
  AOI221xp5_ASAP7_75t_L     g13480(.A1(new_n7334), .A2(\b[21] ), .B1(new_n7322), .B2(new_n2836), .C(new_n13736), .Y(new_n13737));
  XNOR2x2_ASAP7_75t_L       g13481(.A(new_n7316), .B(new_n13737), .Y(new_n13738));
  INVx1_ASAP7_75t_L         g13482(.A(new_n13738), .Y(new_n13739));
  NOR2xp33_ASAP7_75t_L      g13483(.A(new_n13739), .B(new_n13735), .Y(new_n13740));
  NAND2xp33_ASAP7_75t_L     g13484(.A(new_n13739), .B(new_n13735), .Y(new_n13741));
  INVx1_ASAP7_75t_L         g13485(.A(new_n13741), .Y(new_n13742));
  A2O1A1Ixp33_ASAP7_75t_L   g13486(.A1(new_n13395), .A2(new_n13386), .B(new_n13304), .C(new_n13404), .Y(new_n13743));
  INVx1_ASAP7_75t_L         g13487(.A(new_n13743), .Y(new_n13744));
  NOR3xp33_ASAP7_75t_L      g13488(.A(new_n13742), .B(new_n13744), .C(new_n13740), .Y(new_n13745));
  INVx1_ASAP7_75t_L         g13489(.A(new_n13740), .Y(new_n13746));
  AOI21xp33_ASAP7_75t_L     g13490(.A1(new_n13746), .A2(new_n13741), .B(new_n13743), .Y(new_n13747));
  OAI22xp33_ASAP7_75t_L     g13491(.A1(new_n7304), .A2(new_n2188), .B1(new_n2045), .B2(new_n6741), .Y(new_n13748));
  AOI221xp5_ASAP7_75t_L     g13492(.A1(new_n6442), .A2(\b[24] ), .B1(new_n6450), .B2(new_n2216), .C(new_n13748), .Y(new_n13749));
  XNOR2x2_ASAP7_75t_L       g13493(.A(new_n6439), .B(new_n13749), .Y(new_n13750));
  INVx1_ASAP7_75t_L         g13494(.A(new_n13750), .Y(new_n13751));
  OR3x1_ASAP7_75t_L         g13495(.A(new_n13747), .B(new_n13745), .C(new_n13751), .Y(new_n13752));
  OAI21xp33_ASAP7_75t_L     g13496(.A1(new_n13745), .A2(new_n13747), .B(new_n13751), .Y(new_n13753));
  AND2x2_ASAP7_75t_L        g13497(.A(new_n13753), .B(new_n13752), .Y(new_n13754));
  O2A1O1Ixp33_ASAP7_75t_L   g13498(.A1(new_n13116), .A2(new_n13121), .B(new_n13406), .C(new_n13409), .Y(new_n13755));
  NAND2xp33_ASAP7_75t_L     g13499(.A(new_n13755), .B(new_n13754), .Y(new_n13756));
  NAND2xp33_ASAP7_75t_L     g13500(.A(new_n13753), .B(new_n13752), .Y(new_n13757));
  A2O1A1Ixp33_ASAP7_75t_L   g13501(.A1(new_n13411), .A2(new_n13417), .B(new_n13409), .C(new_n13757), .Y(new_n13758));
  OAI22xp33_ASAP7_75t_L     g13502(.A1(new_n5640), .A2(new_n2703), .B1(new_n2377), .B2(new_n5925), .Y(new_n13759));
  AOI221xp5_ASAP7_75t_L     g13503(.A1(new_n5629), .A2(\b[27] ), .B1(new_n5637), .B2(new_n2887), .C(new_n13759), .Y(new_n13760));
  XNOR2x2_ASAP7_75t_L       g13504(.A(new_n5626), .B(new_n13760), .Y(new_n13761));
  NAND3xp33_ASAP7_75t_L     g13505(.A(new_n13756), .B(new_n13758), .C(new_n13761), .Y(new_n13762));
  NOR3xp33_ASAP7_75t_L      g13506(.A(new_n13757), .B(new_n13419), .C(new_n13409), .Y(new_n13763));
  NOR2xp33_ASAP7_75t_L      g13507(.A(new_n13755), .B(new_n13754), .Y(new_n13764));
  INVx1_ASAP7_75t_L         g13508(.A(new_n13761), .Y(new_n13765));
  OAI21xp33_ASAP7_75t_L     g13509(.A1(new_n13763), .A2(new_n13764), .B(new_n13765), .Y(new_n13766));
  NAND4xp25_ASAP7_75t_L     g13510(.A(new_n13766), .B(new_n13762), .C(new_n13663), .D(new_n13424), .Y(new_n13767));
  INVx1_ASAP7_75t_L         g13511(.A(new_n13767), .Y(new_n13768));
  AOI22xp33_ASAP7_75t_L     g13512(.A1(new_n13663), .A2(new_n13424), .B1(new_n13762), .B2(new_n13766), .Y(new_n13769));
  OAI22xp33_ASAP7_75t_L     g13513(.A1(new_n5144), .A2(new_n3079), .B1(new_n3098), .B2(new_n4903), .Y(new_n13770));
  AOI221xp5_ASAP7_75t_L     g13514(.A1(new_n4917), .A2(\b[30] ), .B1(new_n4912), .B2(new_n4813), .C(new_n13770), .Y(new_n13771));
  XNOR2x2_ASAP7_75t_L       g13515(.A(new_n4906), .B(new_n13771), .Y(new_n13772));
  OAI21xp33_ASAP7_75t_L     g13516(.A1(new_n13769), .A2(new_n13768), .B(new_n13772), .Y(new_n13773));
  INVx1_ASAP7_75t_L         g13517(.A(new_n13769), .Y(new_n13774));
  INVx1_ASAP7_75t_L         g13518(.A(new_n13772), .Y(new_n13775));
  NAND3xp33_ASAP7_75t_L     g13519(.A(new_n13774), .B(new_n13767), .C(new_n13775), .Y(new_n13776));
  NAND3xp33_ASAP7_75t_L     g13520(.A(new_n13424), .B(new_n13422), .C(new_n13430), .Y(new_n13777));
  A2O1A1Ixp33_ASAP7_75t_L   g13521(.A1(new_n13428), .A2(new_n13427), .B(new_n13433), .C(new_n13777), .Y(new_n13778));
  NAND3xp33_ASAP7_75t_L     g13522(.A(new_n13776), .B(new_n13773), .C(new_n13778), .Y(new_n13779));
  AO21x2_ASAP7_75t_L        g13523(.A1(new_n13773), .A2(new_n13776), .B(new_n13778), .Y(new_n13780));
  NAND3xp33_ASAP7_75t_L     g13524(.A(new_n13780), .B(new_n13779), .C(new_n13662), .Y(new_n13781));
  NAND2xp33_ASAP7_75t_L     g13525(.A(new_n13779), .B(new_n13780), .Y(new_n13782));
  NOR2xp33_ASAP7_75t_L      g13526(.A(new_n13662), .B(new_n13782), .Y(new_n13783));
  NOR2xp33_ASAP7_75t_L      g13527(.A(new_n4613), .B(new_n3510), .Y(new_n13784));
  AOI221xp5_ASAP7_75t_L     g13528(.A1(\b[34] ), .A2(new_n3708), .B1(\b[35] ), .B2(new_n3499), .C(new_n13784), .Y(new_n13785));
  OA211x2_ASAP7_75t_L       g13529(.A1(new_n3513), .A2(new_n4622), .B(new_n13785), .C(\a[32] ), .Y(new_n13786));
  O2A1O1Ixp33_ASAP7_75t_L   g13530(.A1(new_n3513), .A2(new_n4622), .B(new_n13785), .C(\a[32] ), .Y(new_n13787));
  NAND2xp33_ASAP7_75t_L     g13531(.A(new_n13434), .B(new_n13442), .Y(new_n13788));
  O2A1O1Ixp33_ASAP7_75t_L   g13532(.A1(new_n13435), .A2(new_n13436), .B(new_n13439), .C(new_n13441), .Y(new_n13789));
  INVx1_ASAP7_75t_L         g13533(.A(new_n13789), .Y(new_n13790));
  NOR2xp33_ASAP7_75t_L      g13534(.A(new_n13787), .B(new_n13786), .Y(new_n13791));
  O2A1O1Ixp33_ASAP7_75t_L   g13535(.A1(new_n13788), .A2(new_n13439), .B(new_n13790), .C(new_n13791), .Y(new_n13792));
  INVx1_ASAP7_75t_L         g13536(.A(new_n13792), .Y(new_n13793));
  INVx1_ASAP7_75t_L         g13537(.A(new_n13791), .Y(new_n13794));
  O2A1O1Ixp33_ASAP7_75t_L   g13538(.A1(new_n13788), .A2(new_n13439), .B(new_n13790), .C(new_n13794), .Y(new_n13795));
  O2A1O1Ixp33_ASAP7_75t_L   g13539(.A1(new_n13786), .A2(new_n13787), .B(new_n13793), .C(new_n13795), .Y(new_n13796));
  A2O1A1Ixp33_ASAP7_75t_L   g13540(.A1(new_n13781), .A2(new_n13662), .B(new_n13783), .C(new_n13796), .Y(new_n13797));
  O2A1O1Ixp33_ASAP7_75t_L   g13541(.A1(new_n13659), .A2(new_n13660), .B(new_n13781), .C(new_n13783), .Y(new_n13798));
  A2O1A1Ixp33_ASAP7_75t_L   g13542(.A1(new_n13794), .A2(new_n13793), .B(new_n13795), .C(new_n13798), .Y(new_n13799));
  NAND2xp33_ASAP7_75t_L     g13543(.A(new_n13797), .B(new_n13799), .Y(new_n13800));
  NAND2xp33_ASAP7_75t_L     g13544(.A(new_n13655), .B(new_n13800), .Y(new_n13801));
  INVx1_ASAP7_75t_L         g13545(.A(new_n13795), .Y(new_n13802));
  O2A1O1Ixp33_ASAP7_75t_L   g13546(.A1(new_n13791), .A2(new_n13792), .B(new_n13802), .C(new_n13798), .Y(new_n13803));
  O2A1O1Ixp33_ASAP7_75t_L   g13547(.A1(new_n13798), .A2(new_n13803), .B(new_n13799), .C(new_n13655), .Y(new_n13804));
  AOI21xp33_ASAP7_75t_L     g13548(.A1(new_n13801), .A2(new_n13655), .B(new_n13804), .Y(new_n13805));
  NOR2xp33_ASAP7_75t_L      g13549(.A(new_n13647), .B(new_n13805), .Y(new_n13806));
  NAND2xp33_ASAP7_75t_L     g13550(.A(new_n13647), .B(new_n13805), .Y(new_n13807));
  NAND2xp33_ASAP7_75t_L     g13551(.A(new_n13635), .B(new_n13807), .Y(new_n13808));
  A2O1A1Ixp33_ASAP7_75t_L   g13552(.A1(new_n13634), .A2(new_n13631), .B(new_n13806), .C(new_n13807), .Y(new_n13809));
  A2O1A1O1Ixp25_ASAP7_75t_L g13553(.A1(new_n13801), .A2(new_n13655), .B(new_n13804), .C(new_n13646), .D(new_n13809), .Y(new_n13810));
  O2A1O1Ixp33_ASAP7_75t_L   g13554(.A1(new_n13806), .A2(new_n13808), .B(new_n13635), .C(new_n13810), .Y(new_n13811));
  NOR3xp33_ASAP7_75t_L      g13555(.A(new_n13811), .B(new_n13627), .C(new_n13625), .Y(new_n13812));
  INVx1_ASAP7_75t_L         g13556(.A(new_n13617), .Y(new_n13813));
  OAI21xp33_ASAP7_75t_L     g13557(.A1(new_n13625), .A2(new_n13627), .B(new_n13811), .Y(new_n13814));
  NAND3xp33_ASAP7_75t_L     g13558(.A(new_n13614), .B(new_n13814), .C(new_n13813), .Y(new_n13815));
  NOR2xp33_ASAP7_75t_L      g13559(.A(new_n13627), .B(new_n13625), .Y(new_n13816));
  INVx1_ASAP7_75t_L         g13560(.A(new_n13635), .Y(new_n13817));
  A2O1A1Ixp33_ASAP7_75t_L   g13561(.A1(new_n13801), .A2(new_n13655), .B(new_n13804), .C(new_n13646), .Y(new_n13818));
  O2A1O1Ixp33_ASAP7_75t_L   g13562(.A1(new_n13642), .A2(new_n13645), .B(new_n13805), .C(new_n13817), .Y(new_n13819));
  NAND3xp33_ASAP7_75t_L     g13563(.A(new_n13807), .B(new_n13818), .C(new_n13817), .Y(new_n13820));
  A2O1A1Ixp33_ASAP7_75t_L   g13564(.A1(new_n13818), .A2(new_n13819), .B(new_n13817), .C(new_n13820), .Y(new_n13821));
  NOR2xp33_ASAP7_75t_L      g13565(.A(new_n13821), .B(new_n13816), .Y(new_n13822));
  AOI211xp5_ASAP7_75t_L     g13566(.A1(new_n13813), .A2(new_n13614), .B(new_n13822), .C(new_n13812), .Y(new_n13823));
  O2A1O1Ixp33_ASAP7_75t_L   g13567(.A1(new_n13812), .A2(new_n13815), .B(new_n13618), .C(new_n13823), .Y(new_n13824));
  O2A1O1Ixp33_ASAP7_75t_L   g13568(.A1(new_n13295), .A2(new_n13516), .B(new_n13518), .C(new_n13521), .Y(new_n13825));
  NOR2xp33_ASAP7_75t_L      g13569(.A(new_n9709), .B(new_n869), .Y(new_n13826));
  AOI221xp5_ASAP7_75t_L     g13570(.A1(\b[52] ), .A2(new_n985), .B1(\b[53] ), .B2(new_n885), .C(new_n13826), .Y(new_n13827));
  OA211x2_ASAP7_75t_L       g13571(.A1(new_n872), .A2(new_n9718), .B(new_n13827), .C(\a[14] ), .Y(new_n13828));
  O2A1O1Ixp33_ASAP7_75t_L   g13572(.A1(new_n872), .A2(new_n9718), .B(new_n13827), .C(\a[14] ), .Y(new_n13829));
  NOR2xp33_ASAP7_75t_L      g13573(.A(new_n13829), .B(new_n13828), .Y(new_n13830));
  INVx1_ASAP7_75t_L         g13574(.A(new_n13830), .Y(new_n13831));
  A2O1A1Ixp33_ASAP7_75t_L   g13575(.A1(new_n13522), .A2(new_n13294), .B(new_n13825), .C(new_n13831), .Y(new_n13832));
  AOI211xp5_ASAP7_75t_L     g13576(.A1(new_n13522), .A2(new_n13294), .B(new_n13825), .C(new_n13830), .Y(new_n13833));
  A2O1A1O1Ixp25_ASAP7_75t_L g13577(.A1(new_n13522), .A2(new_n13294), .B(new_n13825), .C(new_n13832), .D(new_n13833), .Y(new_n13834));
  XOR2x2_ASAP7_75t_L        g13578(.A(new_n13834), .B(new_n13824), .Y(new_n13835));
  OR3x1_ASAP7_75t_L         g13579(.A(new_n13835), .B(new_n13608), .C(new_n13609), .Y(new_n13836));
  OAI21xp33_ASAP7_75t_L     g13580(.A1(new_n13609), .A2(new_n13608), .B(new_n13835), .Y(new_n13837));
  NAND2xp33_ASAP7_75t_L     g13581(.A(new_n13837), .B(new_n13836), .Y(new_n13838));
  INVx1_ASAP7_75t_L         g13582(.A(new_n11634), .Y(new_n13839));
  OAI22xp33_ASAP7_75t_L     g13583(.A1(new_n513), .A2(new_n11591), .B1(new_n11303), .B2(new_n506), .Y(new_n13840));
  AOI221xp5_ASAP7_75t_L     g13584(.A1(new_n475), .A2(\b[60] ), .B1(new_n483), .B2(new_n13839), .C(new_n13840), .Y(new_n13841));
  XNOR2x2_ASAP7_75t_L       g13585(.A(\a[8] ), .B(new_n13841), .Y(new_n13842));
  OAI211xp5_ASAP7_75t_L     g13586(.A1(new_n13549), .A2(new_n13551), .B(new_n13546), .C(new_n13842), .Y(new_n13843));
  XNOR2x2_ASAP7_75t_L       g13587(.A(new_n466), .B(new_n13841), .Y(new_n13844));
  A2O1A1Ixp33_ASAP7_75t_L   g13588(.A1(new_n13542), .A2(new_n13553), .B(new_n13552), .C(new_n13844), .Y(new_n13845));
  NAND2xp33_ASAP7_75t_L     g13589(.A(new_n13845), .B(new_n13843), .Y(new_n13846));
  XOR2x2_ASAP7_75t_L        g13590(.A(new_n13838), .B(new_n13846), .Y(new_n13847));
  AOI21xp33_ASAP7_75t_L     g13591(.A1(new_n13600), .A2(new_n13597), .B(new_n13847), .Y(new_n13848));
  INVx1_ASAP7_75t_L         g13592(.A(new_n13597), .Y(new_n13849));
  AOI211xp5_ASAP7_75t_L     g13593(.A1(new_n13556), .A2(new_n13565), .B(new_n13596), .C(new_n13557), .Y(new_n13850));
  A2O1A1Ixp33_ASAP7_75t_L   g13594(.A1(new_n13542), .A2(new_n13553), .B(new_n13552), .C(new_n13842), .Y(new_n13851));
  INVx1_ASAP7_75t_L         g13595(.A(new_n13845), .Y(new_n13852));
  A2O1A1Ixp33_ASAP7_75t_L   g13596(.A1(new_n13851), .A2(new_n13842), .B(new_n13852), .C(new_n13838), .Y(new_n13853));
  O2A1O1Ixp33_ASAP7_75t_L   g13597(.A1(new_n13549), .A2(new_n13551), .B(new_n13546), .C(new_n13844), .Y(new_n13854));
  O2A1O1Ixp33_ASAP7_75t_L   g13598(.A1(new_n13844), .A2(new_n13854), .B(new_n13845), .C(new_n13838), .Y(new_n13855));
  AOI21xp33_ASAP7_75t_L     g13599(.A1(new_n13853), .A2(new_n13838), .B(new_n13855), .Y(new_n13856));
  NOR3xp33_ASAP7_75t_L      g13600(.A(new_n13856), .B(new_n13849), .C(new_n13850), .Y(new_n13857));
  INVx1_ASAP7_75t_L         g13601(.A(new_n13571), .Y(new_n13858));
  A2O1A1Ixp33_ASAP7_75t_L   g13602(.A1(new_n13563), .A2(new_n13566), .B(new_n13575), .C(new_n13858), .Y(new_n13859));
  NOR3xp33_ASAP7_75t_L      g13603(.A(new_n13857), .B(new_n13859), .C(new_n13848), .Y(new_n13860));
  INVx1_ASAP7_75t_L         g13604(.A(new_n13598), .Y(new_n13861));
  A2O1A1Ixp33_ASAP7_75t_L   g13605(.A1(new_n13556), .A2(new_n13565), .B(new_n13557), .C(new_n13599), .Y(new_n13862));
  A2O1A1Ixp33_ASAP7_75t_L   g13606(.A1(new_n13862), .A2(new_n13861), .B(new_n13850), .C(new_n13856), .Y(new_n13863));
  NAND3xp33_ASAP7_75t_L     g13607(.A(new_n13600), .B(new_n13847), .C(new_n13597), .Y(new_n13864));
  O2A1O1Ixp33_ASAP7_75t_L   g13608(.A1(new_n13578), .A2(new_n13579), .B(new_n13576), .C(new_n13571), .Y(new_n13865));
  AOI21xp33_ASAP7_75t_L     g13609(.A1(new_n13863), .A2(new_n13864), .B(new_n13865), .Y(new_n13866));
  NOR2xp33_ASAP7_75t_L      g13610(.A(new_n13866), .B(new_n13860), .Y(new_n13867));
  O2A1O1Ixp33_ASAP7_75t_L   g13611(.A1(new_n13577), .A2(new_n13581), .B(new_n13583), .C(new_n13590), .Y(new_n13868));
  XNOR2x2_ASAP7_75t_L       g13612(.A(new_n13867), .B(new_n13868), .Y(\f[66] ));
  INVx1_ASAP7_75t_L         g13613(.A(new_n13862), .Y(new_n13870));
  O2A1O1Ixp33_ASAP7_75t_L   g13614(.A1(new_n13850), .A2(new_n13861), .B(new_n13847), .C(new_n13870), .Y(new_n13871));
  O2A1O1Ixp33_ASAP7_75t_L   g13615(.A1(new_n13596), .A2(new_n13870), .B(new_n13597), .C(new_n13856), .Y(new_n13872));
  O2A1O1Ixp33_ASAP7_75t_L   g13616(.A1(new_n13842), .A2(new_n13852), .B(new_n13838), .C(new_n13854), .Y(new_n13873));
  INVx1_ASAP7_75t_L         g13617(.A(new_n375), .Y(new_n13874));
  AOI22xp33_ASAP7_75t_L     g13618(.A1(new_n349), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n13874), .Y(new_n13875));
  A2O1A1Ixp33_ASAP7_75t_L   g13619(.A1(new_n12990), .A2(new_n12988), .B(new_n356), .C(new_n13875), .Y(new_n13876));
  NOR2xp33_ASAP7_75t_L      g13620(.A(new_n346), .B(new_n13876), .Y(new_n13877));
  O2A1O1Ixp33_ASAP7_75t_L   g13621(.A1(new_n356), .A2(new_n12993), .B(new_n13875), .C(\a[5] ), .Y(new_n13878));
  NOR2xp33_ASAP7_75t_L      g13622(.A(new_n13878), .B(new_n13877), .Y(new_n13879));
  INVx1_ASAP7_75t_L         g13623(.A(new_n13879), .Y(new_n13880));
  NOR2xp33_ASAP7_75t_L      g13624(.A(new_n13609), .B(new_n13608), .Y(new_n13881));
  OAI22xp33_ASAP7_75t_L     g13625(.A1(new_n513), .A2(new_n11626), .B1(new_n11591), .B2(new_n506), .Y(new_n13882));
  AOI221xp5_ASAP7_75t_L     g13626(.A1(new_n475), .A2(\b[61] ), .B1(new_n483), .B2(new_n12269), .C(new_n13882), .Y(new_n13883));
  XNOR2x2_ASAP7_75t_L       g13627(.A(\a[8] ), .B(new_n13883), .Y(new_n13884));
  A2O1A1Ixp33_ASAP7_75t_L   g13628(.A1(new_n13881), .A2(new_n13835), .B(new_n13609), .C(new_n13884), .Y(new_n13885));
  XNOR2x2_ASAP7_75t_L       g13629(.A(new_n466), .B(new_n13883), .Y(new_n13886));
  AOI211xp5_ASAP7_75t_L     g13630(.A1(new_n13881), .A2(new_n13835), .B(new_n13886), .C(new_n13609), .Y(new_n13887));
  A2O1A1O1Ixp25_ASAP7_75t_L g13631(.A1(new_n13881), .A2(new_n13835), .B(new_n13609), .C(new_n13885), .D(new_n13887), .Y(new_n13888));
  OAI22xp33_ASAP7_75t_L     g13632(.A1(new_n980), .A2(new_n9683), .B1(new_n9709), .B2(new_n864), .Y(new_n13889));
  AOI221xp5_ASAP7_75t_L     g13633(.A1(new_n886), .A2(\b[55] ), .B1(new_n873), .B2(new_n10320), .C(new_n13889), .Y(new_n13890));
  XNOR2x2_ASAP7_75t_L       g13634(.A(new_n867), .B(new_n13890), .Y(new_n13891));
  INVx1_ASAP7_75t_L         g13635(.A(new_n13891), .Y(new_n13892));
  A2O1A1Ixp33_ASAP7_75t_L   g13636(.A1(new_n13816), .A2(new_n13821), .B(new_n13815), .C(new_n13813), .Y(new_n13893));
  NOR2xp33_ASAP7_75t_L      g13637(.A(new_n13892), .B(new_n13893), .Y(new_n13894));
  O2A1O1Ixp33_ASAP7_75t_L   g13638(.A1(new_n13812), .A2(new_n13815), .B(new_n13813), .C(new_n13891), .Y(new_n13895));
  OAI22xp33_ASAP7_75t_L     g13639(.A1(new_n1654), .A2(new_n7552), .B1(new_n7860), .B2(new_n1517), .Y(new_n13896));
  AOI221xp5_ASAP7_75t_L     g13640(.A1(new_n1511), .A2(\b[49] ), .B1(new_n1513), .B2(new_n8438), .C(new_n13896), .Y(new_n13897));
  XNOR2x2_ASAP7_75t_L       g13641(.A(new_n1501), .B(new_n13897), .Y(new_n13898));
  A2O1A1Ixp33_ASAP7_75t_L   g13642(.A1(new_n13489), .A2(new_n13302), .B(new_n13491), .C(new_n13633), .Y(new_n13899));
  INVx1_ASAP7_75t_L         g13643(.A(new_n13899), .Y(new_n13900));
  O2A1O1Ixp33_ASAP7_75t_L   g13644(.A1(new_n13647), .A2(new_n13805), .B(new_n13819), .C(new_n13900), .Y(new_n13901));
  NAND2xp33_ASAP7_75t_L     g13645(.A(new_n13898), .B(new_n13901), .Y(new_n13902));
  O2A1O1Ixp33_ASAP7_75t_L   g13646(.A1(new_n13806), .A2(new_n13808), .B(new_n13899), .C(new_n13898), .Y(new_n13903));
  INVx1_ASAP7_75t_L         g13647(.A(new_n13903), .Y(new_n13904));
  OAI22xp33_ASAP7_75t_L     g13648(.A1(new_n3703), .A2(new_n4581), .B1(new_n4613), .B2(new_n3509), .Y(new_n13905));
  AOI221xp5_ASAP7_75t_L     g13649(.A1(new_n3503), .A2(\b[37] ), .B1(new_n3505), .B2(new_n10229), .C(new_n13905), .Y(new_n13906));
  XNOR2x2_ASAP7_75t_L       g13650(.A(new_n3493), .B(new_n13906), .Y(new_n13907));
  O2A1O1Ixp33_ASAP7_75t_L   g13651(.A1(new_n13661), .A2(new_n13782), .B(new_n13779), .C(new_n13907), .Y(new_n13908));
  AND3x1_ASAP7_75t_L        g13652(.A(new_n13781), .B(new_n13907), .C(new_n13779), .Y(new_n13909));
  OAI22xp33_ASAP7_75t_L     g13653(.A1(new_n4397), .A2(new_n3891), .B1(new_n4101), .B2(new_n4142), .Y(new_n13910));
  AOI221xp5_ASAP7_75t_L     g13654(.A1(new_n4156), .A2(\b[34] ), .B1(new_n4151), .B2(new_n5599), .C(new_n13910), .Y(new_n13911));
  XNOR2x2_ASAP7_75t_L       g13655(.A(new_n4145), .B(new_n13911), .Y(new_n13912));
  AOI21xp33_ASAP7_75t_L     g13656(.A1(new_n13767), .A2(new_n13775), .B(new_n13769), .Y(new_n13913));
  O2A1O1Ixp33_ASAP7_75t_L   g13657(.A1(new_n13727), .A2(new_n13380), .B(new_n13726), .C(new_n13742), .Y(new_n13914));
  INVx1_ASAP7_75t_L         g13658(.A(new_n13914), .Y(new_n13915));
  NOR2xp33_ASAP7_75t_L      g13659(.A(new_n534), .B(new_n11354), .Y(new_n13916));
  AOI221xp5_ASAP7_75t_L     g13660(.A1(\b[10] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[9] ), .C(new_n13916), .Y(new_n13917));
  O2A1O1Ixp33_ASAP7_75t_L   g13661(.A1(new_n11053), .A2(new_n1175), .B(new_n13917), .C(new_n11048), .Y(new_n13918));
  INVx1_ASAP7_75t_L         g13662(.A(new_n13918), .Y(new_n13919));
  O2A1O1Ixp33_ASAP7_75t_L   g13663(.A1(new_n11053), .A2(new_n1175), .B(new_n13917), .C(\a[59] ), .Y(new_n13920));
  NOR2xp33_ASAP7_75t_L      g13664(.A(new_n301), .B(new_n13030), .Y(new_n13921));
  INVx1_ASAP7_75t_L         g13665(.A(new_n13921), .Y(new_n13922));
  A2O1A1Ixp33_ASAP7_75t_L   g13666(.A1(new_n12685), .A2(new_n12686), .B(new_n332), .C(new_n13922), .Y(new_n13923));
  NOR2xp33_ASAP7_75t_L      g13667(.A(new_n257), .B(new_n13923), .Y(new_n13924));
  O2A1O1Ixp33_ASAP7_75t_L   g13668(.A1(new_n332), .A2(new_n12672), .B(new_n13922), .C(\a[2] ), .Y(new_n13925));
  NOR2xp33_ASAP7_75t_L      g13669(.A(new_n427), .B(new_n12318), .Y(new_n13926));
  AOI221xp5_ASAP7_75t_L     g13670(.A1(new_n11995), .A2(\b[7] ), .B1(new_n13314), .B2(\b[5] ), .C(new_n13926), .Y(new_n13927));
  O2A1O1Ixp33_ASAP7_75t_L   g13671(.A1(new_n11998), .A2(new_n456), .B(new_n13927), .C(new_n11987), .Y(new_n13928));
  O2A1O1Ixp33_ASAP7_75t_L   g13672(.A1(new_n11998), .A2(new_n456), .B(new_n13927), .C(\a[62] ), .Y(new_n13929));
  INVx1_ASAP7_75t_L         g13673(.A(new_n13929), .Y(new_n13930));
  O2A1O1Ixp33_ASAP7_75t_L   g13674(.A1(new_n332), .A2(new_n12672), .B(new_n13922), .C(new_n257), .Y(new_n13931));
  INVx1_ASAP7_75t_L         g13675(.A(new_n13931), .Y(new_n13932));
  A2O1A1O1Ixp25_ASAP7_75t_L g13676(.A1(new_n13028), .A2(\b[4] ), .B(new_n13921), .C(new_n13932), .D(new_n13924), .Y(new_n13933));
  O2A1O1Ixp33_ASAP7_75t_L   g13677(.A1(new_n11987), .A2(new_n13928), .B(new_n13930), .C(new_n13933), .Y(new_n13934));
  INVx1_ASAP7_75t_L         g13678(.A(new_n13934), .Y(new_n13935));
  O2A1O1Ixp33_ASAP7_75t_L   g13679(.A1(new_n11987), .A2(new_n13928), .B(new_n13930), .C(new_n13934), .Y(new_n13936));
  O2A1O1Ixp33_ASAP7_75t_L   g13680(.A1(new_n13924), .A2(new_n13925), .B(new_n13935), .C(new_n13936), .Y(new_n13937));
  A2O1A1O1Ixp25_ASAP7_75t_L g13681(.A1(new_n13028), .A2(\b[3] ), .B(new_n13665), .C(\a[2] ), .D(new_n13677), .Y(new_n13938));
  NAND2xp33_ASAP7_75t_L     g13682(.A(new_n13938), .B(new_n13937), .Y(new_n13939));
  INVx1_ASAP7_75t_L         g13683(.A(new_n13677), .Y(new_n13940));
  O2A1O1Ixp33_ASAP7_75t_L   g13684(.A1(new_n257), .A2(new_n13667), .B(new_n13940), .C(new_n13937), .Y(new_n13941));
  INVx1_ASAP7_75t_L         g13685(.A(new_n13941), .Y(new_n13942));
  NAND2xp33_ASAP7_75t_L     g13686(.A(new_n13939), .B(new_n13942), .Y(new_n13943));
  INVx1_ASAP7_75t_L         g13687(.A(new_n13920), .Y(new_n13944));
  O2A1O1Ixp33_ASAP7_75t_L   g13688(.A1(new_n13918), .A2(new_n11048), .B(new_n13944), .C(new_n13943), .Y(new_n13945));
  INVx1_ASAP7_75t_L         g13689(.A(new_n13945), .Y(new_n13946));
  NOR2xp33_ASAP7_75t_L      g13690(.A(new_n13943), .B(new_n13945), .Y(new_n13947));
  A2O1A1O1Ixp25_ASAP7_75t_L g13691(.A1(new_n13919), .A2(\a[59] ), .B(new_n13920), .C(new_n13946), .D(new_n13947), .Y(new_n13948));
  A2O1A1O1Ixp25_ASAP7_75t_L g13692(.A1(new_n13688), .A2(\a[59] ), .B(new_n13689), .C(new_n13684), .D(new_n13681), .Y(new_n13949));
  NAND2xp33_ASAP7_75t_L     g13693(.A(new_n13949), .B(new_n13948), .Y(new_n13950));
  A2O1A1Ixp33_ASAP7_75t_L   g13694(.A1(\a[59] ), .A2(new_n13919), .B(new_n13920), .C(new_n13943), .Y(new_n13951));
  O2A1O1Ixp33_ASAP7_75t_L   g13695(.A1(new_n13943), .A2(new_n13945), .B(new_n13951), .C(new_n13949), .Y(new_n13952));
  INVx1_ASAP7_75t_L         g13696(.A(new_n13952), .Y(new_n13953));
  AND2x2_ASAP7_75t_L        g13697(.A(new_n13953), .B(new_n13950), .Y(new_n13954));
  NOR2xp33_ASAP7_75t_L      g13698(.A(new_n833), .B(new_n10388), .Y(new_n13955));
  AOI221xp5_ASAP7_75t_L     g13699(.A1(new_n10086), .A2(\b[13] ), .B1(new_n11361), .B2(\b[11] ), .C(new_n13955), .Y(new_n13956));
  O2A1O1Ixp33_ASAP7_75t_L   g13700(.A1(new_n10088), .A2(new_n942), .B(new_n13956), .C(new_n10083), .Y(new_n13957));
  O2A1O1Ixp33_ASAP7_75t_L   g13701(.A1(new_n10088), .A2(new_n942), .B(new_n13956), .C(\a[56] ), .Y(new_n13958));
  INVx1_ASAP7_75t_L         g13702(.A(new_n13958), .Y(new_n13959));
  OAI21xp33_ASAP7_75t_L     g13703(.A1(new_n10083), .A2(new_n13957), .B(new_n13959), .Y(new_n13960));
  NOR2xp33_ASAP7_75t_L      g13704(.A(new_n13960), .B(new_n13954), .Y(new_n13961));
  NAND2xp33_ASAP7_75t_L     g13705(.A(new_n13953), .B(new_n13950), .Y(new_n13962));
  O2A1O1Ixp33_ASAP7_75t_L   g13706(.A1(new_n13957), .A2(new_n10083), .B(new_n13959), .C(new_n13962), .Y(new_n13963));
  NOR2xp33_ASAP7_75t_L      g13707(.A(new_n13963), .B(new_n13961), .Y(new_n13964));
  O2A1O1Ixp33_ASAP7_75t_L   g13708(.A1(new_n13330), .A2(new_n13336), .B(new_n13343), .C(new_n13693), .Y(new_n13965));
  O2A1O1Ixp33_ASAP7_75t_L   g13709(.A1(new_n13702), .A2(new_n13706), .B(new_n13705), .C(new_n13965), .Y(new_n13966));
  INVx1_ASAP7_75t_L         g13710(.A(new_n13966), .Y(new_n13967));
  NAND2xp33_ASAP7_75t_L     g13711(.A(new_n13967), .B(new_n13964), .Y(new_n13968));
  OAI21xp33_ASAP7_75t_L     g13712(.A1(new_n13963), .A2(new_n13961), .B(new_n13966), .Y(new_n13969));
  NAND2xp33_ASAP7_75t_L     g13713(.A(new_n13969), .B(new_n13968), .Y(new_n13970));
  NOR2xp33_ASAP7_75t_L      g13714(.A(new_n1043), .B(new_n10400), .Y(new_n13971));
  AOI221xp5_ASAP7_75t_L     g13715(.A1(new_n9102), .A2(\b[16] ), .B1(new_n10398), .B2(\b[14] ), .C(new_n13971), .Y(new_n13972));
  O2A1O1Ixp33_ASAP7_75t_L   g13716(.A1(new_n9104), .A2(new_n1161), .B(new_n13972), .C(new_n9099), .Y(new_n13973));
  O2A1O1Ixp33_ASAP7_75t_L   g13717(.A1(new_n9104), .A2(new_n1161), .B(new_n13972), .C(\a[53] ), .Y(new_n13974));
  INVx1_ASAP7_75t_L         g13718(.A(new_n13974), .Y(new_n13975));
  O2A1O1Ixp33_ASAP7_75t_L   g13719(.A1(new_n13973), .A2(new_n9099), .B(new_n13975), .C(new_n13970), .Y(new_n13976));
  INVx1_ASAP7_75t_L         g13720(.A(new_n13973), .Y(new_n13977));
  A2O1A1Ixp33_ASAP7_75t_L   g13721(.A1(\a[53] ), .A2(new_n13977), .B(new_n13974), .C(new_n13970), .Y(new_n13978));
  OAI21xp33_ASAP7_75t_L     g13722(.A1(new_n13970), .A2(new_n13976), .B(new_n13978), .Y(new_n13979));
  MAJIxp5_ASAP7_75t_L       g13723(.A(new_n13708), .B(new_n13712), .C(new_n13664), .Y(new_n13980));
  XNOR2x2_ASAP7_75t_L       g13724(.A(new_n13980), .B(new_n13979), .Y(new_n13981));
  NOR2xp33_ASAP7_75t_L      g13725(.A(new_n1458), .B(new_n10065), .Y(new_n13982));
  AOI221xp5_ASAP7_75t_L     g13726(.A1(new_n8175), .A2(\b[19] ), .B1(new_n8484), .B2(\b[17] ), .C(new_n13982), .Y(new_n13983));
  O2A1O1Ixp33_ASAP7_75t_L   g13727(.A1(new_n8176), .A2(new_n1628), .B(new_n13983), .C(new_n8172), .Y(new_n13984));
  O2A1O1Ixp33_ASAP7_75t_L   g13728(.A1(new_n8176), .A2(new_n1628), .B(new_n13983), .C(\a[50] ), .Y(new_n13985));
  INVx1_ASAP7_75t_L         g13729(.A(new_n13985), .Y(new_n13986));
  O2A1O1Ixp33_ASAP7_75t_L   g13730(.A1(new_n13984), .A2(new_n8172), .B(new_n13986), .C(new_n13981), .Y(new_n13987));
  INVx1_ASAP7_75t_L         g13731(.A(new_n13984), .Y(new_n13988));
  A2O1A1Ixp33_ASAP7_75t_L   g13732(.A1(\a[50] ), .A2(new_n13988), .B(new_n13985), .C(new_n13981), .Y(new_n13989));
  MAJIxp5_ASAP7_75t_L       g13733(.A(new_n13713), .B(new_n13715), .C(new_n13731), .Y(new_n13990));
  OA211x2_ASAP7_75t_L       g13734(.A1(new_n13981), .A2(new_n13987), .B(new_n13989), .C(new_n13990), .Y(new_n13991));
  O2A1O1Ixp33_ASAP7_75t_L   g13735(.A1(new_n13981), .A2(new_n13987), .B(new_n13989), .C(new_n13990), .Y(new_n13992));
  NOR2xp33_ASAP7_75t_L      g13736(.A(new_n13992), .B(new_n13991), .Y(new_n13993));
  NOR2xp33_ASAP7_75t_L      g13737(.A(new_n1895), .B(new_n7312), .Y(new_n13994));
  AOI221xp5_ASAP7_75t_L     g13738(.A1(\b[20] ), .A2(new_n7609), .B1(\b[22] ), .B2(new_n7334), .C(new_n13994), .Y(new_n13995));
  O2A1O1Ixp33_ASAP7_75t_L   g13739(.A1(new_n7321), .A2(new_n2522), .B(new_n13995), .C(new_n7316), .Y(new_n13996));
  INVx1_ASAP7_75t_L         g13740(.A(new_n13996), .Y(new_n13997));
  O2A1O1Ixp33_ASAP7_75t_L   g13741(.A1(new_n7321), .A2(new_n2522), .B(new_n13995), .C(\a[47] ), .Y(new_n13998));
  A2O1A1Ixp33_ASAP7_75t_L   g13742(.A1(\a[47] ), .A2(new_n13997), .B(new_n13998), .C(new_n13993), .Y(new_n13999));
  A2O1A1Ixp33_ASAP7_75t_L   g13743(.A1(new_n13997), .A2(\a[47] ), .B(new_n13998), .C(new_n13999), .Y(new_n14000));
  INVx1_ASAP7_75t_L         g13744(.A(new_n14000), .Y(new_n14001));
  A2O1A1Ixp33_ASAP7_75t_L   g13745(.A1(new_n13999), .A2(new_n13993), .B(new_n14001), .C(new_n13915), .Y(new_n14002));
  AOI21xp33_ASAP7_75t_L     g13746(.A1(new_n13997), .A2(\a[47] ), .B(new_n13998), .Y(new_n14003));
  NAND2xp33_ASAP7_75t_L     g13747(.A(new_n14003), .B(new_n13993), .Y(new_n14004));
  INVx1_ASAP7_75t_L         g13748(.A(new_n14004), .Y(new_n14005));
  A2O1A1O1Ixp25_ASAP7_75t_L g13749(.A1(new_n13997), .A2(\a[47] ), .B(new_n13998), .C(new_n13999), .D(new_n14005), .Y(new_n14006));
  NOR2xp33_ASAP7_75t_L      g13750(.A(new_n14006), .B(new_n13915), .Y(new_n14007));
  NOR2xp33_ASAP7_75t_L      g13751(.A(new_n2188), .B(new_n6741), .Y(new_n14008));
  AOI221xp5_ASAP7_75t_L     g13752(.A1(\b[25] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[24] ), .C(new_n14008), .Y(new_n14009));
  O2A1O1Ixp33_ASAP7_75t_L   g13753(.A1(new_n6443), .A2(new_n2385), .B(new_n14009), .C(new_n6439), .Y(new_n14010));
  O2A1O1Ixp33_ASAP7_75t_L   g13754(.A1(new_n6443), .A2(new_n2385), .B(new_n14009), .C(\a[44] ), .Y(new_n14011));
  INVx1_ASAP7_75t_L         g13755(.A(new_n14011), .Y(new_n14012));
  OA21x2_ASAP7_75t_L        g13756(.A1(new_n6439), .A2(new_n14010), .B(new_n14012), .Y(new_n14013));
  A2O1A1Ixp33_ASAP7_75t_L   g13757(.A1(new_n14002), .A2(new_n13915), .B(new_n14007), .C(new_n14013), .Y(new_n14014));
  A2O1A1Ixp33_ASAP7_75t_L   g13758(.A1(new_n13999), .A2(new_n13993), .B(new_n14001), .C(new_n13914), .Y(new_n14015));
  A2O1A1Ixp33_ASAP7_75t_L   g13759(.A1(new_n13735), .A2(new_n13739), .B(new_n13734), .C(new_n14006), .Y(new_n14016));
  INVx1_ASAP7_75t_L         g13760(.A(new_n14013), .Y(new_n14017));
  NAND3xp33_ASAP7_75t_L     g13761(.A(new_n14015), .B(new_n14016), .C(new_n14017), .Y(new_n14018));
  OAI21xp33_ASAP7_75t_L     g13762(.A1(new_n13740), .A2(new_n13742), .B(new_n13744), .Y(new_n14019));
  AOI21xp33_ASAP7_75t_L     g13763(.A1(new_n14019), .A2(new_n13751), .B(new_n13745), .Y(new_n14020));
  NAND3xp33_ASAP7_75t_L     g13764(.A(new_n14014), .B(new_n14018), .C(new_n14020), .Y(new_n14021));
  A2O1A1Ixp33_ASAP7_75t_L   g13765(.A1(new_n14002), .A2(new_n13915), .B(new_n14007), .C(new_n14017), .Y(new_n14022));
  O2A1O1Ixp33_ASAP7_75t_L   g13766(.A1(new_n13730), .A2(new_n13738), .B(new_n13733), .C(new_n14006), .Y(new_n14023));
  O2A1O1Ixp33_ASAP7_75t_L   g13767(.A1(new_n14006), .A2(new_n14023), .B(new_n14016), .C(new_n14017), .Y(new_n14024));
  INVx1_ASAP7_75t_L         g13768(.A(new_n14020), .Y(new_n14025));
  A2O1A1Ixp33_ASAP7_75t_L   g13769(.A1(new_n14022), .A2(new_n14017), .B(new_n14024), .C(new_n14025), .Y(new_n14026));
  NAND2xp33_ASAP7_75t_L     g13770(.A(\b[27] ), .B(new_n5623), .Y(new_n14027));
  OAI221xp5_ASAP7_75t_L     g13771(.A1(new_n5641), .A2(new_n3079), .B1(new_n2703), .B2(new_n5925), .C(new_n14027), .Y(new_n14028));
  A2O1A1Ixp33_ASAP7_75t_L   g13772(.A1(new_n3085), .A2(new_n5637), .B(new_n14028), .C(\a[41] ), .Y(new_n14029));
  NAND2xp33_ASAP7_75t_L     g13773(.A(\a[41] ), .B(new_n14029), .Y(new_n14030));
  A2O1A1Ixp33_ASAP7_75t_L   g13774(.A1(new_n3085), .A2(new_n5637), .B(new_n14028), .C(new_n5626), .Y(new_n14031));
  NAND4xp25_ASAP7_75t_L     g13775(.A(new_n14026), .B(new_n14030), .C(new_n14031), .D(new_n14021), .Y(new_n14032));
  AND3x1_ASAP7_75t_L        g13776(.A(new_n14014), .B(new_n14020), .C(new_n14018), .Y(new_n14033));
  O2A1O1Ixp33_ASAP7_75t_L   g13777(.A1(new_n13914), .A2(new_n14023), .B(new_n14015), .C(new_n14013), .Y(new_n14034));
  O2A1O1Ixp33_ASAP7_75t_L   g13778(.A1(new_n14013), .A2(new_n14034), .B(new_n14014), .C(new_n14020), .Y(new_n14035));
  NAND2xp33_ASAP7_75t_L     g13779(.A(new_n14031), .B(new_n14030), .Y(new_n14036));
  OAI21xp33_ASAP7_75t_L     g13780(.A1(new_n14033), .A2(new_n14035), .B(new_n14036), .Y(new_n14037));
  AOI21xp33_ASAP7_75t_L     g13781(.A1(new_n13756), .A2(new_n13765), .B(new_n13764), .Y(new_n14038));
  NAND3xp33_ASAP7_75t_L     g13782(.A(new_n14037), .B(new_n14032), .C(new_n14038), .Y(new_n14039));
  NAND3xp33_ASAP7_75t_L     g13783(.A(new_n14026), .B(new_n14021), .C(new_n14036), .Y(new_n14040));
  NOR3xp33_ASAP7_75t_L      g13784(.A(new_n14035), .B(new_n14033), .C(new_n14036), .Y(new_n14041));
  INVx1_ASAP7_75t_L         g13785(.A(new_n14038), .Y(new_n14042));
  A2O1A1Ixp33_ASAP7_75t_L   g13786(.A1(new_n14040), .A2(new_n14036), .B(new_n14041), .C(new_n14042), .Y(new_n14043));
  OAI22xp33_ASAP7_75t_L     g13787(.A1(new_n5144), .A2(new_n3098), .B1(new_n3456), .B2(new_n4903), .Y(new_n14044));
  AOI221xp5_ASAP7_75t_L     g13788(.A1(new_n4917), .A2(\b[31] ), .B1(new_n4912), .B2(new_n4317), .C(new_n14044), .Y(new_n14045));
  XNOR2x2_ASAP7_75t_L       g13789(.A(new_n4906), .B(new_n14045), .Y(new_n14046));
  INVx1_ASAP7_75t_L         g13790(.A(new_n14046), .Y(new_n14047));
  AO21x2_ASAP7_75t_L        g13791(.A1(new_n14039), .A2(new_n14043), .B(new_n14047), .Y(new_n14048));
  NAND3xp33_ASAP7_75t_L     g13792(.A(new_n14043), .B(new_n14039), .C(new_n14047), .Y(new_n14049));
  AOI21xp33_ASAP7_75t_L     g13793(.A1(new_n14048), .A2(new_n14049), .B(new_n13913), .Y(new_n14050));
  NAND3xp33_ASAP7_75t_L     g13794(.A(new_n14048), .B(new_n13913), .C(new_n14049), .Y(new_n14051));
  INVx1_ASAP7_75t_L         g13795(.A(new_n14051), .Y(new_n14052));
  NOR3xp33_ASAP7_75t_L      g13796(.A(new_n14052), .B(new_n14050), .C(new_n13912), .Y(new_n14053));
  INVx1_ASAP7_75t_L         g13797(.A(new_n13912), .Y(new_n14054));
  INVx1_ASAP7_75t_L         g13798(.A(new_n14050), .Y(new_n14055));
  AOI21xp33_ASAP7_75t_L     g13799(.A1(new_n14055), .A2(new_n14051), .B(new_n14054), .Y(new_n14056));
  NOR2xp33_ASAP7_75t_L      g13800(.A(new_n14053), .B(new_n14056), .Y(new_n14057));
  OA21x2_ASAP7_75t_L        g13801(.A1(new_n13908), .A2(new_n13909), .B(new_n14057), .Y(new_n14058));
  NOR3xp33_ASAP7_75t_L      g13802(.A(new_n14057), .B(new_n13908), .C(new_n13909), .Y(new_n14059));
  NOR2xp33_ASAP7_75t_L      g13803(.A(new_n14059), .B(new_n14058), .Y(new_n14060));
  OAI22xp33_ASAP7_75t_L     g13804(.A1(new_n3133), .A2(new_n5311), .B1(new_n5570), .B2(new_n2925), .Y(new_n14061));
  AOI221xp5_ASAP7_75t_L     g13805(.A1(new_n2938), .A2(\b[40] ), .B1(new_n2932), .B2(new_n6651), .C(new_n14061), .Y(new_n14062));
  XNOR2x2_ASAP7_75t_L       g13806(.A(new_n2928), .B(new_n14062), .Y(new_n14063));
  INVx1_ASAP7_75t_L         g13807(.A(new_n14063), .Y(new_n14064));
  O2A1O1Ixp33_ASAP7_75t_L   g13808(.A1(new_n13796), .A2(new_n13798), .B(new_n13793), .C(new_n14063), .Y(new_n14065));
  INVx1_ASAP7_75t_L         g13809(.A(new_n14065), .Y(new_n14066));
  O2A1O1Ixp33_ASAP7_75t_L   g13810(.A1(new_n13796), .A2(new_n13798), .B(new_n13793), .C(new_n14064), .Y(new_n14067));
  A2O1A1Ixp33_ASAP7_75t_L   g13811(.A1(new_n14066), .A2(new_n14064), .B(new_n14067), .C(new_n14060), .Y(new_n14068));
  INVx1_ASAP7_75t_L         g13812(.A(new_n14067), .Y(new_n14069));
  O2A1O1Ixp33_ASAP7_75t_L   g13813(.A1(new_n14063), .A2(new_n14065), .B(new_n14069), .C(new_n14060), .Y(new_n14070));
  AOI21xp33_ASAP7_75t_L     g13814(.A1(new_n14068), .A2(new_n14060), .B(new_n14070), .Y(new_n14071));
  OAI22xp33_ASAP7_75t_L     g13815(.A1(new_n2572), .A2(new_n6110), .B1(new_n6378), .B2(new_n2410), .Y(new_n14072));
  AOI221xp5_ASAP7_75t_L     g13816(.A1(new_n2423), .A2(\b[43] ), .B1(new_n2417), .B2(new_n6682), .C(new_n14072), .Y(new_n14073));
  XNOR2x2_ASAP7_75t_L       g13817(.A(new_n2413), .B(new_n14073), .Y(new_n14074));
  INVx1_ASAP7_75t_L         g13818(.A(new_n14074), .Y(new_n14075));
  AOI211xp5_ASAP7_75t_L     g13819(.A1(new_n13800), .A2(new_n13655), .B(new_n14075), .C(new_n13653), .Y(new_n14076));
  INVx1_ASAP7_75t_L         g13820(.A(new_n14076), .Y(new_n14077));
  A2O1A1Ixp33_ASAP7_75t_L   g13821(.A1(new_n13800), .A2(new_n13655), .B(new_n13653), .C(new_n14075), .Y(new_n14078));
  NAND2xp33_ASAP7_75t_L     g13822(.A(new_n14078), .B(new_n14077), .Y(new_n14079));
  OR2x4_ASAP7_75t_L         g13823(.A(new_n14059), .B(new_n14058), .Y(new_n14080));
  O2A1O1Ixp33_ASAP7_75t_L   g13824(.A1(new_n14063), .A2(new_n14065), .B(new_n14069), .C(new_n14080), .Y(new_n14081));
  A2O1A1Ixp33_ASAP7_75t_L   g13825(.A1(new_n14064), .A2(new_n14066), .B(new_n14067), .C(new_n14080), .Y(new_n14082));
  O2A1O1Ixp33_ASAP7_75t_L   g13826(.A1(new_n14080), .A2(new_n14081), .B(new_n14082), .C(new_n14079), .Y(new_n14083));
  NAND3xp33_ASAP7_75t_L     g13827(.A(new_n14071), .B(new_n14078), .C(new_n14077), .Y(new_n14084));
  OAI22xp33_ASAP7_75t_L     g13828(.A1(new_n2089), .A2(new_n6944), .B1(new_n7249), .B2(new_n1962), .Y(new_n14085));
  AOI221xp5_ASAP7_75t_L     g13829(.A1(new_n1955), .A2(\b[46] ), .B1(new_n1964), .B2(new_n7278), .C(new_n14085), .Y(new_n14086));
  XNOR2x2_ASAP7_75t_L       g13830(.A(new_n1952), .B(new_n14086), .Y(new_n14087));
  O2A1O1Ixp33_ASAP7_75t_L   g13831(.A1(new_n13647), .A2(new_n13805), .B(new_n13644), .C(new_n14087), .Y(new_n14088));
  INVx1_ASAP7_75t_L         g13832(.A(new_n14087), .Y(new_n14089));
  A2O1A1O1Ixp25_ASAP7_75t_L g13833(.A1(new_n13655), .A2(new_n13801), .B(new_n13804), .C(new_n13646), .D(new_n13645), .Y(new_n14090));
  NAND2xp33_ASAP7_75t_L     g13834(.A(new_n14089), .B(new_n14090), .Y(new_n14091));
  A2O1A1Ixp33_ASAP7_75t_L   g13835(.A1(new_n13818), .A2(new_n13644), .B(new_n14088), .C(new_n14091), .Y(new_n14092));
  O2A1O1Ixp33_ASAP7_75t_L   g13836(.A1(new_n14071), .A2(new_n14083), .B(new_n14084), .C(new_n14092), .Y(new_n14093));
  INVx1_ASAP7_75t_L         g13837(.A(new_n14078), .Y(new_n14094));
  OAI21xp33_ASAP7_75t_L     g13838(.A1(new_n14080), .A2(new_n14081), .B(new_n14082), .Y(new_n14095));
  OAI21xp33_ASAP7_75t_L     g13839(.A1(new_n14076), .A2(new_n14094), .B(new_n14095), .Y(new_n14096));
  NAND2xp33_ASAP7_75t_L     g13840(.A(new_n14084), .B(new_n14096), .Y(new_n14097));
  O2A1O1Ixp33_ASAP7_75t_L   g13841(.A1(new_n14090), .A2(new_n14088), .B(new_n14091), .C(new_n14097), .Y(new_n14098));
  NOR2xp33_ASAP7_75t_L      g13842(.A(new_n14093), .B(new_n14098), .Y(new_n14099));
  NAND3xp33_ASAP7_75t_L     g13843(.A(new_n14099), .B(new_n13904), .C(new_n13902), .Y(new_n14100));
  INVx1_ASAP7_75t_L         g13844(.A(new_n13902), .Y(new_n14101));
  OR2x4_ASAP7_75t_L         g13845(.A(new_n14093), .B(new_n14098), .Y(new_n14102));
  OAI21xp33_ASAP7_75t_L     g13846(.A1(new_n14101), .A2(new_n13903), .B(new_n14102), .Y(new_n14103));
  NAND2xp33_ASAP7_75t_L     g13847(.A(new_n14100), .B(new_n14103), .Y(new_n14104));
  INVx1_ASAP7_75t_L         g13848(.A(new_n13627), .Y(new_n14105));
  NAND2xp33_ASAP7_75t_L     g13849(.A(new_n13818), .B(new_n13819), .Y(new_n14106));
  NAND2xp33_ASAP7_75t_L     g13850(.A(new_n13635), .B(new_n14106), .Y(new_n14107));
  OAI22xp33_ASAP7_75t_L     g13851(.A1(new_n1285), .A2(new_n8755), .B1(new_n8779), .B2(new_n2118), .Y(new_n14108));
  AOI221xp5_ASAP7_75t_L     g13852(.A1(new_n1209), .A2(\b[52] ), .B1(new_n1216), .B2(new_n9367), .C(new_n14108), .Y(new_n14109));
  XNOR2x2_ASAP7_75t_L       g13853(.A(new_n1206), .B(new_n14109), .Y(new_n14110));
  A2O1A1O1Ixp25_ASAP7_75t_L g13854(.A1(new_n13820), .A2(new_n14107), .B(new_n13625), .C(new_n14105), .D(new_n14110), .Y(new_n14111));
  INVx1_ASAP7_75t_L         g13855(.A(new_n14111), .Y(new_n14112));
  A2O1A1Ixp33_ASAP7_75t_L   g13856(.A1(new_n14107), .A2(new_n13820), .B(new_n13625), .C(new_n14105), .Y(new_n14113));
  NOR2xp33_ASAP7_75t_L      g13857(.A(new_n14110), .B(new_n14113), .Y(new_n14114));
  O2A1O1Ixp33_ASAP7_75t_L   g13858(.A1(new_n13627), .A2(new_n13812), .B(new_n14112), .C(new_n14114), .Y(new_n14115));
  NAND2xp33_ASAP7_75t_L     g13859(.A(new_n14115), .B(new_n14104), .Y(new_n14116));
  AND2x2_ASAP7_75t_L        g13860(.A(new_n14100), .B(new_n14103), .Y(new_n14117));
  A2O1A1Ixp33_ASAP7_75t_L   g13861(.A1(new_n14113), .A2(new_n14112), .B(new_n14114), .C(new_n14117), .Y(new_n14118));
  NAND2xp33_ASAP7_75t_L     g13862(.A(new_n14116), .B(new_n14118), .Y(new_n14119));
  NOR3xp33_ASAP7_75t_L      g13863(.A(new_n14119), .B(new_n13895), .C(new_n13894), .Y(new_n14120));
  INVx1_ASAP7_75t_L         g13864(.A(new_n13894), .Y(new_n14121));
  INVx1_ASAP7_75t_L         g13865(.A(new_n13895), .Y(new_n14122));
  AOI22xp33_ASAP7_75t_L     g13866(.A1(new_n14116), .A2(new_n14118), .B1(new_n14122), .B2(new_n14121), .Y(new_n14123));
  NOR2xp33_ASAP7_75t_L      g13867(.A(new_n14120), .B(new_n14123), .Y(new_n14124));
  OAI22xp33_ASAP7_75t_L     g13868(.A1(new_n1550), .A2(new_n10978), .B1(new_n10332), .B2(new_n712), .Y(new_n14125));
  AOI221xp5_ASAP7_75t_L     g13869(.A1(new_n640), .A2(\b[58] ), .B1(new_n718), .B2(new_n11314), .C(new_n14125), .Y(new_n14126));
  XNOR2x2_ASAP7_75t_L       g13870(.A(\a[11] ), .B(new_n14126), .Y(new_n14127));
  INVx1_ASAP7_75t_L         g13871(.A(new_n14127), .Y(new_n14128));
  O2A1O1Ixp33_ASAP7_75t_L   g13872(.A1(new_n13834), .A2(new_n13824), .B(new_n13832), .C(new_n14128), .Y(new_n14129));
  O2A1O1Ixp33_ASAP7_75t_L   g13873(.A1(new_n13834), .A2(new_n13824), .B(new_n13832), .C(new_n14127), .Y(new_n14130));
  INVx1_ASAP7_75t_L         g13874(.A(new_n14130), .Y(new_n14131));
  O2A1O1Ixp33_ASAP7_75t_L   g13875(.A1(new_n14128), .A2(new_n14129), .B(new_n14131), .C(new_n14124), .Y(new_n14132));
  INVx1_ASAP7_75t_L         g13876(.A(new_n14129), .Y(new_n14133));
  A2O1A1Ixp33_ASAP7_75t_L   g13877(.A1(new_n14127), .A2(new_n14133), .B(new_n14130), .C(new_n14124), .Y(new_n14134));
  O2A1O1Ixp33_ASAP7_75t_L   g13878(.A1(new_n14124), .A2(new_n14132), .B(new_n14134), .C(new_n13888), .Y(new_n14135));
  OAI21xp33_ASAP7_75t_L     g13879(.A1(new_n14124), .A2(new_n14132), .B(new_n14134), .Y(new_n14136));
  NAND2xp33_ASAP7_75t_L     g13880(.A(new_n13888), .B(new_n14136), .Y(new_n14137));
  A2O1A1Ixp33_ASAP7_75t_L   g13881(.A1(new_n13846), .A2(new_n13838), .B(new_n13854), .C(new_n13880), .Y(new_n14138));
  A2O1A1Ixp33_ASAP7_75t_L   g13882(.A1(new_n13846), .A2(new_n13838), .B(new_n13854), .C(new_n13879), .Y(new_n14139));
  INVx1_ASAP7_75t_L         g13883(.A(new_n14139), .Y(new_n14140));
  O2A1O1Ixp33_ASAP7_75t_L   g13884(.A1(new_n13877), .A2(new_n13878), .B(new_n14138), .C(new_n14140), .Y(new_n14141));
  O2A1O1Ixp33_ASAP7_75t_L   g13885(.A1(new_n13888), .A2(new_n14135), .B(new_n14137), .C(new_n14141), .Y(new_n14142));
  A2O1A1Ixp33_ASAP7_75t_L   g13886(.A1(new_n13881), .A2(new_n13835), .B(new_n13609), .C(new_n13886), .Y(new_n14143));
  AOI21xp33_ASAP7_75t_L     g13887(.A1(new_n13881), .A2(new_n13835), .B(new_n13609), .Y(new_n14144));
  NAND2xp33_ASAP7_75t_L     g13888(.A(new_n13884), .B(new_n14144), .Y(new_n14145));
  A2O1A1Ixp33_ASAP7_75t_L   g13889(.A1(new_n14145), .A2(new_n14143), .B(new_n14135), .C(new_n14137), .Y(new_n14146));
  O2A1O1Ixp33_ASAP7_75t_L   g13890(.A1(new_n13877), .A2(new_n13878), .B(new_n14138), .C(new_n14146), .Y(new_n14147));
  O2A1O1Ixp33_ASAP7_75t_L   g13891(.A1(new_n13880), .A2(new_n13873), .B(new_n14147), .C(new_n14142), .Y(new_n14148));
  A2O1A1Ixp33_ASAP7_75t_L   g13892(.A1(new_n13599), .A2(new_n13861), .B(new_n13872), .C(new_n14148), .Y(new_n14149));
  INVx1_ASAP7_75t_L         g13893(.A(new_n14149), .Y(new_n14150));
  A2O1A1Ixp33_ASAP7_75t_L   g13894(.A1(new_n13591), .A2(new_n13588), .B(new_n13587), .C(new_n13867), .Y(new_n14151));
  A2O1A1Ixp33_ASAP7_75t_L   g13895(.A1(new_n13880), .A2(new_n14138), .B(new_n14140), .C(new_n14146), .Y(new_n14152));
  NAND2xp33_ASAP7_75t_L     g13896(.A(new_n14143), .B(new_n14145), .Y(new_n14153));
  O2A1O1Ixp33_ASAP7_75t_L   g13897(.A1(new_n14124), .A2(new_n14132), .B(new_n14134), .C(new_n14153), .Y(new_n14154));
  INVx1_ASAP7_75t_L         g13898(.A(new_n13885), .Y(new_n14155));
  O2A1O1Ixp33_ASAP7_75t_L   g13899(.A1(new_n14144), .A2(new_n14155), .B(new_n14145), .C(new_n14136), .Y(new_n14156));
  NOR2xp33_ASAP7_75t_L      g13900(.A(new_n14156), .B(new_n14154), .Y(new_n14157));
  NAND2xp33_ASAP7_75t_L     g13901(.A(new_n13880), .B(new_n13873), .Y(new_n14158));
  NAND2xp33_ASAP7_75t_L     g13902(.A(new_n14158), .B(new_n14157), .Y(new_n14159));
  O2A1O1Ixp33_ASAP7_75t_L   g13903(.A1(new_n14140), .A2(new_n14159), .B(new_n14152), .C(new_n13871), .Y(new_n14160));
  INVx1_ASAP7_75t_L         g13904(.A(new_n13871), .Y(new_n14161));
  AOI211xp5_ASAP7_75t_L     g13905(.A1(new_n13880), .A2(new_n14138), .B(new_n14140), .C(new_n14146), .Y(new_n14162));
  NOR3xp33_ASAP7_75t_L      g13906(.A(new_n14162), .B(new_n14142), .C(new_n14161), .Y(new_n14163));
  NOR2xp33_ASAP7_75t_L      g13907(.A(new_n14160), .B(new_n14163), .Y(new_n14164));
  A2O1A1O1Ixp25_ASAP7_75t_L g13908(.A1(new_n13864), .A2(new_n13863), .B(new_n13865), .C(new_n14151), .D(new_n14164), .Y(new_n14165));
  A2O1A1Ixp33_ASAP7_75t_L   g13909(.A1(new_n13864), .A2(new_n13863), .B(new_n13865), .C(new_n14151), .Y(new_n14166));
  NOR2xp33_ASAP7_75t_L      g13910(.A(new_n14163), .B(new_n14166), .Y(new_n14167));
  O2A1O1Ixp33_ASAP7_75t_L   g13911(.A1(new_n14150), .A2(new_n13871), .B(new_n14167), .C(new_n14165), .Y(\f[67] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13912(.A1(new_n14139), .A2(new_n13879), .B(new_n14157), .C(new_n14138), .Y(new_n14169));
  NOR2xp33_ASAP7_75t_L      g13913(.A(new_n12956), .B(new_n375), .Y(new_n14170));
  A2O1A1Ixp33_ASAP7_75t_L   g13914(.A1(new_n12986), .A2(new_n359), .B(new_n14170), .C(\a[5] ), .Y(new_n14171));
  A2O1A1Ixp33_ASAP7_75t_L   g13915(.A1(new_n12606), .A2(new_n12954), .B(new_n12956), .C(new_n12603), .Y(new_n14172));
  A2O1A1O1Ixp25_ASAP7_75t_L g13916(.A1(new_n359), .A2(new_n14172), .B(new_n13874), .C(\b[63] ), .D(new_n346), .Y(new_n14173));
  A2O1A1O1Ixp25_ASAP7_75t_L g13917(.A1(new_n12986), .A2(new_n359), .B(new_n14170), .C(new_n14171), .D(new_n14173), .Y(new_n14174));
  INVx1_ASAP7_75t_L         g13918(.A(new_n14174), .Y(new_n14175));
  A2O1A1Ixp33_ASAP7_75t_L   g13919(.A1(new_n14153), .A2(new_n14136), .B(new_n14155), .C(new_n14175), .Y(new_n14176));
  INVx1_ASAP7_75t_L         g13920(.A(new_n14176), .Y(new_n14177));
  A2O1A1Ixp33_ASAP7_75t_L   g13921(.A1(new_n14153), .A2(new_n14136), .B(new_n14155), .C(new_n14174), .Y(new_n14178));
  A2O1A1Ixp33_ASAP7_75t_L   g13922(.A1(new_n13231), .A2(new_n13018), .B(new_n13230), .C(new_n13517), .Y(new_n14179));
  O2A1O1Ixp33_ASAP7_75t_L   g13923(.A1(new_n13225), .A2(new_n13230), .B(new_n14179), .C(new_n13525), .Y(new_n14180));
  O2A1O1Ixp33_ASAP7_75t_L   g13924(.A1(new_n14180), .A2(new_n13521), .B(new_n13528), .C(new_n13830), .Y(new_n14181));
  A2O1A1Ixp33_ASAP7_75t_L   g13925(.A1(new_n13522), .A2(new_n13294), .B(new_n13825), .C(new_n13830), .Y(new_n14182));
  O2A1O1Ixp33_ASAP7_75t_L   g13926(.A1(new_n13830), .A2(new_n14181), .B(new_n14182), .C(new_n13824), .Y(new_n14183));
  O2A1O1Ixp33_ASAP7_75t_L   g13927(.A1(new_n14181), .A2(new_n14183), .B(new_n14127), .C(new_n14132), .Y(new_n14184));
  INVx1_ASAP7_75t_L         g13928(.A(new_n14184), .Y(new_n14185));
  OAI22xp33_ASAP7_75t_L     g13929(.A1(new_n513), .A2(new_n12258), .B1(new_n11626), .B2(new_n506), .Y(new_n14186));
  AOI221xp5_ASAP7_75t_L     g13930(.A1(new_n475), .A2(\b[62] ), .B1(new_n483), .B2(new_n13559), .C(new_n14186), .Y(new_n14187));
  XNOR2x2_ASAP7_75t_L       g13931(.A(new_n466), .B(new_n14187), .Y(new_n14188));
  OAI22xp33_ASAP7_75t_L     g13932(.A1(new_n980), .A2(new_n9709), .B1(new_n10309), .B2(new_n864), .Y(new_n14189));
  AOI221xp5_ASAP7_75t_L     g13933(.A1(new_n886), .A2(\b[56] ), .B1(new_n873), .B2(new_n11579), .C(new_n14189), .Y(new_n14190));
  XNOR2x2_ASAP7_75t_L       g13934(.A(\a[14] ), .B(new_n14190), .Y(new_n14191));
  INVx1_ASAP7_75t_L         g13935(.A(new_n14191), .Y(new_n14192));
  A2O1A1O1Ixp25_ASAP7_75t_L g13936(.A1(new_n14103), .A2(new_n14100), .B(new_n14115), .C(new_n14112), .D(new_n14192), .Y(new_n14193));
  INVx1_ASAP7_75t_L         g13937(.A(new_n14193), .Y(new_n14194));
  A2O1A1O1Ixp25_ASAP7_75t_L g13938(.A1(new_n14103), .A2(new_n14100), .B(new_n14115), .C(new_n14112), .D(new_n14191), .Y(new_n14195));
  OAI22xp33_ASAP7_75t_L     g13939(.A1(new_n1285), .A2(new_n8779), .B1(new_n9355), .B2(new_n2118), .Y(new_n14196));
  AOI221xp5_ASAP7_75t_L     g13940(.A1(new_n1209), .A2(\b[53] ), .B1(new_n1216), .B2(new_n9690), .C(new_n14196), .Y(new_n14197));
  XNOR2x2_ASAP7_75t_L       g13941(.A(new_n1206), .B(new_n14197), .Y(new_n14198));
  O2A1O1Ixp33_ASAP7_75t_L   g13942(.A1(new_n14101), .A2(new_n14099), .B(new_n13904), .C(new_n14198), .Y(new_n14199));
  INVx1_ASAP7_75t_L         g13943(.A(new_n14199), .Y(new_n14200));
  O2A1O1Ixp33_ASAP7_75t_L   g13944(.A1(new_n14093), .A2(new_n14098), .B(new_n13902), .C(new_n13903), .Y(new_n14201));
  NAND2xp33_ASAP7_75t_L     g13945(.A(new_n14198), .B(new_n14201), .Y(new_n14202));
  NAND2xp33_ASAP7_75t_L     g13946(.A(new_n14202), .B(new_n14200), .Y(new_n14203));
  NOR2xp33_ASAP7_75t_L      g13947(.A(new_n8427), .B(new_n1517), .Y(new_n14204));
  AOI221xp5_ASAP7_75t_L     g13948(.A1(\b[48] ), .A2(new_n1659), .B1(\b[50] ), .B2(new_n1511), .C(new_n14204), .Y(new_n14205));
  INVx1_ASAP7_75t_L         g13949(.A(new_n14205), .Y(new_n14206));
  A2O1A1Ixp33_ASAP7_75t_L   g13950(.A1(new_n8763), .A2(new_n1513), .B(new_n14206), .C(\a[20] ), .Y(new_n14207));
  O2A1O1Ixp33_ASAP7_75t_L   g13951(.A1(new_n1521), .A2(new_n8764), .B(new_n14205), .C(\a[20] ), .Y(new_n14208));
  AO21x2_ASAP7_75t_L        g13952(.A1(\a[20] ), .A2(new_n14207), .B(new_n14208), .Y(new_n14209));
  A2O1A1Ixp33_ASAP7_75t_L   g13953(.A1(new_n14097), .A2(new_n14092), .B(new_n14088), .C(new_n14209), .Y(new_n14210));
  A2O1A1Ixp33_ASAP7_75t_L   g13954(.A1(new_n13641), .A2(new_n13639), .B(new_n13806), .C(new_n14089), .Y(new_n14211));
  O2A1O1Ixp33_ASAP7_75t_L   g13955(.A1(new_n13647), .A2(new_n13805), .B(new_n13644), .C(new_n14089), .Y(new_n14212));
  A2O1A1Ixp33_ASAP7_75t_L   g13956(.A1(new_n14089), .A2(new_n14211), .B(new_n14212), .C(new_n14097), .Y(new_n14213));
  O2A1O1Ixp33_ASAP7_75t_L   g13957(.A1(new_n14090), .A2(new_n14087), .B(new_n14213), .C(new_n14209), .Y(new_n14214));
  A2O1A1O1Ixp25_ASAP7_75t_L g13958(.A1(new_n14207), .A2(\a[20] ), .B(new_n14208), .C(new_n14210), .D(new_n14214), .Y(new_n14215));
  NOR2xp33_ASAP7_75t_L      g13959(.A(new_n7270), .B(new_n1962), .Y(new_n14216));
  AOI221xp5_ASAP7_75t_L     g13960(.A1(new_n1955), .A2(\b[47] ), .B1(new_n2093), .B2(\b[45] ), .C(new_n14216), .Y(new_n14217));
  O2A1O1Ixp33_ASAP7_75t_L   g13961(.A1(new_n1956), .A2(new_n7560), .B(new_n14217), .C(new_n1952), .Y(new_n14218));
  INVx1_ASAP7_75t_L         g13962(.A(new_n14218), .Y(new_n14219));
  O2A1O1Ixp33_ASAP7_75t_L   g13963(.A1(new_n1956), .A2(new_n7560), .B(new_n14217), .C(\a[23] ), .Y(new_n14220));
  AOI21xp33_ASAP7_75t_L     g13964(.A1(new_n14219), .A2(\a[23] ), .B(new_n14220), .Y(new_n14221));
  A2O1A1O1Ixp25_ASAP7_75t_L g13965(.A1(new_n14068), .A2(new_n14060), .B(new_n14070), .C(new_n14077), .D(new_n14094), .Y(new_n14222));
  NAND2xp33_ASAP7_75t_L     g13966(.A(new_n14221), .B(new_n14222), .Y(new_n14223));
  INVx1_ASAP7_75t_L         g13967(.A(new_n14221), .Y(new_n14224));
  A2O1A1Ixp33_ASAP7_75t_L   g13968(.A1(new_n14095), .A2(new_n14077), .B(new_n14094), .C(new_n14224), .Y(new_n14225));
  NAND2xp33_ASAP7_75t_L     g13969(.A(new_n14225), .B(new_n14223), .Y(new_n14226));
  NOR2xp33_ASAP7_75t_L      g13970(.A(new_n332), .B(new_n13030), .Y(new_n14227));
  INVx1_ASAP7_75t_L         g13971(.A(new_n14227), .Y(new_n14228));
  O2A1O1Ixp33_ASAP7_75t_L   g13972(.A1(new_n384), .A2(new_n12672), .B(new_n14228), .C(new_n257), .Y(new_n14229));
  NOR2xp33_ASAP7_75t_L      g13973(.A(new_n257), .B(new_n14229), .Y(new_n14230));
  O2A1O1Ixp33_ASAP7_75t_L   g13974(.A1(new_n384), .A2(new_n12672), .B(new_n14228), .C(\a[2] ), .Y(new_n14231));
  NOR2xp33_ASAP7_75t_L      g13975(.A(new_n448), .B(new_n12318), .Y(new_n14232));
  AOI221xp5_ASAP7_75t_L     g13976(.A1(new_n11995), .A2(\b[8] ), .B1(new_n13314), .B2(\b[6] ), .C(new_n14232), .Y(new_n14233));
  INVx1_ASAP7_75t_L         g13977(.A(new_n14233), .Y(new_n14234));
  A2O1A1Ixp33_ASAP7_75t_L   g13978(.A1(new_n1684), .A2(new_n11997), .B(new_n14234), .C(\a[62] ), .Y(new_n14235));
  O2A1O1Ixp33_ASAP7_75t_L   g13979(.A1(new_n11998), .A2(new_n540), .B(new_n14233), .C(\a[62] ), .Y(new_n14236));
  INVx1_ASAP7_75t_L         g13980(.A(new_n14229), .Y(new_n14237));
  A2O1A1O1Ixp25_ASAP7_75t_L g13981(.A1(new_n13028), .A2(\b[5] ), .B(new_n14227), .C(new_n14237), .D(new_n14230), .Y(new_n14238));
  INVx1_ASAP7_75t_L         g13982(.A(new_n14238), .Y(new_n14239));
  A2O1A1Ixp33_ASAP7_75t_L   g13983(.A1(new_n14235), .A2(\a[62] ), .B(new_n14236), .C(new_n14239), .Y(new_n14240));
  O2A1O1Ixp33_ASAP7_75t_L   g13984(.A1(new_n11998), .A2(new_n540), .B(new_n14233), .C(new_n11987), .Y(new_n14241));
  INVx1_ASAP7_75t_L         g13985(.A(new_n14236), .Y(new_n14242));
  O2A1O1Ixp33_ASAP7_75t_L   g13986(.A1(new_n11987), .A2(new_n14241), .B(new_n14242), .C(new_n14239), .Y(new_n14243));
  O2A1O1Ixp33_ASAP7_75t_L   g13987(.A1(new_n14230), .A2(new_n14231), .B(new_n14240), .C(new_n14243), .Y(new_n14244));
  A2O1A1O1Ixp25_ASAP7_75t_L g13988(.A1(new_n13028), .A2(\b[4] ), .B(new_n13921), .C(\a[2] ), .D(new_n13934), .Y(new_n14245));
  NAND2xp33_ASAP7_75t_L     g13989(.A(new_n14245), .B(new_n14244), .Y(new_n14246));
  O2A1O1Ixp33_ASAP7_75t_L   g13990(.A1(new_n11987), .A2(new_n14241), .B(new_n14242), .C(new_n14238), .Y(new_n14247));
  A2O1A1Ixp33_ASAP7_75t_L   g13991(.A1(new_n14235), .A2(\a[62] ), .B(new_n14236), .C(new_n14238), .Y(new_n14248));
  O2A1O1Ixp33_ASAP7_75t_L   g13992(.A1(new_n14238), .A2(new_n14247), .B(new_n14248), .C(new_n14245), .Y(new_n14249));
  INVx1_ASAP7_75t_L         g13993(.A(new_n14249), .Y(new_n14250));
  NAND2xp33_ASAP7_75t_L     g13994(.A(new_n14246), .B(new_n14250), .Y(new_n14251));
  NOR2xp33_ASAP7_75t_L      g13995(.A(new_n590), .B(new_n11354), .Y(new_n14252));
  AOI221xp5_ASAP7_75t_L     g13996(.A1(\b[11] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[10] ), .C(new_n14252), .Y(new_n14253));
  O2A1O1Ixp33_ASAP7_75t_L   g13997(.A1(new_n11053), .A2(new_n754), .B(new_n14253), .C(new_n11048), .Y(new_n14254));
  O2A1O1Ixp33_ASAP7_75t_L   g13998(.A1(new_n11053), .A2(new_n754), .B(new_n14253), .C(\a[59] ), .Y(new_n14255));
  INVx1_ASAP7_75t_L         g13999(.A(new_n14255), .Y(new_n14256));
  OAI211xp5_ASAP7_75t_L     g14000(.A1(new_n11048), .A2(new_n14254), .B(new_n14251), .C(new_n14256), .Y(new_n14257));
  O2A1O1Ixp33_ASAP7_75t_L   g14001(.A1(new_n14254), .A2(new_n11048), .B(new_n14256), .C(new_n14251), .Y(new_n14258));
  INVx1_ASAP7_75t_L         g14002(.A(new_n14258), .Y(new_n14259));
  AND2x2_ASAP7_75t_L        g14003(.A(new_n14257), .B(new_n14259), .Y(new_n14260));
  INVx1_ASAP7_75t_L         g14004(.A(new_n14260), .Y(new_n14261));
  O2A1O1Ixp33_ASAP7_75t_L   g14005(.A1(new_n13937), .A2(new_n13938), .B(new_n13946), .C(new_n14261), .Y(new_n14262));
  NOR3xp33_ASAP7_75t_L      g14006(.A(new_n14260), .B(new_n13945), .C(new_n13941), .Y(new_n14263));
  NOR2xp33_ASAP7_75t_L      g14007(.A(new_n14263), .B(new_n14262), .Y(new_n14264));
  NOR2xp33_ASAP7_75t_L      g14008(.A(new_n936), .B(new_n10388), .Y(new_n14265));
  AOI221xp5_ASAP7_75t_L     g14009(.A1(new_n10086), .A2(\b[14] ), .B1(new_n11361), .B2(\b[12] ), .C(new_n14265), .Y(new_n14266));
  O2A1O1Ixp33_ASAP7_75t_L   g14010(.A1(new_n10088), .A2(new_n1268), .B(new_n14266), .C(new_n10083), .Y(new_n14267));
  INVx1_ASAP7_75t_L         g14011(.A(new_n14267), .Y(new_n14268));
  O2A1O1Ixp33_ASAP7_75t_L   g14012(.A1(new_n10088), .A2(new_n1268), .B(new_n14266), .C(\a[56] ), .Y(new_n14269));
  A2O1A1Ixp33_ASAP7_75t_L   g14013(.A1(\a[56] ), .A2(new_n14268), .B(new_n14269), .C(new_n14264), .Y(new_n14270));
  INVx1_ASAP7_75t_L         g14014(.A(new_n14269), .Y(new_n14271));
  O2A1O1Ixp33_ASAP7_75t_L   g14015(.A1(new_n14267), .A2(new_n10083), .B(new_n14271), .C(new_n14264), .Y(new_n14272));
  INVx1_ASAP7_75t_L         g14016(.A(new_n13957), .Y(new_n14273));
  A2O1A1O1Ixp25_ASAP7_75t_L g14017(.A1(new_n14273), .A2(\a[56] ), .B(new_n13958), .C(new_n13950), .D(new_n13952), .Y(new_n14274));
  A2O1A1Ixp33_ASAP7_75t_L   g14018(.A1(new_n14270), .A2(new_n14264), .B(new_n14272), .C(new_n14274), .Y(new_n14275));
  AOI21xp33_ASAP7_75t_L     g14019(.A1(new_n14270), .A2(new_n14264), .B(new_n14272), .Y(new_n14276));
  A2O1A1Ixp33_ASAP7_75t_L   g14020(.A1(new_n13954), .A2(new_n13960), .B(new_n13952), .C(new_n14276), .Y(new_n14277));
  AND2x2_ASAP7_75t_L        g14021(.A(new_n14275), .B(new_n14277), .Y(new_n14278));
  NOR2xp33_ASAP7_75t_L      g14022(.A(new_n1150), .B(new_n10400), .Y(new_n14279));
  AOI221xp5_ASAP7_75t_L     g14023(.A1(new_n9102), .A2(\b[17] ), .B1(new_n10398), .B2(\b[15] ), .C(new_n14279), .Y(new_n14280));
  O2A1O1Ixp33_ASAP7_75t_L   g14024(.A1(new_n9104), .A2(new_n1356), .B(new_n14280), .C(new_n9099), .Y(new_n14281));
  O2A1O1Ixp33_ASAP7_75t_L   g14025(.A1(new_n9104), .A2(new_n1356), .B(new_n14280), .C(\a[53] ), .Y(new_n14282));
  INVx1_ASAP7_75t_L         g14026(.A(new_n14282), .Y(new_n14283));
  O2A1O1Ixp33_ASAP7_75t_L   g14027(.A1(new_n14281), .A2(new_n9099), .B(new_n14283), .C(new_n14278), .Y(new_n14284));
  INVx1_ASAP7_75t_L         g14028(.A(new_n14281), .Y(new_n14285));
  A2O1A1Ixp33_ASAP7_75t_L   g14029(.A1(\a[53] ), .A2(new_n14285), .B(new_n14282), .C(new_n14278), .Y(new_n14286));
  INVx1_ASAP7_75t_L         g14030(.A(new_n13968), .Y(new_n14287));
  A2O1A1O1Ixp25_ASAP7_75t_L g14031(.A1(new_n13977), .A2(\a[53] ), .B(new_n13974), .C(new_n13969), .D(new_n14287), .Y(new_n14288));
  OAI211xp5_ASAP7_75t_L     g14032(.A1(new_n14278), .A2(new_n14284), .B(new_n14286), .C(new_n14288), .Y(new_n14289));
  O2A1O1Ixp33_ASAP7_75t_L   g14033(.A1(new_n14278), .A2(new_n14284), .B(new_n14286), .C(new_n14288), .Y(new_n14290));
  INVx1_ASAP7_75t_L         g14034(.A(new_n14290), .Y(new_n14291));
  NAND2xp33_ASAP7_75t_L     g14035(.A(new_n14289), .B(new_n14291), .Y(new_n14292));
  NOR2xp33_ASAP7_75t_L      g14036(.A(new_n1599), .B(new_n10065), .Y(new_n14293));
  AOI221xp5_ASAP7_75t_L     g14037(.A1(new_n8175), .A2(\b[20] ), .B1(new_n8484), .B2(\b[18] ), .C(new_n14293), .Y(new_n14294));
  O2A1O1Ixp33_ASAP7_75t_L   g14038(.A1(new_n8176), .A2(new_n1754), .B(new_n14294), .C(new_n8172), .Y(new_n14295));
  INVx1_ASAP7_75t_L         g14039(.A(new_n14295), .Y(new_n14296));
  O2A1O1Ixp33_ASAP7_75t_L   g14040(.A1(new_n8176), .A2(new_n1754), .B(new_n14294), .C(\a[50] ), .Y(new_n14297));
  AOI21xp33_ASAP7_75t_L     g14041(.A1(new_n14296), .A2(\a[50] ), .B(new_n14297), .Y(new_n14298));
  NAND2xp33_ASAP7_75t_L     g14042(.A(new_n14298), .B(new_n14292), .Y(new_n14299));
  AND2x2_ASAP7_75t_L        g14043(.A(new_n14289), .B(new_n14291), .Y(new_n14300));
  A2O1A1Ixp33_ASAP7_75t_L   g14044(.A1(\a[50] ), .A2(new_n14296), .B(new_n14297), .C(new_n14300), .Y(new_n14301));
  NAND2xp33_ASAP7_75t_L     g14045(.A(new_n14299), .B(new_n14301), .Y(new_n14302));
  AOI21xp33_ASAP7_75t_L     g14046(.A1(new_n13980), .A2(new_n13979), .B(new_n13987), .Y(new_n14303));
  XNOR2x2_ASAP7_75t_L       g14047(.A(new_n14303), .B(new_n14302), .Y(new_n14304));
  NOR2xp33_ASAP7_75t_L      g14048(.A(new_n2188), .B(new_n7318), .Y(new_n14305));
  AOI221xp5_ASAP7_75t_L     g14049(.A1(new_n7333), .A2(\b[22] ), .B1(new_n7609), .B2(\b[21] ), .C(new_n14305), .Y(new_n14306));
  O2A1O1Ixp33_ASAP7_75t_L   g14050(.A1(new_n7321), .A2(new_n2194), .B(new_n14306), .C(new_n7316), .Y(new_n14307));
  O2A1O1Ixp33_ASAP7_75t_L   g14051(.A1(new_n7321), .A2(new_n2194), .B(new_n14306), .C(\a[47] ), .Y(new_n14308));
  INVx1_ASAP7_75t_L         g14052(.A(new_n14308), .Y(new_n14309));
  O2A1O1Ixp33_ASAP7_75t_L   g14053(.A1(new_n14307), .A2(new_n7316), .B(new_n14309), .C(new_n14304), .Y(new_n14310));
  INVx1_ASAP7_75t_L         g14054(.A(new_n14307), .Y(new_n14311));
  A2O1A1Ixp33_ASAP7_75t_L   g14055(.A1(\a[47] ), .A2(new_n14311), .B(new_n14308), .C(new_n14304), .Y(new_n14312));
  OAI21xp33_ASAP7_75t_L     g14056(.A1(new_n14304), .A2(new_n14310), .B(new_n14312), .Y(new_n14313));
  INVx1_ASAP7_75t_L         g14057(.A(new_n13992), .Y(new_n14314));
  NAND2xp33_ASAP7_75t_L     g14058(.A(new_n14314), .B(new_n13999), .Y(new_n14315));
  XOR2x2_ASAP7_75t_L        g14059(.A(new_n14315), .B(new_n14313), .Y(new_n14316));
  NOR2xp33_ASAP7_75t_L      g14060(.A(new_n2205), .B(new_n6741), .Y(new_n14317));
  AOI221xp5_ASAP7_75t_L     g14061(.A1(\b[26] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[25] ), .C(new_n14317), .Y(new_n14318));
  O2A1O1Ixp33_ASAP7_75t_L   g14062(.A1(new_n6443), .A2(new_n2708), .B(new_n14318), .C(new_n6439), .Y(new_n14319));
  INVx1_ASAP7_75t_L         g14063(.A(new_n14319), .Y(new_n14320));
  O2A1O1Ixp33_ASAP7_75t_L   g14064(.A1(new_n6443), .A2(new_n2708), .B(new_n14318), .C(\a[44] ), .Y(new_n14321));
  AOI21xp33_ASAP7_75t_L     g14065(.A1(new_n14320), .A2(\a[44] ), .B(new_n14321), .Y(new_n14322));
  XOR2x2_ASAP7_75t_L        g14066(.A(new_n14322), .B(new_n14316), .Y(new_n14323));
  O2A1O1Ixp33_ASAP7_75t_L   g14067(.A1(new_n13915), .A2(new_n14007), .B(new_n14017), .C(new_n14023), .Y(new_n14324));
  NAND2xp33_ASAP7_75t_L     g14068(.A(new_n14324), .B(new_n14323), .Y(new_n14325));
  A2O1A1Ixp33_ASAP7_75t_L   g14069(.A1(new_n13741), .A2(new_n13733), .B(new_n14023), .C(new_n14015), .Y(new_n14326));
  INVx1_ASAP7_75t_L         g14070(.A(new_n14323), .Y(new_n14327));
  A2O1A1Ixp33_ASAP7_75t_L   g14071(.A1(new_n14326), .A2(new_n14017), .B(new_n14023), .C(new_n14327), .Y(new_n14328));
  NOR2xp33_ASAP7_75t_L      g14072(.A(new_n3098), .B(new_n5641), .Y(new_n14329));
  AOI221xp5_ASAP7_75t_L     g14073(.A1(\b[27] ), .A2(new_n5920), .B1(\b[28] ), .B2(new_n5623), .C(new_n14329), .Y(new_n14330));
  O2A1O1Ixp33_ASAP7_75t_L   g14074(.A1(new_n5630), .A2(new_n3104), .B(new_n14330), .C(new_n5626), .Y(new_n14331));
  NOR2xp33_ASAP7_75t_L      g14075(.A(new_n5626), .B(new_n14331), .Y(new_n14332));
  O2A1O1Ixp33_ASAP7_75t_L   g14076(.A1(new_n5630), .A2(new_n3104), .B(new_n14330), .C(\a[41] ), .Y(new_n14333));
  NOR2xp33_ASAP7_75t_L      g14077(.A(new_n14333), .B(new_n14332), .Y(new_n14334));
  NAND3xp33_ASAP7_75t_L     g14078(.A(new_n14328), .B(new_n14325), .C(new_n14334), .Y(new_n14335));
  INVx1_ASAP7_75t_L         g14079(.A(new_n14325), .Y(new_n14336));
  O2A1O1Ixp33_ASAP7_75t_L   g14080(.A1(new_n13734), .A2(new_n13742), .B(new_n14002), .C(new_n14007), .Y(new_n14337));
  O2A1O1Ixp33_ASAP7_75t_L   g14081(.A1(new_n14337), .A2(new_n14013), .B(new_n14002), .C(new_n14323), .Y(new_n14338));
  INVx1_ASAP7_75t_L         g14082(.A(new_n14334), .Y(new_n14339));
  OAI21xp33_ASAP7_75t_L     g14083(.A1(new_n14338), .A2(new_n14336), .B(new_n14339), .Y(new_n14340));
  NAND4xp25_ASAP7_75t_L     g14084(.A(new_n14340), .B(new_n14026), .C(new_n14335), .D(new_n14040), .Y(new_n14341));
  NOR3xp33_ASAP7_75t_L      g14085(.A(new_n14336), .B(new_n14338), .C(new_n14339), .Y(new_n14342));
  AOI21xp33_ASAP7_75t_L     g14086(.A1(new_n14328), .A2(new_n14325), .B(new_n14334), .Y(new_n14343));
  A2O1A1Ixp33_ASAP7_75t_L   g14087(.A1(new_n14030), .A2(new_n14031), .B(new_n14033), .C(new_n14026), .Y(new_n14344));
  OAI21xp33_ASAP7_75t_L     g14088(.A1(new_n14342), .A2(new_n14343), .B(new_n14344), .Y(new_n14345));
  NOR2xp33_ASAP7_75t_L      g14089(.A(new_n3891), .B(new_n4908), .Y(new_n14346));
  AOI221xp5_ASAP7_75t_L     g14090(.A1(\b[30] ), .A2(new_n5139), .B1(\b[31] ), .B2(new_n4916), .C(new_n14346), .Y(new_n14347));
  O2A1O1Ixp33_ASAP7_75t_L   g14091(.A1(new_n4911), .A2(new_n3897), .B(new_n14347), .C(new_n4906), .Y(new_n14348));
  NOR2xp33_ASAP7_75t_L      g14092(.A(new_n4906), .B(new_n14348), .Y(new_n14349));
  O2A1O1Ixp33_ASAP7_75t_L   g14093(.A1(new_n4911), .A2(new_n3897), .B(new_n14347), .C(\a[38] ), .Y(new_n14350));
  NOR2xp33_ASAP7_75t_L      g14094(.A(new_n14350), .B(new_n14349), .Y(new_n14351));
  INVx1_ASAP7_75t_L         g14095(.A(new_n14351), .Y(new_n14352));
  AO21x2_ASAP7_75t_L        g14096(.A1(new_n14345), .A2(new_n14341), .B(new_n14352), .Y(new_n14353));
  NAND3xp33_ASAP7_75t_L     g14097(.A(new_n14341), .B(new_n14345), .C(new_n14352), .Y(new_n14354));
  A2O1A1Ixp33_ASAP7_75t_L   g14098(.A1(new_n14037), .A2(new_n14032), .B(new_n14038), .C(new_n14049), .Y(new_n14355));
  NAND3xp33_ASAP7_75t_L     g14099(.A(new_n14353), .B(new_n14355), .C(new_n14354), .Y(new_n14356));
  AOI21xp33_ASAP7_75t_L     g14100(.A1(new_n14341), .A2(new_n14345), .B(new_n14352), .Y(new_n14357));
  AND3x1_ASAP7_75t_L        g14101(.A(new_n14341), .B(new_n14345), .C(new_n14352), .Y(new_n14358));
  INVx1_ASAP7_75t_L         g14102(.A(new_n14355), .Y(new_n14359));
  OAI21xp33_ASAP7_75t_L     g14103(.A1(new_n14357), .A2(new_n14358), .B(new_n14359), .Y(new_n14360));
  NOR2xp33_ASAP7_75t_L      g14104(.A(new_n4581), .B(new_n4147), .Y(new_n14361));
  AOI221xp5_ASAP7_75t_L     g14105(.A1(\b[33] ), .A2(new_n4402), .B1(\b[34] ), .B2(new_n4155), .C(new_n14361), .Y(new_n14362));
  O2A1O1Ixp33_ASAP7_75t_L   g14106(.A1(new_n4150), .A2(new_n4589), .B(new_n14362), .C(new_n4145), .Y(new_n14363));
  INVx1_ASAP7_75t_L         g14107(.A(new_n14363), .Y(new_n14364));
  O2A1O1Ixp33_ASAP7_75t_L   g14108(.A1(new_n4150), .A2(new_n4589), .B(new_n14362), .C(\a[35] ), .Y(new_n14365));
  AOI21xp33_ASAP7_75t_L     g14109(.A1(new_n14364), .A2(\a[35] ), .B(new_n14365), .Y(new_n14366));
  NAND3xp33_ASAP7_75t_L     g14110(.A(new_n14360), .B(new_n14356), .C(new_n14366), .Y(new_n14367));
  AO21x2_ASAP7_75t_L        g14111(.A1(new_n14356), .A2(new_n14360), .B(new_n14366), .Y(new_n14368));
  NAND2xp33_ASAP7_75t_L     g14112(.A(new_n14367), .B(new_n14368), .Y(new_n14369));
  NAND2xp33_ASAP7_75t_L     g14113(.A(new_n14049), .B(new_n14048), .Y(new_n14370));
  MAJIxp5_ASAP7_75t_L       g14114(.A(new_n14370), .B(new_n13912), .C(new_n13913), .Y(new_n14371));
  NAND2xp33_ASAP7_75t_L     g14115(.A(\b[37] ), .B(new_n3499), .Y(new_n14372));
  OAI221xp5_ASAP7_75t_L     g14116(.A1(new_n3510), .A2(new_n5311), .B1(new_n4613), .B2(new_n3703), .C(new_n14372), .Y(new_n14373));
  AOI21xp33_ASAP7_75t_L     g14117(.A1(new_n6083), .A2(new_n3505), .B(new_n14373), .Y(new_n14374));
  NAND2xp33_ASAP7_75t_L     g14118(.A(\a[32] ), .B(new_n14374), .Y(new_n14375));
  A2O1A1Ixp33_ASAP7_75t_L   g14119(.A1(new_n6083), .A2(new_n3505), .B(new_n14373), .C(new_n3493), .Y(new_n14376));
  NAND2xp33_ASAP7_75t_L     g14120(.A(new_n14376), .B(new_n14375), .Y(new_n14377));
  XNOR2x2_ASAP7_75t_L       g14121(.A(new_n14377), .B(new_n14371), .Y(new_n14378));
  AOI21xp33_ASAP7_75t_L     g14122(.A1(new_n14368), .A2(new_n14367), .B(new_n14378), .Y(new_n14379));
  INVx1_ASAP7_75t_L         g14123(.A(new_n14379), .Y(new_n14380));
  NOR2xp33_ASAP7_75t_L      g14124(.A(new_n14378), .B(new_n14369), .Y(new_n14381));
  NAND2xp33_ASAP7_75t_L     g14125(.A(\b[40] ), .B(new_n2936), .Y(new_n14382));
  OAI221xp5_ASAP7_75t_L     g14126(.A1(new_n2930), .A2(new_n6110), .B1(new_n5570), .B2(new_n3133), .C(new_n14382), .Y(new_n14383));
  A2O1A1Ixp33_ASAP7_75t_L   g14127(.A1(new_n6118), .A2(new_n2932), .B(new_n14383), .C(\a[29] ), .Y(new_n14384));
  NAND2xp33_ASAP7_75t_L     g14128(.A(\a[29] ), .B(new_n14384), .Y(new_n14385));
  A2O1A1Ixp33_ASAP7_75t_L   g14129(.A1(new_n6118), .A2(new_n2932), .B(new_n14383), .C(new_n2928), .Y(new_n14386));
  INVx1_ASAP7_75t_L         g14130(.A(new_n13779), .Y(new_n14387));
  O2A1O1Ixp33_ASAP7_75t_L   g14131(.A1(new_n13659), .A2(new_n13660), .B(new_n13780), .C(new_n14387), .Y(new_n14388));
  NAND2xp33_ASAP7_75t_L     g14132(.A(new_n13907), .B(new_n14388), .Y(new_n14389));
  O2A1O1Ixp33_ASAP7_75t_L   g14133(.A1(new_n14053), .A2(new_n14056), .B(new_n14389), .C(new_n13908), .Y(new_n14390));
  NAND3xp33_ASAP7_75t_L     g14134(.A(new_n14390), .B(new_n14386), .C(new_n14385), .Y(new_n14391));
  AOI21xp33_ASAP7_75t_L     g14135(.A1(new_n14386), .A2(new_n14385), .B(new_n14390), .Y(new_n14392));
  INVx1_ASAP7_75t_L         g14136(.A(new_n14392), .Y(new_n14393));
  NAND2xp33_ASAP7_75t_L     g14137(.A(new_n14378), .B(new_n14369), .Y(new_n14394));
  OAI21xp33_ASAP7_75t_L     g14138(.A1(new_n14378), .A2(new_n14379), .B(new_n14394), .Y(new_n14395));
  NAND3xp33_ASAP7_75t_L     g14139(.A(new_n14395), .B(new_n14393), .C(new_n14391), .Y(new_n14396));
  INVx1_ASAP7_75t_L         g14140(.A(new_n14391), .Y(new_n14397));
  NOR3xp33_ASAP7_75t_L      g14141(.A(new_n14395), .B(new_n14392), .C(new_n14397), .Y(new_n14398));
  A2O1A1O1Ixp25_ASAP7_75t_L g14142(.A1(new_n14380), .A2(new_n14369), .B(new_n14381), .C(new_n14396), .D(new_n14398), .Y(new_n14399));
  NAND2xp33_ASAP7_75t_L     g14143(.A(\b[43] ), .B(new_n2421), .Y(new_n14400));
  OAI221xp5_ASAP7_75t_L     g14144(.A1(new_n2415), .A2(new_n6944), .B1(new_n6378), .B2(new_n2572), .C(new_n14400), .Y(new_n14401));
  AOI21xp33_ASAP7_75t_L     g14145(.A1(new_n7824), .A2(new_n2417), .B(new_n14401), .Y(new_n14402));
  NAND2xp33_ASAP7_75t_L     g14146(.A(\a[26] ), .B(new_n14402), .Y(new_n14403));
  A2O1A1Ixp33_ASAP7_75t_L   g14147(.A1(new_n7824), .A2(new_n2417), .B(new_n14401), .C(new_n2413), .Y(new_n14404));
  NAND2xp33_ASAP7_75t_L     g14148(.A(new_n14404), .B(new_n14403), .Y(new_n14405));
  INVx1_ASAP7_75t_L         g14149(.A(new_n14405), .Y(new_n14406));
  A2O1A1O1Ixp25_ASAP7_75t_L g14150(.A1(new_n14069), .A2(new_n14063), .B(new_n14080), .C(new_n14066), .D(new_n14406), .Y(new_n14407));
  A2O1A1O1Ixp25_ASAP7_75t_L g14151(.A1(new_n14069), .A2(new_n14063), .B(new_n14080), .C(new_n14066), .D(new_n14405), .Y(new_n14408));
  INVx1_ASAP7_75t_L         g14152(.A(new_n14408), .Y(new_n14409));
  O2A1O1Ixp33_ASAP7_75t_L   g14153(.A1(new_n14406), .A2(new_n14407), .B(new_n14409), .C(new_n14399), .Y(new_n14410));
  INVx1_ASAP7_75t_L         g14154(.A(new_n14407), .Y(new_n14411));
  A2O1A1Ixp33_ASAP7_75t_L   g14155(.A1(new_n14411), .A2(new_n14405), .B(new_n14408), .C(new_n14399), .Y(new_n14412));
  OAI21xp33_ASAP7_75t_L     g14156(.A1(new_n14399), .A2(new_n14410), .B(new_n14412), .Y(new_n14413));
  XOR2x2_ASAP7_75t_L        g14157(.A(new_n14226), .B(new_n14413), .Y(new_n14414));
  XNOR2x2_ASAP7_75t_L       g14158(.A(new_n14414), .B(new_n14215), .Y(new_n14415));
  XNOR2x2_ASAP7_75t_L       g14159(.A(new_n14203), .B(new_n14415), .Y(new_n14416));
  A2O1A1Ixp33_ASAP7_75t_L   g14160(.A1(new_n14194), .A2(new_n14191), .B(new_n14195), .C(new_n14416), .Y(new_n14417));
  O2A1O1Ixp33_ASAP7_75t_L   g14161(.A1(new_n13625), .A2(new_n13811), .B(new_n14105), .C(new_n14111), .Y(new_n14418));
  O2A1O1Ixp33_ASAP7_75t_L   g14162(.A1(new_n14114), .A2(new_n14418), .B(new_n14104), .C(new_n14111), .Y(new_n14419));
  NAND2xp33_ASAP7_75t_L     g14163(.A(new_n14191), .B(new_n14419), .Y(new_n14420));
  INVx1_ASAP7_75t_L         g14164(.A(new_n14195), .Y(new_n14421));
  XOR2x2_ASAP7_75t_L        g14165(.A(new_n14203), .B(new_n14415), .Y(new_n14422));
  NAND3xp33_ASAP7_75t_L     g14166(.A(new_n14422), .B(new_n14421), .C(new_n14420), .Y(new_n14423));
  NAND2xp33_ASAP7_75t_L     g14167(.A(new_n14423), .B(new_n14417), .Y(new_n14424));
  OAI22xp33_ASAP7_75t_L     g14168(.A1(new_n1550), .A2(new_n11303), .B1(new_n10978), .B2(new_n712), .Y(new_n14425));
  AOI221xp5_ASAP7_75t_L     g14169(.A1(new_n640), .A2(\b[59] ), .B1(new_n718), .B2(new_n12577), .C(new_n14425), .Y(new_n14426));
  XNOR2x2_ASAP7_75t_L       g14170(.A(\a[11] ), .B(new_n14426), .Y(new_n14427));
  A2O1A1Ixp33_ASAP7_75t_L   g14171(.A1(new_n14118), .A2(new_n14116), .B(new_n13894), .C(new_n14122), .Y(new_n14428));
  NOR2xp33_ASAP7_75t_L      g14172(.A(new_n14427), .B(new_n14428), .Y(new_n14429));
  INVx1_ASAP7_75t_L         g14173(.A(new_n14429), .Y(new_n14430));
  A2O1A1Ixp33_ASAP7_75t_L   g14174(.A1(new_n14119), .A2(new_n14121), .B(new_n13895), .C(new_n14427), .Y(new_n14431));
  NAND3xp33_ASAP7_75t_L     g14175(.A(new_n14424), .B(new_n14431), .C(new_n14430), .Y(new_n14432));
  INVx1_ASAP7_75t_L         g14176(.A(new_n14431), .Y(new_n14433));
  NOR3xp33_ASAP7_75t_L      g14177(.A(new_n14424), .B(new_n14433), .C(new_n14429), .Y(new_n14434));
  AOI21xp33_ASAP7_75t_L     g14178(.A1(new_n14432), .A2(new_n14424), .B(new_n14434), .Y(new_n14435));
  A2O1A1O1Ixp25_ASAP7_75t_L g14179(.A1(new_n14131), .A2(new_n14128), .B(new_n14124), .C(new_n14133), .D(new_n14188), .Y(new_n14436));
  A2O1A1Ixp33_ASAP7_75t_L   g14180(.A1(new_n14182), .A2(new_n13830), .B(new_n13824), .C(new_n13832), .Y(new_n14437));
  A2O1A1Ixp33_ASAP7_75t_L   g14181(.A1(new_n14127), .A2(new_n14437), .B(new_n14132), .C(new_n14188), .Y(new_n14438));
  O2A1O1Ixp33_ASAP7_75t_L   g14182(.A1(new_n14188), .A2(new_n14436), .B(new_n14438), .C(new_n14435), .Y(new_n14439));
  INVx1_ASAP7_75t_L         g14183(.A(new_n14439), .Y(new_n14440));
  OAI21xp33_ASAP7_75t_L     g14184(.A1(new_n14188), .A2(new_n14436), .B(new_n14435), .Y(new_n14441));
  A2O1A1Ixp33_ASAP7_75t_L   g14185(.A1(new_n14185), .A2(new_n14188), .B(new_n14441), .C(new_n14440), .Y(new_n14442));
  O2A1O1Ixp33_ASAP7_75t_L   g14186(.A1(new_n14174), .A2(new_n14177), .B(new_n14178), .C(new_n14442), .Y(new_n14443));
  A2O1A1O1Ixp25_ASAP7_75t_L g14187(.A1(new_n12263), .A2(new_n12267), .B(new_n12262), .C(new_n12605), .D(new_n12604), .Y(new_n14444));
  A2O1A1O1Ixp25_ASAP7_75t_L g14188(.A1(new_n12603), .A2(new_n14444), .B(new_n356), .C(new_n375), .D(new_n12956), .Y(new_n14445));
  OAI221xp5_ASAP7_75t_L     g14189(.A1(new_n14128), .A2(new_n14129), .B1(new_n14120), .B2(new_n14123), .C(new_n14131), .Y(new_n14446));
  A2O1A1O1Ixp25_ASAP7_75t_L g14190(.A1(new_n14134), .A2(new_n14446), .B(new_n13888), .C(new_n13885), .D(new_n14175), .Y(new_n14447));
  A2O1A1O1Ixp25_ASAP7_75t_L g14191(.A1(new_n14171), .A2(new_n14445), .B(new_n14173), .C(new_n14176), .D(new_n14447), .Y(new_n14448));
  INVx1_ASAP7_75t_L         g14192(.A(new_n14441), .Y(new_n14449));
  A2O1A1Ixp33_ASAP7_75t_L   g14193(.A1(new_n14449), .A2(new_n14438), .B(new_n14439), .C(new_n14448), .Y(new_n14450));
  INVx1_ASAP7_75t_L         g14194(.A(new_n14450), .Y(new_n14451));
  OAI21xp33_ASAP7_75t_L     g14195(.A1(new_n14443), .A2(new_n14451), .B(new_n14169), .Y(new_n14452));
  A2O1A1Ixp33_ASAP7_75t_L   g14196(.A1(new_n14446), .A2(new_n14134), .B(new_n13888), .C(new_n13885), .Y(new_n14453));
  INVx1_ASAP7_75t_L         g14197(.A(new_n14171), .Y(new_n14454));
  A2O1A1Ixp33_ASAP7_75t_L   g14198(.A1(new_n12986), .A2(new_n359), .B(new_n14170), .C(new_n346), .Y(new_n14455));
  O2A1O1Ixp33_ASAP7_75t_L   g14199(.A1(new_n14454), .A2(new_n346), .B(new_n14455), .C(new_n14453), .Y(new_n14456));
  INVx1_ASAP7_75t_L         g14200(.A(new_n14188), .Y(new_n14457));
  O2A1O1Ixp33_ASAP7_75t_L   g14201(.A1(new_n14457), .A2(new_n14184), .B(new_n14449), .C(new_n14439), .Y(new_n14458));
  A2O1A1Ixp33_ASAP7_75t_L   g14202(.A1(new_n14176), .A2(new_n14453), .B(new_n14456), .C(new_n14458), .Y(new_n14459));
  NAND4xp25_ASAP7_75t_L     g14203(.A(new_n14459), .B(new_n14138), .C(new_n14152), .D(new_n14450), .Y(new_n14460));
  NAND2xp33_ASAP7_75t_L     g14204(.A(new_n14460), .B(new_n14452), .Y(new_n14461));
  A2O1A1Ixp33_ASAP7_75t_L   g14205(.A1(new_n14148), .A2(new_n14149), .B(new_n14160), .C(new_n14166), .Y(new_n14462));
  NAND3xp33_ASAP7_75t_L     g14206(.A(new_n14462), .B(new_n14149), .C(new_n14460), .Y(new_n14463));
  O2A1O1Ixp33_ASAP7_75t_L   g14207(.A1(new_n14443), .A2(new_n14451), .B(new_n14169), .C(new_n14463), .Y(new_n14464));
  O2A1O1Ixp33_ASAP7_75t_L   g14208(.A1(new_n14150), .A2(new_n14165), .B(new_n14461), .C(new_n14464), .Y(\f[68] ));
  INVx1_ASAP7_75t_L         g14209(.A(new_n13866), .Y(new_n14466));
  A2O1A1Ixp33_ASAP7_75t_L   g14210(.A1(new_n14151), .A2(new_n14466), .B(new_n14164), .C(new_n14149), .Y(new_n14467));
  NAND2xp33_ASAP7_75t_L     g14211(.A(new_n14450), .B(new_n14459), .Y(new_n14468));
  O2A1O1Ixp33_ASAP7_75t_L   g14212(.A1(new_n13873), .A2(new_n13879), .B(new_n14152), .C(new_n14468), .Y(new_n14469));
  O2A1O1Ixp33_ASAP7_75t_L   g14213(.A1(new_n14456), .A2(new_n14453), .B(new_n14458), .C(new_n14177), .Y(new_n14470));
  OAI22xp33_ASAP7_75t_L     g14214(.A1(new_n513), .A2(new_n12603), .B1(new_n12258), .B2(new_n506), .Y(new_n14471));
  AOI221xp5_ASAP7_75t_L     g14215(.A1(new_n475), .A2(\b[63] ), .B1(new_n483), .B2(new_n12961), .C(new_n14471), .Y(new_n14472));
  XNOR2x2_ASAP7_75t_L       g14216(.A(new_n466), .B(new_n14472), .Y(new_n14473));
  INVx1_ASAP7_75t_L         g14217(.A(new_n14473), .Y(new_n14474));
  INVx1_ASAP7_75t_L         g14218(.A(new_n14436), .Y(new_n14475));
  A2O1A1O1Ixp25_ASAP7_75t_L g14219(.A1(new_n14438), .A2(new_n14188), .B(new_n14435), .C(new_n14475), .D(new_n14473), .Y(new_n14476));
  INVx1_ASAP7_75t_L         g14220(.A(new_n14476), .Y(new_n14477));
  A2O1A1O1Ixp25_ASAP7_75t_L g14221(.A1(new_n14438), .A2(new_n14188), .B(new_n14435), .C(new_n14475), .D(new_n14474), .Y(new_n14478));
  OAI22xp33_ASAP7_75t_L     g14222(.A1(new_n1550), .A2(new_n11591), .B1(new_n11303), .B2(new_n712), .Y(new_n14479));
  AOI221xp5_ASAP7_75t_L     g14223(.A1(new_n640), .A2(\b[60] ), .B1(new_n718), .B2(new_n13839), .C(new_n14479), .Y(new_n14480));
  XNOR2x2_ASAP7_75t_L       g14224(.A(new_n637), .B(new_n14480), .Y(new_n14481));
  INVx1_ASAP7_75t_L         g14225(.A(new_n14481), .Y(new_n14482));
  A2O1A1Ixp33_ASAP7_75t_L   g14226(.A1(new_n14417), .A2(new_n14423), .B(new_n14429), .C(new_n14431), .Y(new_n14483));
  NOR2xp33_ASAP7_75t_L      g14227(.A(new_n14482), .B(new_n14483), .Y(new_n14484));
  A2O1A1O1Ixp25_ASAP7_75t_L g14228(.A1(new_n14423), .A2(new_n14417), .B(new_n14429), .C(new_n14431), .D(new_n14481), .Y(new_n14485));
  NAND2xp33_ASAP7_75t_L     g14229(.A(\b[48] ), .B(new_n1955), .Y(new_n14486));
  OAI221xp5_ASAP7_75t_L     g14230(.A1(new_n1962), .A2(new_n7552), .B1(new_n7270), .B2(new_n2089), .C(new_n14486), .Y(new_n14487));
  A2O1A1Ixp33_ASAP7_75t_L   g14231(.A1(new_n11656), .A2(new_n1964), .B(new_n14487), .C(\a[23] ), .Y(new_n14488));
  NAND2xp33_ASAP7_75t_L     g14232(.A(\a[23] ), .B(new_n14488), .Y(new_n14489));
  A2O1A1Ixp33_ASAP7_75t_L   g14233(.A1(new_n11656), .A2(new_n1964), .B(new_n14487), .C(new_n1952), .Y(new_n14490));
  INVx1_ASAP7_75t_L         g14234(.A(new_n14225), .Y(new_n14491));
  AO21x2_ASAP7_75t_L        g14235(.A1(new_n14395), .A2(new_n14396), .B(new_n14398), .Y(new_n14492));
  A2O1A1Ixp33_ASAP7_75t_L   g14236(.A1(new_n14405), .A2(new_n14411), .B(new_n14408), .C(new_n14492), .Y(new_n14493));
  INVx1_ASAP7_75t_L         g14237(.A(new_n14412), .Y(new_n14494));
  A2O1A1O1Ixp25_ASAP7_75t_L g14238(.A1(new_n14492), .A2(new_n14493), .B(new_n14494), .C(new_n14223), .D(new_n14491), .Y(new_n14495));
  NAND3xp33_ASAP7_75t_L     g14239(.A(new_n14495), .B(new_n14490), .C(new_n14489), .Y(new_n14496));
  NAND2xp33_ASAP7_75t_L     g14240(.A(new_n14490), .B(new_n14489), .Y(new_n14497));
  A2O1A1Ixp33_ASAP7_75t_L   g14241(.A1(new_n14413), .A2(new_n14223), .B(new_n14491), .C(new_n14497), .Y(new_n14498));
  AND2x2_ASAP7_75t_L        g14242(.A(new_n14498), .B(new_n14496), .Y(new_n14499));
  OAI22xp33_ASAP7_75t_L     g14243(.A1(new_n2572), .A2(new_n6671), .B1(new_n6944), .B2(new_n2410), .Y(new_n14500));
  AOI221xp5_ASAP7_75t_L     g14244(.A1(new_n2423), .A2(\b[45] ), .B1(new_n2417), .B2(new_n7256), .C(new_n14500), .Y(new_n14501));
  XNOR2x2_ASAP7_75t_L       g14245(.A(new_n2413), .B(new_n14501), .Y(new_n14502));
  INVx1_ASAP7_75t_L         g14246(.A(new_n14502), .Y(new_n14503));
  A2O1A1O1Ixp25_ASAP7_75t_L g14247(.A1(new_n14409), .A2(new_n14406), .B(new_n14399), .C(new_n14411), .D(new_n14502), .Y(new_n14504));
  INVx1_ASAP7_75t_L         g14248(.A(new_n14504), .Y(new_n14505));
  O2A1O1Ixp33_ASAP7_75t_L   g14249(.A1(new_n14067), .A2(new_n14064), .B(new_n14060), .C(new_n14065), .Y(new_n14506));
  NAND2xp33_ASAP7_75t_L     g14250(.A(new_n14405), .B(new_n14506), .Y(new_n14507));
  A2O1A1O1Ixp25_ASAP7_75t_L g14251(.A1(new_n14507), .A2(new_n14506), .B(new_n14399), .C(new_n14411), .D(new_n14503), .Y(new_n14508));
  OAI22xp33_ASAP7_75t_L     g14252(.A1(new_n3133), .A2(new_n5855), .B1(new_n6110), .B2(new_n2925), .Y(new_n14509));
  AOI221xp5_ASAP7_75t_L     g14253(.A1(new_n2938), .A2(\b[42] ), .B1(new_n2932), .B2(new_n6389), .C(new_n14509), .Y(new_n14510));
  XNOR2x2_ASAP7_75t_L       g14254(.A(new_n2928), .B(new_n14510), .Y(new_n14511));
  A2O1A1O1Ixp25_ASAP7_75t_L g14255(.A1(new_n14369), .A2(new_n14380), .B(new_n14381), .C(new_n14391), .D(new_n14392), .Y(new_n14512));
  NAND2xp33_ASAP7_75t_L     g14256(.A(new_n14511), .B(new_n14512), .Y(new_n14513));
  INVx1_ASAP7_75t_L         g14257(.A(new_n14511), .Y(new_n14514));
  A2O1A1Ixp33_ASAP7_75t_L   g14258(.A1(new_n14395), .A2(new_n14391), .B(new_n14392), .C(new_n14514), .Y(new_n14515));
  NOR3xp33_ASAP7_75t_L      g14259(.A(new_n14358), .B(new_n14359), .C(new_n14357), .Y(new_n14516));
  A2O1A1O1Ixp25_ASAP7_75t_L g14260(.A1(new_n14364), .A2(\a[35] ), .B(new_n14365), .C(new_n14360), .D(new_n14516), .Y(new_n14517));
  INVx1_ASAP7_75t_L         g14261(.A(new_n14517), .Y(new_n14518));
  NOR2xp33_ASAP7_75t_L      g14262(.A(new_n4101), .B(new_n4908), .Y(new_n14519));
  AOI221xp5_ASAP7_75t_L     g14263(.A1(\b[31] ), .A2(new_n5139), .B1(\b[32] ), .B2(new_n4916), .C(new_n14519), .Y(new_n14520));
  O2A1O1Ixp33_ASAP7_75t_L   g14264(.A1(new_n4911), .A2(new_n4108), .B(new_n14520), .C(new_n4906), .Y(new_n14521));
  O2A1O1Ixp33_ASAP7_75t_L   g14265(.A1(new_n4911), .A2(new_n4108), .B(new_n14520), .C(\a[38] ), .Y(new_n14522));
  INVx1_ASAP7_75t_L         g14266(.A(new_n14522), .Y(new_n14523));
  OAI21xp33_ASAP7_75t_L     g14267(.A1(new_n4906), .A2(new_n14521), .B(new_n14523), .Y(new_n14524));
  INVx1_ASAP7_75t_L         g14268(.A(new_n14302), .Y(new_n14525));
  A2O1A1O1Ixp25_ASAP7_75t_L g14269(.A1(new_n13980), .A2(new_n13979), .B(new_n13987), .C(new_n14525), .D(new_n14310), .Y(new_n14526));
  INVx1_ASAP7_75t_L         g14270(.A(new_n14254), .Y(new_n14527));
  A2O1A1O1Ixp25_ASAP7_75t_L g14271(.A1(\a[59] ), .A2(new_n14527), .B(new_n14255), .C(new_n14246), .D(new_n14249), .Y(new_n14528));
  NOR2xp33_ASAP7_75t_L      g14272(.A(new_n384), .B(new_n13030), .Y(new_n14529));
  INVx1_ASAP7_75t_L         g14273(.A(new_n14529), .Y(new_n14530));
  XNOR2x2_ASAP7_75t_L       g14274(.A(\a[5] ), .B(\a[2] ), .Y(new_n14531));
  O2A1O1Ixp33_ASAP7_75t_L   g14275(.A1(new_n427), .A2(new_n12672), .B(new_n14530), .C(new_n14531), .Y(new_n14532));
  O2A1O1Ixp33_ASAP7_75t_L   g14276(.A1(new_n12669), .A2(new_n12671), .B(\b[6] ), .C(new_n14529), .Y(new_n14533));
  AND2x2_ASAP7_75t_L        g14277(.A(new_n14531), .B(new_n14533), .Y(new_n14534));
  NOR2xp33_ASAP7_75t_L      g14278(.A(new_n14532), .B(new_n14534), .Y(new_n14535));
  NOR3xp33_ASAP7_75t_L      g14279(.A(new_n14247), .B(new_n14535), .C(new_n14229), .Y(new_n14536));
  O2A1O1Ixp33_ASAP7_75t_L   g14280(.A1(new_n12669), .A2(new_n12671), .B(\b[5] ), .C(new_n14227), .Y(new_n14537));
  INVx1_ASAP7_75t_L         g14281(.A(new_n14535), .Y(new_n14538));
  O2A1O1Ixp33_ASAP7_75t_L   g14282(.A1(new_n257), .A2(new_n14537), .B(new_n14240), .C(new_n14538), .Y(new_n14539));
  OAI22xp33_ASAP7_75t_L     g14283(.A1(new_n12320), .A2(new_n448), .B1(new_n534), .B2(new_n12318), .Y(new_n14540));
  AOI221xp5_ASAP7_75t_L     g14284(.A1(new_n11995), .A2(\b[9] ), .B1(new_n11997), .B2(new_n602), .C(new_n14540), .Y(new_n14541));
  XNOR2x2_ASAP7_75t_L       g14285(.A(new_n11987), .B(new_n14541), .Y(new_n14542));
  OAI21xp33_ASAP7_75t_L     g14286(.A1(new_n14536), .A2(new_n14539), .B(new_n14542), .Y(new_n14543));
  NOR2xp33_ASAP7_75t_L      g14287(.A(new_n14539), .B(new_n14536), .Y(new_n14544));
  INVx1_ASAP7_75t_L         g14288(.A(new_n14542), .Y(new_n14545));
  NAND2xp33_ASAP7_75t_L     g14289(.A(new_n14544), .B(new_n14545), .Y(new_n14546));
  NAND2xp33_ASAP7_75t_L     g14290(.A(new_n14543), .B(new_n14546), .Y(new_n14547));
  NOR2xp33_ASAP7_75t_L      g14291(.A(new_n680), .B(new_n11354), .Y(new_n14548));
  AOI221xp5_ASAP7_75t_L     g14292(.A1(\b[12] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[11] ), .C(new_n14548), .Y(new_n14549));
  O2A1O1Ixp33_ASAP7_75t_L   g14293(.A1(new_n11053), .A2(new_n841), .B(new_n14549), .C(new_n11048), .Y(new_n14550));
  INVx1_ASAP7_75t_L         g14294(.A(new_n14550), .Y(new_n14551));
  O2A1O1Ixp33_ASAP7_75t_L   g14295(.A1(new_n11053), .A2(new_n841), .B(new_n14549), .C(\a[59] ), .Y(new_n14552));
  INVx1_ASAP7_75t_L         g14296(.A(new_n14547), .Y(new_n14553));
  A2O1A1Ixp33_ASAP7_75t_L   g14297(.A1(new_n14551), .A2(\a[59] ), .B(new_n14552), .C(new_n14553), .Y(new_n14554));
  INVx1_ASAP7_75t_L         g14298(.A(new_n14554), .Y(new_n14555));
  A2O1A1Ixp33_ASAP7_75t_L   g14299(.A1(new_n14551), .A2(\a[59] ), .B(new_n14552), .C(new_n14547), .Y(new_n14556));
  O2A1O1Ixp33_ASAP7_75t_L   g14300(.A1(new_n14547), .A2(new_n14555), .B(new_n14556), .C(new_n14528), .Y(new_n14557));
  O2A1O1Ixp33_ASAP7_75t_L   g14301(.A1(new_n14244), .A2(new_n14245), .B(new_n14259), .C(new_n14557), .Y(new_n14558));
  INVx1_ASAP7_75t_L         g14302(.A(new_n14528), .Y(new_n14559));
  O2A1O1Ixp33_ASAP7_75t_L   g14303(.A1(new_n14547), .A2(new_n14555), .B(new_n14556), .C(new_n14559), .Y(new_n14560));
  INVx1_ASAP7_75t_L         g14304(.A(new_n14560), .Y(new_n14561));
  A2O1A1Ixp33_ASAP7_75t_L   g14305(.A1(new_n14259), .A2(new_n14250), .B(new_n14557), .C(new_n14561), .Y(new_n14562));
  NOR2xp33_ASAP7_75t_L      g14306(.A(new_n960), .B(new_n10388), .Y(new_n14563));
  AOI221xp5_ASAP7_75t_L     g14307(.A1(new_n10086), .A2(\b[15] ), .B1(new_n11361), .B2(\b[13] ), .C(new_n14563), .Y(new_n14564));
  O2A1O1Ixp33_ASAP7_75t_L   g14308(.A1(new_n10088), .A2(new_n1774), .B(new_n14564), .C(new_n10083), .Y(new_n14565));
  INVx1_ASAP7_75t_L         g14309(.A(new_n14565), .Y(new_n14566));
  O2A1O1Ixp33_ASAP7_75t_L   g14310(.A1(new_n10088), .A2(new_n1774), .B(new_n14564), .C(\a[56] ), .Y(new_n14567));
  A2O1A1Ixp33_ASAP7_75t_L   g14311(.A1(\a[56] ), .A2(new_n14566), .B(new_n14567), .C(new_n14562), .Y(new_n14568));
  INVx1_ASAP7_75t_L         g14312(.A(new_n14567), .Y(new_n14569));
  O2A1O1Ixp33_ASAP7_75t_L   g14313(.A1(new_n14565), .A2(new_n10083), .B(new_n14569), .C(new_n14562), .Y(new_n14570));
  O2A1O1Ixp33_ASAP7_75t_L   g14314(.A1(new_n14558), .A2(new_n14560), .B(new_n14568), .C(new_n14570), .Y(new_n14571));
  A2O1A1O1Ixp25_ASAP7_75t_L g14315(.A1(new_n14268), .A2(\a[56] ), .B(new_n14269), .C(new_n14264), .D(new_n14262), .Y(new_n14572));
  NAND2xp33_ASAP7_75t_L     g14316(.A(new_n14572), .B(new_n14571), .Y(new_n14573));
  INVx1_ASAP7_75t_L         g14317(.A(new_n14572), .Y(new_n14574));
  A2O1A1Ixp33_ASAP7_75t_L   g14318(.A1(new_n14568), .A2(new_n14562), .B(new_n14570), .C(new_n14574), .Y(new_n14575));
  AND2x2_ASAP7_75t_L        g14319(.A(new_n14575), .B(new_n14573), .Y(new_n14576));
  NOR2xp33_ASAP7_75t_L      g14320(.A(new_n1349), .B(new_n10400), .Y(new_n14577));
  AOI221xp5_ASAP7_75t_L     g14321(.A1(new_n9102), .A2(\b[18] ), .B1(new_n10398), .B2(\b[16] ), .C(new_n14577), .Y(new_n14578));
  O2A1O1Ixp33_ASAP7_75t_L   g14322(.A1(new_n9104), .A2(new_n1464), .B(new_n14578), .C(new_n9099), .Y(new_n14579));
  INVx1_ASAP7_75t_L         g14323(.A(new_n14579), .Y(new_n14580));
  O2A1O1Ixp33_ASAP7_75t_L   g14324(.A1(new_n9104), .A2(new_n1464), .B(new_n14578), .C(\a[53] ), .Y(new_n14581));
  A2O1A1Ixp33_ASAP7_75t_L   g14325(.A1(\a[53] ), .A2(new_n14580), .B(new_n14581), .C(new_n14576), .Y(new_n14582));
  INVx1_ASAP7_75t_L         g14326(.A(new_n14581), .Y(new_n14583));
  O2A1O1Ixp33_ASAP7_75t_L   g14327(.A1(new_n14579), .A2(new_n9099), .B(new_n14583), .C(new_n14576), .Y(new_n14584));
  AOI21xp33_ASAP7_75t_L     g14328(.A1(new_n14582), .A2(new_n14576), .B(new_n14584), .Y(new_n14585));
  A2O1A1Ixp33_ASAP7_75t_L   g14329(.A1(\a[56] ), .A2(new_n14273), .B(new_n13958), .C(new_n13954), .Y(new_n14586));
  O2A1O1Ixp33_ASAP7_75t_L   g14330(.A1(new_n13948), .A2(new_n13949), .B(new_n14586), .C(new_n14276), .Y(new_n14587));
  A2O1A1Ixp33_ASAP7_75t_L   g14331(.A1(new_n14586), .A2(new_n13953), .B(new_n14587), .C(new_n14275), .Y(new_n14588));
  A2O1A1O1Ixp25_ASAP7_75t_L g14332(.A1(new_n14285), .A2(\a[53] ), .B(new_n14282), .C(new_n14588), .D(new_n14587), .Y(new_n14589));
  NAND2xp33_ASAP7_75t_L     g14333(.A(new_n14589), .B(new_n14585), .Y(new_n14590));
  INVx1_ASAP7_75t_L         g14334(.A(new_n14589), .Y(new_n14591));
  A2O1A1Ixp33_ASAP7_75t_L   g14335(.A1(new_n14582), .A2(new_n14576), .B(new_n14584), .C(new_n14591), .Y(new_n14592));
  NAND2xp33_ASAP7_75t_L     g14336(.A(new_n14592), .B(new_n14590), .Y(new_n14593));
  NOR2xp33_ASAP7_75t_L      g14337(.A(new_n1745), .B(new_n10065), .Y(new_n14594));
  AOI221xp5_ASAP7_75t_L     g14338(.A1(new_n8175), .A2(\b[21] ), .B1(new_n8484), .B2(\b[19] ), .C(new_n14594), .Y(new_n14595));
  O2A1O1Ixp33_ASAP7_75t_L   g14339(.A1(new_n8176), .A2(new_n1901), .B(new_n14595), .C(new_n8172), .Y(new_n14596));
  O2A1O1Ixp33_ASAP7_75t_L   g14340(.A1(new_n8176), .A2(new_n1901), .B(new_n14595), .C(\a[50] ), .Y(new_n14597));
  INVx1_ASAP7_75t_L         g14341(.A(new_n14597), .Y(new_n14598));
  O2A1O1Ixp33_ASAP7_75t_L   g14342(.A1(new_n14596), .A2(new_n8172), .B(new_n14598), .C(new_n14593), .Y(new_n14599));
  INVx1_ASAP7_75t_L         g14343(.A(new_n14596), .Y(new_n14600));
  A2O1A1Ixp33_ASAP7_75t_L   g14344(.A1(\a[50] ), .A2(new_n14600), .B(new_n14597), .C(new_n14593), .Y(new_n14601));
  OAI21xp33_ASAP7_75t_L     g14345(.A1(new_n14593), .A2(new_n14599), .B(new_n14601), .Y(new_n14602));
  O2A1O1Ixp33_ASAP7_75t_L   g14346(.A1(new_n14292), .A2(new_n14298), .B(new_n14291), .C(new_n14602), .Y(new_n14603));
  A2O1A1O1Ixp25_ASAP7_75t_L g14347(.A1(new_n14296), .A2(\a[50] ), .B(new_n14297), .C(new_n14289), .D(new_n14290), .Y(new_n14604));
  INVx1_ASAP7_75t_L         g14348(.A(new_n14604), .Y(new_n14605));
  O2A1O1Ixp33_ASAP7_75t_L   g14349(.A1(new_n14593), .A2(new_n14599), .B(new_n14601), .C(new_n14605), .Y(new_n14606));
  NOR2xp33_ASAP7_75t_L      g14350(.A(new_n14606), .B(new_n14603), .Y(new_n14607));
  NOR2xp33_ASAP7_75t_L      g14351(.A(new_n2205), .B(new_n7318), .Y(new_n14608));
  AOI221xp5_ASAP7_75t_L     g14352(.A1(new_n7333), .A2(\b[23] ), .B1(new_n7609), .B2(\b[22] ), .C(new_n14608), .Y(new_n14609));
  O2A1O1Ixp33_ASAP7_75t_L   g14353(.A1(new_n7321), .A2(new_n2853), .B(new_n14609), .C(new_n7316), .Y(new_n14610));
  INVx1_ASAP7_75t_L         g14354(.A(new_n14610), .Y(new_n14611));
  O2A1O1Ixp33_ASAP7_75t_L   g14355(.A1(new_n7321), .A2(new_n2853), .B(new_n14609), .C(\a[47] ), .Y(new_n14612));
  AOI21xp33_ASAP7_75t_L     g14356(.A1(new_n14611), .A2(\a[47] ), .B(new_n14612), .Y(new_n14613));
  XNOR2x2_ASAP7_75t_L       g14357(.A(new_n14613), .B(new_n14607), .Y(new_n14614));
  XOR2x2_ASAP7_75t_L        g14358(.A(new_n14526), .B(new_n14614), .Y(new_n14615));
  NOR2xp33_ASAP7_75t_L      g14359(.A(new_n2377), .B(new_n6741), .Y(new_n14616));
  AOI221xp5_ASAP7_75t_L     g14360(.A1(\b[27] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[26] ), .C(new_n14616), .Y(new_n14617));
  O2A1O1Ixp33_ASAP7_75t_L   g14361(.A1(new_n6443), .A2(new_n2889), .B(new_n14617), .C(new_n6439), .Y(new_n14618));
  INVx1_ASAP7_75t_L         g14362(.A(new_n14618), .Y(new_n14619));
  O2A1O1Ixp33_ASAP7_75t_L   g14363(.A1(new_n6443), .A2(new_n2889), .B(new_n14617), .C(\a[44] ), .Y(new_n14620));
  AOI21xp33_ASAP7_75t_L     g14364(.A1(new_n14619), .A2(\a[44] ), .B(new_n14620), .Y(new_n14621));
  XNOR2x2_ASAP7_75t_L       g14365(.A(new_n14621), .B(new_n14615), .Y(new_n14622));
  INVx1_ASAP7_75t_L         g14366(.A(new_n14313), .Y(new_n14623));
  A2O1A1Ixp33_ASAP7_75t_L   g14367(.A1(\a[44] ), .A2(new_n14320), .B(new_n14321), .C(new_n14316), .Y(new_n14624));
  A2O1A1Ixp33_ASAP7_75t_L   g14368(.A1(new_n13999), .A2(new_n14314), .B(new_n14623), .C(new_n14624), .Y(new_n14625));
  XNOR2x2_ASAP7_75t_L       g14369(.A(new_n14625), .B(new_n14622), .Y(new_n14626));
  NOR2xp33_ASAP7_75t_L      g14370(.A(new_n3456), .B(new_n5641), .Y(new_n14627));
  AOI221xp5_ASAP7_75t_L     g14371(.A1(\b[28] ), .A2(new_n5920), .B1(\b[29] ), .B2(new_n5623), .C(new_n14627), .Y(new_n14628));
  O2A1O1Ixp33_ASAP7_75t_L   g14372(.A1(new_n5630), .A2(new_n3464), .B(new_n14628), .C(new_n5626), .Y(new_n14629));
  O2A1O1Ixp33_ASAP7_75t_L   g14373(.A1(new_n5630), .A2(new_n3464), .B(new_n14628), .C(\a[41] ), .Y(new_n14630));
  INVx1_ASAP7_75t_L         g14374(.A(new_n14630), .Y(new_n14631));
  OAI21xp33_ASAP7_75t_L     g14375(.A1(new_n5626), .A2(new_n14629), .B(new_n14631), .Y(new_n14632));
  INVx1_ASAP7_75t_L         g14376(.A(new_n14632), .Y(new_n14633));
  NAND2xp33_ASAP7_75t_L     g14377(.A(new_n14633), .B(new_n14626), .Y(new_n14634));
  O2A1O1Ixp33_ASAP7_75t_L   g14378(.A1(new_n14332), .A2(new_n14333), .B(new_n14325), .C(new_n14338), .Y(new_n14635));
  OR2x4_ASAP7_75t_L         g14379(.A(new_n14625), .B(new_n14622), .Y(new_n14636));
  A2O1A1Ixp33_ASAP7_75t_L   g14380(.A1(\a[44] ), .A2(new_n14619), .B(new_n14620), .C(new_n14615), .Y(new_n14637));
  INVx1_ASAP7_75t_L         g14381(.A(new_n14620), .Y(new_n14638));
  O2A1O1Ixp33_ASAP7_75t_L   g14382(.A1(new_n14618), .A2(new_n6439), .B(new_n14638), .C(new_n14615), .Y(new_n14639));
  A2O1A1Ixp33_ASAP7_75t_L   g14383(.A1(new_n14637), .A2(new_n14615), .B(new_n14639), .C(new_n14625), .Y(new_n14640));
  NAND3xp33_ASAP7_75t_L     g14384(.A(new_n14636), .B(new_n14640), .C(new_n14632), .Y(new_n14641));
  AOI21xp33_ASAP7_75t_L     g14385(.A1(new_n14634), .A2(new_n14641), .B(new_n14635), .Y(new_n14642));
  O2A1O1Ixp33_ASAP7_75t_L   g14386(.A1(new_n14629), .A2(new_n5626), .B(new_n14631), .C(new_n14626), .Y(new_n14643));
  A2O1A1O1Ixp25_ASAP7_75t_L g14387(.A1(new_n14325), .A2(new_n14339), .B(new_n14338), .C(new_n14634), .D(new_n14643), .Y(new_n14644));
  A2O1A1Ixp33_ASAP7_75t_L   g14388(.A1(new_n14644), .A2(new_n14634), .B(new_n14642), .C(new_n14524), .Y(new_n14645));
  AND3x1_ASAP7_75t_L        g14389(.A(new_n14634), .B(new_n14641), .C(new_n14635), .Y(new_n14646));
  INVx1_ASAP7_75t_L         g14390(.A(new_n14524), .Y(new_n14647));
  OA21x2_ASAP7_75t_L        g14391(.A1(new_n14642), .A2(new_n14646), .B(new_n14647), .Y(new_n14648));
  AO221x2_ASAP7_75t_L       g14392(.A1(new_n14354), .A2(new_n14345), .B1(new_n14645), .B2(new_n14524), .C(new_n14648), .Y(new_n14649));
  O2A1O1Ixp33_ASAP7_75t_L   g14393(.A1(new_n14342), .A2(new_n14343), .B(new_n14344), .C(new_n14358), .Y(new_n14650));
  A2O1A1Ixp33_ASAP7_75t_L   g14394(.A1(new_n14645), .A2(new_n14524), .B(new_n14648), .C(new_n14650), .Y(new_n14651));
  NOR2xp33_ASAP7_75t_L      g14395(.A(new_n4613), .B(new_n4147), .Y(new_n14652));
  AOI221xp5_ASAP7_75t_L     g14396(.A1(\b[34] ), .A2(new_n4402), .B1(\b[35] ), .B2(new_n4155), .C(new_n14652), .Y(new_n14653));
  O2A1O1Ixp33_ASAP7_75t_L   g14397(.A1(new_n4150), .A2(new_n4622), .B(new_n14653), .C(new_n4145), .Y(new_n14654));
  NOR2xp33_ASAP7_75t_L      g14398(.A(new_n4145), .B(new_n14654), .Y(new_n14655));
  O2A1O1Ixp33_ASAP7_75t_L   g14399(.A1(new_n4150), .A2(new_n4622), .B(new_n14653), .C(\a[35] ), .Y(new_n14656));
  NOR2xp33_ASAP7_75t_L      g14400(.A(new_n14656), .B(new_n14655), .Y(new_n14657));
  AO21x2_ASAP7_75t_L        g14401(.A1(new_n14649), .A2(new_n14651), .B(new_n14657), .Y(new_n14658));
  NAND3xp33_ASAP7_75t_L     g14402(.A(new_n14651), .B(new_n14649), .C(new_n14657), .Y(new_n14659));
  AOI21xp33_ASAP7_75t_L     g14403(.A1(new_n14658), .A2(new_n14659), .B(new_n14518), .Y(new_n14660));
  AOI21xp33_ASAP7_75t_L     g14404(.A1(new_n14651), .A2(new_n14649), .B(new_n14657), .Y(new_n14661));
  AND3x1_ASAP7_75t_L        g14405(.A(new_n14651), .B(new_n14649), .C(new_n14657), .Y(new_n14662));
  NOR3xp33_ASAP7_75t_L      g14406(.A(new_n14662), .B(new_n14661), .C(new_n14517), .Y(new_n14663));
  NOR2xp33_ASAP7_75t_L      g14407(.A(new_n14660), .B(new_n14663), .Y(new_n14664));
  OAI22xp33_ASAP7_75t_L     g14408(.A1(new_n3703), .A2(new_n5074), .B1(new_n5311), .B2(new_n3509), .Y(new_n14665));
  AOI221xp5_ASAP7_75t_L     g14409(.A1(new_n3503), .A2(\b[39] ), .B1(new_n3505), .B2(new_n11869), .C(new_n14665), .Y(new_n14666));
  XNOR2x2_ASAP7_75t_L       g14410(.A(new_n3493), .B(new_n14666), .Y(new_n14667));
  INVx1_ASAP7_75t_L         g14411(.A(new_n14667), .Y(new_n14668));
  O2A1O1Ixp33_ASAP7_75t_L   g14412(.A1(new_n13768), .A2(new_n13772), .B(new_n13774), .C(new_n14370), .Y(new_n14669));
  A2O1A1Ixp33_ASAP7_75t_L   g14413(.A1(new_n13776), .A2(new_n13774), .B(new_n14669), .C(new_n14051), .Y(new_n14670));
  A2O1A1Ixp33_ASAP7_75t_L   g14414(.A1(new_n14670), .A2(new_n14054), .B(new_n14669), .C(new_n14377), .Y(new_n14671));
  A2O1A1Ixp33_ASAP7_75t_L   g14415(.A1(new_n14367), .A2(new_n14368), .B(new_n14378), .C(new_n14671), .Y(new_n14672));
  NOR2xp33_ASAP7_75t_L      g14416(.A(new_n14668), .B(new_n14672), .Y(new_n14673));
  INVx1_ASAP7_75t_L         g14417(.A(new_n14673), .Y(new_n14674));
  A2O1A1O1Ixp25_ASAP7_75t_L g14418(.A1(new_n14368), .A2(new_n14367), .B(new_n14378), .C(new_n14671), .D(new_n14667), .Y(new_n14675));
  INVx1_ASAP7_75t_L         g14419(.A(new_n14675), .Y(new_n14676));
  NAND3xp33_ASAP7_75t_L     g14420(.A(new_n14674), .B(new_n14664), .C(new_n14676), .Y(new_n14677));
  OAI21xp33_ASAP7_75t_L     g14421(.A1(new_n14661), .A2(new_n14662), .B(new_n14517), .Y(new_n14678));
  NAND3xp33_ASAP7_75t_L     g14422(.A(new_n14658), .B(new_n14518), .C(new_n14659), .Y(new_n14679));
  NAND2xp33_ASAP7_75t_L     g14423(.A(new_n14679), .B(new_n14678), .Y(new_n14680));
  OAI21xp33_ASAP7_75t_L     g14424(.A1(new_n14673), .A2(new_n14675), .B(new_n14680), .Y(new_n14681));
  AND2x2_ASAP7_75t_L        g14425(.A(new_n14681), .B(new_n14677), .Y(new_n14682));
  NAND3xp33_ASAP7_75t_L     g14426(.A(new_n14682), .B(new_n14515), .C(new_n14513), .Y(new_n14683));
  INVx1_ASAP7_75t_L         g14427(.A(new_n14513), .Y(new_n14684));
  INVx1_ASAP7_75t_L         g14428(.A(new_n14515), .Y(new_n14685));
  NAND2xp33_ASAP7_75t_L     g14429(.A(new_n14681), .B(new_n14677), .Y(new_n14686));
  OAI21xp33_ASAP7_75t_L     g14430(.A1(new_n14684), .A2(new_n14685), .B(new_n14686), .Y(new_n14687));
  NAND2xp33_ASAP7_75t_L     g14431(.A(new_n14687), .B(new_n14683), .Y(new_n14688));
  A2O1A1Ixp33_ASAP7_75t_L   g14432(.A1(new_n14505), .A2(new_n14503), .B(new_n14508), .C(new_n14688), .Y(new_n14689));
  INVx1_ASAP7_75t_L         g14433(.A(new_n14508), .Y(new_n14690));
  O2A1O1Ixp33_ASAP7_75t_L   g14434(.A1(new_n14408), .A2(new_n14405), .B(new_n14492), .C(new_n14407), .Y(new_n14691));
  NAND2xp33_ASAP7_75t_L     g14435(.A(new_n14503), .B(new_n14691), .Y(new_n14692));
  NOR3xp33_ASAP7_75t_L      g14436(.A(new_n14686), .B(new_n14685), .C(new_n14684), .Y(new_n14693));
  AOI21xp33_ASAP7_75t_L     g14437(.A1(new_n14515), .A2(new_n14513), .B(new_n14682), .Y(new_n14694));
  NOR2xp33_ASAP7_75t_L      g14438(.A(new_n14693), .B(new_n14694), .Y(new_n14695));
  NAND3xp33_ASAP7_75t_L     g14439(.A(new_n14695), .B(new_n14692), .C(new_n14690), .Y(new_n14696));
  NAND2xp33_ASAP7_75t_L     g14440(.A(new_n14696), .B(new_n14689), .Y(new_n14697));
  NAND3xp33_ASAP7_75t_L     g14441(.A(new_n14697), .B(new_n14498), .C(new_n14496), .Y(new_n14698));
  AOI22xp33_ASAP7_75t_L     g14442(.A1(new_n14689), .A2(new_n14696), .B1(new_n14498), .B2(new_n14496), .Y(new_n14699));
  AOI21xp33_ASAP7_75t_L     g14443(.A1(new_n14499), .A2(new_n14698), .B(new_n14699), .Y(new_n14700));
  O2A1O1Ixp33_ASAP7_75t_L   g14444(.A1(new_n14212), .A2(new_n14089), .B(new_n14097), .C(new_n14088), .Y(new_n14701));
  A2O1A1Ixp33_ASAP7_75t_L   g14445(.A1(new_n14207), .A2(\a[20] ), .B(new_n14208), .C(new_n14701), .Y(new_n14702));
  A2O1A1Ixp33_ASAP7_75t_L   g14446(.A1(new_n14092), .A2(new_n14097), .B(new_n14088), .C(new_n14210), .Y(new_n14703));
  OAI22xp33_ASAP7_75t_L     g14447(.A1(new_n1654), .A2(new_n8427), .B1(new_n8755), .B2(new_n1517), .Y(new_n14704));
  AOI221xp5_ASAP7_75t_L     g14448(.A1(new_n1511), .A2(\b[51] ), .B1(new_n1513), .B2(new_n8790), .C(new_n14704), .Y(new_n14705));
  XNOR2x2_ASAP7_75t_L       g14449(.A(new_n1501), .B(new_n14705), .Y(new_n14706));
  A2O1A1O1Ixp25_ASAP7_75t_L g14450(.A1(new_n14702), .A2(new_n14703), .B(new_n14414), .C(new_n14210), .D(new_n14706), .Y(new_n14707));
  INVx1_ASAP7_75t_L         g14451(.A(new_n14706), .Y(new_n14708));
  A2O1A1Ixp33_ASAP7_75t_L   g14452(.A1(new_n14703), .A2(new_n14702), .B(new_n14414), .C(new_n14210), .Y(new_n14709));
  NOR2xp33_ASAP7_75t_L      g14453(.A(new_n14708), .B(new_n14709), .Y(new_n14710));
  NOR2xp33_ASAP7_75t_L      g14454(.A(new_n14707), .B(new_n14710), .Y(new_n14711));
  XOR2x2_ASAP7_75t_L        g14455(.A(new_n14700), .B(new_n14711), .Y(new_n14712));
  XOR2x2_ASAP7_75t_L        g14456(.A(new_n14414), .B(new_n14215), .Y(new_n14713));
  AOI21xp33_ASAP7_75t_L     g14457(.A1(new_n14713), .A2(new_n14202), .B(new_n14199), .Y(new_n14714));
  OAI22xp33_ASAP7_75t_L     g14458(.A1(new_n1285), .A2(new_n9355), .B1(new_n9683), .B2(new_n2118), .Y(new_n14715));
  AOI221xp5_ASAP7_75t_L     g14459(.A1(new_n1209), .A2(\b[54] ), .B1(new_n1216), .B2(new_n9717), .C(new_n14715), .Y(new_n14716));
  XNOR2x2_ASAP7_75t_L       g14460(.A(new_n1206), .B(new_n14716), .Y(new_n14717));
  INVx1_ASAP7_75t_L         g14461(.A(new_n14717), .Y(new_n14718));
  A2O1A1Ixp33_ASAP7_75t_L   g14462(.A1(new_n14713), .A2(new_n14202), .B(new_n14199), .C(new_n14718), .Y(new_n14719));
  INVx1_ASAP7_75t_L         g14463(.A(new_n14719), .Y(new_n14720));
  NAND2xp33_ASAP7_75t_L     g14464(.A(new_n14718), .B(new_n14714), .Y(new_n14721));
  O2A1O1Ixp33_ASAP7_75t_L   g14465(.A1(new_n14714), .A2(new_n14720), .B(new_n14721), .C(new_n14712), .Y(new_n14722));
  O2A1O1Ixp33_ASAP7_75t_L   g14466(.A1(new_n14203), .A2(new_n14415), .B(new_n14200), .C(new_n14718), .Y(new_n14723));
  A2O1A1Ixp33_ASAP7_75t_L   g14467(.A1(new_n14719), .A2(new_n14718), .B(new_n14723), .C(new_n14712), .Y(new_n14724));
  OAI21xp33_ASAP7_75t_L     g14468(.A1(new_n14712), .A2(new_n14722), .B(new_n14724), .Y(new_n14725));
  OAI22xp33_ASAP7_75t_L     g14469(.A1(new_n980), .A2(new_n10309), .B1(new_n10332), .B2(new_n864), .Y(new_n14726));
  AOI221xp5_ASAP7_75t_L     g14470(.A1(new_n886), .A2(\b[57] ), .B1(new_n873), .B2(new_n10991), .C(new_n14726), .Y(new_n14727));
  XNOR2x2_ASAP7_75t_L       g14471(.A(new_n867), .B(new_n14727), .Y(new_n14728));
  A2O1A1O1Ixp25_ASAP7_75t_L g14472(.A1(new_n14421), .A2(new_n14192), .B(new_n14416), .C(new_n14194), .D(new_n14728), .Y(new_n14729));
  INVx1_ASAP7_75t_L         g14473(.A(new_n14728), .Y(new_n14730));
  A2O1A1Ixp33_ASAP7_75t_L   g14474(.A1(new_n14192), .A2(new_n14421), .B(new_n14416), .C(new_n14194), .Y(new_n14731));
  NOR2xp33_ASAP7_75t_L      g14475(.A(new_n14730), .B(new_n14731), .Y(new_n14732));
  OAI21xp33_ASAP7_75t_L     g14476(.A1(new_n14732), .A2(new_n14729), .B(new_n14725), .Y(new_n14733));
  XNOR2x2_ASAP7_75t_L       g14477(.A(new_n14700), .B(new_n14711), .Y(new_n14734));
  A2O1A1Ixp33_ASAP7_75t_L   g14478(.A1(new_n14719), .A2(new_n14718), .B(new_n14723), .C(new_n14734), .Y(new_n14735));
  INVx1_ASAP7_75t_L         g14479(.A(new_n14723), .Y(new_n14736));
  O2A1O1Ixp33_ASAP7_75t_L   g14480(.A1(new_n14717), .A2(new_n14720), .B(new_n14736), .C(new_n14734), .Y(new_n14737));
  AOI21xp33_ASAP7_75t_L     g14481(.A1(new_n14735), .A2(new_n14734), .B(new_n14737), .Y(new_n14738));
  INVx1_ASAP7_75t_L         g14482(.A(new_n14729), .Y(new_n14739));
  O2A1O1Ixp33_ASAP7_75t_L   g14483(.A1(new_n14195), .A2(new_n14191), .B(new_n14422), .C(new_n14193), .Y(new_n14740));
  NAND2xp33_ASAP7_75t_L     g14484(.A(new_n14728), .B(new_n14740), .Y(new_n14741));
  NAND3xp33_ASAP7_75t_L     g14485(.A(new_n14738), .B(new_n14741), .C(new_n14739), .Y(new_n14742));
  NAND2xp33_ASAP7_75t_L     g14486(.A(new_n14733), .B(new_n14742), .Y(new_n14743));
  NOR3xp33_ASAP7_75t_L      g14487(.A(new_n14743), .B(new_n14485), .C(new_n14484), .Y(new_n14744));
  NOR2xp33_ASAP7_75t_L      g14488(.A(new_n14485), .B(new_n14484), .Y(new_n14745));
  NAND2xp33_ASAP7_75t_L     g14489(.A(new_n14741), .B(new_n14739), .Y(new_n14746));
  O2A1O1Ixp33_ASAP7_75t_L   g14490(.A1(new_n14712), .A2(new_n14722), .B(new_n14724), .C(new_n14746), .Y(new_n14747));
  O2A1O1Ixp33_ASAP7_75t_L   g14491(.A1(new_n14738), .A2(new_n14747), .B(new_n14742), .C(new_n14745), .Y(new_n14748));
  NOR2xp33_ASAP7_75t_L      g14492(.A(new_n14748), .B(new_n14744), .Y(new_n14749));
  A2O1A1Ixp33_ASAP7_75t_L   g14493(.A1(new_n14477), .A2(new_n14474), .B(new_n14478), .C(new_n14749), .Y(new_n14750));
  AO21x2_ASAP7_75t_L        g14494(.A1(new_n14424), .A2(new_n14432), .B(new_n14434), .Y(new_n14751));
  A2O1A1O1Ixp25_ASAP7_75t_L g14495(.A1(new_n14131), .A2(new_n14128), .B(new_n14124), .C(new_n14133), .D(new_n14457), .Y(new_n14752));
  O2A1O1Ixp33_ASAP7_75t_L   g14496(.A1(new_n14457), .A2(new_n14752), .B(new_n14751), .C(new_n14436), .Y(new_n14753));
  NAND2xp33_ASAP7_75t_L     g14497(.A(new_n14474), .B(new_n14753), .Y(new_n14754));
  OAI221xp5_ASAP7_75t_L     g14498(.A1(new_n14476), .A2(new_n14753), .B1(new_n14744), .B2(new_n14748), .C(new_n14754), .Y(new_n14755));
  NAND2xp33_ASAP7_75t_L     g14499(.A(new_n14750), .B(new_n14755), .Y(new_n14756));
  XNOR2x2_ASAP7_75t_L       g14500(.A(new_n14470), .B(new_n14756), .Y(new_n14757));
  A2O1A1Ixp33_ASAP7_75t_L   g14501(.A1(new_n14467), .A2(new_n14461), .B(new_n14469), .C(new_n14757), .Y(new_n14758));
  INVx1_ASAP7_75t_L         g14502(.A(new_n14758), .Y(new_n14759));
  A2O1A1Ixp33_ASAP7_75t_L   g14503(.A1(new_n14148), .A2(new_n14161), .B(new_n14165), .C(new_n14461), .Y(new_n14760));
  A2O1A1Ixp33_ASAP7_75t_L   g14504(.A1(new_n14152), .A2(new_n14138), .B(new_n14468), .C(new_n14760), .Y(new_n14761));
  NOR2xp33_ASAP7_75t_L      g14505(.A(new_n14757), .B(new_n14761), .Y(new_n14762));
  NOR2xp33_ASAP7_75t_L      g14506(.A(new_n14759), .B(new_n14762), .Y(\f[69] ));
  INVx1_ASAP7_75t_L         g14507(.A(new_n12269), .Y(new_n14764));
  NOR2xp33_ASAP7_75t_L      g14508(.A(new_n11591), .B(new_n712), .Y(new_n14765));
  AOI221xp5_ASAP7_75t_L     g14509(.A1(\b[61] ), .A2(new_n640), .B1(new_n635), .B2(\b[60] ), .C(new_n14765), .Y(new_n14766));
  O2A1O1Ixp33_ASAP7_75t_L   g14510(.A1(new_n641), .A2(new_n14764), .B(new_n14766), .C(new_n637), .Y(new_n14767));
  O2A1O1Ixp33_ASAP7_75t_L   g14511(.A1(new_n641), .A2(new_n14764), .B(new_n14766), .C(\a[11] ), .Y(new_n14768));
  INVx1_ASAP7_75t_L         g14512(.A(new_n14768), .Y(new_n14769));
  A2O1A1O1Ixp25_ASAP7_75t_L g14513(.A1(new_n14735), .A2(new_n14734), .B(new_n14737), .C(new_n14741), .D(new_n14729), .Y(new_n14770));
  OAI211xp5_ASAP7_75t_L     g14514(.A1(new_n637), .A2(new_n14767), .B(new_n14770), .C(new_n14769), .Y(new_n14771));
  OAI21xp33_ASAP7_75t_L     g14515(.A1(new_n637), .A2(new_n14767), .B(new_n14769), .Y(new_n14772));
  A2O1A1Ixp33_ASAP7_75t_L   g14516(.A1(new_n14725), .A2(new_n14741), .B(new_n14729), .C(new_n14772), .Y(new_n14773));
  NAND2xp33_ASAP7_75t_L     g14517(.A(\b[57] ), .B(new_n885), .Y(new_n14774));
  OAI221xp5_ASAP7_75t_L     g14518(.A1(new_n869), .A2(new_n11303), .B1(new_n10332), .B2(new_n980), .C(new_n14774), .Y(new_n14775));
  AOI21xp33_ASAP7_75t_L     g14519(.A1(new_n11314), .A2(new_n873), .B(new_n14775), .Y(new_n14776));
  NAND2xp33_ASAP7_75t_L     g14520(.A(\a[14] ), .B(new_n14776), .Y(new_n14777));
  A2O1A1Ixp33_ASAP7_75t_L   g14521(.A1(new_n11314), .A2(new_n873), .B(new_n14775), .C(new_n867), .Y(new_n14778));
  AND2x2_ASAP7_75t_L        g14522(.A(new_n14778), .B(new_n14777), .Y(new_n14779));
  A2O1A1O1Ixp25_ASAP7_75t_L g14523(.A1(new_n14714), .A2(new_n14721), .B(new_n14712), .C(new_n14719), .D(new_n14779), .Y(new_n14780));
  INVx1_ASAP7_75t_L         g14524(.A(new_n14780), .Y(new_n14781));
  NAND3xp33_ASAP7_75t_L     g14525(.A(new_n14735), .B(new_n14719), .C(new_n14779), .Y(new_n14782));
  NAND2xp33_ASAP7_75t_L     g14526(.A(new_n14782), .B(new_n14781), .Y(new_n14783));
  NAND2xp33_ASAP7_75t_L     g14527(.A(\b[54] ), .B(new_n1204), .Y(new_n14784));
  OAI221xp5_ASAP7_75t_L     g14528(.A1(new_n1284), .A2(new_n10309), .B1(new_n9683), .B2(new_n1285), .C(new_n14784), .Y(new_n14785));
  A2O1A1Ixp33_ASAP7_75t_L   g14529(.A1(new_n10320), .A2(new_n1216), .B(new_n14785), .C(\a[17] ), .Y(new_n14786));
  NAND2xp33_ASAP7_75t_L     g14530(.A(\a[17] ), .B(new_n14786), .Y(new_n14787));
  A2O1A1Ixp33_ASAP7_75t_L   g14531(.A1(new_n10320), .A2(new_n1216), .B(new_n14785), .C(new_n1206), .Y(new_n14788));
  NAND2xp33_ASAP7_75t_L     g14532(.A(new_n14788), .B(new_n14787), .Y(new_n14789));
  A2O1A1O1Ixp25_ASAP7_75t_L g14533(.A1(new_n14698), .A2(new_n14499), .B(new_n14699), .C(new_n14711), .D(new_n14707), .Y(new_n14790));
  XNOR2x2_ASAP7_75t_L       g14534(.A(new_n14789), .B(new_n14790), .Y(new_n14791));
  NAND2xp33_ASAP7_75t_L     g14535(.A(\b[51] ), .B(new_n1507), .Y(new_n14792));
  OAI221xp5_ASAP7_75t_L     g14536(.A1(new_n1518), .A2(new_n9355), .B1(new_n8755), .B2(new_n1654), .C(new_n14792), .Y(new_n14793));
  A2O1A1Ixp33_ASAP7_75t_L   g14537(.A1(new_n9367), .A2(new_n1513), .B(new_n14793), .C(\a[20] ), .Y(new_n14794));
  NAND2xp33_ASAP7_75t_L     g14538(.A(\a[20] ), .B(new_n14794), .Y(new_n14795));
  A2O1A1Ixp33_ASAP7_75t_L   g14539(.A1(new_n9367), .A2(new_n1513), .B(new_n14793), .C(new_n1501), .Y(new_n14796));
  NAND2xp33_ASAP7_75t_L     g14540(.A(new_n14796), .B(new_n14795), .Y(new_n14797));
  A2O1A1Ixp33_ASAP7_75t_L   g14541(.A1(new_n14490), .A2(new_n14489), .B(new_n14495), .C(new_n14698), .Y(new_n14798));
  XOR2x2_ASAP7_75t_L        g14542(.A(new_n14797), .B(new_n14798), .Y(new_n14799));
  O2A1O1Ixp33_ASAP7_75t_L   g14543(.A1(new_n14502), .A2(new_n14504), .B(new_n14690), .C(new_n14688), .Y(new_n14800));
  INVx1_ASAP7_75t_L         g14544(.A(new_n14800), .Y(new_n14801));
  INVx1_ASAP7_75t_L         g14545(.A(new_n8438), .Y(new_n14802));
  NOR2xp33_ASAP7_75t_L      g14546(.A(new_n7860), .B(new_n1962), .Y(new_n14803));
  AOI221xp5_ASAP7_75t_L     g14547(.A1(new_n1955), .A2(\b[49] ), .B1(new_n2093), .B2(\b[47] ), .C(new_n14803), .Y(new_n14804));
  O2A1O1Ixp33_ASAP7_75t_L   g14548(.A1(new_n1956), .A2(new_n14802), .B(new_n14804), .C(new_n1952), .Y(new_n14805));
  O2A1O1Ixp33_ASAP7_75t_L   g14549(.A1(new_n1956), .A2(new_n14802), .B(new_n14804), .C(\a[23] ), .Y(new_n14806));
  INVx1_ASAP7_75t_L         g14550(.A(new_n14806), .Y(new_n14807));
  O2A1O1Ixp33_ASAP7_75t_L   g14551(.A1(new_n14508), .A2(new_n14503), .B(new_n14695), .C(new_n14504), .Y(new_n14808));
  O2A1O1Ixp33_ASAP7_75t_L   g14552(.A1(new_n1952), .A2(new_n14805), .B(new_n14807), .C(new_n14808), .Y(new_n14809));
  INVx1_ASAP7_75t_L         g14553(.A(new_n14805), .Y(new_n14810));
  A2O1A1Ixp33_ASAP7_75t_L   g14554(.A1(new_n14810), .A2(\a[23] ), .B(new_n14806), .C(new_n14808), .Y(new_n14811));
  A2O1A1Ixp33_ASAP7_75t_L   g14555(.A1(new_n14801), .A2(new_n14505), .B(new_n14809), .C(new_n14811), .Y(new_n14812));
  NAND2xp33_ASAP7_75t_L     g14556(.A(\b[45] ), .B(new_n2421), .Y(new_n14813));
  OAI221xp5_ASAP7_75t_L     g14557(.A1(new_n2415), .A2(new_n7270), .B1(new_n6944), .B2(new_n2572), .C(new_n14813), .Y(new_n14814));
  AOI21xp33_ASAP7_75t_L     g14558(.A1(new_n7278), .A2(new_n2417), .B(new_n14814), .Y(new_n14815));
  NAND2xp33_ASAP7_75t_L     g14559(.A(\a[26] ), .B(new_n14815), .Y(new_n14816));
  A2O1A1Ixp33_ASAP7_75t_L   g14560(.A1(new_n7278), .A2(new_n2417), .B(new_n14814), .C(new_n2413), .Y(new_n14817));
  AND2x2_ASAP7_75t_L        g14561(.A(new_n14817), .B(new_n14816), .Y(new_n14818));
  O2A1O1Ixp33_ASAP7_75t_L   g14562(.A1(new_n14684), .A2(new_n14686), .B(new_n14515), .C(new_n14818), .Y(new_n14819));
  INVx1_ASAP7_75t_L         g14563(.A(new_n14819), .Y(new_n14820));
  NAND3xp33_ASAP7_75t_L     g14564(.A(new_n14683), .B(new_n14515), .C(new_n14818), .Y(new_n14821));
  NAND2xp33_ASAP7_75t_L     g14565(.A(new_n14820), .B(new_n14821), .Y(new_n14822));
  NOR2xp33_ASAP7_75t_L      g14566(.A(new_n6671), .B(new_n2930), .Y(new_n14823));
  AOI221xp5_ASAP7_75t_L     g14567(.A1(\b[41] ), .A2(new_n3129), .B1(\b[42] ), .B2(new_n2936), .C(new_n14823), .Y(new_n14824));
  O2A1O1Ixp33_ASAP7_75t_L   g14568(.A1(new_n2940), .A2(new_n6679), .B(new_n14824), .C(new_n2928), .Y(new_n14825));
  O2A1O1Ixp33_ASAP7_75t_L   g14569(.A1(new_n2940), .A2(new_n6679), .B(new_n14824), .C(\a[29] ), .Y(new_n14826));
  INVx1_ASAP7_75t_L         g14570(.A(new_n14826), .Y(new_n14827));
  AOI21xp33_ASAP7_75t_L     g14571(.A1(new_n14674), .A2(new_n14664), .B(new_n14675), .Y(new_n14828));
  O2A1O1Ixp33_ASAP7_75t_L   g14572(.A1(new_n2928), .A2(new_n14825), .B(new_n14827), .C(new_n14828), .Y(new_n14829));
  INVx1_ASAP7_75t_L         g14573(.A(new_n14825), .Y(new_n14830));
  A2O1A1Ixp33_ASAP7_75t_L   g14574(.A1(new_n14830), .A2(\a[29] ), .B(new_n14826), .C(new_n14828), .Y(new_n14831));
  A2O1A1Ixp33_ASAP7_75t_L   g14575(.A1(new_n14677), .A2(new_n14676), .B(new_n14829), .C(new_n14831), .Y(new_n14832));
  NOR2xp33_ASAP7_75t_L      g14576(.A(new_n5855), .B(new_n3510), .Y(new_n14833));
  AOI221xp5_ASAP7_75t_L     g14577(.A1(\b[38] ), .A2(new_n3708), .B1(\b[39] ), .B2(new_n3499), .C(new_n14833), .Y(new_n14834));
  O2A1O1Ixp33_ASAP7_75t_L   g14578(.A1(new_n3513), .A2(new_n5862), .B(new_n14834), .C(new_n3493), .Y(new_n14835));
  NOR2xp33_ASAP7_75t_L      g14579(.A(new_n3493), .B(new_n14835), .Y(new_n14836));
  O2A1O1Ixp33_ASAP7_75t_L   g14580(.A1(new_n3513), .A2(new_n5862), .B(new_n14834), .C(\a[32] ), .Y(new_n14837));
  NOR2xp33_ASAP7_75t_L      g14581(.A(new_n14837), .B(new_n14836), .Y(new_n14838));
  INVx1_ASAP7_75t_L         g14582(.A(new_n14838), .Y(new_n14839));
  A2O1A1Ixp33_ASAP7_75t_L   g14583(.A1(new_n14651), .A2(new_n14649), .B(new_n14657), .C(new_n14679), .Y(new_n14840));
  NOR2xp33_ASAP7_75t_L      g14584(.A(new_n14839), .B(new_n14840), .Y(new_n14841));
  O2A1O1Ixp33_ASAP7_75t_L   g14585(.A1(new_n14517), .A2(new_n14662), .B(new_n14658), .C(new_n14838), .Y(new_n14842));
  NOR2xp33_ASAP7_75t_L      g14586(.A(new_n14842), .B(new_n14841), .Y(new_n14843));
  NOR2xp33_ASAP7_75t_L      g14587(.A(new_n5074), .B(new_n4147), .Y(new_n14844));
  AOI221xp5_ASAP7_75t_L     g14588(.A1(\b[35] ), .A2(new_n4402), .B1(\b[36] ), .B2(new_n4155), .C(new_n14844), .Y(new_n14845));
  O2A1O1Ixp33_ASAP7_75t_L   g14589(.A1(new_n4150), .A2(new_n5083), .B(new_n14845), .C(new_n4145), .Y(new_n14846));
  NOR2xp33_ASAP7_75t_L      g14590(.A(new_n4145), .B(new_n14846), .Y(new_n14847));
  O2A1O1Ixp33_ASAP7_75t_L   g14591(.A1(new_n4150), .A2(new_n5083), .B(new_n14845), .C(\a[35] ), .Y(new_n14848));
  NOR2xp33_ASAP7_75t_L      g14592(.A(new_n14848), .B(new_n14847), .Y(new_n14849));
  INVx1_ASAP7_75t_L         g14593(.A(new_n14849), .Y(new_n14850));
  INVx1_ASAP7_75t_L         g14594(.A(new_n14648), .Y(new_n14851));
  A2O1A1Ixp33_ASAP7_75t_L   g14595(.A1(new_n14851), .A2(new_n14647), .B(new_n14650), .C(new_n14645), .Y(new_n14852));
  NOR2xp33_ASAP7_75t_L      g14596(.A(new_n4344), .B(new_n4908), .Y(new_n14853));
  AOI221xp5_ASAP7_75t_L     g14597(.A1(\b[32] ), .A2(new_n5139), .B1(\b[33] ), .B2(new_n4916), .C(new_n14853), .Y(new_n14854));
  O2A1O1Ixp33_ASAP7_75t_L   g14598(.A1(new_n4911), .A2(new_n4352), .B(new_n14854), .C(new_n4906), .Y(new_n14855));
  INVx1_ASAP7_75t_L         g14599(.A(new_n14855), .Y(new_n14856));
  O2A1O1Ixp33_ASAP7_75t_L   g14600(.A1(new_n4911), .A2(new_n4352), .B(new_n14854), .C(\a[38] ), .Y(new_n14857));
  NOR2xp33_ASAP7_75t_L      g14601(.A(new_n1043), .B(new_n10388), .Y(new_n14858));
  AOI221xp5_ASAP7_75t_L     g14602(.A1(new_n10086), .A2(\b[16] ), .B1(new_n11361), .B2(\b[14] ), .C(new_n14858), .Y(new_n14859));
  O2A1O1Ixp33_ASAP7_75t_L   g14603(.A1(new_n10088), .A2(new_n1161), .B(new_n14859), .C(new_n10083), .Y(new_n14860));
  INVx1_ASAP7_75t_L         g14604(.A(new_n14860), .Y(new_n14861));
  O2A1O1Ixp33_ASAP7_75t_L   g14605(.A1(new_n10088), .A2(new_n1161), .B(new_n14859), .C(\a[56] ), .Y(new_n14862));
  A2O1A1O1Ixp25_ASAP7_75t_L g14606(.A1(\a[62] ), .A2(new_n14235), .B(new_n14236), .C(new_n14239), .D(new_n14229), .Y(new_n14863));
  INVx1_ASAP7_75t_L         g14607(.A(new_n14532), .Y(new_n14864));
  NOR2xp33_ASAP7_75t_L      g14608(.A(new_n427), .B(new_n13030), .Y(new_n14865));
  O2A1O1Ixp33_ASAP7_75t_L   g14609(.A1(new_n12669), .A2(new_n12671), .B(\b[7] ), .C(new_n14865), .Y(new_n14866));
  INVx1_ASAP7_75t_L         g14610(.A(new_n14866), .Y(new_n14867));
  O2A1O1Ixp33_ASAP7_75t_L   g14611(.A1(\a[2] ), .A2(\a[5] ), .B(new_n14864), .C(new_n14867), .Y(new_n14868));
  INVx1_ASAP7_75t_L         g14612(.A(new_n14868), .Y(new_n14869));
  AOI21xp33_ASAP7_75t_L     g14613(.A1(new_n346), .A2(new_n257), .B(new_n14532), .Y(new_n14870));
  A2O1A1Ixp33_ASAP7_75t_L   g14614(.A1(\b[7] ), .A2(new_n13028), .B(new_n14865), .C(new_n14870), .Y(new_n14871));
  NAND2xp33_ASAP7_75t_L     g14615(.A(new_n14871), .B(new_n14869), .Y(new_n14872));
  NAND2xp33_ASAP7_75t_L     g14616(.A(\b[10] ), .B(new_n11995), .Y(new_n14873));
  OAI221xp5_ASAP7_75t_L     g14617(.A1(new_n12318), .A2(new_n590), .B1(new_n534), .B2(new_n12320), .C(new_n14873), .Y(new_n14874));
  AOI21xp33_ASAP7_75t_L     g14618(.A1(new_n690), .A2(new_n11997), .B(new_n14874), .Y(new_n14875));
  NAND2xp33_ASAP7_75t_L     g14619(.A(\a[62] ), .B(new_n14875), .Y(new_n14876));
  A2O1A1Ixp33_ASAP7_75t_L   g14620(.A1(new_n690), .A2(new_n11997), .B(new_n14874), .C(new_n11987), .Y(new_n14877));
  NAND2xp33_ASAP7_75t_L     g14621(.A(new_n14877), .B(new_n14876), .Y(new_n14878));
  XNOR2x2_ASAP7_75t_L       g14622(.A(new_n14872), .B(new_n14878), .Y(new_n14879));
  INVx1_ASAP7_75t_L         g14623(.A(new_n14879), .Y(new_n14880));
  O2A1O1Ixp33_ASAP7_75t_L   g14624(.A1(new_n14863), .A2(new_n14538), .B(new_n14546), .C(new_n14880), .Y(new_n14881));
  A2O1A1Ixp33_ASAP7_75t_L   g14625(.A1(new_n14240), .A2(new_n14237), .B(new_n14538), .C(new_n14546), .Y(new_n14882));
  NOR2xp33_ASAP7_75t_L      g14626(.A(new_n14879), .B(new_n14882), .Y(new_n14883));
  NOR2xp33_ASAP7_75t_L      g14627(.A(new_n14883), .B(new_n14881), .Y(new_n14884));
  NOR2xp33_ASAP7_75t_L      g14628(.A(new_n748), .B(new_n11354), .Y(new_n14885));
  AOI221xp5_ASAP7_75t_L     g14629(.A1(\b[13] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[12] ), .C(new_n14885), .Y(new_n14886));
  O2A1O1Ixp33_ASAP7_75t_L   g14630(.A1(new_n11053), .A2(new_n942), .B(new_n14886), .C(new_n11048), .Y(new_n14887));
  INVx1_ASAP7_75t_L         g14631(.A(new_n14887), .Y(new_n14888));
  O2A1O1Ixp33_ASAP7_75t_L   g14632(.A1(new_n11053), .A2(new_n942), .B(new_n14886), .C(\a[59] ), .Y(new_n14889));
  A2O1A1Ixp33_ASAP7_75t_L   g14633(.A1(\a[59] ), .A2(new_n14888), .B(new_n14889), .C(new_n14884), .Y(new_n14890));
  INVx1_ASAP7_75t_L         g14634(.A(new_n14889), .Y(new_n14891));
  O2A1O1Ixp33_ASAP7_75t_L   g14635(.A1(new_n14887), .A2(new_n11048), .B(new_n14891), .C(new_n14884), .Y(new_n14892));
  AOI21xp33_ASAP7_75t_L     g14636(.A1(new_n14890), .A2(new_n14884), .B(new_n14892), .Y(new_n14893));
  INVx1_ASAP7_75t_L         g14637(.A(new_n14556), .Y(new_n14894));
  O2A1O1Ixp33_ASAP7_75t_L   g14638(.A1(new_n14894), .A2(new_n14553), .B(new_n14559), .C(new_n14555), .Y(new_n14895));
  NAND2xp33_ASAP7_75t_L     g14639(.A(new_n14895), .B(new_n14893), .Y(new_n14896));
  A2O1A1O1Ixp25_ASAP7_75t_L g14640(.A1(new_n14556), .A2(new_n14547), .B(new_n14528), .C(new_n14554), .D(new_n14893), .Y(new_n14897));
  INVx1_ASAP7_75t_L         g14641(.A(new_n14897), .Y(new_n14898));
  NAND2xp33_ASAP7_75t_L     g14642(.A(new_n14896), .B(new_n14898), .Y(new_n14899));
  INVx1_ASAP7_75t_L         g14643(.A(new_n14862), .Y(new_n14900));
  O2A1O1Ixp33_ASAP7_75t_L   g14644(.A1(new_n14860), .A2(new_n10083), .B(new_n14900), .C(new_n14899), .Y(new_n14901));
  INVx1_ASAP7_75t_L         g14645(.A(new_n14901), .Y(new_n14902));
  NOR2xp33_ASAP7_75t_L      g14646(.A(new_n14899), .B(new_n14901), .Y(new_n14903));
  A2O1A1O1Ixp25_ASAP7_75t_L g14647(.A1(new_n14861), .A2(\a[56] ), .B(new_n14862), .C(new_n14902), .D(new_n14903), .Y(new_n14904));
  INVx1_ASAP7_75t_L         g14648(.A(new_n14568), .Y(new_n14905));
  O2A1O1Ixp33_ASAP7_75t_L   g14649(.A1(new_n14570), .A2(new_n14562), .B(new_n14574), .C(new_n14905), .Y(new_n14906));
  NAND2xp33_ASAP7_75t_L     g14650(.A(new_n14906), .B(new_n14904), .Y(new_n14907));
  A2O1A1Ixp33_ASAP7_75t_L   g14651(.A1(\a[56] ), .A2(new_n14861), .B(new_n14862), .C(new_n14899), .Y(new_n14908));
  O2A1O1Ixp33_ASAP7_75t_L   g14652(.A1(new_n14899), .A2(new_n14901), .B(new_n14908), .C(new_n14906), .Y(new_n14909));
  INVx1_ASAP7_75t_L         g14653(.A(new_n14909), .Y(new_n14910));
  NAND2xp33_ASAP7_75t_L     g14654(.A(new_n14910), .B(new_n14907), .Y(new_n14911));
  NOR2xp33_ASAP7_75t_L      g14655(.A(new_n1458), .B(new_n10400), .Y(new_n14912));
  AOI221xp5_ASAP7_75t_L     g14656(.A1(new_n9102), .A2(\b[19] ), .B1(new_n10398), .B2(\b[17] ), .C(new_n14912), .Y(new_n14913));
  O2A1O1Ixp33_ASAP7_75t_L   g14657(.A1(new_n9104), .A2(new_n1628), .B(new_n14913), .C(new_n9099), .Y(new_n14914));
  O2A1O1Ixp33_ASAP7_75t_L   g14658(.A1(new_n9104), .A2(new_n1628), .B(new_n14913), .C(\a[53] ), .Y(new_n14915));
  INVx1_ASAP7_75t_L         g14659(.A(new_n14915), .Y(new_n14916));
  O2A1O1Ixp33_ASAP7_75t_L   g14660(.A1(new_n14914), .A2(new_n9099), .B(new_n14916), .C(new_n14911), .Y(new_n14917));
  INVx1_ASAP7_75t_L         g14661(.A(new_n14914), .Y(new_n14918));
  A2O1A1Ixp33_ASAP7_75t_L   g14662(.A1(\a[53] ), .A2(new_n14918), .B(new_n14915), .C(new_n14911), .Y(new_n14919));
  INVx1_ASAP7_75t_L         g14663(.A(new_n14587), .Y(new_n14920));
  A2O1A1Ixp33_ASAP7_75t_L   g14664(.A1(\a[53] ), .A2(new_n14285), .B(new_n14282), .C(new_n14588), .Y(new_n14921));
  A2O1A1Ixp33_ASAP7_75t_L   g14665(.A1(new_n14920), .A2(new_n14921), .B(new_n14585), .C(new_n14582), .Y(new_n14922));
  INVx1_ASAP7_75t_L         g14666(.A(new_n14922), .Y(new_n14923));
  OAI211xp5_ASAP7_75t_L     g14667(.A1(new_n14911), .A2(new_n14917), .B(new_n14923), .C(new_n14919), .Y(new_n14924));
  OAI21xp33_ASAP7_75t_L     g14668(.A1(new_n9099), .A2(new_n14914), .B(new_n14916), .Y(new_n14925));
  INVx1_ASAP7_75t_L         g14669(.A(new_n14917), .Y(new_n14926));
  NOR2xp33_ASAP7_75t_L      g14670(.A(new_n14925), .B(new_n14911), .Y(new_n14927));
  A2O1A1Ixp33_ASAP7_75t_L   g14671(.A1(new_n14926), .A2(new_n14925), .B(new_n14927), .C(new_n14922), .Y(new_n14928));
  NAND2xp33_ASAP7_75t_L     g14672(.A(new_n14924), .B(new_n14928), .Y(new_n14929));
  NOR2xp33_ASAP7_75t_L      g14673(.A(new_n1895), .B(new_n10065), .Y(new_n14930));
  AOI221xp5_ASAP7_75t_L     g14674(.A1(new_n8175), .A2(\b[22] ), .B1(new_n8484), .B2(\b[20] ), .C(new_n14930), .Y(new_n14931));
  O2A1O1Ixp33_ASAP7_75t_L   g14675(.A1(new_n8176), .A2(new_n2522), .B(new_n14931), .C(new_n8172), .Y(new_n14932));
  O2A1O1Ixp33_ASAP7_75t_L   g14676(.A1(new_n8176), .A2(new_n2522), .B(new_n14931), .C(\a[50] ), .Y(new_n14933));
  INVx1_ASAP7_75t_L         g14677(.A(new_n14933), .Y(new_n14934));
  O2A1O1Ixp33_ASAP7_75t_L   g14678(.A1(new_n14932), .A2(new_n8172), .B(new_n14934), .C(new_n14929), .Y(new_n14935));
  INVx1_ASAP7_75t_L         g14679(.A(new_n14932), .Y(new_n14936));
  A2O1A1Ixp33_ASAP7_75t_L   g14680(.A1(\a[50] ), .A2(new_n14936), .B(new_n14933), .C(new_n14929), .Y(new_n14937));
  INVx1_ASAP7_75t_L         g14681(.A(new_n14601), .Y(new_n14938));
  A2O1A1O1Ixp25_ASAP7_75t_L g14682(.A1(new_n14590), .A2(new_n14592), .B(new_n14938), .C(new_n14605), .D(new_n14599), .Y(new_n14939));
  OA211x2_ASAP7_75t_L       g14683(.A1(new_n14929), .A2(new_n14935), .B(new_n14937), .C(new_n14939), .Y(new_n14940));
  O2A1O1Ixp33_ASAP7_75t_L   g14684(.A1(new_n14929), .A2(new_n14935), .B(new_n14937), .C(new_n14939), .Y(new_n14941));
  NOR2xp33_ASAP7_75t_L      g14685(.A(new_n14941), .B(new_n14940), .Y(new_n14942));
  NOR2xp33_ASAP7_75t_L      g14686(.A(new_n2205), .B(new_n7312), .Y(new_n14943));
  AOI221xp5_ASAP7_75t_L     g14687(.A1(\b[23] ), .A2(new_n7609), .B1(\b[25] ), .B2(new_n7334), .C(new_n14943), .Y(new_n14944));
  O2A1O1Ixp33_ASAP7_75t_L   g14688(.A1(new_n7321), .A2(new_n2385), .B(new_n14944), .C(new_n7316), .Y(new_n14945));
  INVx1_ASAP7_75t_L         g14689(.A(new_n14945), .Y(new_n14946));
  O2A1O1Ixp33_ASAP7_75t_L   g14690(.A1(new_n7321), .A2(new_n2385), .B(new_n14944), .C(\a[47] ), .Y(new_n14947));
  A2O1A1Ixp33_ASAP7_75t_L   g14691(.A1(\a[47] ), .A2(new_n14946), .B(new_n14947), .C(new_n14942), .Y(new_n14948));
  INVx1_ASAP7_75t_L         g14692(.A(new_n14947), .Y(new_n14949));
  O2A1O1Ixp33_ASAP7_75t_L   g14693(.A1(new_n14945), .A2(new_n7316), .B(new_n14949), .C(new_n14942), .Y(new_n14950));
  AOI21xp33_ASAP7_75t_L     g14694(.A1(new_n14948), .A2(new_n14942), .B(new_n14950), .Y(new_n14951));
  INVx1_ASAP7_75t_L         g14695(.A(new_n14613), .Y(new_n14952));
  INVx1_ASAP7_75t_L         g14696(.A(new_n14310), .Y(new_n14953));
  O2A1O1Ixp33_ASAP7_75t_L   g14697(.A1(new_n14302), .A2(new_n14303), .B(new_n14953), .C(new_n14614), .Y(new_n14954));
  O2A1O1Ixp33_ASAP7_75t_L   g14698(.A1(new_n14603), .A2(new_n14606), .B(new_n14952), .C(new_n14954), .Y(new_n14955));
  XNOR2x2_ASAP7_75t_L       g14699(.A(new_n14955), .B(new_n14951), .Y(new_n14956));
  NOR2xp33_ASAP7_75t_L      g14700(.A(new_n2703), .B(new_n6741), .Y(new_n14957));
  AOI221xp5_ASAP7_75t_L     g14701(.A1(\b[28] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[27] ), .C(new_n14957), .Y(new_n14958));
  O2A1O1Ixp33_ASAP7_75t_L   g14702(.A1(new_n6443), .A2(new_n3087), .B(new_n14958), .C(new_n6439), .Y(new_n14959));
  O2A1O1Ixp33_ASAP7_75t_L   g14703(.A1(new_n6443), .A2(new_n3087), .B(new_n14958), .C(\a[44] ), .Y(new_n14960));
  INVx1_ASAP7_75t_L         g14704(.A(new_n14960), .Y(new_n14961));
  O2A1O1Ixp33_ASAP7_75t_L   g14705(.A1(new_n14959), .A2(new_n6439), .B(new_n14961), .C(new_n14956), .Y(new_n14962));
  INVx1_ASAP7_75t_L         g14706(.A(new_n14959), .Y(new_n14963));
  A2O1A1Ixp33_ASAP7_75t_L   g14707(.A1(\a[44] ), .A2(new_n14963), .B(new_n14960), .C(new_n14956), .Y(new_n14964));
  OAI21xp33_ASAP7_75t_L     g14708(.A1(new_n14956), .A2(new_n14962), .B(new_n14964), .Y(new_n14965));
  NAND2xp33_ASAP7_75t_L     g14709(.A(new_n14637), .B(new_n14640), .Y(new_n14966));
  XOR2x2_ASAP7_75t_L        g14710(.A(new_n14966), .B(new_n14965), .Y(new_n14967));
  NOR2xp33_ASAP7_75t_L      g14711(.A(new_n3674), .B(new_n5641), .Y(new_n14968));
  AOI221xp5_ASAP7_75t_L     g14712(.A1(\b[29] ), .A2(new_n5920), .B1(\b[30] ), .B2(new_n5623), .C(new_n14968), .Y(new_n14969));
  O2A1O1Ixp33_ASAP7_75t_L   g14713(.A1(new_n5630), .A2(new_n3681), .B(new_n14969), .C(new_n5626), .Y(new_n14970));
  INVx1_ASAP7_75t_L         g14714(.A(new_n14970), .Y(new_n14971));
  O2A1O1Ixp33_ASAP7_75t_L   g14715(.A1(new_n5630), .A2(new_n3681), .B(new_n14969), .C(\a[41] ), .Y(new_n14972));
  AOI21xp33_ASAP7_75t_L     g14716(.A1(new_n14971), .A2(\a[41] ), .B(new_n14972), .Y(new_n14973));
  XOR2x2_ASAP7_75t_L        g14717(.A(new_n14973), .B(new_n14967), .Y(new_n14974));
  XOR2x2_ASAP7_75t_L        g14718(.A(new_n14644), .B(new_n14974), .Y(new_n14975));
  A2O1A1Ixp33_ASAP7_75t_L   g14719(.A1(new_n14856), .A2(\a[38] ), .B(new_n14857), .C(new_n14975), .Y(new_n14976));
  AOI21xp33_ASAP7_75t_L     g14720(.A1(new_n14856), .A2(\a[38] ), .B(new_n14857), .Y(new_n14977));
  XNOR2x2_ASAP7_75t_L       g14721(.A(new_n14644), .B(new_n14974), .Y(new_n14978));
  NAND2xp33_ASAP7_75t_L     g14722(.A(new_n14977), .B(new_n14978), .Y(new_n14979));
  NAND3xp33_ASAP7_75t_L     g14723(.A(new_n14976), .B(new_n14852), .C(new_n14979), .Y(new_n14980));
  INVx1_ASAP7_75t_L         g14724(.A(new_n14852), .Y(new_n14981));
  INVx1_ASAP7_75t_L         g14725(.A(new_n14857), .Y(new_n14982));
  O2A1O1Ixp33_ASAP7_75t_L   g14726(.A1(new_n4906), .A2(new_n14855), .B(new_n14982), .C(new_n14978), .Y(new_n14983));
  INVx1_ASAP7_75t_L         g14727(.A(new_n14977), .Y(new_n14984));
  NOR2xp33_ASAP7_75t_L      g14728(.A(new_n14984), .B(new_n14975), .Y(new_n14985));
  OAI21xp33_ASAP7_75t_L     g14729(.A1(new_n14985), .A2(new_n14983), .B(new_n14981), .Y(new_n14986));
  NAND3xp33_ASAP7_75t_L     g14730(.A(new_n14986), .B(new_n14980), .C(new_n14850), .Y(new_n14987));
  AND3x1_ASAP7_75t_L        g14731(.A(new_n14986), .B(new_n14980), .C(new_n14849), .Y(new_n14988));
  O2A1O1Ixp33_ASAP7_75t_L   g14732(.A1(new_n14847), .A2(new_n14848), .B(new_n14987), .C(new_n14988), .Y(new_n14989));
  XNOR2x2_ASAP7_75t_L       g14733(.A(new_n14843), .B(new_n14989), .Y(new_n14990));
  XNOR2x2_ASAP7_75t_L       g14734(.A(new_n14832), .B(new_n14990), .Y(new_n14991));
  XNOR2x2_ASAP7_75t_L       g14735(.A(new_n14822), .B(new_n14991), .Y(new_n14992));
  XNOR2x2_ASAP7_75t_L       g14736(.A(new_n14812), .B(new_n14992), .Y(new_n14993));
  XOR2x2_ASAP7_75t_L        g14737(.A(new_n14993), .B(new_n14799), .Y(new_n14994));
  NAND2xp33_ASAP7_75t_L     g14738(.A(new_n14791), .B(new_n14994), .Y(new_n14995));
  NOR2xp33_ASAP7_75t_L      g14739(.A(new_n14791), .B(new_n14994), .Y(new_n14996));
  NOR2xp33_ASAP7_75t_L      g14740(.A(new_n14996), .B(new_n14783), .Y(new_n14997));
  INVx1_ASAP7_75t_L         g14741(.A(new_n14996), .Y(new_n14998));
  NAND3xp33_ASAP7_75t_L     g14742(.A(new_n14783), .B(new_n14995), .C(new_n14998), .Y(new_n14999));
  A2O1A1Ixp33_ASAP7_75t_L   g14743(.A1(new_n14997), .A2(new_n14995), .B(new_n14783), .C(new_n14999), .Y(new_n15000));
  NAND3xp33_ASAP7_75t_L     g14744(.A(new_n15000), .B(new_n14773), .C(new_n14771), .Y(new_n15001));
  INVx1_ASAP7_75t_L         g14745(.A(new_n15001), .Y(new_n15002));
  INVx1_ASAP7_75t_L         g14746(.A(new_n14485), .Y(new_n15003));
  AOI22xp33_ASAP7_75t_L     g14747(.A1(new_n470), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n560), .Y(new_n15004));
  A2O1A1Ixp33_ASAP7_75t_L   g14748(.A1(new_n12990), .A2(new_n12988), .B(new_n477), .C(new_n15004), .Y(new_n15005));
  NOR2xp33_ASAP7_75t_L      g14749(.A(new_n466), .B(new_n15005), .Y(new_n15006));
  O2A1O1Ixp33_ASAP7_75t_L   g14750(.A1(new_n477), .A2(new_n12993), .B(new_n15004), .C(\a[8] ), .Y(new_n15007));
  NOR2xp33_ASAP7_75t_L      g14751(.A(new_n15007), .B(new_n15006), .Y(new_n15008));
  A2O1A1O1Ixp25_ASAP7_75t_L g14752(.A1(new_n14733), .A2(new_n14742), .B(new_n14484), .C(new_n15003), .D(new_n15008), .Y(new_n15009));
  A2O1A1Ixp33_ASAP7_75t_L   g14753(.A1(new_n14742), .A2(new_n14733), .B(new_n14484), .C(new_n15003), .Y(new_n15010));
  INVx1_ASAP7_75t_L         g14754(.A(new_n15008), .Y(new_n15011));
  NOR2xp33_ASAP7_75t_L      g14755(.A(new_n15011), .B(new_n15010), .Y(new_n15012));
  NOR2xp33_ASAP7_75t_L      g14756(.A(new_n15009), .B(new_n15012), .Y(new_n15013));
  NAND2xp33_ASAP7_75t_L     g14757(.A(new_n14773), .B(new_n14771), .Y(new_n15014));
  AND4x1_ASAP7_75t_L        g14758(.A(new_n14998), .B(new_n14995), .C(new_n14782), .D(new_n14781), .Y(new_n15015));
  OAI211xp5_ASAP7_75t_L     g14759(.A1(new_n14783), .A2(new_n15015), .B(new_n15014), .C(new_n14999), .Y(new_n15016));
  NAND3xp33_ASAP7_75t_L     g14760(.A(new_n15013), .B(new_n15001), .C(new_n15016), .Y(new_n15017));
  NAND2xp33_ASAP7_75t_L     g14761(.A(new_n15013), .B(new_n15017), .Y(new_n15018));
  A2O1A1Ixp33_ASAP7_75t_L   g14762(.A1(new_n14773), .A2(new_n14771), .B(new_n15000), .C(new_n15017), .Y(new_n15019));
  A2O1A1Ixp33_ASAP7_75t_L   g14763(.A1(new_n14754), .A2(new_n14753), .B(new_n14749), .C(new_n14477), .Y(new_n15020));
  O2A1O1Ixp33_ASAP7_75t_L   g14764(.A1(new_n15002), .A2(new_n15019), .B(new_n15018), .C(new_n15020), .Y(new_n15021));
  NAND3xp33_ASAP7_75t_L     g14765(.A(new_n15017), .B(new_n15016), .C(new_n15001), .Y(new_n15022));
  NAND2xp33_ASAP7_75t_L     g14766(.A(new_n15018), .B(new_n15022), .Y(new_n15023));
  O2A1O1Ixp33_ASAP7_75t_L   g14767(.A1(new_n14753), .A2(new_n14476), .B(new_n14754), .C(new_n14749), .Y(new_n15024));
  INVx1_ASAP7_75t_L         g14768(.A(new_n15024), .Y(new_n15025));
  O2A1O1Ixp33_ASAP7_75t_L   g14769(.A1(new_n14473), .A2(new_n14753), .B(new_n15025), .C(new_n15023), .Y(new_n15026));
  NOR2xp33_ASAP7_75t_L      g14770(.A(new_n15021), .B(new_n15026), .Y(new_n15027));
  A2O1A1O1Ixp25_ASAP7_75t_L g14771(.A1(new_n14750), .A2(new_n14755), .B(new_n14470), .C(new_n14758), .D(new_n15027), .Y(new_n15028));
  A2O1A1Ixp33_ASAP7_75t_L   g14772(.A1(new_n14175), .A2(new_n14453), .B(new_n14443), .C(new_n14756), .Y(new_n15029));
  AND3x1_ASAP7_75t_L        g14773(.A(new_n15027), .B(new_n14758), .C(new_n15029), .Y(new_n15030));
  NOR2xp33_ASAP7_75t_L      g14774(.A(new_n15028), .B(new_n15030), .Y(\f[70] ));
  NAND2xp33_ASAP7_75t_L     g14775(.A(new_n14745), .B(new_n14743), .Y(new_n15032));
  A2O1A1Ixp33_ASAP7_75t_L   g14776(.A1(new_n15032), .A2(new_n15003), .B(new_n15008), .C(new_n15017), .Y(new_n15033));
  INVx1_ASAP7_75t_L         g14777(.A(new_n14773), .Y(new_n15034));
  NOR2xp33_ASAP7_75t_L      g14778(.A(new_n12956), .B(new_n506), .Y(new_n15035));
  A2O1A1Ixp33_ASAP7_75t_L   g14779(.A1(new_n12986), .A2(new_n483), .B(new_n15035), .C(\a[8] ), .Y(new_n15036));
  A2O1A1O1Ixp25_ASAP7_75t_L g14780(.A1(new_n483), .A2(new_n14172), .B(new_n560), .C(\b[63] ), .D(new_n466), .Y(new_n15037));
  A2O1A1O1Ixp25_ASAP7_75t_L g14781(.A1(new_n12986), .A2(new_n483), .B(new_n15035), .C(new_n15036), .D(new_n15037), .Y(new_n15038));
  INVx1_ASAP7_75t_L         g14782(.A(new_n15038), .Y(new_n15039));
  A2O1A1Ixp33_ASAP7_75t_L   g14783(.A1(new_n15000), .A2(new_n14771), .B(new_n15034), .C(new_n15039), .Y(new_n15040));
  INVx1_ASAP7_75t_L         g14784(.A(new_n15040), .Y(new_n15041));
  A2O1A1O1Ixp25_ASAP7_75t_L g14785(.A1(new_n12603), .A2(new_n14444), .B(new_n477), .C(new_n506), .D(new_n12956), .Y(new_n15042));
  A2O1A1Ixp33_ASAP7_75t_L   g14786(.A1(new_n15036), .A2(new_n15042), .B(new_n15037), .C(new_n15040), .Y(new_n15043));
  A2O1A1Ixp33_ASAP7_75t_L   g14787(.A1(new_n15001), .A2(new_n14773), .B(new_n15041), .C(new_n15043), .Y(new_n15044));
  NOR2xp33_ASAP7_75t_L      g14788(.A(new_n8427), .B(new_n1962), .Y(new_n15045));
  AOI221xp5_ASAP7_75t_L     g14789(.A1(new_n1955), .A2(\b[50] ), .B1(new_n2093), .B2(\b[48] ), .C(new_n15045), .Y(new_n15046));
  INVx1_ASAP7_75t_L         g14790(.A(new_n15046), .Y(new_n15047));
  O2A1O1Ixp33_ASAP7_75t_L   g14791(.A1(new_n1956), .A2(new_n8764), .B(new_n15046), .C(new_n1952), .Y(new_n15048));
  INVx1_ASAP7_75t_L         g14792(.A(new_n15048), .Y(new_n15049));
  NOR2xp33_ASAP7_75t_L      g14793(.A(new_n1952), .B(new_n15048), .Y(new_n15050));
  A2O1A1O1Ixp25_ASAP7_75t_L g14794(.A1(new_n8763), .A2(new_n1964), .B(new_n15047), .C(new_n15049), .D(new_n15050), .Y(new_n15051));
  INVx1_ASAP7_75t_L         g14795(.A(new_n15051), .Y(new_n15052));
  OAI21xp33_ASAP7_75t_L     g14796(.A1(new_n2928), .A2(new_n14825), .B(new_n14827), .Y(new_n15053));
  INVx1_ASAP7_75t_L         g14797(.A(new_n14829), .Y(new_n15054));
  O2A1O1Ixp33_ASAP7_75t_L   g14798(.A1(new_n14673), .A2(new_n14680), .B(new_n14676), .C(new_n15053), .Y(new_n15055));
  INVx1_ASAP7_75t_L         g14799(.A(new_n14990), .Y(new_n15056));
  A2O1A1Ixp33_ASAP7_75t_L   g14800(.A1(new_n15054), .A2(new_n15053), .B(new_n15055), .C(new_n15056), .Y(new_n15057));
  INVx1_ASAP7_75t_L         g14801(.A(new_n14832), .Y(new_n15058));
  NAND2xp33_ASAP7_75t_L     g14802(.A(new_n15058), .B(new_n14990), .Y(new_n15059));
  A2O1A1Ixp33_ASAP7_75t_L   g14803(.A1(new_n15057), .A2(new_n15059), .B(new_n14822), .C(new_n14820), .Y(new_n15060));
  NOR2xp33_ASAP7_75t_L      g14804(.A(new_n15052), .B(new_n15060), .Y(new_n15061));
  O2A1O1Ixp33_ASAP7_75t_L   g14805(.A1(new_n14822), .A2(new_n14991), .B(new_n14820), .C(new_n15051), .Y(new_n15062));
  NOR2xp33_ASAP7_75t_L      g14806(.A(new_n7270), .B(new_n2410), .Y(new_n15063));
  AOI221xp5_ASAP7_75t_L     g14807(.A1(\b[45] ), .A2(new_n2577), .B1(\b[47] ), .B2(new_n2423), .C(new_n15063), .Y(new_n15064));
  O2A1O1Ixp33_ASAP7_75t_L   g14808(.A1(new_n2425), .A2(new_n7560), .B(new_n15064), .C(new_n2413), .Y(new_n15065));
  O2A1O1Ixp33_ASAP7_75t_L   g14809(.A1(new_n2425), .A2(new_n7560), .B(new_n15064), .C(\a[26] ), .Y(new_n15066));
  INVx1_ASAP7_75t_L         g14810(.A(new_n15066), .Y(new_n15067));
  OAI21xp33_ASAP7_75t_L     g14811(.A1(new_n2413), .A2(new_n15065), .B(new_n15067), .Y(new_n15068));
  A2O1A1Ixp33_ASAP7_75t_L   g14812(.A1(new_n14990), .A2(new_n14832), .B(new_n14829), .C(new_n15068), .Y(new_n15069));
  O2A1O1Ixp33_ASAP7_75t_L   g14813(.A1(new_n15058), .A2(new_n15056), .B(new_n15054), .C(new_n15068), .Y(new_n15070));
  NOR2xp33_ASAP7_75t_L      g14814(.A(new_n6671), .B(new_n2925), .Y(new_n15071));
  AOI221xp5_ASAP7_75t_L     g14815(.A1(\b[42] ), .A2(new_n3129), .B1(\b[44] ), .B2(new_n2938), .C(new_n15071), .Y(new_n15072));
  INVx1_ASAP7_75t_L         g14816(.A(new_n15072), .Y(new_n15073));
  A2O1A1Ixp33_ASAP7_75t_L   g14817(.A1(new_n2927), .A2(new_n2929), .B(new_n2739), .C(new_n15072), .Y(new_n15074));
  A2O1A1O1Ixp25_ASAP7_75t_L g14818(.A1(new_n6950), .A2(new_n6947), .B(new_n15073), .C(new_n15074), .D(new_n2928), .Y(new_n15075));
  O2A1O1Ixp33_ASAP7_75t_L   g14819(.A1(new_n2940), .A2(new_n6951), .B(new_n15072), .C(\a[29] ), .Y(new_n15076));
  NOR2xp33_ASAP7_75t_L      g14820(.A(new_n15075), .B(new_n15076), .Y(new_n15077));
  INVx1_ASAP7_75t_L         g14821(.A(new_n15077), .Y(new_n15078));
  INVx1_ASAP7_75t_L         g14822(.A(new_n14842), .Y(new_n15079));
  O2A1O1Ixp33_ASAP7_75t_L   g14823(.A1(new_n14841), .A2(new_n14989), .B(new_n15079), .C(new_n15077), .Y(new_n15080));
  INVx1_ASAP7_75t_L         g14824(.A(new_n15080), .Y(new_n15081));
  O2A1O1Ixp33_ASAP7_75t_L   g14825(.A1(new_n14841), .A2(new_n14989), .B(new_n15079), .C(new_n15078), .Y(new_n15082));
  NOR2xp33_ASAP7_75t_L      g14826(.A(new_n6110), .B(new_n3510), .Y(new_n15083));
  AOI221xp5_ASAP7_75t_L     g14827(.A1(\b[39] ), .A2(new_n3708), .B1(\b[40] ), .B2(new_n3499), .C(new_n15083), .Y(new_n15084));
  O2A1O1Ixp33_ASAP7_75t_L   g14828(.A1(new_n3513), .A2(new_n6117), .B(new_n15084), .C(new_n3493), .Y(new_n15085));
  INVx1_ASAP7_75t_L         g14829(.A(new_n15085), .Y(new_n15086));
  O2A1O1Ixp33_ASAP7_75t_L   g14830(.A1(new_n3513), .A2(new_n6117), .B(new_n15084), .C(\a[32] ), .Y(new_n15087));
  AOI21xp33_ASAP7_75t_L     g14831(.A1(new_n15086), .A2(\a[32] ), .B(new_n15087), .Y(new_n15088));
  NAND3xp33_ASAP7_75t_L     g14832(.A(new_n14987), .B(new_n14980), .C(new_n15088), .Y(new_n15089));
  NAND2xp33_ASAP7_75t_L     g14833(.A(new_n14979), .B(new_n14976), .Y(new_n15090));
  MAJIxp5_ASAP7_75t_L       g14834(.A(new_n15090), .B(new_n14849), .C(new_n14981), .Y(new_n15091));
  A2O1A1Ixp33_ASAP7_75t_L   g14835(.A1(new_n15086), .A2(\a[32] ), .B(new_n15087), .C(new_n15091), .Y(new_n15092));
  NAND2xp33_ASAP7_75t_L     g14836(.A(new_n15092), .B(new_n15089), .Y(new_n15093));
  O2A1O1Ixp33_ASAP7_75t_L   g14837(.A1(new_n9099), .A2(new_n14914), .B(new_n14916), .C(new_n14917), .Y(new_n15094));
  O2A1O1Ixp33_ASAP7_75t_L   g14838(.A1(new_n14927), .A2(new_n15094), .B(new_n14922), .C(new_n14935), .Y(new_n15095));
  INVx1_ASAP7_75t_L         g14839(.A(new_n15095), .Y(new_n15096));
  NOR2xp33_ASAP7_75t_L      g14840(.A(new_n2045), .B(new_n10065), .Y(new_n15097));
  AOI221xp5_ASAP7_75t_L     g14841(.A1(new_n8175), .A2(\b[23] ), .B1(new_n8484), .B2(\b[21] ), .C(new_n15097), .Y(new_n15098));
  O2A1O1Ixp33_ASAP7_75t_L   g14842(.A1(new_n8176), .A2(new_n2194), .B(new_n15098), .C(new_n8172), .Y(new_n15099));
  INVx1_ASAP7_75t_L         g14843(.A(new_n15099), .Y(new_n15100));
  O2A1O1Ixp33_ASAP7_75t_L   g14844(.A1(new_n8176), .A2(new_n2194), .B(new_n15098), .C(\a[50] ), .Y(new_n15101));
  INVx1_ASAP7_75t_L         g14845(.A(new_n14904), .Y(new_n15102));
  INVx1_ASAP7_75t_L         g14846(.A(new_n14906), .Y(new_n15103));
  A2O1A1O1Ixp25_ASAP7_75t_L g14847(.A1(new_n14888), .A2(\a[59] ), .B(new_n14889), .C(new_n14884), .D(new_n14881), .Y(new_n15104));
  A2O1A1Ixp33_ASAP7_75t_L   g14848(.A1(new_n14876), .A2(new_n14877), .B(new_n14872), .C(new_n14869), .Y(new_n15105));
  NOR2xp33_ASAP7_75t_L      g14849(.A(new_n448), .B(new_n13030), .Y(new_n15106));
  INVx1_ASAP7_75t_L         g14850(.A(new_n15106), .Y(new_n15107));
  O2A1O1Ixp33_ASAP7_75t_L   g14851(.A1(new_n12672), .A2(new_n534), .B(new_n15107), .C(new_n14867), .Y(new_n15108));
  INVx1_ASAP7_75t_L         g14852(.A(new_n15108), .Y(new_n15109));
  O2A1O1Ixp33_ASAP7_75t_L   g14853(.A1(new_n12669), .A2(new_n12671), .B(\b[8] ), .C(new_n15106), .Y(new_n15110));
  A2O1A1Ixp33_ASAP7_75t_L   g14854(.A1(new_n13028), .A2(\b[7] ), .B(new_n14865), .C(new_n15110), .Y(new_n15111));
  INVx1_ASAP7_75t_L         g14855(.A(new_n15111), .Y(new_n15112));
  A2O1A1O1Ixp25_ASAP7_75t_L g14856(.A1(new_n14877), .A2(new_n14876), .B(new_n14872), .C(new_n14869), .D(new_n15112), .Y(new_n15113));
  NAND2xp33_ASAP7_75t_L     g14857(.A(new_n15109), .B(new_n15113), .Y(new_n15114));
  NAND3xp33_ASAP7_75t_L     g14858(.A(new_n14878), .B(new_n14871), .C(new_n14869), .Y(new_n15115));
  A2O1A1Ixp33_ASAP7_75t_L   g14859(.A1(new_n15115), .A2(new_n14869), .B(new_n15108), .C(new_n15111), .Y(new_n15116));
  A2O1A1O1Ixp25_ASAP7_75t_L g14860(.A1(new_n13028), .A2(\b[8] ), .B(new_n15106), .C(new_n14866), .D(new_n15116), .Y(new_n15117));
  OAI22xp33_ASAP7_75t_L     g14861(.A1(new_n12320), .A2(new_n590), .B1(new_n680), .B2(new_n12318), .Y(new_n15118));
  AOI221xp5_ASAP7_75t_L     g14862(.A1(new_n11995), .A2(\b[11] ), .B1(new_n11997), .B2(new_n976), .C(new_n15118), .Y(new_n15119));
  XNOR2x2_ASAP7_75t_L       g14863(.A(new_n11987), .B(new_n15119), .Y(new_n15120));
  A2O1A1Ixp33_ASAP7_75t_L   g14864(.A1(new_n15114), .A2(new_n15105), .B(new_n15117), .C(new_n15120), .Y(new_n15121));
  A2O1A1Ixp33_ASAP7_75t_L   g14865(.A1(new_n14871), .A2(new_n14878), .B(new_n14868), .C(new_n15114), .Y(new_n15122));
  INVx1_ASAP7_75t_L         g14866(.A(new_n15120), .Y(new_n15123));
  OAI211xp5_ASAP7_75t_L     g14867(.A1(new_n15108), .A2(new_n15116), .B(new_n15122), .C(new_n15123), .Y(new_n15124));
  NAND2xp33_ASAP7_75t_L     g14868(.A(new_n15124), .B(new_n15121), .Y(new_n15125));
  NOR2xp33_ASAP7_75t_L      g14869(.A(new_n833), .B(new_n11354), .Y(new_n15126));
  AOI221xp5_ASAP7_75t_L     g14870(.A1(\b[14] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[13] ), .C(new_n15126), .Y(new_n15127));
  O2A1O1Ixp33_ASAP7_75t_L   g14871(.A1(new_n11053), .A2(new_n1268), .B(new_n15127), .C(new_n11048), .Y(new_n15128));
  NOR2xp33_ASAP7_75t_L      g14872(.A(new_n11048), .B(new_n15128), .Y(new_n15129));
  O2A1O1Ixp33_ASAP7_75t_L   g14873(.A1(new_n11053), .A2(new_n1268), .B(new_n15127), .C(\a[59] ), .Y(new_n15130));
  NOR2xp33_ASAP7_75t_L      g14874(.A(new_n15130), .B(new_n15129), .Y(new_n15131));
  XOR2x2_ASAP7_75t_L        g14875(.A(new_n15131), .B(new_n15125), .Y(new_n15132));
  AND2x2_ASAP7_75t_L        g14876(.A(new_n15104), .B(new_n15132), .Y(new_n15133));
  INVx1_ASAP7_75t_L         g14877(.A(new_n14882), .Y(new_n15134));
  O2A1O1Ixp33_ASAP7_75t_L   g14878(.A1(new_n15134), .A2(new_n14880), .B(new_n14890), .C(new_n15132), .Y(new_n15135));
  NOR2xp33_ASAP7_75t_L      g14879(.A(new_n15135), .B(new_n15133), .Y(new_n15136));
  NOR2xp33_ASAP7_75t_L      g14880(.A(new_n1150), .B(new_n10388), .Y(new_n15137));
  AOI221xp5_ASAP7_75t_L     g14881(.A1(new_n10086), .A2(\b[17] ), .B1(new_n11361), .B2(\b[15] ), .C(new_n15137), .Y(new_n15138));
  O2A1O1Ixp33_ASAP7_75t_L   g14882(.A1(new_n10088), .A2(new_n1356), .B(new_n15138), .C(new_n10083), .Y(new_n15139));
  INVx1_ASAP7_75t_L         g14883(.A(new_n15139), .Y(new_n15140));
  O2A1O1Ixp33_ASAP7_75t_L   g14884(.A1(new_n10088), .A2(new_n1356), .B(new_n15138), .C(\a[56] ), .Y(new_n15141));
  A2O1A1Ixp33_ASAP7_75t_L   g14885(.A1(\a[56] ), .A2(new_n15140), .B(new_n15141), .C(new_n15136), .Y(new_n15142));
  INVx1_ASAP7_75t_L         g14886(.A(new_n15141), .Y(new_n15143));
  O2A1O1Ixp33_ASAP7_75t_L   g14887(.A1(new_n15139), .A2(new_n10083), .B(new_n15143), .C(new_n15136), .Y(new_n15144));
  AOI21xp33_ASAP7_75t_L     g14888(.A1(new_n15142), .A2(new_n15136), .B(new_n15144), .Y(new_n15145));
  A2O1A1O1Ixp25_ASAP7_75t_L g14889(.A1(new_n14861), .A2(\a[56] ), .B(new_n14862), .C(new_n14896), .D(new_n14897), .Y(new_n15146));
  AND2x2_ASAP7_75t_L        g14890(.A(new_n15146), .B(new_n15145), .Y(new_n15147));
  O2A1O1Ixp33_ASAP7_75t_L   g14891(.A1(new_n14893), .A2(new_n14895), .B(new_n14902), .C(new_n15145), .Y(new_n15148));
  NOR2xp33_ASAP7_75t_L      g14892(.A(new_n15148), .B(new_n15147), .Y(new_n15149));
  NOR2xp33_ASAP7_75t_L      g14893(.A(new_n1599), .B(new_n10400), .Y(new_n15150));
  AOI221xp5_ASAP7_75t_L     g14894(.A1(new_n9102), .A2(\b[20] ), .B1(new_n10398), .B2(\b[18] ), .C(new_n15150), .Y(new_n15151));
  O2A1O1Ixp33_ASAP7_75t_L   g14895(.A1(new_n9104), .A2(new_n1754), .B(new_n15151), .C(new_n9099), .Y(new_n15152));
  NOR2xp33_ASAP7_75t_L      g14896(.A(new_n9099), .B(new_n15152), .Y(new_n15153));
  O2A1O1Ixp33_ASAP7_75t_L   g14897(.A1(new_n9104), .A2(new_n1754), .B(new_n15151), .C(\a[53] ), .Y(new_n15154));
  OR3x1_ASAP7_75t_L         g14898(.A(new_n15149), .B(new_n15153), .C(new_n15154), .Y(new_n15155));
  INVx1_ASAP7_75t_L         g14899(.A(new_n15152), .Y(new_n15156));
  A2O1A1Ixp33_ASAP7_75t_L   g14900(.A1(\a[53] ), .A2(new_n15156), .B(new_n15154), .C(new_n15149), .Y(new_n15157));
  AND2x2_ASAP7_75t_L        g14901(.A(new_n15157), .B(new_n15155), .Y(new_n15158));
  A2O1A1Ixp33_ASAP7_75t_L   g14902(.A1(new_n15103), .A2(new_n15102), .B(new_n14917), .C(new_n15158), .Y(new_n15159));
  A2O1A1Ixp33_ASAP7_75t_L   g14903(.A1(new_n15103), .A2(new_n15102), .B(new_n14917), .C(new_n15159), .Y(new_n15160));
  A2O1A1O1Ixp25_ASAP7_75t_L g14904(.A1(new_n14918), .A2(\a[53] ), .B(new_n14915), .C(new_n14907), .D(new_n14909), .Y(new_n15161));
  NAND2xp33_ASAP7_75t_L     g14905(.A(new_n15161), .B(new_n15158), .Y(new_n15162));
  NAND2xp33_ASAP7_75t_L     g14906(.A(new_n15162), .B(new_n15160), .Y(new_n15163));
  AOI21xp33_ASAP7_75t_L     g14907(.A1(new_n15100), .A2(\a[50] ), .B(new_n15101), .Y(new_n15164));
  NAND2xp33_ASAP7_75t_L     g14908(.A(new_n15164), .B(new_n15162), .Y(new_n15165));
  O2A1O1Ixp33_ASAP7_75t_L   g14909(.A1(new_n14909), .A2(new_n14917), .B(new_n15159), .C(new_n15165), .Y(new_n15166));
  A2O1A1O1Ixp25_ASAP7_75t_L g14910(.A1(new_n15100), .A2(\a[50] ), .B(new_n15101), .C(new_n15163), .D(new_n15166), .Y(new_n15167));
  NAND2xp33_ASAP7_75t_L     g14911(.A(new_n15167), .B(new_n15096), .Y(new_n15168));
  AO21x2_ASAP7_75t_L        g14912(.A1(\a[50] ), .A2(new_n15100), .B(new_n15101), .Y(new_n15169));
  A2O1A1Ixp33_ASAP7_75t_L   g14913(.A1(new_n15163), .A2(new_n15169), .B(new_n15166), .C(new_n15095), .Y(new_n15170));
  NAND2xp33_ASAP7_75t_L     g14914(.A(new_n15170), .B(new_n15168), .Y(new_n15171));
  NOR2xp33_ASAP7_75t_L      g14915(.A(new_n2377), .B(new_n7312), .Y(new_n15172));
  AOI221xp5_ASAP7_75t_L     g14916(.A1(\b[24] ), .A2(new_n7609), .B1(\b[26] ), .B2(new_n7334), .C(new_n15172), .Y(new_n15173));
  O2A1O1Ixp33_ASAP7_75t_L   g14917(.A1(new_n7321), .A2(new_n2708), .B(new_n15173), .C(new_n7316), .Y(new_n15174));
  O2A1O1Ixp33_ASAP7_75t_L   g14918(.A1(new_n7321), .A2(new_n2708), .B(new_n15173), .C(\a[47] ), .Y(new_n15175));
  INVx1_ASAP7_75t_L         g14919(.A(new_n15175), .Y(new_n15176));
  O2A1O1Ixp33_ASAP7_75t_L   g14920(.A1(new_n15174), .A2(new_n7316), .B(new_n15176), .C(new_n15171), .Y(new_n15177));
  INVx1_ASAP7_75t_L         g14921(.A(new_n15174), .Y(new_n15178));
  A2O1A1Ixp33_ASAP7_75t_L   g14922(.A1(\a[47] ), .A2(new_n15178), .B(new_n15175), .C(new_n15171), .Y(new_n15179));
  OAI21xp33_ASAP7_75t_L     g14923(.A1(new_n15171), .A2(new_n15177), .B(new_n15179), .Y(new_n15180));
  A2O1A1O1Ixp25_ASAP7_75t_L g14924(.A1(new_n14946), .A2(\a[47] ), .B(new_n14947), .C(new_n14942), .D(new_n14941), .Y(new_n15181));
  XNOR2x2_ASAP7_75t_L       g14925(.A(new_n15181), .B(new_n15180), .Y(new_n15182));
  NOR2xp33_ASAP7_75t_L      g14926(.A(new_n3079), .B(new_n7304), .Y(new_n15183));
  AOI221xp5_ASAP7_75t_L     g14927(.A1(\b[27] ), .A2(new_n6742), .B1(\b[29] ), .B2(new_n6442), .C(new_n15183), .Y(new_n15184));
  O2A1O1Ixp33_ASAP7_75t_L   g14928(.A1(new_n6443), .A2(new_n3104), .B(new_n15184), .C(new_n6439), .Y(new_n15185));
  INVx1_ASAP7_75t_L         g14929(.A(new_n15185), .Y(new_n15186));
  O2A1O1Ixp33_ASAP7_75t_L   g14930(.A1(new_n6443), .A2(new_n3104), .B(new_n15184), .C(\a[44] ), .Y(new_n15187));
  AO21x2_ASAP7_75t_L        g14931(.A1(\a[44] ), .A2(new_n15186), .B(new_n15187), .Y(new_n15188));
  XNOR2x2_ASAP7_75t_L       g14932(.A(new_n15188), .B(new_n15182), .Y(new_n15189));
  INVx1_ASAP7_75t_L         g14933(.A(new_n14954), .Y(new_n15190));
  O2A1O1Ixp33_ASAP7_75t_L   g14934(.A1(new_n14607), .A2(new_n14613), .B(new_n15190), .C(new_n14951), .Y(new_n15191));
  INVx1_ASAP7_75t_L         g14935(.A(new_n14956), .Y(new_n15192));
  A2O1A1O1Ixp25_ASAP7_75t_L g14936(.A1(new_n14963), .A2(\a[44] ), .B(new_n14960), .C(new_n15192), .D(new_n15191), .Y(new_n15193));
  XNOR2x2_ASAP7_75t_L       g14937(.A(new_n15193), .B(new_n15189), .Y(new_n15194));
  NOR2xp33_ASAP7_75t_L      g14938(.A(new_n3891), .B(new_n5641), .Y(new_n15195));
  AOI221xp5_ASAP7_75t_L     g14939(.A1(\b[30] ), .A2(new_n5920), .B1(\b[31] ), .B2(new_n5623), .C(new_n15195), .Y(new_n15196));
  O2A1O1Ixp33_ASAP7_75t_L   g14940(.A1(new_n5630), .A2(new_n3897), .B(new_n15196), .C(new_n5626), .Y(new_n15197));
  O2A1O1Ixp33_ASAP7_75t_L   g14941(.A1(new_n5630), .A2(new_n3897), .B(new_n15196), .C(\a[41] ), .Y(new_n15198));
  INVx1_ASAP7_75t_L         g14942(.A(new_n15198), .Y(new_n15199));
  OAI21xp33_ASAP7_75t_L     g14943(.A1(new_n5626), .A2(new_n15197), .B(new_n15199), .Y(new_n15200));
  XNOR2x2_ASAP7_75t_L       g14944(.A(new_n15200), .B(new_n15194), .Y(new_n15201));
  INVx1_ASAP7_75t_L         g14945(.A(new_n14962), .Y(new_n15202));
  O2A1O1Ixp33_ASAP7_75t_L   g14946(.A1(new_n14959), .A2(new_n6439), .B(new_n14961), .C(new_n15192), .Y(new_n15203));
  A2O1A1Ixp33_ASAP7_75t_L   g14947(.A1(new_n15202), .A2(new_n15192), .B(new_n15203), .C(new_n14966), .Y(new_n15204));
  A2O1A1Ixp33_ASAP7_75t_L   g14948(.A1(\a[41] ), .A2(new_n14971), .B(new_n14972), .C(new_n14967), .Y(new_n15205));
  NAND2xp33_ASAP7_75t_L     g14949(.A(new_n15204), .B(new_n15205), .Y(new_n15206));
  XNOR2x2_ASAP7_75t_L       g14950(.A(new_n15206), .B(new_n15201), .Y(new_n15207));
  NOR2xp33_ASAP7_75t_L      g14951(.A(new_n4581), .B(new_n4908), .Y(new_n15208));
  AOI221xp5_ASAP7_75t_L     g14952(.A1(\b[33] ), .A2(new_n5139), .B1(\b[34] ), .B2(new_n4916), .C(new_n15208), .Y(new_n15209));
  O2A1O1Ixp33_ASAP7_75t_L   g14953(.A1(new_n4911), .A2(new_n4589), .B(new_n15209), .C(new_n4906), .Y(new_n15210));
  INVx1_ASAP7_75t_L         g14954(.A(new_n15210), .Y(new_n15211));
  NAND2xp33_ASAP7_75t_L     g14955(.A(\a[38] ), .B(new_n15211), .Y(new_n15212));
  O2A1O1Ixp33_ASAP7_75t_L   g14956(.A1(new_n4911), .A2(new_n4589), .B(new_n15209), .C(\a[38] ), .Y(new_n15213));
  INVx1_ASAP7_75t_L         g14957(.A(new_n15213), .Y(new_n15214));
  NAND2xp33_ASAP7_75t_L     g14958(.A(new_n15214), .B(new_n15212), .Y(new_n15215));
  XNOR2x2_ASAP7_75t_L       g14959(.A(new_n15215), .B(new_n15207), .Y(new_n15216));
  A2O1A1Ixp33_ASAP7_75t_L   g14960(.A1(new_n14339), .A2(new_n14325), .B(new_n14338), .C(new_n14634), .Y(new_n15217));
  O2A1O1Ixp33_ASAP7_75t_L   g14961(.A1(new_n14626), .A2(new_n14633), .B(new_n15217), .C(new_n14974), .Y(new_n15218));
  A2O1A1O1Ixp25_ASAP7_75t_L g14962(.A1(new_n14856), .A2(\a[38] ), .B(new_n14857), .C(new_n14975), .D(new_n15218), .Y(new_n15219));
  INVx1_ASAP7_75t_L         g14963(.A(new_n15219), .Y(new_n15220));
  NOR2xp33_ASAP7_75t_L      g14964(.A(new_n15220), .B(new_n15216), .Y(new_n15221));
  O2A1O1Ixp33_ASAP7_75t_L   g14965(.A1(new_n15210), .A2(new_n4906), .B(new_n15214), .C(new_n15207), .Y(new_n15222));
  A2O1A1Ixp33_ASAP7_75t_L   g14966(.A1(\a[38] ), .A2(new_n15211), .B(new_n15213), .C(new_n15207), .Y(new_n15223));
  O2A1O1Ixp33_ASAP7_75t_L   g14967(.A1(new_n15207), .A2(new_n15222), .B(new_n15223), .C(new_n15219), .Y(new_n15224));
  NOR2xp33_ASAP7_75t_L      g14968(.A(new_n5311), .B(new_n4147), .Y(new_n15225));
  AOI221xp5_ASAP7_75t_L     g14969(.A1(\b[36] ), .A2(new_n4402), .B1(\b[37] ), .B2(new_n4155), .C(new_n15225), .Y(new_n15226));
  O2A1O1Ixp33_ASAP7_75t_L   g14970(.A1(new_n4150), .A2(new_n5318), .B(new_n15226), .C(new_n4145), .Y(new_n15227));
  NOR2xp33_ASAP7_75t_L      g14971(.A(new_n4145), .B(new_n15227), .Y(new_n15228));
  O2A1O1Ixp33_ASAP7_75t_L   g14972(.A1(new_n4150), .A2(new_n5318), .B(new_n15226), .C(\a[35] ), .Y(new_n15229));
  NOR2xp33_ASAP7_75t_L      g14973(.A(new_n15229), .B(new_n15228), .Y(new_n15230));
  NOR3xp33_ASAP7_75t_L      g14974(.A(new_n15221), .B(new_n15224), .C(new_n15230), .Y(new_n15231));
  OA21x2_ASAP7_75t_L        g14975(.A1(new_n15224), .A2(new_n15221), .B(new_n15230), .Y(new_n15232));
  NOR3xp33_ASAP7_75t_L      g14976(.A(new_n15093), .B(new_n15231), .C(new_n15232), .Y(new_n15233));
  AO211x2_ASAP7_75t_L       g14977(.A1(new_n15092), .A2(new_n15089), .B(new_n15231), .C(new_n15232), .Y(new_n15234));
  OAI21xp33_ASAP7_75t_L     g14978(.A1(new_n15093), .A2(new_n15233), .B(new_n15234), .Y(new_n15235));
  A2O1A1Ixp33_ASAP7_75t_L   g14979(.A1(new_n15078), .A2(new_n15081), .B(new_n15082), .C(new_n15235), .Y(new_n15236));
  A2O1A1Ixp33_ASAP7_75t_L   g14980(.A1(new_n14850), .A2(new_n14987), .B(new_n14988), .C(new_n14843), .Y(new_n15237));
  A2O1A1O1Ixp25_ASAP7_75t_L g14981(.A1(new_n14987), .A2(new_n14850), .B(new_n14988), .C(new_n14843), .D(new_n14842), .Y(new_n15238));
  NAND2xp33_ASAP7_75t_L     g14982(.A(new_n15078), .B(new_n15238), .Y(new_n15239));
  A2O1A1Ixp33_ASAP7_75t_L   g14983(.A1(new_n15237), .A2(new_n15079), .B(new_n15080), .C(new_n15239), .Y(new_n15240));
  O2A1O1Ixp33_ASAP7_75t_L   g14984(.A1(new_n15093), .A2(new_n15233), .B(new_n15234), .C(new_n15240), .Y(new_n15241));
  A2O1A1O1Ixp25_ASAP7_75t_L g14985(.A1(new_n15081), .A2(new_n15078), .B(new_n15082), .C(new_n15236), .D(new_n15241), .Y(new_n15242));
  A2O1A1Ixp33_ASAP7_75t_L   g14986(.A1(new_n15069), .A2(new_n15068), .B(new_n15070), .C(new_n15242), .Y(new_n15243));
  INVx1_ASAP7_75t_L         g14987(.A(new_n15065), .Y(new_n15244));
  A2O1A1O1Ixp25_ASAP7_75t_L g14988(.A1(new_n15244), .A2(\a[26] ), .B(new_n15066), .C(new_n15069), .D(new_n15070), .Y(new_n15245));
  O2A1O1Ixp33_ASAP7_75t_L   g14989(.A1(new_n15238), .A2(new_n15080), .B(new_n15239), .C(new_n15235), .Y(new_n15246));
  A2O1A1Ixp33_ASAP7_75t_L   g14990(.A1(new_n15235), .A2(new_n15236), .B(new_n15246), .C(new_n15245), .Y(new_n15247));
  OAI211xp5_ASAP7_75t_L     g14991(.A1(new_n15062), .A2(new_n15061), .B(new_n15243), .C(new_n15247), .Y(new_n15248));
  NOR2xp33_ASAP7_75t_L      g14992(.A(new_n15062), .B(new_n15061), .Y(new_n15249));
  O2A1O1Ixp33_ASAP7_75t_L   g14993(.A1(new_n15055), .A2(new_n15053), .B(new_n14990), .C(new_n14829), .Y(new_n15250));
  A2O1A1Ixp33_ASAP7_75t_L   g14994(.A1(new_n15244), .A2(\a[26] ), .B(new_n15066), .C(new_n15250), .Y(new_n15251));
  A2O1A1Ixp33_ASAP7_75t_L   g14995(.A1(new_n14832), .A2(new_n14990), .B(new_n14829), .C(new_n15069), .Y(new_n15252));
  NAND2xp33_ASAP7_75t_L     g14996(.A(new_n15251), .B(new_n15252), .Y(new_n15253));
  AO21x2_ASAP7_75t_L        g14997(.A1(new_n15235), .A2(new_n15236), .B(new_n15246), .Y(new_n15254));
  NAND2xp33_ASAP7_75t_L     g14998(.A(new_n15254), .B(new_n15253), .Y(new_n15255));
  NOR2xp33_ASAP7_75t_L      g14999(.A(new_n15253), .B(new_n15242), .Y(new_n15256));
  A2O1A1Ixp33_ASAP7_75t_L   g15000(.A1(new_n15253), .A2(new_n15255), .B(new_n15256), .C(new_n15249), .Y(new_n15257));
  NAND2xp33_ASAP7_75t_L     g15001(.A(new_n15248), .B(new_n15257), .Y(new_n15258));
  NOR2xp33_ASAP7_75t_L      g15002(.A(new_n9355), .B(new_n1517), .Y(new_n15259));
  AOI221xp5_ASAP7_75t_L     g15003(.A1(\b[51] ), .A2(new_n1659), .B1(\b[53] ), .B2(new_n1511), .C(new_n15259), .Y(new_n15260));
  INVx1_ASAP7_75t_L         g15004(.A(new_n15260), .Y(new_n15261));
  A2O1A1Ixp33_ASAP7_75t_L   g15005(.A1(new_n1508), .A2(new_n1509), .B(new_n1389), .C(new_n15260), .Y(new_n15262));
  A2O1A1O1Ixp25_ASAP7_75t_L g15006(.A1(new_n9689), .A2(new_n9686), .B(new_n15261), .C(new_n15262), .D(new_n1501), .Y(new_n15263));
  O2A1O1Ixp33_ASAP7_75t_L   g15007(.A1(new_n1521), .A2(new_n9691), .B(new_n15260), .C(\a[20] ), .Y(new_n15264));
  NOR2xp33_ASAP7_75t_L      g15008(.A(new_n15263), .B(new_n15264), .Y(new_n15265));
  INVx1_ASAP7_75t_L         g15009(.A(new_n14809), .Y(new_n15266));
  A2O1A1O1Ixp25_ASAP7_75t_L g15010(.A1(new_n14811), .A2(new_n14808), .B(new_n14992), .C(new_n15266), .D(new_n15265), .Y(new_n15267));
  INVx1_ASAP7_75t_L         g15011(.A(new_n15265), .Y(new_n15268));
  A2O1A1O1Ixp25_ASAP7_75t_L g15012(.A1(new_n14811), .A2(new_n14808), .B(new_n14992), .C(new_n15266), .D(new_n15268), .Y(new_n15269));
  INVx1_ASAP7_75t_L         g15013(.A(new_n15269), .Y(new_n15270));
  O2A1O1Ixp33_ASAP7_75t_L   g15014(.A1(new_n15265), .A2(new_n15267), .B(new_n15270), .C(new_n15258), .Y(new_n15271));
  INVx1_ASAP7_75t_L         g15015(.A(new_n15267), .Y(new_n15272));
  A2O1A1Ixp33_ASAP7_75t_L   g15016(.A1(new_n15268), .A2(new_n15272), .B(new_n15269), .C(new_n15258), .Y(new_n15273));
  OAI21xp33_ASAP7_75t_L     g15017(.A1(new_n15258), .A2(new_n15271), .B(new_n15273), .Y(new_n15274));
  NAND2xp33_ASAP7_75t_L     g15018(.A(\b[55] ), .B(new_n1204), .Y(new_n15275));
  OAI221xp5_ASAP7_75t_L     g15019(.A1(new_n1284), .A2(new_n10332), .B1(new_n9709), .B2(new_n1285), .C(new_n15275), .Y(new_n15276));
  A2O1A1Ixp33_ASAP7_75t_L   g15020(.A1(new_n11579), .A2(new_n1216), .B(new_n15276), .C(\a[17] ), .Y(new_n15277));
  NAND2xp33_ASAP7_75t_L     g15021(.A(\a[17] ), .B(new_n15277), .Y(new_n15278));
  A2O1A1Ixp33_ASAP7_75t_L   g15022(.A1(new_n11579), .A2(new_n1216), .B(new_n15276), .C(new_n1206), .Y(new_n15279));
  NAND2xp33_ASAP7_75t_L     g15023(.A(new_n15279), .B(new_n15278), .Y(new_n15280));
  MAJx2_ASAP7_75t_L         g15024(.A(new_n14993), .B(new_n14798), .C(new_n14797), .Y(new_n15281));
  NOR2xp33_ASAP7_75t_L      g15025(.A(new_n15280), .B(new_n15281), .Y(new_n15282));
  INVx1_ASAP7_75t_L         g15026(.A(new_n15282), .Y(new_n15283));
  NAND2xp33_ASAP7_75t_L     g15027(.A(new_n15280), .B(new_n15281), .Y(new_n15284));
  NAND3xp33_ASAP7_75t_L     g15028(.A(new_n15274), .B(new_n15284), .C(new_n15283), .Y(new_n15285));
  INVx1_ASAP7_75t_L         g15029(.A(new_n15284), .Y(new_n15286));
  NOR3xp33_ASAP7_75t_L      g15030(.A(new_n15274), .B(new_n15286), .C(new_n15282), .Y(new_n15287));
  NOR2xp33_ASAP7_75t_L      g15031(.A(new_n11303), .B(new_n864), .Y(new_n15288));
  AOI221xp5_ASAP7_75t_L     g15032(.A1(\b[57] ), .A2(new_n985), .B1(\b[59] ), .B2(new_n886), .C(new_n15288), .Y(new_n15289));
  INVx1_ASAP7_75t_L         g15033(.A(new_n15289), .Y(new_n15290));
  A2O1A1Ixp33_ASAP7_75t_L   g15034(.A1(new_n12577), .A2(new_n873), .B(new_n15290), .C(\a[14] ), .Y(new_n15291));
  O2A1O1Ixp33_ASAP7_75t_L   g15035(.A1(new_n872), .A2(new_n11597), .B(new_n15289), .C(\a[14] ), .Y(new_n15292));
  AOI21xp33_ASAP7_75t_L     g15036(.A1(new_n14788), .A2(new_n14787), .B(new_n14790), .Y(new_n15293));
  AO21x2_ASAP7_75t_L        g15037(.A1(\a[14] ), .A2(new_n15291), .B(new_n15292), .Y(new_n15294));
  A2O1A1Ixp33_ASAP7_75t_L   g15038(.A1(new_n14994), .A2(new_n14791), .B(new_n15293), .C(new_n15294), .Y(new_n15295));
  A2O1A1O1Ixp25_ASAP7_75t_L g15039(.A1(new_n14788), .A2(new_n14787), .B(new_n14790), .C(new_n14995), .D(new_n15294), .Y(new_n15296));
  A2O1A1O1Ixp25_ASAP7_75t_L g15040(.A1(new_n15291), .A2(\a[14] ), .B(new_n15292), .C(new_n15295), .D(new_n15296), .Y(new_n15297));
  A2O1A1Ixp33_ASAP7_75t_L   g15041(.A1(new_n15285), .A2(new_n15274), .B(new_n15287), .C(new_n15297), .Y(new_n15298));
  AOI21xp33_ASAP7_75t_L     g15042(.A1(new_n15285), .A2(new_n15274), .B(new_n15287), .Y(new_n15299));
  A2O1A1Ixp33_ASAP7_75t_L   g15043(.A1(new_n15294), .A2(new_n15295), .B(new_n15296), .C(new_n15299), .Y(new_n15300));
  NAND2xp33_ASAP7_75t_L     g15044(.A(new_n15300), .B(new_n15298), .Y(new_n15301));
  NAND2xp33_ASAP7_75t_L     g15045(.A(\b[61] ), .B(new_n635), .Y(new_n15302));
  OAI221xp5_ASAP7_75t_L     g15046(.A1(new_n710), .A2(new_n12603), .B1(new_n11626), .B2(new_n712), .C(new_n15302), .Y(new_n15303));
  AOI21xp33_ASAP7_75t_L     g15047(.A1(new_n13559), .A2(new_n718), .B(new_n15303), .Y(new_n15304));
  NAND2xp33_ASAP7_75t_L     g15048(.A(\a[11] ), .B(new_n15304), .Y(new_n15305));
  A2O1A1Ixp33_ASAP7_75t_L   g15049(.A1(new_n13559), .A2(new_n718), .B(new_n15303), .C(new_n637), .Y(new_n15306));
  NAND2xp33_ASAP7_75t_L     g15050(.A(new_n15306), .B(new_n15305), .Y(new_n15307));
  INVx1_ASAP7_75t_L         g15051(.A(new_n15015), .Y(new_n15308));
  INVx1_ASAP7_75t_L         g15052(.A(new_n15307), .Y(new_n15309));
  A2O1A1O1Ixp25_ASAP7_75t_L g15053(.A1(new_n14735), .A2(new_n14719), .B(new_n14779), .C(new_n15308), .D(new_n15309), .Y(new_n15310));
  INVx1_ASAP7_75t_L         g15054(.A(new_n15310), .Y(new_n15311));
  A2O1A1O1Ixp25_ASAP7_75t_L g15055(.A1(new_n14735), .A2(new_n14719), .B(new_n14779), .C(new_n15308), .D(new_n15307), .Y(new_n15312));
  A2O1A1Ixp33_ASAP7_75t_L   g15056(.A1(new_n15311), .A2(new_n15307), .B(new_n15312), .C(new_n15301), .Y(new_n15313));
  AND2x2_ASAP7_75t_L        g15057(.A(new_n15300), .B(new_n15298), .Y(new_n15314));
  INVx1_ASAP7_75t_L         g15058(.A(new_n15312), .Y(new_n15315));
  INVx1_ASAP7_75t_L         g15059(.A(new_n14779), .Y(new_n15316));
  O2A1O1Ixp33_ASAP7_75t_L   g15060(.A1(new_n14720), .A2(new_n14722), .B(new_n15316), .C(new_n15015), .Y(new_n15317));
  NAND2xp33_ASAP7_75t_L     g15061(.A(new_n15307), .B(new_n15317), .Y(new_n15318));
  NAND3xp33_ASAP7_75t_L     g15062(.A(new_n15314), .B(new_n15315), .C(new_n15318), .Y(new_n15319));
  NAND3xp33_ASAP7_75t_L     g15063(.A(new_n15044), .B(new_n15313), .C(new_n15319), .Y(new_n15320));
  INVx1_ASAP7_75t_L         g15064(.A(new_n15320), .Y(new_n15321));
  INVx1_ASAP7_75t_L         g15065(.A(new_n15317), .Y(new_n15322));
  A2O1A1Ixp33_ASAP7_75t_L   g15066(.A1(new_n15305), .A2(new_n15306), .B(new_n15322), .C(new_n15314), .Y(new_n15323));
  O2A1O1Ixp33_ASAP7_75t_L   g15067(.A1(new_n15323), .A2(new_n15312), .B(new_n15313), .C(new_n15044), .Y(new_n15324));
  OAI21xp33_ASAP7_75t_L     g15068(.A1(new_n15324), .A2(new_n15321), .B(new_n15033), .Y(new_n15325));
  INVx1_ASAP7_75t_L         g15069(.A(new_n15033), .Y(new_n15326));
  INVx1_ASAP7_75t_L         g15070(.A(new_n15324), .Y(new_n15327));
  NAND3xp33_ASAP7_75t_L     g15071(.A(new_n15327), .B(new_n15320), .C(new_n15326), .Y(new_n15328));
  NAND2xp33_ASAP7_75t_L     g15072(.A(new_n15325), .B(new_n15328), .Y(new_n15329));
  A2O1A1Ixp33_ASAP7_75t_L   g15073(.A1(new_n14438), .A2(new_n14188), .B(new_n14435), .C(new_n14475), .Y(new_n15330));
  A2O1A1Ixp33_ASAP7_75t_L   g15074(.A1(new_n15330), .A2(new_n14474), .B(new_n15024), .C(new_n15023), .Y(new_n15331));
  A2O1A1Ixp33_ASAP7_75t_L   g15075(.A1(new_n14758), .A2(new_n15029), .B(new_n15027), .C(new_n15331), .Y(new_n15332));
  INVx1_ASAP7_75t_L         g15076(.A(new_n15332), .Y(new_n15333));
  NAND2xp33_ASAP7_75t_L     g15077(.A(new_n15328), .B(new_n15333), .Y(new_n15334));
  O2A1O1Ixp33_ASAP7_75t_L   g15078(.A1(new_n15321), .A2(new_n15324), .B(new_n15033), .C(new_n15334), .Y(new_n15335));
  A2O1A1O1Ixp25_ASAP7_75t_L g15079(.A1(new_n15020), .A2(new_n15023), .B(new_n15028), .C(new_n15329), .D(new_n15335), .Y(\f[71] ));
  NAND2xp33_ASAP7_75t_L     g15080(.A(new_n15320), .B(new_n15327), .Y(new_n15337));
  A2O1A1O1Ixp25_ASAP7_75t_L g15081(.A1(new_n15032), .A2(new_n15003), .B(new_n15008), .C(new_n15017), .D(new_n15337), .Y(new_n15338));
  O2A1O1Ixp33_ASAP7_75t_L   g15082(.A1(new_n15337), .A2(new_n15338), .B(new_n15325), .C(new_n15333), .Y(new_n15339));
  AOI31xp33_ASAP7_75t_L     g15083(.A1(new_n15044), .A2(new_n15313), .A3(new_n15319), .B(new_n15041), .Y(new_n15340));
  INVx1_ASAP7_75t_L         g15084(.A(new_n15340), .Y(new_n15341));
  OAI22xp33_ASAP7_75t_L     g15085(.A1(new_n1550), .A2(new_n12603), .B1(new_n12258), .B2(new_n712), .Y(new_n15342));
  AOI221xp5_ASAP7_75t_L     g15086(.A1(new_n640), .A2(\b[63] ), .B1(new_n718), .B2(new_n12961), .C(new_n15342), .Y(new_n15343));
  XNOR2x2_ASAP7_75t_L       g15087(.A(new_n637), .B(new_n15343), .Y(new_n15344));
  INVx1_ASAP7_75t_L         g15088(.A(new_n15344), .Y(new_n15345));
  A2O1A1O1Ixp25_ASAP7_75t_L g15089(.A1(new_n15318), .A2(new_n15317), .B(new_n15314), .C(new_n15311), .D(new_n15344), .Y(new_n15346));
  INVx1_ASAP7_75t_L         g15090(.A(new_n15346), .Y(new_n15347));
  A2O1A1O1Ixp25_ASAP7_75t_L g15091(.A1(new_n15318), .A2(new_n15317), .B(new_n15314), .C(new_n15311), .D(new_n15345), .Y(new_n15348));
  A2O1A1Ixp33_ASAP7_75t_L   g15092(.A1(new_n14788), .A2(new_n14787), .B(new_n14790), .C(new_n14995), .Y(new_n15349));
  O2A1O1Ixp33_ASAP7_75t_L   g15093(.A1(new_n872), .A2(new_n11597), .B(new_n15289), .C(new_n867), .Y(new_n15350));
  NOR2xp33_ASAP7_75t_L      g15094(.A(new_n867), .B(new_n15350), .Y(new_n15351));
  A2O1A1O1Ixp25_ASAP7_75t_L g15095(.A1(new_n12577), .A2(new_n873), .B(new_n15290), .C(new_n15291), .D(new_n15351), .Y(new_n15352));
  A2O1A1O1Ixp25_ASAP7_75t_L g15096(.A1(new_n14788), .A2(new_n14787), .B(new_n14790), .C(new_n14995), .D(new_n15352), .Y(new_n15353));
  A2O1A1Ixp33_ASAP7_75t_L   g15097(.A1(new_n14791), .A2(new_n14994), .B(new_n15293), .C(new_n15295), .Y(new_n15354));
  O2A1O1Ixp33_ASAP7_75t_L   g15098(.A1(new_n15352), .A2(new_n15353), .B(new_n15354), .C(new_n15299), .Y(new_n15355));
  OAI22xp33_ASAP7_75t_L     g15099(.A1(new_n980), .A2(new_n11303), .B1(new_n11591), .B2(new_n864), .Y(new_n15356));
  AOI221xp5_ASAP7_75t_L     g15100(.A1(new_n886), .A2(\b[60] ), .B1(new_n873), .B2(new_n13839), .C(new_n15356), .Y(new_n15357));
  XNOR2x2_ASAP7_75t_L       g15101(.A(new_n867), .B(new_n15357), .Y(new_n15358));
  A2O1A1Ixp33_ASAP7_75t_L   g15102(.A1(new_n15349), .A2(new_n15294), .B(new_n15355), .C(new_n15358), .Y(new_n15359));
  A2O1A1Ixp33_ASAP7_75t_L   g15103(.A1(new_n15291), .A2(\a[14] ), .B(new_n15292), .C(new_n15295), .Y(new_n15360));
  NAND2xp33_ASAP7_75t_L     g15104(.A(new_n15360), .B(new_n15354), .Y(new_n15361));
  A2O1A1O1Ixp25_ASAP7_75t_L g15105(.A1(new_n15285), .A2(new_n15274), .B(new_n15287), .C(new_n15361), .D(new_n15353), .Y(new_n15362));
  INVx1_ASAP7_75t_L         g15106(.A(new_n15358), .Y(new_n15363));
  NAND2xp33_ASAP7_75t_L     g15107(.A(new_n15363), .B(new_n15362), .Y(new_n15364));
  OAI22xp33_ASAP7_75t_L     g15108(.A1(new_n1285), .A2(new_n10309), .B1(new_n10332), .B2(new_n2118), .Y(new_n15365));
  AOI221xp5_ASAP7_75t_L     g15109(.A1(new_n1209), .A2(\b[57] ), .B1(new_n1216), .B2(new_n10991), .C(new_n15365), .Y(new_n15366));
  XNOR2x2_ASAP7_75t_L       g15110(.A(new_n1206), .B(new_n15366), .Y(new_n15367));
  INVx1_ASAP7_75t_L         g15111(.A(new_n15367), .Y(new_n15368));
  AOI211xp5_ASAP7_75t_L     g15112(.A1(new_n15274), .A2(new_n15283), .B(new_n15368), .C(new_n15286), .Y(new_n15369));
  A2O1A1Ixp33_ASAP7_75t_L   g15113(.A1(new_n15274), .A2(new_n15283), .B(new_n15286), .C(new_n15368), .Y(new_n15370));
  INVx1_ASAP7_75t_L         g15114(.A(new_n15370), .Y(new_n15371));
  NOR2xp33_ASAP7_75t_L      g15115(.A(new_n15369), .B(new_n15371), .Y(new_n15372));
  OAI22xp33_ASAP7_75t_L     g15116(.A1(new_n1654), .A2(new_n9355), .B1(new_n9683), .B2(new_n1517), .Y(new_n15373));
  AOI221xp5_ASAP7_75t_L     g15117(.A1(new_n1511), .A2(\b[54] ), .B1(new_n1513), .B2(new_n9717), .C(new_n15373), .Y(new_n15374));
  XNOR2x2_ASAP7_75t_L       g15118(.A(new_n1501), .B(new_n15374), .Y(new_n15375));
  A2O1A1O1Ixp25_ASAP7_75t_L g15119(.A1(new_n15270), .A2(new_n15265), .B(new_n15258), .C(new_n15272), .D(new_n15375), .Y(new_n15376));
  INVx1_ASAP7_75t_L         g15120(.A(new_n15376), .Y(new_n15377));
  A2O1A1Ixp33_ASAP7_75t_L   g15121(.A1(new_n15270), .A2(new_n15265), .B(new_n15258), .C(new_n15272), .Y(new_n15378));
  NOR2xp33_ASAP7_75t_L      g15122(.A(new_n15375), .B(new_n15378), .Y(new_n15379));
  O2A1O1Ixp33_ASAP7_75t_L   g15123(.A1(new_n15267), .A2(new_n15271), .B(new_n15377), .C(new_n15379), .Y(new_n15380));
  INVx1_ASAP7_75t_L         g15124(.A(new_n15380), .Y(new_n15381));
  INVx1_ASAP7_75t_L         g15125(.A(new_n15062), .Y(new_n15382));
  OAI22xp33_ASAP7_75t_L     g15126(.A1(new_n2089), .A2(new_n8427), .B1(new_n8755), .B2(new_n1962), .Y(new_n15383));
  AOI221xp5_ASAP7_75t_L     g15127(.A1(new_n1955), .A2(\b[51] ), .B1(new_n1964), .B2(new_n8790), .C(new_n15383), .Y(new_n15384));
  XNOR2x2_ASAP7_75t_L       g15128(.A(new_n1952), .B(new_n15384), .Y(new_n15385));
  A2O1A1O1Ixp25_ASAP7_75t_L g15129(.A1(new_n15247), .A2(new_n15243), .B(new_n15061), .C(new_n15382), .D(new_n15385), .Y(new_n15386));
  INVx1_ASAP7_75t_L         g15130(.A(new_n15386), .Y(new_n15387));
  INVx1_ASAP7_75t_L         g15131(.A(new_n15069), .Y(new_n15388));
  O2A1O1Ixp33_ASAP7_75t_L   g15132(.A1(new_n15250), .A2(new_n15388), .B(new_n15251), .C(new_n15254), .Y(new_n15389));
  O2A1O1Ixp33_ASAP7_75t_L   g15133(.A1(new_n15389), .A2(new_n15256), .B(new_n15249), .C(new_n15062), .Y(new_n15390));
  NAND2xp33_ASAP7_75t_L     g15134(.A(new_n15385), .B(new_n15390), .Y(new_n15391));
  AND2x2_ASAP7_75t_L        g15135(.A(new_n15387), .B(new_n15391), .Y(new_n15392));
  OAI22xp33_ASAP7_75t_L     g15136(.A1(new_n3133), .A2(new_n6671), .B1(new_n6944), .B2(new_n2925), .Y(new_n15393));
  AOI221xp5_ASAP7_75t_L     g15137(.A1(new_n2938), .A2(\b[45] ), .B1(new_n2932), .B2(new_n7256), .C(new_n15393), .Y(new_n15394));
  XNOR2x2_ASAP7_75t_L       g15138(.A(new_n2928), .B(new_n15394), .Y(new_n15395));
  INVx1_ASAP7_75t_L         g15139(.A(new_n15395), .Y(new_n15396));
  A2O1A1Ixp33_ASAP7_75t_L   g15140(.A1(new_n15240), .A2(new_n15235), .B(new_n15080), .C(new_n15396), .Y(new_n15397));
  O2A1O1Ixp33_ASAP7_75t_L   g15141(.A1(new_n15238), .A2(new_n15077), .B(new_n15236), .C(new_n15396), .Y(new_n15398));
  INVx1_ASAP7_75t_L         g15142(.A(new_n15205), .Y(new_n15399));
  A2O1A1Ixp33_ASAP7_75t_L   g15143(.A1(new_n14966), .A2(new_n14965), .B(new_n15399), .C(new_n15201), .Y(new_n15400));
  A2O1A1Ixp33_ASAP7_75t_L   g15144(.A1(new_n15212), .A2(new_n15214), .B(new_n15207), .C(new_n15400), .Y(new_n15401));
  INVx1_ASAP7_75t_L         g15145(.A(new_n15401), .Y(new_n15402));
  INVx1_ASAP7_75t_L         g15146(.A(new_n15189), .Y(new_n15403));
  INVx1_ASAP7_75t_L         g15147(.A(new_n15193), .Y(new_n15404));
  O2A1O1Ixp33_ASAP7_75t_L   g15148(.A1(new_n15197), .A2(new_n5626), .B(new_n15199), .C(new_n15194), .Y(new_n15405));
  NOR2xp33_ASAP7_75t_L      g15149(.A(new_n3891), .B(new_n5640), .Y(new_n15406));
  AOI221xp5_ASAP7_75t_L     g15150(.A1(\b[31] ), .A2(new_n5920), .B1(\b[33] ), .B2(new_n5629), .C(new_n15406), .Y(new_n15407));
  INVx1_ASAP7_75t_L         g15151(.A(new_n15407), .Y(new_n15408));
  A2O1A1Ixp33_ASAP7_75t_L   g15152(.A1(new_n4831), .A2(new_n5637), .B(new_n15408), .C(\a[41] ), .Y(new_n15409));
  O2A1O1Ixp33_ASAP7_75t_L   g15153(.A1(new_n5630), .A2(new_n4108), .B(new_n15407), .C(\a[41] ), .Y(new_n15410));
  O2A1O1Ixp33_ASAP7_75t_L   g15154(.A1(new_n15171), .A2(new_n15177), .B(new_n15179), .C(new_n15181), .Y(new_n15411));
  INVx1_ASAP7_75t_L         g15155(.A(new_n15411), .Y(new_n15412));
  A2O1A1Ixp33_ASAP7_75t_L   g15156(.A1(\a[44] ), .A2(new_n15186), .B(new_n15187), .C(new_n15182), .Y(new_n15413));
  A2O1A1Ixp33_ASAP7_75t_L   g15157(.A1(new_n15162), .A2(new_n15161), .B(new_n15164), .C(new_n15159), .Y(new_n15414));
  O2A1O1Ixp33_ASAP7_75t_L   g15158(.A1(new_n15108), .A2(new_n15116), .B(new_n15122), .C(new_n15120), .Y(new_n15415));
  O2A1O1Ixp33_ASAP7_75t_L   g15159(.A1(new_n15129), .A2(new_n15130), .B(new_n15125), .C(new_n15415), .Y(new_n15416));
  INVx1_ASAP7_75t_L         g15160(.A(new_n15416), .Y(new_n15417));
  NAND2xp33_ASAP7_75t_L     g15161(.A(\b[12] ), .B(new_n11995), .Y(new_n15418));
  OAI221xp5_ASAP7_75t_L     g15162(.A1(new_n12318), .A2(new_n748), .B1(new_n680), .B2(new_n12320), .C(new_n15418), .Y(new_n15419));
  A2O1A1Ixp33_ASAP7_75t_L   g15163(.A1(new_n1057), .A2(new_n11997), .B(new_n15419), .C(\a[62] ), .Y(new_n15420));
  NAND2xp33_ASAP7_75t_L     g15164(.A(\a[62] ), .B(new_n15420), .Y(new_n15421));
  A2O1A1Ixp33_ASAP7_75t_L   g15165(.A1(new_n1057), .A2(new_n11997), .B(new_n15419), .C(new_n11987), .Y(new_n15422));
  NAND2xp33_ASAP7_75t_L     g15166(.A(new_n15422), .B(new_n15421), .Y(new_n15423));
  NOR2xp33_ASAP7_75t_L      g15167(.A(new_n534), .B(new_n13030), .Y(new_n15424));
  O2A1O1Ixp33_ASAP7_75t_L   g15168(.A1(new_n534), .A2(new_n12672), .B(new_n15107), .C(new_n466), .Y(new_n15425));
  AOI211xp5_ASAP7_75t_L     g15169(.A1(new_n13028), .A2(\b[8] ), .B(new_n15106), .C(\a[8] ), .Y(new_n15426));
  NOR2xp33_ASAP7_75t_L      g15170(.A(new_n15426), .B(new_n15425), .Y(new_n15427));
  INVx1_ASAP7_75t_L         g15171(.A(new_n15427), .Y(new_n15428));
  A2O1A1Ixp33_ASAP7_75t_L   g15172(.A1(new_n13028), .A2(\b[9] ), .B(new_n15424), .C(new_n15428), .Y(new_n15429));
  O2A1O1Ixp33_ASAP7_75t_L   g15173(.A1(new_n12669), .A2(new_n12671), .B(\b[9] ), .C(new_n15424), .Y(new_n15430));
  NAND2xp33_ASAP7_75t_L     g15174(.A(new_n15430), .B(new_n15427), .Y(new_n15431));
  AND2x2_ASAP7_75t_L        g15175(.A(new_n15431), .B(new_n15429), .Y(new_n15432));
  A2O1A1Ixp33_ASAP7_75t_L   g15176(.A1(new_n15105), .A2(new_n15109), .B(new_n15112), .C(new_n15432), .Y(new_n15433));
  A2O1A1O1Ixp25_ASAP7_75t_L g15177(.A1(new_n14871), .A2(new_n14878), .B(new_n14868), .C(new_n15109), .D(new_n15112), .Y(new_n15434));
  INVx1_ASAP7_75t_L         g15178(.A(new_n15432), .Y(new_n15435));
  NAND2xp33_ASAP7_75t_L     g15179(.A(new_n15435), .B(new_n15434), .Y(new_n15436));
  NAND2xp33_ASAP7_75t_L     g15180(.A(new_n15433), .B(new_n15436), .Y(new_n15437));
  XNOR2x2_ASAP7_75t_L       g15181(.A(new_n15423), .B(new_n15437), .Y(new_n15438));
  NOR2xp33_ASAP7_75t_L      g15182(.A(new_n936), .B(new_n11354), .Y(new_n15439));
  AOI221xp5_ASAP7_75t_L     g15183(.A1(\b[15] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[14] ), .C(new_n15439), .Y(new_n15440));
  O2A1O1Ixp33_ASAP7_75t_L   g15184(.A1(new_n11053), .A2(new_n1774), .B(new_n15440), .C(new_n11048), .Y(new_n15441));
  INVx1_ASAP7_75t_L         g15185(.A(new_n15441), .Y(new_n15442));
  O2A1O1Ixp33_ASAP7_75t_L   g15186(.A1(new_n11053), .A2(new_n1774), .B(new_n15440), .C(\a[59] ), .Y(new_n15443));
  AOI21xp33_ASAP7_75t_L     g15187(.A1(new_n15442), .A2(\a[59] ), .B(new_n15443), .Y(new_n15444));
  XNOR2x2_ASAP7_75t_L       g15188(.A(new_n15438), .B(new_n15444), .Y(new_n15445));
  NAND2xp33_ASAP7_75t_L     g15189(.A(new_n15417), .B(new_n15445), .Y(new_n15446));
  INVx1_ASAP7_75t_L         g15190(.A(new_n15445), .Y(new_n15447));
  NAND2xp33_ASAP7_75t_L     g15191(.A(new_n15416), .B(new_n15447), .Y(new_n15448));
  NAND2xp33_ASAP7_75t_L     g15192(.A(new_n15446), .B(new_n15448), .Y(new_n15449));
  INVx1_ASAP7_75t_L         g15193(.A(new_n15449), .Y(new_n15450));
  NOR2xp33_ASAP7_75t_L      g15194(.A(new_n1349), .B(new_n10388), .Y(new_n15451));
  AOI221xp5_ASAP7_75t_L     g15195(.A1(new_n10086), .A2(\b[18] ), .B1(new_n11361), .B2(\b[16] ), .C(new_n15451), .Y(new_n15452));
  O2A1O1Ixp33_ASAP7_75t_L   g15196(.A1(new_n10088), .A2(new_n1464), .B(new_n15452), .C(new_n10083), .Y(new_n15453));
  INVx1_ASAP7_75t_L         g15197(.A(new_n15453), .Y(new_n15454));
  O2A1O1Ixp33_ASAP7_75t_L   g15198(.A1(new_n10088), .A2(new_n1464), .B(new_n15452), .C(\a[56] ), .Y(new_n15455));
  A2O1A1Ixp33_ASAP7_75t_L   g15199(.A1(\a[56] ), .A2(new_n15454), .B(new_n15455), .C(new_n15450), .Y(new_n15456));
  INVx1_ASAP7_75t_L         g15200(.A(new_n15456), .Y(new_n15457));
  A2O1A1Ixp33_ASAP7_75t_L   g15201(.A1(\a[56] ), .A2(new_n15454), .B(new_n15455), .C(new_n15449), .Y(new_n15458));
  A2O1A1O1Ixp25_ASAP7_75t_L g15202(.A1(new_n15140), .A2(\a[56] ), .B(new_n15141), .C(new_n15136), .D(new_n15135), .Y(new_n15459));
  OAI211xp5_ASAP7_75t_L     g15203(.A1(new_n15449), .A2(new_n15457), .B(new_n15458), .C(new_n15459), .Y(new_n15460));
  INVx1_ASAP7_75t_L         g15204(.A(new_n15458), .Y(new_n15461));
  INVx1_ASAP7_75t_L         g15205(.A(new_n15459), .Y(new_n15462));
  A2O1A1Ixp33_ASAP7_75t_L   g15206(.A1(new_n15456), .A2(new_n15450), .B(new_n15461), .C(new_n15462), .Y(new_n15463));
  AND2x2_ASAP7_75t_L        g15207(.A(new_n15463), .B(new_n15460), .Y(new_n15464));
  NOR2xp33_ASAP7_75t_L      g15208(.A(new_n1745), .B(new_n10400), .Y(new_n15465));
  AOI221xp5_ASAP7_75t_L     g15209(.A1(new_n9102), .A2(\b[21] ), .B1(new_n10398), .B2(\b[19] ), .C(new_n15465), .Y(new_n15466));
  O2A1O1Ixp33_ASAP7_75t_L   g15210(.A1(new_n9104), .A2(new_n1901), .B(new_n15466), .C(new_n9099), .Y(new_n15467));
  INVx1_ASAP7_75t_L         g15211(.A(new_n15467), .Y(new_n15468));
  O2A1O1Ixp33_ASAP7_75t_L   g15212(.A1(new_n9104), .A2(new_n1901), .B(new_n15466), .C(\a[53] ), .Y(new_n15469));
  A2O1A1Ixp33_ASAP7_75t_L   g15213(.A1(\a[53] ), .A2(new_n15468), .B(new_n15469), .C(new_n15464), .Y(new_n15470));
  INVx1_ASAP7_75t_L         g15214(.A(new_n15469), .Y(new_n15471));
  O2A1O1Ixp33_ASAP7_75t_L   g15215(.A1(new_n15467), .A2(new_n9099), .B(new_n15471), .C(new_n15464), .Y(new_n15472));
  AO21x2_ASAP7_75t_L        g15216(.A1(new_n15464), .A2(new_n15470), .B(new_n15472), .Y(new_n15473));
  O2A1O1Ixp33_ASAP7_75t_L   g15217(.A1(new_n15153), .A2(new_n15154), .B(new_n15149), .C(new_n15148), .Y(new_n15474));
  XNOR2x2_ASAP7_75t_L       g15218(.A(new_n15474), .B(new_n15473), .Y(new_n15475));
  NOR2xp33_ASAP7_75t_L      g15219(.A(new_n2188), .B(new_n10065), .Y(new_n15476));
  AOI221xp5_ASAP7_75t_L     g15220(.A1(new_n8175), .A2(\b[24] ), .B1(new_n8484), .B2(\b[22] ), .C(new_n15476), .Y(new_n15477));
  O2A1O1Ixp33_ASAP7_75t_L   g15221(.A1(new_n8176), .A2(new_n2853), .B(new_n15477), .C(new_n8172), .Y(new_n15478));
  INVx1_ASAP7_75t_L         g15222(.A(new_n15478), .Y(new_n15479));
  O2A1O1Ixp33_ASAP7_75t_L   g15223(.A1(new_n8176), .A2(new_n2853), .B(new_n15477), .C(\a[50] ), .Y(new_n15480));
  A2O1A1Ixp33_ASAP7_75t_L   g15224(.A1(new_n15479), .A2(\a[50] ), .B(new_n15480), .C(new_n15475), .Y(new_n15481));
  INVx1_ASAP7_75t_L         g15225(.A(new_n15480), .Y(new_n15482));
  O2A1O1Ixp33_ASAP7_75t_L   g15226(.A1(new_n8172), .A2(new_n15478), .B(new_n15482), .C(new_n15475), .Y(new_n15483));
  A2O1A1Ixp33_ASAP7_75t_L   g15227(.A1(new_n15481), .A2(new_n15475), .B(new_n15483), .C(new_n15414), .Y(new_n15484));
  AOI21xp33_ASAP7_75t_L     g15228(.A1(new_n15479), .A2(\a[50] ), .B(new_n15480), .Y(new_n15485));
  NOR2xp33_ASAP7_75t_L      g15229(.A(new_n8172), .B(new_n15478), .Y(new_n15486));
  OA21x2_ASAP7_75t_L        g15230(.A1(new_n15486), .A2(new_n15480), .B(new_n15475), .Y(new_n15487));
  NAND2xp33_ASAP7_75t_L     g15231(.A(new_n15485), .B(new_n15475), .Y(new_n15488));
  O2A1O1Ixp33_ASAP7_75t_L   g15232(.A1(new_n15485), .A2(new_n15487), .B(new_n15488), .C(new_n15414), .Y(new_n15489));
  NOR2xp33_ASAP7_75t_L      g15233(.A(new_n2703), .B(new_n7312), .Y(new_n15490));
  AOI221xp5_ASAP7_75t_L     g15234(.A1(\b[25] ), .A2(new_n7609), .B1(\b[27] ), .B2(new_n7334), .C(new_n15490), .Y(new_n15491));
  INVx1_ASAP7_75t_L         g15235(.A(new_n15491), .Y(new_n15492));
  A2O1A1Ixp33_ASAP7_75t_L   g15236(.A1(new_n2887), .A2(new_n7322), .B(new_n15492), .C(\a[47] ), .Y(new_n15493));
  O2A1O1Ixp33_ASAP7_75t_L   g15237(.A1(new_n7321), .A2(new_n2889), .B(new_n15491), .C(\a[47] ), .Y(new_n15494));
  AO21x2_ASAP7_75t_L        g15238(.A1(\a[47] ), .A2(new_n15493), .B(new_n15494), .Y(new_n15495));
  A2O1A1Ixp33_ASAP7_75t_L   g15239(.A1(new_n15484), .A2(new_n15414), .B(new_n15489), .C(new_n15495), .Y(new_n15496));
  A2O1A1Ixp33_ASAP7_75t_L   g15240(.A1(new_n15484), .A2(new_n15414), .B(new_n15489), .C(new_n15496), .Y(new_n15497));
  A2O1A1Ixp33_ASAP7_75t_L   g15241(.A1(new_n15493), .A2(\a[47] ), .B(new_n15494), .C(new_n15496), .Y(new_n15498));
  INVx1_ASAP7_75t_L         g15242(.A(new_n15168), .Y(new_n15499));
  A2O1A1O1Ixp25_ASAP7_75t_L g15243(.A1(new_n15178), .A2(\a[47] ), .B(new_n15175), .C(new_n15170), .D(new_n15499), .Y(new_n15500));
  NAND3xp33_ASAP7_75t_L     g15244(.A(new_n15500), .B(new_n15498), .C(new_n15497), .Y(new_n15501));
  NAND2xp33_ASAP7_75t_L     g15245(.A(new_n15498), .B(new_n15497), .Y(new_n15502));
  A2O1A1Ixp33_ASAP7_75t_L   g15246(.A1(new_n15167), .A2(new_n15096), .B(new_n15177), .C(new_n15502), .Y(new_n15503));
  NAND2xp33_ASAP7_75t_L     g15247(.A(new_n15501), .B(new_n15503), .Y(new_n15504));
  NOR2xp33_ASAP7_75t_L      g15248(.A(new_n3098), .B(new_n7304), .Y(new_n15505));
  AOI221xp5_ASAP7_75t_L     g15249(.A1(\b[28] ), .A2(new_n6742), .B1(\b[30] ), .B2(new_n6442), .C(new_n15505), .Y(new_n15506));
  O2A1O1Ixp33_ASAP7_75t_L   g15250(.A1(new_n6443), .A2(new_n3464), .B(new_n15506), .C(new_n6439), .Y(new_n15507));
  INVx1_ASAP7_75t_L         g15251(.A(new_n15506), .Y(new_n15508));
  A2O1A1Ixp33_ASAP7_75t_L   g15252(.A1(new_n4813), .A2(new_n6450), .B(new_n15508), .C(new_n6439), .Y(new_n15509));
  O2A1O1Ixp33_ASAP7_75t_L   g15253(.A1(new_n15507), .A2(new_n6439), .B(new_n15509), .C(new_n15504), .Y(new_n15510));
  OAI211xp5_ASAP7_75t_L     g15254(.A1(new_n6443), .A2(new_n3464), .B(\a[44] ), .C(new_n15506), .Y(new_n15511));
  AND3x1_ASAP7_75t_L        g15255(.A(new_n15504), .B(new_n15509), .C(new_n15511), .Y(new_n15512));
  INVx1_ASAP7_75t_L         g15256(.A(new_n15512), .Y(new_n15513));
  A2O1A1Ixp33_ASAP7_75t_L   g15257(.A1(new_n15182), .A2(new_n15188), .B(new_n15411), .C(new_n15513), .Y(new_n15514));
  NOR2xp33_ASAP7_75t_L      g15258(.A(new_n15510), .B(new_n15514), .Y(new_n15515));
  A2O1A1O1Ixp25_ASAP7_75t_L g15259(.A1(new_n15182), .A2(new_n15188), .B(new_n15411), .C(new_n15513), .D(new_n15510), .Y(new_n15516));
  NAND2xp33_ASAP7_75t_L     g15260(.A(new_n15513), .B(new_n15516), .Y(new_n15517));
  A2O1A1Ixp33_ASAP7_75t_L   g15261(.A1(new_n15413), .A2(new_n15412), .B(new_n15515), .C(new_n15517), .Y(new_n15518));
  A2O1A1Ixp33_ASAP7_75t_L   g15262(.A1(\a[41] ), .A2(new_n15409), .B(new_n15410), .C(new_n15518), .Y(new_n15519));
  A2O1A1O1Ixp25_ASAP7_75t_L g15263(.A1(new_n15186), .A2(\a[44] ), .B(new_n15187), .C(new_n15182), .D(new_n15411), .Y(new_n15520));
  AO21x2_ASAP7_75t_L        g15264(.A1(\a[41] ), .A2(new_n15409), .B(new_n15410), .Y(new_n15521));
  O2A1O1Ixp33_ASAP7_75t_L   g15265(.A1(new_n15520), .A2(new_n15515), .B(new_n15517), .C(new_n15521), .Y(new_n15522));
  A2O1A1O1Ixp25_ASAP7_75t_L g15266(.A1(new_n15409), .A2(\a[41] ), .B(new_n15410), .C(new_n15519), .D(new_n15522), .Y(new_n15523));
  A2O1A1Ixp33_ASAP7_75t_L   g15267(.A1(new_n15404), .A2(new_n15403), .B(new_n15405), .C(new_n15523), .Y(new_n15524));
  O2A1O1Ixp33_ASAP7_75t_L   g15268(.A1(new_n15191), .A2(new_n14962), .B(new_n15403), .C(new_n15405), .Y(new_n15525));
  A2O1A1Ixp33_ASAP7_75t_L   g15269(.A1(new_n15519), .A2(new_n15521), .B(new_n15522), .C(new_n15525), .Y(new_n15526));
  NOR2xp33_ASAP7_75t_L      g15270(.A(new_n4613), .B(new_n4908), .Y(new_n15527));
  AOI221xp5_ASAP7_75t_L     g15271(.A1(\b[34] ), .A2(new_n5139), .B1(\b[35] ), .B2(new_n4916), .C(new_n15527), .Y(new_n15528));
  O2A1O1Ixp33_ASAP7_75t_L   g15272(.A1(new_n4911), .A2(new_n4622), .B(new_n15528), .C(new_n4906), .Y(new_n15529));
  INVx1_ASAP7_75t_L         g15273(.A(new_n15529), .Y(new_n15530));
  O2A1O1Ixp33_ASAP7_75t_L   g15274(.A1(new_n4911), .A2(new_n4622), .B(new_n15528), .C(\a[38] ), .Y(new_n15531));
  AOI21xp33_ASAP7_75t_L     g15275(.A1(new_n15530), .A2(\a[38] ), .B(new_n15531), .Y(new_n15532));
  AOI21xp33_ASAP7_75t_L     g15276(.A1(new_n15524), .A2(new_n15526), .B(new_n15532), .Y(new_n15533));
  NAND3xp33_ASAP7_75t_L     g15277(.A(new_n15524), .B(new_n15526), .C(new_n15532), .Y(new_n15534));
  INVx1_ASAP7_75t_L         g15278(.A(new_n15534), .Y(new_n15535));
  OAI21xp33_ASAP7_75t_L     g15279(.A1(new_n15533), .A2(new_n15535), .B(new_n15402), .Y(new_n15536));
  INVx1_ASAP7_75t_L         g15280(.A(new_n15533), .Y(new_n15537));
  NAND3xp33_ASAP7_75t_L     g15281(.A(new_n15537), .B(new_n15401), .C(new_n15534), .Y(new_n15538));
  NOR2xp33_ASAP7_75t_L      g15282(.A(new_n5570), .B(new_n4147), .Y(new_n15539));
  AOI221xp5_ASAP7_75t_L     g15283(.A1(\b[37] ), .A2(new_n4402), .B1(\b[38] ), .B2(new_n4155), .C(new_n15539), .Y(new_n15540));
  O2A1O1Ixp33_ASAP7_75t_L   g15284(.A1(new_n4150), .A2(new_n5578), .B(new_n15540), .C(new_n4145), .Y(new_n15541));
  NOR2xp33_ASAP7_75t_L      g15285(.A(new_n4145), .B(new_n15541), .Y(new_n15542));
  O2A1O1Ixp33_ASAP7_75t_L   g15286(.A1(new_n4150), .A2(new_n5578), .B(new_n15540), .C(\a[35] ), .Y(new_n15543));
  NOR2xp33_ASAP7_75t_L      g15287(.A(new_n15543), .B(new_n15542), .Y(new_n15544));
  AND3x1_ASAP7_75t_L        g15288(.A(new_n15538), .B(new_n15536), .C(new_n15544), .Y(new_n15545));
  AOI21xp33_ASAP7_75t_L     g15289(.A1(new_n15538), .A2(new_n15536), .B(new_n15544), .Y(new_n15546));
  O2A1O1Ixp33_ASAP7_75t_L   g15290(.A1(new_n15218), .A2(new_n14983), .B(new_n15216), .C(new_n15231), .Y(new_n15547));
  OA21x2_ASAP7_75t_L        g15291(.A1(new_n15546), .A2(new_n15545), .B(new_n15547), .Y(new_n15548));
  NOR3xp33_ASAP7_75t_L      g15292(.A(new_n15547), .B(new_n15546), .C(new_n15545), .Y(new_n15549));
  NOR2xp33_ASAP7_75t_L      g15293(.A(new_n15549), .B(new_n15548), .Y(new_n15550));
  OAI22xp33_ASAP7_75t_L     g15294(.A1(new_n3703), .A2(new_n5855), .B1(new_n6110), .B2(new_n3509), .Y(new_n15551));
  AOI221xp5_ASAP7_75t_L     g15295(.A1(new_n3503), .A2(\b[42] ), .B1(new_n3505), .B2(new_n6389), .C(new_n15551), .Y(new_n15552));
  XNOR2x2_ASAP7_75t_L       g15296(.A(new_n3493), .B(new_n15552), .Y(new_n15553));
  INVx1_ASAP7_75t_L         g15297(.A(new_n15088), .Y(new_n15554));
  INVx1_ASAP7_75t_L         g15298(.A(new_n15553), .Y(new_n15555));
  A2O1A1Ixp33_ASAP7_75t_L   g15299(.A1(new_n15091), .A2(new_n15554), .B(new_n15233), .C(new_n15555), .Y(new_n15556));
  INVx1_ASAP7_75t_L         g15300(.A(new_n15556), .Y(new_n15557));
  A2O1A1Ixp33_ASAP7_75t_L   g15301(.A1(new_n15091), .A2(new_n15554), .B(new_n15233), .C(new_n15553), .Y(new_n15558));
  O2A1O1Ixp33_ASAP7_75t_L   g15302(.A1(new_n15553), .A2(new_n15557), .B(new_n15558), .C(new_n15550), .Y(new_n15559));
  OAI31xp33_ASAP7_75t_L     g15303(.A1(new_n15093), .A2(new_n15232), .A3(new_n15231), .B(new_n15092), .Y(new_n15560));
  NOR2xp33_ASAP7_75t_L      g15304(.A(new_n15553), .B(new_n15560), .Y(new_n15561));
  A2O1A1Ixp33_ASAP7_75t_L   g15305(.A1(new_n15556), .A2(new_n15560), .B(new_n15561), .C(new_n15550), .Y(new_n15562));
  OA21x2_ASAP7_75t_L        g15306(.A1(new_n15550), .A2(new_n15559), .B(new_n15562), .Y(new_n15563));
  A2O1A1Ixp33_ASAP7_75t_L   g15307(.A1(new_n15397), .A2(new_n15396), .B(new_n15398), .C(new_n15563), .Y(new_n15564));
  INVx1_ASAP7_75t_L         g15308(.A(new_n15398), .Y(new_n15565));
  O2A1O1Ixp33_ASAP7_75t_L   g15309(.A1(new_n15082), .A2(new_n15078), .B(new_n15235), .C(new_n15080), .Y(new_n15566));
  NAND2xp33_ASAP7_75t_L     g15310(.A(new_n15396), .B(new_n15566), .Y(new_n15567));
  OAI21xp33_ASAP7_75t_L     g15311(.A1(new_n15550), .A2(new_n15559), .B(new_n15562), .Y(new_n15568));
  NAND3xp33_ASAP7_75t_L     g15312(.A(new_n15568), .B(new_n15567), .C(new_n15565), .Y(new_n15569));
  NAND2xp33_ASAP7_75t_L     g15313(.A(new_n15569), .B(new_n15564), .Y(new_n15570));
  OAI22xp33_ASAP7_75t_L     g15314(.A1(new_n2572), .A2(new_n7270), .B1(new_n7552), .B2(new_n2410), .Y(new_n15571));
  AOI221xp5_ASAP7_75t_L     g15315(.A1(new_n2423), .A2(\b[48] ), .B1(new_n2417), .B2(new_n11656), .C(new_n15571), .Y(new_n15572));
  XNOR2x2_ASAP7_75t_L       g15316(.A(new_n2413), .B(new_n15572), .Y(new_n15573));
  INVx1_ASAP7_75t_L         g15317(.A(new_n15573), .Y(new_n15574));
  INVx1_ASAP7_75t_L         g15318(.A(new_n15241), .Y(new_n15575));
  INVx1_ASAP7_75t_L         g15319(.A(new_n15246), .Y(new_n15576));
  A2O1A1Ixp33_ASAP7_75t_L   g15320(.A1(new_n15575), .A2(new_n15576), .B(new_n15245), .C(new_n15069), .Y(new_n15577));
  NOR2xp33_ASAP7_75t_L      g15321(.A(new_n15574), .B(new_n15577), .Y(new_n15578));
  INVx1_ASAP7_75t_L         g15322(.A(new_n15578), .Y(new_n15579));
  A2O1A1O1Ixp25_ASAP7_75t_L g15323(.A1(new_n15576), .A2(new_n15575), .B(new_n15245), .C(new_n15069), .D(new_n15573), .Y(new_n15580));
  INVx1_ASAP7_75t_L         g15324(.A(new_n15580), .Y(new_n15581));
  NAND3xp33_ASAP7_75t_L     g15325(.A(new_n15570), .B(new_n15581), .C(new_n15579), .Y(new_n15582));
  NOR3xp33_ASAP7_75t_L      g15326(.A(new_n15570), .B(new_n15580), .C(new_n15578), .Y(new_n15583));
  A2O1A1Ixp33_ASAP7_75t_L   g15327(.A1(new_n15582), .A2(new_n15570), .B(new_n15583), .C(new_n15392), .Y(new_n15584));
  INVx1_ASAP7_75t_L         g15328(.A(new_n15564), .Y(new_n15585));
  INVx1_ASAP7_75t_L         g15329(.A(new_n15569), .Y(new_n15586));
  O2A1O1Ixp33_ASAP7_75t_L   g15330(.A1(new_n15585), .A2(new_n15586), .B(new_n15582), .C(new_n15583), .Y(new_n15587));
  NOR2xp33_ASAP7_75t_L      g15331(.A(new_n15392), .B(new_n15587), .Y(new_n15588));
  A2O1A1Ixp33_ASAP7_75t_L   g15332(.A1(new_n15392), .A2(new_n15584), .B(new_n15588), .C(new_n15381), .Y(new_n15589));
  AOI21xp33_ASAP7_75t_L     g15333(.A1(new_n15584), .A2(new_n15392), .B(new_n15588), .Y(new_n15590));
  NOR2xp33_ASAP7_75t_L      g15334(.A(new_n15590), .B(new_n15381), .Y(new_n15591));
  A2O1A1Ixp33_ASAP7_75t_L   g15335(.A1(new_n15589), .A2(new_n15381), .B(new_n15591), .C(new_n15372), .Y(new_n15592));
  INVx1_ASAP7_75t_L         g15336(.A(new_n15375), .Y(new_n15593));
  A2O1A1O1Ixp25_ASAP7_75t_L g15337(.A1(new_n15270), .A2(new_n15265), .B(new_n15258), .C(new_n15272), .D(new_n15593), .Y(new_n15594));
  A2O1A1Ixp33_ASAP7_75t_L   g15338(.A1(new_n15377), .A2(new_n15593), .B(new_n15594), .C(new_n15590), .Y(new_n15595));
  A2O1A1Ixp33_ASAP7_75t_L   g15339(.A1(new_n15392), .A2(new_n15584), .B(new_n15588), .C(new_n15380), .Y(new_n15596));
  OAI211xp5_ASAP7_75t_L     g15340(.A1(new_n15371), .A2(new_n15369), .B(new_n15595), .C(new_n15596), .Y(new_n15597));
  AOI22xp33_ASAP7_75t_L     g15341(.A1(new_n15592), .A2(new_n15597), .B1(new_n15359), .B2(new_n15364), .Y(new_n15598));
  NAND4xp25_ASAP7_75t_L     g15342(.A(new_n15364), .B(new_n15359), .C(new_n15592), .D(new_n15597), .Y(new_n15599));
  INVx1_ASAP7_75t_L         g15343(.A(new_n15599), .Y(new_n15600));
  NOR2xp33_ASAP7_75t_L      g15344(.A(new_n15598), .B(new_n15600), .Y(new_n15601));
  A2O1A1Ixp33_ASAP7_75t_L   g15345(.A1(new_n15347), .A2(new_n15345), .B(new_n15348), .C(new_n15601), .Y(new_n15602));
  INVx1_ASAP7_75t_L         g15346(.A(new_n15348), .Y(new_n15603));
  O2A1O1Ixp33_ASAP7_75t_L   g15347(.A1(new_n15307), .A2(new_n15312), .B(new_n15301), .C(new_n15310), .Y(new_n15604));
  NAND2xp33_ASAP7_75t_L     g15348(.A(new_n15345), .B(new_n15604), .Y(new_n15605));
  INVx1_ASAP7_75t_L         g15349(.A(new_n15598), .Y(new_n15606));
  NAND2xp33_ASAP7_75t_L     g15350(.A(new_n15599), .B(new_n15606), .Y(new_n15607));
  NAND3xp33_ASAP7_75t_L     g15351(.A(new_n15607), .B(new_n15605), .C(new_n15603), .Y(new_n15608));
  NAND3xp33_ASAP7_75t_L     g15352(.A(new_n15341), .B(new_n15602), .C(new_n15608), .Y(new_n15609));
  O2A1O1Ixp33_ASAP7_75t_L   g15353(.A1(new_n15344), .A2(new_n15346), .B(new_n15603), .C(new_n15607), .Y(new_n15610));
  A2O1A1Ixp33_ASAP7_75t_L   g15354(.A1(new_n15313), .A2(new_n15311), .B(new_n15346), .C(new_n15605), .Y(new_n15611));
  NOR2xp33_ASAP7_75t_L      g15355(.A(new_n15601), .B(new_n15611), .Y(new_n15612));
  OAI21xp33_ASAP7_75t_L     g15356(.A1(new_n15610), .A2(new_n15612), .B(new_n15340), .Y(new_n15613));
  NAND2xp33_ASAP7_75t_L     g15357(.A(new_n15609), .B(new_n15613), .Y(new_n15614));
  NOR2xp33_ASAP7_75t_L      g15358(.A(new_n15610), .B(new_n15612), .Y(new_n15615));
  A2O1A1O1Ixp25_ASAP7_75t_L g15359(.A1(new_n15020), .A2(new_n15023), .B(new_n15028), .C(new_n15329), .D(new_n15338), .Y(new_n15616));
  A2O1A1Ixp33_ASAP7_75t_L   g15360(.A1(new_n15602), .A2(new_n15608), .B(new_n15341), .C(new_n15616), .Y(new_n15617));
  O2A1O1Ixp33_ASAP7_75t_L   g15361(.A1(new_n15041), .A2(new_n15321), .B(new_n15615), .C(new_n15617), .Y(new_n15618));
  O2A1O1Ixp33_ASAP7_75t_L   g15362(.A1(new_n15338), .A2(new_n15339), .B(new_n15614), .C(new_n15618), .Y(\f[72] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15363(.A1(new_n15348), .A2(new_n15345), .B(new_n15607), .C(new_n15346), .Y(new_n15620));
  NOR2xp33_ASAP7_75t_L      g15364(.A(new_n12258), .B(new_n869), .Y(new_n15621));
  AOI221xp5_ASAP7_75t_L     g15365(.A1(\b[59] ), .A2(new_n985), .B1(\b[60] ), .B2(new_n885), .C(new_n15621), .Y(new_n15622));
  O2A1O1Ixp33_ASAP7_75t_L   g15366(.A1(new_n872), .A2(new_n14764), .B(new_n15622), .C(new_n867), .Y(new_n15623));
  NOR2xp33_ASAP7_75t_L      g15367(.A(new_n867), .B(new_n15623), .Y(new_n15624));
  O2A1O1Ixp33_ASAP7_75t_L   g15368(.A1(new_n872), .A2(new_n14764), .B(new_n15622), .C(\a[14] ), .Y(new_n15625));
  NOR2xp33_ASAP7_75t_L      g15369(.A(new_n15625), .B(new_n15624), .Y(new_n15626));
  A2O1A1O1Ixp25_ASAP7_75t_L g15370(.A1(new_n15596), .A2(new_n15595), .B(new_n15369), .C(new_n15370), .D(new_n15626), .Y(new_n15627));
  INVx1_ASAP7_75t_L         g15371(.A(new_n15626), .Y(new_n15628));
  A2O1A1O1Ixp25_ASAP7_75t_L g15372(.A1(new_n15596), .A2(new_n15595), .B(new_n15369), .C(new_n15370), .D(new_n15628), .Y(new_n15629));
  INVx1_ASAP7_75t_L         g15373(.A(new_n15629), .Y(new_n15630));
  NAND2xp33_ASAP7_75t_L     g15374(.A(\b[52] ), .B(new_n1955), .Y(new_n15631));
  OAI221xp5_ASAP7_75t_L     g15375(.A1(new_n1962), .A2(new_n8779), .B1(new_n8755), .B2(new_n2089), .C(new_n15631), .Y(new_n15632));
  A2O1A1Ixp33_ASAP7_75t_L   g15376(.A1(new_n9367), .A2(new_n1964), .B(new_n15632), .C(\a[23] ), .Y(new_n15633));
  NAND2xp33_ASAP7_75t_L     g15377(.A(\a[23] ), .B(new_n15633), .Y(new_n15634));
  A2O1A1Ixp33_ASAP7_75t_L   g15378(.A1(new_n9367), .A2(new_n1964), .B(new_n15632), .C(new_n1952), .Y(new_n15635));
  O2A1O1Ixp33_ASAP7_75t_L   g15379(.A1(new_n15586), .A2(new_n15585), .B(new_n15579), .C(new_n15580), .Y(new_n15636));
  NAND3xp33_ASAP7_75t_L     g15380(.A(new_n15636), .B(new_n15635), .C(new_n15634), .Y(new_n15637));
  NAND2xp33_ASAP7_75t_L     g15381(.A(new_n15635), .B(new_n15634), .Y(new_n15638));
  A2O1A1Ixp33_ASAP7_75t_L   g15382(.A1(new_n15570), .A2(new_n15579), .B(new_n15580), .C(new_n15638), .Y(new_n15639));
  NAND2xp33_ASAP7_75t_L     g15383(.A(new_n15639), .B(new_n15637), .Y(new_n15640));
  NOR2xp33_ASAP7_75t_L      g15384(.A(new_n5855), .B(new_n4147), .Y(new_n15641));
  AOI221xp5_ASAP7_75t_L     g15385(.A1(\b[38] ), .A2(new_n4402), .B1(\b[39] ), .B2(new_n4155), .C(new_n15641), .Y(new_n15642));
  O2A1O1Ixp33_ASAP7_75t_L   g15386(.A1(new_n4150), .A2(new_n5862), .B(new_n15642), .C(new_n4145), .Y(new_n15643));
  NOR2xp33_ASAP7_75t_L      g15387(.A(new_n4145), .B(new_n15643), .Y(new_n15644));
  O2A1O1Ixp33_ASAP7_75t_L   g15388(.A1(new_n4150), .A2(new_n5862), .B(new_n15642), .C(\a[35] ), .Y(new_n15645));
  NOR2xp33_ASAP7_75t_L      g15389(.A(new_n15645), .B(new_n15644), .Y(new_n15646));
  INVx1_ASAP7_75t_L         g15390(.A(new_n15646), .Y(new_n15647));
  NOR2xp33_ASAP7_75t_L      g15391(.A(new_n15525), .B(new_n15523), .Y(new_n15648));
  A2O1A1O1Ixp25_ASAP7_75t_L g15392(.A1(new_n15409), .A2(\a[41] ), .B(new_n15410), .C(new_n15518), .D(new_n15648), .Y(new_n15649));
  NOR2xp33_ASAP7_75t_L      g15393(.A(new_n4344), .B(new_n5641), .Y(new_n15650));
  AOI221xp5_ASAP7_75t_L     g15394(.A1(\b[32] ), .A2(new_n5920), .B1(\b[33] ), .B2(new_n5623), .C(new_n15650), .Y(new_n15651));
  O2A1O1Ixp33_ASAP7_75t_L   g15395(.A1(new_n5630), .A2(new_n4352), .B(new_n15651), .C(new_n5626), .Y(new_n15652));
  INVx1_ASAP7_75t_L         g15396(.A(new_n15652), .Y(new_n15653));
  O2A1O1Ixp33_ASAP7_75t_L   g15397(.A1(new_n5630), .A2(new_n4352), .B(new_n15651), .C(\a[41] ), .Y(new_n15654));
  NOR2xp33_ASAP7_75t_L      g15398(.A(new_n590), .B(new_n13030), .Y(new_n15655));
  O2A1O1Ixp33_ASAP7_75t_L   g15399(.A1(new_n12669), .A2(new_n12671), .B(\b[10] ), .C(new_n15655), .Y(new_n15656));
  INVx1_ASAP7_75t_L         g15400(.A(new_n15656), .Y(new_n15657));
  O2A1O1Ixp33_ASAP7_75t_L   g15401(.A1(new_n534), .A2(new_n12672), .B(new_n15107), .C(\a[8] ), .Y(new_n15658));
  INVx1_ASAP7_75t_L         g15402(.A(new_n15658), .Y(new_n15659));
  O2A1O1Ixp33_ASAP7_75t_L   g15403(.A1(new_n15430), .A2(new_n15427), .B(new_n15659), .C(new_n15657), .Y(new_n15660));
  NOR2xp33_ASAP7_75t_L      g15404(.A(new_n15657), .B(new_n15660), .Y(new_n15661));
  O2A1O1Ixp33_ASAP7_75t_L   g15405(.A1(new_n15430), .A2(new_n15427), .B(new_n15659), .C(new_n15656), .Y(new_n15662));
  NOR2xp33_ASAP7_75t_L      g15406(.A(new_n833), .B(new_n12318), .Y(new_n15663));
  AOI221xp5_ASAP7_75t_L     g15407(.A1(new_n11995), .A2(\b[13] ), .B1(new_n13314), .B2(\b[11] ), .C(new_n15663), .Y(new_n15664));
  O2A1O1Ixp33_ASAP7_75t_L   g15408(.A1(new_n11998), .A2(new_n942), .B(new_n15664), .C(new_n11987), .Y(new_n15665));
  INVx1_ASAP7_75t_L         g15409(.A(new_n15664), .Y(new_n15666));
  A2O1A1Ixp33_ASAP7_75t_L   g15410(.A1(new_n1166), .A2(new_n11997), .B(new_n15666), .C(new_n11987), .Y(new_n15667));
  INVx1_ASAP7_75t_L         g15411(.A(new_n15429), .Y(new_n15668));
  INVx1_ASAP7_75t_L         g15412(.A(new_n15660), .Y(new_n15669));
  O2A1O1Ixp33_ASAP7_75t_L   g15413(.A1(new_n15658), .A2(new_n15668), .B(new_n15669), .C(new_n15661), .Y(new_n15670));
  O2A1O1Ixp33_ASAP7_75t_L   g15414(.A1(new_n11987), .A2(new_n15665), .B(new_n15667), .C(new_n15670), .Y(new_n15671));
  INVx1_ASAP7_75t_L         g15415(.A(new_n15671), .Y(new_n15672));
  O2A1O1Ixp33_ASAP7_75t_L   g15416(.A1(new_n11987), .A2(new_n15665), .B(new_n15667), .C(new_n15671), .Y(new_n15673));
  O2A1O1Ixp33_ASAP7_75t_L   g15417(.A1(new_n15661), .A2(new_n15662), .B(new_n15672), .C(new_n15673), .Y(new_n15674));
  INVx1_ASAP7_75t_L         g15418(.A(new_n15674), .Y(new_n15675));
  A2O1A1O1Ixp25_ASAP7_75t_L g15419(.A1(new_n15422), .A2(new_n15421), .B(new_n15437), .C(new_n15433), .D(new_n15674), .Y(new_n15676));
  INVx1_ASAP7_75t_L         g15420(.A(new_n15676), .Y(new_n15677));
  A2O1A1O1Ixp25_ASAP7_75t_L g15421(.A1(new_n15422), .A2(new_n15421), .B(new_n15437), .C(new_n15433), .D(new_n15675), .Y(new_n15678));
  AO21x2_ASAP7_75t_L        g15422(.A1(new_n15675), .A2(new_n15677), .B(new_n15678), .Y(new_n15679));
  NOR2xp33_ASAP7_75t_L      g15423(.A(new_n960), .B(new_n11354), .Y(new_n15680));
  AOI221xp5_ASAP7_75t_L     g15424(.A1(\b[16] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[15] ), .C(new_n15680), .Y(new_n15681));
  O2A1O1Ixp33_ASAP7_75t_L   g15425(.A1(new_n11053), .A2(new_n1161), .B(new_n15681), .C(new_n11048), .Y(new_n15682));
  INVx1_ASAP7_75t_L         g15426(.A(new_n15682), .Y(new_n15683));
  O2A1O1Ixp33_ASAP7_75t_L   g15427(.A1(new_n11053), .A2(new_n1161), .B(new_n15681), .C(\a[59] ), .Y(new_n15684));
  A2O1A1Ixp33_ASAP7_75t_L   g15428(.A1(\a[59] ), .A2(new_n15683), .B(new_n15684), .C(new_n15679), .Y(new_n15685));
  INVx1_ASAP7_75t_L         g15429(.A(new_n15684), .Y(new_n15686));
  O2A1O1Ixp33_ASAP7_75t_L   g15430(.A1(new_n15682), .A2(new_n11048), .B(new_n15686), .C(new_n15679), .Y(new_n15687));
  A2O1A1O1Ixp25_ASAP7_75t_L g15431(.A1(new_n15677), .A2(new_n15675), .B(new_n15678), .C(new_n15685), .D(new_n15687), .Y(new_n15688));
  INVx1_ASAP7_75t_L         g15432(.A(new_n15446), .Y(new_n15689));
  A2O1A1O1Ixp25_ASAP7_75t_L g15433(.A1(new_n15442), .A2(\a[59] ), .B(new_n15443), .C(new_n15438), .D(new_n15689), .Y(new_n15690));
  NAND2xp33_ASAP7_75t_L     g15434(.A(new_n15690), .B(new_n15688), .Y(new_n15691));
  INVx1_ASAP7_75t_L         g15435(.A(new_n15690), .Y(new_n15692));
  A2O1A1Ixp33_ASAP7_75t_L   g15436(.A1(new_n15685), .A2(new_n15679), .B(new_n15687), .C(new_n15692), .Y(new_n15693));
  AND2x2_ASAP7_75t_L        g15437(.A(new_n15691), .B(new_n15693), .Y(new_n15694));
  NOR2xp33_ASAP7_75t_L      g15438(.A(new_n1458), .B(new_n10388), .Y(new_n15695));
  AOI221xp5_ASAP7_75t_L     g15439(.A1(new_n10086), .A2(\b[19] ), .B1(new_n11361), .B2(\b[17] ), .C(new_n15695), .Y(new_n15696));
  O2A1O1Ixp33_ASAP7_75t_L   g15440(.A1(new_n10088), .A2(new_n1628), .B(new_n15696), .C(new_n10083), .Y(new_n15697));
  INVx1_ASAP7_75t_L         g15441(.A(new_n15697), .Y(new_n15698));
  O2A1O1Ixp33_ASAP7_75t_L   g15442(.A1(new_n10088), .A2(new_n1628), .B(new_n15696), .C(\a[56] ), .Y(new_n15699));
  A2O1A1Ixp33_ASAP7_75t_L   g15443(.A1(\a[56] ), .A2(new_n15698), .B(new_n15699), .C(new_n15694), .Y(new_n15700));
  INVx1_ASAP7_75t_L         g15444(.A(new_n15699), .Y(new_n15701));
  O2A1O1Ixp33_ASAP7_75t_L   g15445(.A1(new_n15697), .A2(new_n10083), .B(new_n15701), .C(new_n15694), .Y(new_n15702));
  AOI21xp33_ASAP7_75t_L     g15446(.A1(new_n15700), .A2(new_n15694), .B(new_n15702), .Y(new_n15703));
  O2A1O1Ixp33_ASAP7_75t_L   g15447(.A1(new_n15461), .A2(new_n15450), .B(new_n15462), .C(new_n15457), .Y(new_n15704));
  AND2x2_ASAP7_75t_L        g15448(.A(new_n15704), .B(new_n15703), .Y(new_n15705));
  A2O1A1O1Ixp25_ASAP7_75t_L g15449(.A1(new_n15458), .A2(new_n15449), .B(new_n15459), .C(new_n15456), .D(new_n15703), .Y(new_n15706));
  NOR2xp33_ASAP7_75t_L      g15450(.A(new_n15706), .B(new_n15705), .Y(new_n15707));
  NOR2xp33_ASAP7_75t_L      g15451(.A(new_n1895), .B(new_n10400), .Y(new_n15708));
  AOI221xp5_ASAP7_75t_L     g15452(.A1(new_n9102), .A2(\b[22] ), .B1(new_n10398), .B2(\b[20] ), .C(new_n15708), .Y(new_n15709));
  O2A1O1Ixp33_ASAP7_75t_L   g15453(.A1(new_n9104), .A2(new_n2522), .B(new_n15709), .C(new_n9099), .Y(new_n15710));
  INVx1_ASAP7_75t_L         g15454(.A(new_n15710), .Y(new_n15711));
  O2A1O1Ixp33_ASAP7_75t_L   g15455(.A1(new_n9104), .A2(new_n2522), .B(new_n15709), .C(\a[53] ), .Y(new_n15712));
  A2O1A1Ixp33_ASAP7_75t_L   g15456(.A1(\a[53] ), .A2(new_n15711), .B(new_n15712), .C(new_n15707), .Y(new_n15713));
  INVx1_ASAP7_75t_L         g15457(.A(new_n15712), .Y(new_n15714));
  O2A1O1Ixp33_ASAP7_75t_L   g15458(.A1(new_n15710), .A2(new_n9099), .B(new_n15714), .C(new_n15707), .Y(new_n15715));
  AOI21xp33_ASAP7_75t_L     g15459(.A1(new_n15713), .A2(new_n15707), .B(new_n15715), .Y(new_n15716));
  INVx1_ASAP7_75t_L         g15460(.A(new_n15474), .Y(new_n15717));
  A2O1A1Ixp33_ASAP7_75t_L   g15461(.A1(new_n15470), .A2(new_n15464), .B(new_n15472), .C(new_n15717), .Y(new_n15718));
  NAND2xp33_ASAP7_75t_L     g15462(.A(new_n15470), .B(new_n15718), .Y(new_n15719));
  INVx1_ASAP7_75t_L         g15463(.A(new_n15719), .Y(new_n15720));
  NAND2xp33_ASAP7_75t_L     g15464(.A(new_n15720), .B(new_n15716), .Y(new_n15721));
  A2O1A1Ixp33_ASAP7_75t_L   g15465(.A1(new_n15713), .A2(new_n15707), .B(new_n15715), .C(new_n15719), .Y(new_n15722));
  NAND2xp33_ASAP7_75t_L     g15466(.A(new_n15722), .B(new_n15721), .Y(new_n15723));
  NOR2xp33_ASAP7_75t_L      g15467(.A(new_n2205), .B(new_n10065), .Y(new_n15724));
  AOI221xp5_ASAP7_75t_L     g15468(.A1(new_n8175), .A2(\b[25] ), .B1(new_n8484), .B2(\b[23] ), .C(new_n15724), .Y(new_n15725));
  O2A1O1Ixp33_ASAP7_75t_L   g15469(.A1(new_n8176), .A2(new_n2385), .B(new_n15725), .C(new_n8172), .Y(new_n15726));
  INVx1_ASAP7_75t_L         g15470(.A(new_n15726), .Y(new_n15727));
  O2A1O1Ixp33_ASAP7_75t_L   g15471(.A1(new_n8176), .A2(new_n2385), .B(new_n15725), .C(\a[50] ), .Y(new_n15728));
  AO21x2_ASAP7_75t_L        g15472(.A1(\a[50] ), .A2(new_n15727), .B(new_n15728), .Y(new_n15729));
  NAND3xp33_ASAP7_75t_L     g15473(.A(new_n15721), .B(new_n15722), .C(new_n15729), .Y(new_n15730));
  INVx1_ASAP7_75t_L         g15474(.A(new_n15730), .Y(new_n15731));
  A2O1A1Ixp33_ASAP7_75t_L   g15475(.A1(\a[50] ), .A2(new_n15727), .B(new_n15728), .C(new_n15723), .Y(new_n15732));
  O2A1O1Ixp33_ASAP7_75t_L   g15476(.A1(new_n15475), .A2(new_n15483), .B(new_n15414), .C(new_n15487), .Y(new_n15733));
  OAI211xp5_ASAP7_75t_L     g15477(.A1(new_n15731), .A2(new_n15723), .B(new_n15732), .C(new_n15733), .Y(new_n15734));
  NOR2xp33_ASAP7_75t_L      g15478(.A(new_n15729), .B(new_n15723), .Y(new_n15735));
  INVx1_ASAP7_75t_L         g15479(.A(new_n15733), .Y(new_n15736));
  A2O1A1Ixp33_ASAP7_75t_L   g15480(.A1(new_n15730), .A2(new_n15729), .B(new_n15735), .C(new_n15736), .Y(new_n15737));
  NAND2xp33_ASAP7_75t_L     g15481(.A(new_n15737), .B(new_n15734), .Y(new_n15738));
  NOR2xp33_ASAP7_75t_L      g15482(.A(new_n2879), .B(new_n7312), .Y(new_n15739));
  AOI221xp5_ASAP7_75t_L     g15483(.A1(\b[26] ), .A2(new_n7609), .B1(\b[28] ), .B2(new_n7334), .C(new_n15739), .Y(new_n15740));
  O2A1O1Ixp33_ASAP7_75t_L   g15484(.A1(new_n7321), .A2(new_n3087), .B(new_n15740), .C(new_n7316), .Y(new_n15741));
  O2A1O1Ixp33_ASAP7_75t_L   g15485(.A1(new_n7321), .A2(new_n3087), .B(new_n15740), .C(\a[47] ), .Y(new_n15742));
  INVx1_ASAP7_75t_L         g15486(.A(new_n15742), .Y(new_n15743));
  O2A1O1Ixp33_ASAP7_75t_L   g15487(.A1(new_n15741), .A2(new_n7316), .B(new_n15743), .C(new_n15738), .Y(new_n15744));
  INVx1_ASAP7_75t_L         g15488(.A(new_n15740), .Y(new_n15745));
  A2O1A1Ixp33_ASAP7_75t_L   g15489(.A1(new_n3085), .A2(new_n7322), .B(new_n15745), .C(\a[47] ), .Y(new_n15746));
  A2O1A1Ixp33_ASAP7_75t_L   g15490(.A1(\a[47] ), .A2(new_n15746), .B(new_n15742), .C(new_n15738), .Y(new_n15747));
  OA21x2_ASAP7_75t_L        g15491(.A1(new_n15738), .A2(new_n15744), .B(new_n15747), .Y(new_n15748));
  A2O1A1Ixp33_ASAP7_75t_L   g15492(.A1(new_n15497), .A2(new_n15498), .B(new_n15500), .C(new_n15496), .Y(new_n15749));
  INVx1_ASAP7_75t_L         g15493(.A(new_n15749), .Y(new_n15750));
  NAND2xp33_ASAP7_75t_L     g15494(.A(new_n15750), .B(new_n15748), .Y(new_n15751));
  O2A1O1Ixp33_ASAP7_75t_L   g15495(.A1(new_n15738), .A2(new_n15744), .B(new_n15747), .C(new_n15750), .Y(new_n15752));
  INVx1_ASAP7_75t_L         g15496(.A(new_n15752), .Y(new_n15753));
  NAND2xp33_ASAP7_75t_L     g15497(.A(new_n15753), .B(new_n15751), .Y(new_n15754));
  INVx1_ASAP7_75t_L         g15498(.A(new_n15754), .Y(new_n15755));
  NOR2xp33_ASAP7_75t_L      g15499(.A(new_n3098), .B(new_n6741), .Y(new_n15756));
  AOI221xp5_ASAP7_75t_L     g15500(.A1(\b[31] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[30] ), .C(new_n15756), .Y(new_n15757));
  O2A1O1Ixp33_ASAP7_75t_L   g15501(.A1(new_n6443), .A2(new_n3681), .B(new_n15757), .C(new_n6439), .Y(new_n15758));
  INVx1_ASAP7_75t_L         g15502(.A(new_n15758), .Y(new_n15759));
  O2A1O1Ixp33_ASAP7_75t_L   g15503(.A1(new_n6443), .A2(new_n3681), .B(new_n15757), .C(\a[44] ), .Y(new_n15760));
  AOI211xp5_ASAP7_75t_L     g15504(.A1(new_n15759), .A2(\a[44] ), .B(new_n15760), .C(new_n15755), .Y(new_n15761));
  A2O1A1Ixp33_ASAP7_75t_L   g15505(.A1(\a[44] ), .A2(new_n15759), .B(new_n15760), .C(new_n15755), .Y(new_n15762));
  INVx1_ASAP7_75t_L         g15506(.A(new_n15762), .Y(new_n15763));
  NOR2xp33_ASAP7_75t_L      g15507(.A(new_n15761), .B(new_n15763), .Y(new_n15764));
  XNOR2x2_ASAP7_75t_L       g15508(.A(new_n15516), .B(new_n15764), .Y(new_n15765));
  A2O1A1Ixp33_ASAP7_75t_L   g15509(.A1(new_n15653), .A2(\a[41] ), .B(new_n15654), .C(new_n15765), .Y(new_n15766));
  NOR2xp33_ASAP7_75t_L      g15510(.A(new_n5626), .B(new_n15652), .Y(new_n15767));
  OR3x1_ASAP7_75t_L         g15511(.A(new_n15765), .B(new_n15767), .C(new_n15654), .Y(new_n15768));
  NAND2xp33_ASAP7_75t_L     g15512(.A(new_n15766), .B(new_n15768), .Y(new_n15769));
  O2A1O1Ixp33_ASAP7_75t_L   g15513(.A1(new_n15525), .A2(new_n15523), .B(new_n15519), .C(new_n15769), .Y(new_n15770));
  NOR2xp33_ASAP7_75t_L      g15514(.A(new_n5074), .B(new_n4908), .Y(new_n15771));
  AOI221xp5_ASAP7_75t_L     g15515(.A1(\b[35] ), .A2(new_n5139), .B1(\b[36] ), .B2(new_n4916), .C(new_n15771), .Y(new_n15772));
  O2A1O1Ixp33_ASAP7_75t_L   g15516(.A1(new_n4911), .A2(new_n5083), .B(new_n15772), .C(new_n4906), .Y(new_n15773));
  NOR2xp33_ASAP7_75t_L      g15517(.A(new_n4906), .B(new_n15773), .Y(new_n15774));
  O2A1O1Ixp33_ASAP7_75t_L   g15518(.A1(new_n4911), .A2(new_n5083), .B(new_n15772), .C(\a[38] ), .Y(new_n15775));
  NOR2xp33_ASAP7_75t_L      g15519(.A(new_n15775), .B(new_n15774), .Y(new_n15776));
  NAND3xp33_ASAP7_75t_L     g15520(.A(new_n15649), .B(new_n15766), .C(new_n15768), .Y(new_n15777));
  O2A1O1Ixp33_ASAP7_75t_L   g15521(.A1(new_n15649), .A2(new_n15770), .B(new_n15777), .C(new_n15776), .Y(new_n15778));
  AND2x2_ASAP7_75t_L        g15522(.A(new_n15776), .B(new_n15777), .Y(new_n15779));
  O2A1O1Ixp33_ASAP7_75t_L   g15523(.A1(new_n15770), .A2(new_n15649), .B(new_n15779), .C(new_n15778), .Y(new_n15780));
  A2O1A1Ixp33_ASAP7_75t_L   g15524(.A1(new_n15534), .A2(new_n15401), .B(new_n15533), .C(new_n15780), .Y(new_n15781));
  O2A1O1Ixp33_ASAP7_75t_L   g15525(.A1(new_n15402), .A2(new_n15535), .B(new_n15537), .C(new_n15780), .Y(new_n15782));
  A2O1A1Ixp33_ASAP7_75t_L   g15526(.A1(new_n15781), .A2(new_n15780), .B(new_n15782), .C(new_n15647), .Y(new_n15783));
  A2O1A1Ixp33_ASAP7_75t_L   g15527(.A1(new_n15521), .A2(new_n15518), .B(new_n15648), .C(new_n15769), .Y(new_n15784));
  AO21x2_ASAP7_75t_L        g15528(.A1(new_n15779), .A2(new_n15784), .B(new_n15778), .Y(new_n15785));
  O2A1O1Ixp33_ASAP7_75t_L   g15529(.A1(new_n15402), .A2(new_n15535), .B(new_n15537), .C(new_n15785), .Y(new_n15786));
  A2O1A1Ixp33_ASAP7_75t_L   g15530(.A1(new_n15534), .A2(new_n15401), .B(new_n15533), .C(new_n15785), .Y(new_n15787));
  O2A1O1Ixp33_ASAP7_75t_L   g15531(.A1(new_n15785), .A2(new_n15786), .B(new_n15787), .C(new_n15647), .Y(new_n15788));
  O2A1O1Ixp33_ASAP7_75t_L   g15532(.A1(new_n15644), .A2(new_n15645), .B(new_n15783), .C(new_n15788), .Y(new_n15789));
  NOR2xp33_ASAP7_75t_L      g15533(.A(new_n6378), .B(new_n3509), .Y(new_n15790));
  AOI221xp5_ASAP7_75t_L     g15534(.A1(\b[41] ), .A2(new_n3708), .B1(\b[43] ), .B2(new_n3503), .C(new_n15790), .Y(new_n15791));
  O2A1O1Ixp33_ASAP7_75t_L   g15535(.A1(new_n3513), .A2(new_n6679), .B(new_n15791), .C(new_n3493), .Y(new_n15792));
  INVx1_ASAP7_75t_L         g15536(.A(new_n15791), .Y(new_n15793));
  A2O1A1Ixp33_ASAP7_75t_L   g15537(.A1(new_n6682), .A2(new_n3505), .B(new_n15793), .C(new_n3493), .Y(new_n15794));
  OAI21xp33_ASAP7_75t_L     g15538(.A1(new_n3493), .A2(new_n15792), .B(new_n15794), .Y(new_n15795));
  NAND2xp33_ASAP7_75t_L     g15539(.A(new_n15536), .B(new_n15538), .Y(new_n15796));
  MAJIxp5_ASAP7_75t_L       g15540(.A(new_n15547), .B(new_n15544), .C(new_n15796), .Y(new_n15797));
  NOR2xp33_ASAP7_75t_L      g15541(.A(new_n15795), .B(new_n15797), .Y(new_n15798));
  AND2x2_ASAP7_75t_L        g15542(.A(new_n15795), .B(new_n15797), .Y(new_n15799));
  NOR2xp33_ASAP7_75t_L      g15543(.A(new_n15798), .B(new_n15799), .Y(new_n15800));
  A2O1A1Ixp33_ASAP7_75t_L   g15544(.A1(new_n15647), .A2(new_n15783), .B(new_n15788), .C(new_n15800), .Y(new_n15801));
  INVx1_ASAP7_75t_L         g15545(.A(new_n15801), .Y(new_n15802));
  NAND2xp33_ASAP7_75t_L     g15546(.A(new_n15800), .B(new_n15789), .Y(new_n15803));
  NAND2xp33_ASAP7_75t_L     g15547(.A(\b[45] ), .B(new_n2936), .Y(new_n15804));
  OAI221xp5_ASAP7_75t_L     g15548(.A1(new_n2930), .A2(new_n7270), .B1(new_n6944), .B2(new_n3133), .C(new_n15804), .Y(new_n15805));
  AOI21xp33_ASAP7_75t_L     g15549(.A1(new_n7278), .A2(new_n2932), .B(new_n15805), .Y(new_n15806));
  NAND2xp33_ASAP7_75t_L     g15550(.A(\a[29] ), .B(new_n15806), .Y(new_n15807));
  A2O1A1Ixp33_ASAP7_75t_L   g15551(.A1(new_n7278), .A2(new_n2932), .B(new_n15805), .C(new_n2928), .Y(new_n15808));
  NAND2xp33_ASAP7_75t_L     g15552(.A(new_n15808), .B(new_n15807), .Y(new_n15809));
  INVx1_ASAP7_75t_L         g15553(.A(new_n15809), .Y(new_n15810));
  A2O1A1O1Ixp25_ASAP7_75t_L g15554(.A1(new_n15558), .A2(new_n15553), .B(new_n15550), .C(new_n15556), .D(new_n15810), .Y(new_n15811));
  A2O1A1Ixp33_ASAP7_75t_L   g15555(.A1(new_n15555), .A2(new_n15560), .B(new_n15559), .C(new_n15810), .Y(new_n15812));
  A2O1A1Ixp33_ASAP7_75t_L   g15556(.A1(new_n15808), .A2(new_n15807), .B(new_n15811), .C(new_n15812), .Y(new_n15813));
  O2A1O1Ixp33_ASAP7_75t_L   g15557(.A1(new_n15789), .A2(new_n15802), .B(new_n15803), .C(new_n15813), .Y(new_n15814));
  O2A1O1Ixp33_ASAP7_75t_L   g15558(.A1(new_n15785), .A2(new_n15786), .B(new_n15787), .C(new_n15646), .Y(new_n15815));
  A2O1A1Ixp33_ASAP7_75t_L   g15559(.A1(new_n15781), .A2(new_n15780), .B(new_n15782), .C(new_n15646), .Y(new_n15816));
  O2A1O1Ixp33_ASAP7_75t_L   g15560(.A1(new_n15646), .A2(new_n15815), .B(new_n15816), .C(new_n15800), .Y(new_n15817));
  AO21x2_ASAP7_75t_L        g15561(.A1(new_n15800), .A2(new_n15801), .B(new_n15817), .Y(new_n15818));
  O2A1O1Ixp33_ASAP7_75t_L   g15562(.A1(new_n15810), .A2(new_n15811), .B(new_n15812), .C(new_n15818), .Y(new_n15819));
  NOR2xp33_ASAP7_75t_L      g15563(.A(new_n15819), .B(new_n15814), .Y(new_n15820));
  NOR2xp33_ASAP7_75t_L      g15564(.A(new_n8427), .B(new_n2415), .Y(new_n15821));
  AOI221xp5_ASAP7_75t_L     g15565(.A1(\b[47] ), .A2(new_n2577), .B1(\b[48] ), .B2(new_n2421), .C(new_n15821), .Y(new_n15822));
  O2A1O1Ixp33_ASAP7_75t_L   g15566(.A1(new_n2425), .A2(new_n14802), .B(new_n15822), .C(new_n2413), .Y(new_n15823));
  INVx1_ASAP7_75t_L         g15567(.A(new_n15823), .Y(new_n15824));
  O2A1O1Ixp33_ASAP7_75t_L   g15568(.A1(new_n2425), .A2(new_n14802), .B(new_n15822), .C(\a[26] ), .Y(new_n15825));
  AOI21xp33_ASAP7_75t_L     g15569(.A1(new_n15824), .A2(\a[26] ), .B(new_n15825), .Y(new_n15826));
  A2O1A1O1Ixp25_ASAP7_75t_L g15570(.A1(new_n15565), .A2(new_n15395), .B(new_n15563), .C(new_n15397), .D(new_n15826), .Y(new_n15827));
  INVx1_ASAP7_75t_L         g15571(.A(new_n15397), .Y(new_n15828));
  A2O1A1Ixp33_ASAP7_75t_L   g15572(.A1(new_n15236), .A2(new_n15081), .B(new_n15828), .C(new_n15567), .Y(new_n15829));
  A2O1A1Ixp33_ASAP7_75t_L   g15573(.A1(new_n15829), .A2(new_n15568), .B(new_n15828), .C(new_n15826), .Y(new_n15830));
  O2A1O1Ixp33_ASAP7_75t_L   g15574(.A1(new_n15826), .A2(new_n15827), .B(new_n15830), .C(new_n15820), .Y(new_n15831));
  O2A1O1Ixp33_ASAP7_75t_L   g15575(.A1(new_n15398), .A2(new_n15396), .B(new_n15568), .C(new_n15828), .Y(new_n15832));
  INVx1_ASAP7_75t_L         g15576(.A(new_n15832), .Y(new_n15833));
  INVx1_ASAP7_75t_L         g15577(.A(new_n15827), .Y(new_n15834));
  INVx1_ASAP7_75t_L         g15578(.A(new_n15825), .Y(new_n15835));
  O2A1O1Ixp33_ASAP7_75t_L   g15579(.A1(new_n2413), .A2(new_n15823), .B(new_n15835), .C(new_n15827), .Y(new_n15836));
  A2O1A1Ixp33_ASAP7_75t_L   g15580(.A1(new_n15834), .A2(new_n15833), .B(new_n15836), .C(new_n15820), .Y(new_n15837));
  O2A1O1Ixp33_ASAP7_75t_L   g15581(.A1(new_n15820), .A2(new_n15831), .B(new_n15837), .C(new_n15640), .Y(new_n15838));
  INVx1_ASAP7_75t_L         g15582(.A(new_n15811), .Y(new_n15839));
  A2O1A1Ixp33_ASAP7_75t_L   g15583(.A1(new_n15553), .A2(new_n15558), .B(new_n15550), .C(new_n15556), .Y(new_n15840));
  NOR2xp33_ASAP7_75t_L      g15584(.A(new_n15810), .B(new_n15840), .Y(new_n15841));
  O2A1O1Ixp33_ASAP7_75t_L   g15585(.A1(new_n15557), .A2(new_n15559), .B(new_n15839), .C(new_n15841), .Y(new_n15842));
  A2O1A1Ixp33_ASAP7_75t_L   g15586(.A1(new_n15801), .A2(new_n15800), .B(new_n15817), .C(new_n15842), .Y(new_n15843));
  O2A1O1Ixp33_ASAP7_75t_L   g15587(.A1(new_n15789), .A2(new_n15802), .B(new_n15803), .C(new_n15842), .Y(new_n15844));
  INVx1_ASAP7_75t_L         g15588(.A(new_n15844), .Y(new_n15845));
  A2O1A1Ixp33_ASAP7_75t_L   g15589(.A1(new_n15839), .A2(new_n15840), .B(new_n15841), .C(new_n15845), .Y(new_n15846));
  A2O1A1Ixp33_ASAP7_75t_L   g15590(.A1(new_n15846), .A2(new_n15843), .B(new_n15831), .C(new_n15837), .Y(new_n15847));
  AOI21xp33_ASAP7_75t_L     g15591(.A1(new_n15639), .A2(new_n15637), .B(new_n15847), .Y(new_n15848));
  INVx1_ASAP7_75t_L         g15592(.A(new_n10320), .Y(new_n15849));
  NOR2xp33_ASAP7_75t_L      g15593(.A(new_n10309), .B(new_n1518), .Y(new_n15850));
  AOI221xp5_ASAP7_75t_L     g15594(.A1(\b[53] ), .A2(new_n1659), .B1(\b[54] ), .B2(new_n1507), .C(new_n15850), .Y(new_n15851));
  O2A1O1Ixp33_ASAP7_75t_L   g15595(.A1(new_n1521), .A2(new_n15849), .B(new_n15851), .C(new_n1501), .Y(new_n15852));
  INVx1_ASAP7_75t_L         g15596(.A(new_n15852), .Y(new_n15853));
  O2A1O1Ixp33_ASAP7_75t_L   g15597(.A1(new_n1521), .A2(new_n15849), .B(new_n15851), .C(\a[20] ), .Y(new_n15854));
  AOI21xp33_ASAP7_75t_L     g15598(.A1(new_n15853), .A2(\a[20] ), .B(new_n15854), .Y(new_n15855));
  A2O1A1O1Ixp25_ASAP7_75t_L g15599(.A1(new_n15570), .A2(new_n15582), .B(new_n15583), .C(new_n15391), .D(new_n15386), .Y(new_n15856));
  AND2x2_ASAP7_75t_L        g15600(.A(new_n15855), .B(new_n15856), .Y(new_n15857));
  O2A1O1Ixp33_ASAP7_75t_L   g15601(.A1(new_n15385), .A2(new_n15390), .B(new_n15584), .C(new_n15855), .Y(new_n15858));
  NOR4xp25_ASAP7_75t_L      g15602(.A(new_n15858), .B(new_n15838), .C(new_n15848), .D(new_n15857), .Y(new_n15859));
  NOR2xp33_ASAP7_75t_L      g15603(.A(new_n15857), .B(new_n15858), .Y(new_n15860));
  OAI21xp33_ASAP7_75t_L     g15604(.A1(new_n15838), .A2(new_n15848), .B(new_n15860), .Y(new_n15861));
  OAI31xp33_ASAP7_75t_L     g15605(.A1(new_n15838), .A2(new_n15859), .A3(new_n15848), .B(new_n15861), .Y(new_n15862));
  NAND2xp33_ASAP7_75t_L     g15606(.A(\b[57] ), .B(new_n1204), .Y(new_n15863));
  OAI221xp5_ASAP7_75t_L     g15607(.A1(new_n1284), .A2(new_n11303), .B1(new_n10332), .B2(new_n1285), .C(new_n15863), .Y(new_n15864));
  AOI21xp33_ASAP7_75t_L     g15608(.A1(new_n11314), .A2(new_n1216), .B(new_n15864), .Y(new_n15865));
  NAND2xp33_ASAP7_75t_L     g15609(.A(\a[17] ), .B(new_n15865), .Y(new_n15866));
  A2O1A1Ixp33_ASAP7_75t_L   g15610(.A1(new_n11314), .A2(new_n1216), .B(new_n15864), .C(new_n1206), .Y(new_n15867));
  NAND2xp33_ASAP7_75t_L     g15611(.A(new_n15867), .B(new_n15866), .Y(new_n15868));
  O2A1O1Ixp33_ASAP7_75t_L   g15612(.A1(new_n15380), .A2(new_n15590), .B(new_n15377), .C(new_n15868), .Y(new_n15869));
  INVx1_ASAP7_75t_L         g15613(.A(new_n15594), .Y(new_n15870));
  A2O1A1Ixp33_ASAP7_75t_L   g15614(.A1(new_n15375), .A2(new_n15870), .B(new_n15590), .C(new_n15377), .Y(new_n15871));
  INVx1_ASAP7_75t_L         g15615(.A(new_n15868), .Y(new_n15872));
  NOR2xp33_ASAP7_75t_L      g15616(.A(new_n15872), .B(new_n15871), .Y(new_n15873));
  NOR2xp33_ASAP7_75t_L      g15617(.A(new_n15869), .B(new_n15873), .Y(new_n15874));
  XNOR2x2_ASAP7_75t_L       g15618(.A(new_n15862), .B(new_n15874), .Y(new_n15875));
  O2A1O1Ixp33_ASAP7_75t_L   g15619(.A1(new_n15626), .A2(new_n15627), .B(new_n15630), .C(new_n15875), .Y(new_n15876));
  INVx1_ASAP7_75t_L         g15620(.A(new_n15625), .Y(new_n15877));
  A2O1A1Ixp33_ASAP7_75t_L   g15621(.A1(new_n15595), .A2(new_n15596), .B(new_n15369), .C(new_n15370), .Y(new_n15878));
  O2A1O1Ixp33_ASAP7_75t_L   g15622(.A1(new_n867), .A2(new_n15623), .B(new_n15877), .C(new_n15878), .Y(new_n15879));
  XOR2x2_ASAP7_75t_L        g15623(.A(new_n15862), .B(new_n15874), .Y(new_n15880));
  NOR3xp33_ASAP7_75t_L      g15624(.A(new_n15880), .B(new_n15629), .C(new_n15879), .Y(new_n15881));
  NAND2xp33_ASAP7_75t_L     g15625(.A(new_n15359), .B(new_n15364), .Y(new_n15882));
  NAND3xp33_ASAP7_75t_L     g15626(.A(new_n15882), .B(new_n15592), .C(new_n15597), .Y(new_n15883));
  A2O1A1O1Ixp25_ASAP7_75t_L g15627(.A1(new_n15360), .A2(new_n15354), .B(new_n15299), .C(new_n15295), .D(new_n15358), .Y(new_n15884));
  INVx1_ASAP7_75t_L         g15628(.A(new_n15884), .Y(new_n15885));
  AOI22xp33_ASAP7_75t_L     g15629(.A1(new_n635), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n713), .Y(new_n15886));
  A2O1A1Ixp33_ASAP7_75t_L   g15630(.A1(new_n12990), .A2(new_n12988), .B(new_n641), .C(new_n15886), .Y(new_n15887));
  NOR2xp33_ASAP7_75t_L      g15631(.A(new_n637), .B(new_n15887), .Y(new_n15888));
  O2A1O1Ixp33_ASAP7_75t_L   g15632(.A1(new_n641), .A2(new_n12993), .B(new_n15886), .C(\a[11] ), .Y(new_n15889));
  NOR2xp33_ASAP7_75t_L      g15633(.A(new_n15889), .B(new_n15888), .Y(new_n15890));
  O2A1O1Ixp33_ASAP7_75t_L   g15634(.A1(new_n15362), .A2(new_n15358), .B(new_n15883), .C(new_n15890), .Y(new_n15891));
  INVx1_ASAP7_75t_L         g15635(.A(new_n15890), .Y(new_n15892));
  NAND3xp33_ASAP7_75t_L     g15636(.A(new_n15883), .B(new_n15885), .C(new_n15892), .Y(new_n15893));
  A2O1A1Ixp33_ASAP7_75t_L   g15637(.A1(new_n15885), .A2(new_n15883), .B(new_n15891), .C(new_n15893), .Y(new_n15894));
  INVx1_ASAP7_75t_L         g15638(.A(new_n15627), .Y(new_n15895));
  A2O1A1Ixp33_ASAP7_75t_L   g15639(.A1(new_n15895), .A2(new_n15878), .B(new_n15879), .C(new_n15880), .Y(new_n15896));
  O2A1O1Ixp33_ASAP7_75t_L   g15640(.A1(new_n15624), .A2(new_n15625), .B(new_n15895), .C(new_n15629), .Y(new_n15897));
  O2A1O1Ixp33_ASAP7_75t_L   g15641(.A1(new_n15375), .A2(new_n15376), .B(new_n15870), .C(new_n15590), .Y(new_n15898));
  A2O1A1Ixp33_ASAP7_75t_L   g15642(.A1(new_n15593), .A2(new_n15378), .B(new_n15898), .C(new_n15868), .Y(new_n15899));
  A2O1A1Ixp33_ASAP7_75t_L   g15643(.A1(new_n15871), .A2(new_n15899), .B(new_n15873), .C(new_n15862), .Y(new_n15900));
  O2A1O1Ixp33_ASAP7_75t_L   g15644(.A1(new_n15380), .A2(new_n15590), .B(new_n15377), .C(new_n15872), .Y(new_n15901));
  A2O1A1Ixp33_ASAP7_75t_L   g15645(.A1(new_n15593), .A2(new_n15378), .B(new_n15898), .C(new_n15872), .Y(new_n15902));
  O2A1O1Ixp33_ASAP7_75t_L   g15646(.A1(new_n15872), .A2(new_n15901), .B(new_n15902), .C(new_n15862), .Y(new_n15903));
  A2O1A1Ixp33_ASAP7_75t_L   g15647(.A1(new_n15862), .A2(new_n15900), .B(new_n15903), .C(new_n15897), .Y(new_n15904));
  NAND2xp33_ASAP7_75t_L     g15648(.A(new_n15904), .B(new_n15896), .Y(new_n15905));
  AND2x2_ASAP7_75t_L        g15649(.A(new_n15597), .B(new_n15882), .Y(new_n15906));
  A2O1A1Ixp33_ASAP7_75t_L   g15650(.A1(new_n15906), .A2(new_n15592), .B(new_n15884), .C(new_n15892), .Y(new_n15907));
  O2A1O1Ixp33_ASAP7_75t_L   g15651(.A1(new_n15362), .A2(new_n15358), .B(new_n15883), .C(new_n15892), .Y(new_n15908));
  AOI211xp5_ASAP7_75t_L     g15652(.A1(new_n15892), .A2(new_n15907), .B(new_n15908), .C(new_n15905), .Y(new_n15909));
  O2A1O1Ixp33_ASAP7_75t_L   g15653(.A1(new_n15876), .A2(new_n15881), .B(new_n15894), .C(new_n15909), .Y(new_n15910));
  A2O1A1Ixp33_ASAP7_75t_L   g15654(.A1(new_n15332), .A2(new_n15329), .B(new_n15338), .C(new_n15614), .Y(new_n15911));
  A2O1A1Ixp33_ASAP7_75t_L   g15655(.A1(new_n15895), .A2(new_n15878), .B(new_n15879), .C(new_n15875), .Y(new_n15912));
  O2A1O1Ixp33_ASAP7_75t_L   g15656(.A1(new_n15879), .A2(new_n15629), .B(new_n15912), .C(new_n15881), .Y(new_n15913));
  INVx1_ASAP7_75t_L         g15657(.A(new_n15894), .Y(new_n15914));
  INVx1_ASAP7_75t_L         g15658(.A(new_n15908), .Y(new_n15915));
  NAND3xp33_ASAP7_75t_L     g15659(.A(new_n15913), .B(new_n15915), .C(new_n15893), .Y(new_n15916));
  O2A1O1Ixp33_ASAP7_75t_L   g15660(.A1(new_n15913), .A2(new_n15914), .B(new_n15916), .C(new_n15620), .Y(new_n15917));
  INVx1_ASAP7_75t_L         g15661(.A(new_n15620), .Y(new_n15918));
  AOI21xp33_ASAP7_75t_L     g15662(.A1(new_n15893), .A2(new_n15915), .B(new_n15913), .Y(new_n15919));
  NOR3xp33_ASAP7_75t_L      g15663(.A(new_n15919), .B(new_n15909), .C(new_n15918), .Y(new_n15920));
  NOR2xp33_ASAP7_75t_L      g15664(.A(new_n15920), .B(new_n15917), .Y(new_n15921));
  O2A1O1Ixp33_ASAP7_75t_L   g15665(.A1(new_n15340), .A2(new_n15615), .B(new_n15911), .C(new_n15921), .Y(new_n15922));
  A2O1A1Ixp33_ASAP7_75t_L   g15666(.A1(new_n15602), .A2(new_n15608), .B(new_n15340), .C(new_n15911), .Y(new_n15923));
  NOR2xp33_ASAP7_75t_L      g15667(.A(new_n15920), .B(new_n15923), .Y(new_n15924));
  O2A1O1Ixp33_ASAP7_75t_L   g15668(.A1(new_n15910), .A2(new_n15620), .B(new_n15924), .C(new_n15922), .Y(\f[73] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15669(.A1(new_n15908), .A2(new_n15892), .B(new_n15905), .C(new_n15891), .Y(new_n15926));
  NOR2xp33_ASAP7_75t_L      g15670(.A(new_n12956), .B(new_n712), .Y(new_n15927));
  A2O1A1Ixp33_ASAP7_75t_L   g15671(.A1(new_n12986), .A2(new_n718), .B(new_n15927), .C(\a[11] ), .Y(new_n15928));
  A2O1A1O1Ixp25_ASAP7_75t_L g15672(.A1(new_n718), .A2(new_n14172), .B(new_n713), .C(\b[63] ), .D(new_n637), .Y(new_n15929));
  A2O1A1O1Ixp25_ASAP7_75t_L g15673(.A1(new_n12986), .A2(new_n718), .B(new_n15927), .C(new_n15928), .D(new_n15929), .Y(new_n15930));
  O2A1O1Ixp33_ASAP7_75t_L   g15674(.A1(new_n15897), .A2(new_n15880), .B(new_n15895), .C(new_n15930), .Y(new_n15931));
  O2A1O1Ixp33_ASAP7_75t_L   g15675(.A1(new_n15626), .A2(new_n15627), .B(new_n15630), .C(new_n15880), .Y(new_n15932));
  A2O1A1Ixp33_ASAP7_75t_L   g15676(.A1(new_n15878), .A2(new_n15628), .B(new_n15932), .C(new_n15930), .Y(new_n15933));
  A2O1A1Ixp33_ASAP7_75t_L   g15677(.A1(new_n15867), .A2(new_n15866), .B(new_n15901), .C(new_n15902), .Y(new_n15934));
  NAND2xp33_ASAP7_75t_L     g15678(.A(\b[61] ), .B(new_n885), .Y(new_n15935));
  OAI221xp5_ASAP7_75t_L     g15679(.A1(new_n869), .A2(new_n12603), .B1(new_n11626), .B2(new_n980), .C(new_n15935), .Y(new_n15936));
  AOI21xp33_ASAP7_75t_L     g15680(.A1(new_n13559), .A2(new_n873), .B(new_n15936), .Y(new_n15937));
  NAND2xp33_ASAP7_75t_L     g15681(.A(\a[14] ), .B(new_n15937), .Y(new_n15938));
  A2O1A1Ixp33_ASAP7_75t_L   g15682(.A1(new_n13559), .A2(new_n873), .B(new_n15936), .C(new_n867), .Y(new_n15939));
  AND2x2_ASAP7_75t_L        g15683(.A(new_n15939), .B(new_n15938), .Y(new_n15940));
  INVx1_ASAP7_75t_L         g15684(.A(new_n15940), .Y(new_n15941));
  A2O1A1Ixp33_ASAP7_75t_L   g15685(.A1(new_n15934), .A2(new_n15862), .B(new_n15901), .C(new_n15941), .Y(new_n15942));
  O2A1O1Ixp33_ASAP7_75t_L   g15686(.A1(new_n15869), .A2(new_n15873), .B(new_n15862), .C(new_n15901), .Y(new_n15943));
  NAND2xp33_ASAP7_75t_L     g15687(.A(new_n15940), .B(new_n15943), .Y(new_n15944));
  NAND2xp33_ASAP7_75t_L     g15688(.A(new_n15942), .B(new_n15944), .Y(new_n15945));
  INVx1_ASAP7_75t_L         g15689(.A(new_n15858), .Y(new_n15946));
  INVx1_ASAP7_75t_L         g15690(.A(new_n15859), .Y(new_n15947));
  NOR2xp33_ASAP7_75t_L      g15691(.A(new_n11591), .B(new_n1284), .Y(new_n15948));
  AOI221xp5_ASAP7_75t_L     g15692(.A1(\b[57] ), .A2(new_n1290), .B1(\b[58] ), .B2(new_n1204), .C(new_n15948), .Y(new_n15949));
  O2A1O1Ixp33_ASAP7_75t_L   g15693(.A1(new_n1210), .A2(new_n11597), .B(new_n15949), .C(new_n1206), .Y(new_n15950));
  INVx1_ASAP7_75t_L         g15694(.A(new_n15950), .Y(new_n15951));
  O2A1O1Ixp33_ASAP7_75t_L   g15695(.A1(new_n1210), .A2(new_n11597), .B(new_n15949), .C(\a[17] ), .Y(new_n15952));
  AOI21xp33_ASAP7_75t_L     g15696(.A1(new_n15951), .A2(\a[17] ), .B(new_n15952), .Y(new_n15953));
  NAND3xp33_ASAP7_75t_L     g15697(.A(new_n15947), .B(new_n15946), .C(new_n15953), .Y(new_n15954));
  INVx1_ASAP7_75t_L         g15698(.A(new_n15954), .Y(new_n15955));
  O2A1O1Ixp33_ASAP7_75t_L   g15699(.A1(new_n15855), .A2(new_n15856), .B(new_n15947), .C(new_n15953), .Y(new_n15956));
  NOR2xp33_ASAP7_75t_L      g15700(.A(new_n15956), .B(new_n15955), .Y(new_n15957));
  NAND2xp33_ASAP7_75t_L     g15701(.A(\b[49] ), .B(new_n2421), .Y(new_n15958));
  OAI221xp5_ASAP7_75t_L     g15702(.A1(new_n2415), .A2(new_n8755), .B1(new_n7860), .B2(new_n2572), .C(new_n15958), .Y(new_n15959));
  AOI21xp33_ASAP7_75t_L     g15703(.A1(new_n8763), .A2(new_n2417), .B(new_n15959), .Y(new_n15960));
  NAND2xp33_ASAP7_75t_L     g15704(.A(\a[26] ), .B(new_n15960), .Y(new_n15961));
  A2O1A1Ixp33_ASAP7_75t_L   g15705(.A1(new_n8763), .A2(new_n2417), .B(new_n15959), .C(new_n2413), .Y(new_n15962));
  AND2x2_ASAP7_75t_L        g15706(.A(new_n15962), .B(new_n15961), .Y(new_n15963));
  INVx1_ASAP7_75t_L         g15707(.A(new_n15963), .Y(new_n15964));
  A2O1A1Ixp33_ASAP7_75t_L   g15708(.A1(new_n15813), .A2(new_n15818), .B(new_n15811), .C(new_n15964), .Y(new_n15965));
  O2A1O1Ixp33_ASAP7_75t_L   g15709(.A1(new_n15841), .A2(new_n15840), .B(new_n15818), .C(new_n15811), .Y(new_n15966));
  NAND2xp33_ASAP7_75t_L     g15710(.A(new_n15963), .B(new_n15966), .Y(new_n15967));
  NAND2xp33_ASAP7_75t_L     g15711(.A(new_n15965), .B(new_n15967), .Y(new_n15968));
  NOR2xp33_ASAP7_75t_L      g15712(.A(new_n7552), .B(new_n2930), .Y(new_n15969));
  AOI221xp5_ASAP7_75t_L     g15713(.A1(\b[45] ), .A2(new_n3129), .B1(\b[46] ), .B2(new_n2936), .C(new_n15969), .Y(new_n15970));
  O2A1O1Ixp33_ASAP7_75t_L   g15714(.A1(new_n2940), .A2(new_n7560), .B(new_n15970), .C(new_n2928), .Y(new_n15971));
  O2A1O1Ixp33_ASAP7_75t_L   g15715(.A1(new_n2940), .A2(new_n7560), .B(new_n15970), .C(\a[29] ), .Y(new_n15972));
  INVx1_ASAP7_75t_L         g15716(.A(new_n15972), .Y(new_n15973));
  A2O1A1O1Ixp25_ASAP7_75t_L g15717(.A1(new_n15783), .A2(new_n15647), .B(new_n15788), .C(new_n15800), .D(new_n15799), .Y(new_n15974));
  OA211x2_ASAP7_75t_L       g15718(.A1(new_n15971), .A2(new_n2928), .B(new_n15974), .C(new_n15973), .Y(new_n15975));
  O2A1O1Ixp33_ASAP7_75t_L   g15719(.A1(new_n2928), .A2(new_n15971), .B(new_n15973), .C(new_n15974), .Y(new_n15976));
  NOR2xp33_ASAP7_75t_L      g15720(.A(new_n15976), .B(new_n15975), .Y(new_n15977));
  NAND2xp33_ASAP7_75t_L     g15721(.A(\b[43] ), .B(new_n3499), .Y(new_n15978));
  OAI221xp5_ASAP7_75t_L     g15722(.A1(new_n3510), .A2(new_n6944), .B1(new_n6378), .B2(new_n3703), .C(new_n15978), .Y(new_n15979));
  AOI21xp33_ASAP7_75t_L     g15723(.A1(new_n7824), .A2(new_n3505), .B(new_n15979), .Y(new_n15980));
  NAND2xp33_ASAP7_75t_L     g15724(.A(\a[32] ), .B(new_n15980), .Y(new_n15981));
  A2O1A1Ixp33_ASAP7_75t_L   g15725(.A1(new_n7824), .A2(new_n3505), .B(new_n15979), .C(new_n3493), .Y(new_n15982));
  NAND2xp33_ASAP7_75t_L     g15726(.A(new_n15982), .B(new_n15981), .Y(new_n15983));
  INVx1_ASAP7_75t_L         g15727(.A(new_n15983), .Y(new_n15984));
  A2O1A1O1Ixp25_ASAP7_75t_L g15728(.A1(new_n15785), .A2(new_n15787), .B(new_n15646), .C(new_n15781), .D(new_n15984), .Y(new_n15985));
  INVx1_ASAP7_75t_L         g15729(.A(new_n15985), .Y(new_n15986));
  O2A1O1Ixp33_ASAP7_75t_L   g15730(.A1(new_n15780), .A2(new_n15782), .B(new_n15647), .C(new_n15786), .Y(new_n15987));
  NAND2xp33_ASAP7_75t_L     g15731(.A(new_n15984), .B(new_n15987), .Y(new_n15988));
  NAND2xp33_ASAP7_75t_L     g15732(.A(new_n15988), .B(new_n15986), .Y(new_n15989));
  NAND2xp33_ASAP7_75t_L     g15733(.A(new_n15777), .B(new_n15784), .Y(new_n15990));
  O2A1O1Ixp33_ASAP7_75t_L   g15734(.A1(new_n15775), .A2(new_n15774), .B(new_n15990), .C(new_n15770), .Y(new_n15991));
  NAND2xp33_ASAP7_75t_L     g15735(.A(new_n15412), .B(new_n15413), .Y(new_n15992));
  A2O1A1Ixp33_ASAP7_75t_L   g15736(.A1(new_n15513), .A2(new_n15992), .B(new_n15510), .C(new_n15764), .Y(new_n15993));
  A2O1A1Ixp33_ASAP7_75t_L   g15737(.A1(new_n15718), .A2(new_n15470), .B(new_n15716), .C(new_n15730), .Y(new_n15994));
  NOR2xp33_ASAP7_75t_L      g15738(.A(new_n2377), .B(new_n10065), .Y(new_n15995));
  AOI221xp5_ASAP7_75t_L     g15739(.A1(new_n8175), .A2(\b[26] ), .B1(new_n8484), .B2(\b[24] ), .C(new_n15995), .Y(new_n15996));
  INVx1_ASAP7_75t_L         g15740(.A(new_n15996), .Y(new_n15997));
  A2O1A1Ixp33_ASAP7_75t_L   g15741(.A1(new_n2709), .A2(new_n8490), .B(new_n15997), .C(\a[50] ), .Y(new_n15998));
  O2A1O1Ixp33_ASAP7_75t_L   g15742(.A1(new_n8176), .A2(new_n2708), .B(new_n15996), .C(\a[50] ), .Y(new_n15999));
  A2O1A1O1Ixp25_ASAP7_75t_L g15743(.A1(new_n15711), .A2(\a[53] ), .B(new_n15712), .C(new_n15707), .D(new_n15706), .Y(new_n16000));
  NOR2xp33_ASAP7_75t_L      g15744(.A(new_n2045), .B(new_n10400), .Y(new_n16001));
  AOI221xp5_ASAP7_75t_L     g15745(.A1(new_n9102), .A2(\b[23] ), .B1(new_n10398), .B2(\b[21] ), .C(new_n16001), .Y(new_n16002));
  O2A1O1Ixp33_ASAP7_75t_L   g15746(.A1(new_n9104), .A2(new_n2194), .B(new_n16002), .C(new_n9099), .Y(new_n16003));
  INVx1_ASAP7_75t_L         g15747(.A(new_n16003), .Y(new_n16004));
  O2A1O1Ixp33_ASAP7_75t_L   g15748(.A1(new_n9104), .A2(new_n2194), .B(new_n16002), .C(\a[53] ), .Y(new_n16005));
  AOI21xp33_ASAP7_75t_L     g15749(.A1(new_n16004), .A2(\a[53] ), .B(new_n16005), .Y(new_n16006));
  A2O1A1Ixp33_ASAP7_75t_L   g15750(.A1(\a[59] ), .A2(new_n15442), .B(new_n15443), .C(new_n15438), .Y(new_n16007));
  A2O1A1Ixp33_ASAP7_75t_L   g15751(.A1(new_n15446), .A2(new_n16007), .B(new_n15688), .C(new_n15700), .Y(new_n16008));
  INVx1_ASAP7_75t_L         g15752(.A(new_n16008), .Y(new_n16009));
  OAI22xp33_ASAP7_75t_L     g15753(.A1(new_n12320), .A2(new_n833), .B1(new_n936), .B2(new_n12318), .Y(new_n16010));
  AOI221xp5_ASAP7_75t_L     g15754(.A1(new_n11995), .A2(\b[14] ), .B1(new_n11997), .B2(new_n971), .C(new_n16010), .Y(new_n16011));
  XNOR2x2_ASAP7_75t_L       g15755(.A(new_n11987), .B(new_n16011), .Y(new_n16012));
  INVx1_ASAP7_75t_L         g15756(.A(new_n16012), .Y(new_n16013));
  O2A1O1Ixp33_ASAP7_75t_L   g15757(.A1(new_n15668), .A2(new_n15658), .B(new_n15656), .C(new_n15671), .Y(new_n16014));
  NOR2xp33_ASAP7_75t_L      g15758(.A(new_n680), .B(new_n13030), .Y(new_n16015));
  INVx1_ASAP7_75t_L         g15759(.A(new_n16015), .Y(new_n16016));
  O2A1O1Ixp33_ASAP7_75t_L   g15760(.A1(new_n12672), .A2(new_n748), .B(new_n16016), .C(new_n15657), .Y(new_n16017));
  O2A1O1Ixp33_ASAP7_75t_L   g15761(.A1(new_n12672), .A2(new_n748), .B(new_n16016), .C(new_n15656), .Y(new_n16018));
  INVx1_ASAP7_75t_L         g15762(.A(new_n16018), .Y(new_n16019));
  O2A1O1Ixp33_ASAP7_75t_L   g15763(.A1(new_n16017), .A2(new_n15657), .B(new_n16019), .C(new_n16014), .Y(new_n16020));
  INVx1_ASAP7_75t_L         g15764(.A(new_n16014), .Y(new_n16021));
  O2A1O1Ixp33_ASAP7_75t_L   g15765(.A1(new_n16017), .A2(new_n15657), .B(new_n16019), .C(new_n16021), .Y(new_n16022));
  INVx1_ASAP7_75t_L         g15766(.A(new_n16022), .Y(new_n16023));
  O2A1O1Ixp33_ASAP7_75t_L   g15767(.A1(new_n16014), .A2(new_n16020), .B(new_n16023), .C(new_n16012), .Y(new_n16024));
  INVx1_ASAP7_75t_L         g15768(.A(new_n16024), .Y(new_n16025));
  O2A1O1Ixp33_ASAP7_75t_L   g15769(.A1(new_n16014), .A2(new_n16020), .B(new_n16023), .C(new_n16013), .Y(new_n16026));
  NOR2xp33_ASAP7_75t_L      g15770(.A(new_n1043), .B(new_n11354), .Y(new_n16027));
  AOI221xp5_ASAP7_75t_L     g15771(.A1(\b[17] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[16] ), .C(new_n16027), .Y(new_n16028));
  O2A1O1Ixp33_ASAP7_75t_L   g15772(.A1(new_n11053), .A2(new_n1356), .B(new_n16028), .C(new_n11048), .Y(new_n16029));
  O2A1O1Ixp33_ASAP7_75t_L   g15773(.A1(new_n11053), .A2(new_n1356), .B(new_n16028), .C(\a[59] ), .Y(new_n16030));
  INVx1_ASAP7_75t_L         g15774(.A(new_n16030), .Y(new_n16031));
  OAI21xp33_ASAP7_75t_L     g15775(.A1(new_n11048), .A2(new_n16029), .B(new_n16031), .Y(new_n16032));
  A2O1A1Ixp33_ASAP7_75t_L   g15776(.A1(new_n16025), .A2(new_n16013), .B(new_n16026), .C(new_n16032), .Y(new_n16033));
  A2O1A1Ixp33_ASAP7_75t_L   g15777(.A1(new_n16025), .A2(new_n16013), .B(new_n16026), .C(new_n16033), .Y(new_n16034));
  INVx1_ASAP7_75t_L         g15778(.A(new_n16034), .Y(new_n16035));
  INVx1_ASAP7_75t_L         g15779(.A(new_n16029), .Y(new_n16036));
  A2O1A1Ixp33_ASAP7_75t_L   g15780(.A1(new_n16036), .A2(\a[59] ), .B(new_n16030), .C(new_n16033), .Y(new_n16037));
  INVx1_ASAP7_75t_L         g15781(.A(new_n16037), .Y(new_n16038));
  A2O1A1O1Ixp25_ASAP7_75t_L g15782(.A1(new_n15683), .A2(\a[59] ), .B(new_n15684), .C(new_n15679), .D(new_n15676), .Y(new_n16039));
  INVx1_ASAP7_75t_L         g15783(.A(new_n16039), .Y(new_n16040));
  NOR3xp33_ASAP7_75t_L      g15784(.A(new_n16035), .B(new_n16038), .C(new_n16040), .Y(new_n16041));
  AOI21xp33_ASAP7_75t_L     g15785(.A1(new_n16037), .A2(new_n16034), .B(new_n16039), .Y(new_n16042));
  NOR2xp33_ASAP7_75t_L      g15786(.A(new_n16042), .B(new_n16041), .Y(new_n16043));
  NOR2xp33_ASAP7_75t_L      g15787(.A(new_n1599), .B(new_n10388), .Y(new_n16044));
  AOI221xp5_ASAP7_75t_L     g15788(.A1(new_n10086), .A2(\b[20] ), .B1(new_n11361), .B2(\b[18] ), .C(new_n16044), .Y(new_n16045));
  O2A1O1Ixp33_ASAP7_75t_L   g15789(.A1(new_n10088), .A2(new_n1754), .B(new_n16045), .C(new_n10083), .Y(new_n16046));
  INVx1_ASAP7_75t_L         g15790(.A(new_n16046), .Y(new_n16047));
  O2A1O1Ixp33_ASAP7_75t_L   g15791(.A1(new_n10088), .A2(new_n1754), .B(new_n16045), .C(\a[56] ), .Y(new_n16048));
  AOI211xp5_ASAP7_75t_L     g15792(.A1(new_n16047), .A2(\a[56] ), .B(new_n16048), .C(new_n16043), .Y(new_n16049));
  AOI21xp33_ASAP7_75t_L     g15793(.A1(new_n16047), .A2(\a[56] ), .B(new_n16048), .Y(new_n16050));
  NOR3xp33_ASAP7_75t_L      g15794(.A(new_n16041), .B(new_n16042), .C(new_n16050), .Y(new_n16051));
  NOR3xp33_ASAP7_75t_L      g15795(.A(new_n16009), .B(new_n16049), .C(new_n16051), .Y(new_n16052));
  NOR2xp33_ASAP7_75t_L      g15796(.A(new_n16051), .B(new_n16049), .Y(new_n16053));
  NAND2xp33_ASAP7_75t_L     g15797(.A(new_n16053), .B(new_n16009), .Y(new_n16054));
  O2A1O1Ixp33_ASAP7_75t_L   g15798(.A1(new_n16009), .A2(new_n16052), .B(new_n16054), .C(new_n16006), .Y(new_n16055));
  NAND2xp33_ASAP7_75t_L     g15799(.A(new_n16006), .B(new_n16054), .Y(new_n16056));
  O2A1O1Ixp33_ASAP7_75t_L   g15800(.A1(new_n16049), .A2(new_n16051), .B(new_n16008), .C(new_n16056), .Y(new_n16057));
  OR3x1_ASAP7_75t_L         g15801(.A(new_n16057), .B(new_n16000), .C(new_n16055), .Y(new_n16058));
  INVx1_ASAP7_75t_L         g15802(.A(new_n16058), .Y(new_n16059));
  INVx1_ASAP7_75t_L         g15803(.A(new_n16000), .Y(new_n16060));
  O2A1O1Ixp33_ASAP7_75t_L   g15804(.A1(new_n15688), .A2(new_n15690), .B(new_n15700), .C(new_n16053), .Y(new_n16061));
  A2O1A1Ixp33_ASAP7_75t_L   g15805(.A1(new_n15700), .A2(new_n15693), .B(new_n16052), .C(new_n16054), .Y(new_n16062));
  A2O1A1Ixp33_ASAP7_75t_L   g15806(.A1(new_n16004), .A2(\a[53] ), .B(new_n16005), .C(new_n16062), .Y(new_n16063));
  O2A1O1Ixp33_ASAP7_75t_L   g15807(.A1(new_n16056), .A2(new_n16061), .B(new_n16063), .C(new_n16060), .Y(new_n16064));
  NOR2xp33_ASAP7_75t_L      g15808(.A(new_n16064), .B(new_n16059), .Y(new_n16065));
  A2O1A1Ixp33_ASAP7_75t_L   g15809(.A1(new_n15998), .A2(\a[50] ), .B(new_n15999), .C(new_n16065), .Y(new_n16066));
  AO21x2_ASAP7_75t_L        g15810(.A1(\a[50] ), .A2(new_n15998), .B(new_n15999), .Y(new_n16067));
  INVx1_ASAP7_75t_L         g15811(.A(new_n16064), .Y(new_n16068));
  AO21x2_ASAP7_75t_L        g15812(.A1(new_n16058), .A2(new_n16068), .B(new_n16067), .Y(new_n16069));
  NAND2xp33_ASAP7_75t_L     g15813(.A(new_n16069), .B(new_n16066), .Y(new_n16070));
  XOR2x2_ASAP7_75t_L        g15814(.A(new_n15994), .B(new_n16070), .Y(new_n16071));
  NOR2xp33_ASAP7_75t_L      g15815(.A(new_n3079), .B(new_n7312), .Y(new_n16072));
  AOI221xp5_ASAP7_75t_L     g15816(.A1(\b[27] ), .A2(new_n7609), .B1(\b[29] ), .B2(new_n7334), .C(new_n16072), .Y(new_n16073));
  O2A1O1Ixp33_ASAP7_75t_L   g15817(.A1(new_n7321), .A2(new_n3104), .B(new_n16073), .C(new_n7316), .Y(new_n16074));
  O2A1O1Ixp33_ASAP7_75t_L   g15818(.A1(new_n7321), .A2(new_n3104), .B(new_n16073), .C(\a[47] ), .Y(new_n16075));
  INVx1_ASAP7_75t_L         g15819(.A(new_n16075), .Y(new_n16076));
  O2A1O1Ixp33_ASAP7_75t_L   g15820(.A1(new_n16074), .A2(new_n7316), .B(new_n16076), .C(new_n16071), .Y(new_n16077));
  INVx1_ASAP7_75t_L         g15821(.A(new_n16074), .Y(new_n16078));
  A2O1A1Ixp33_ASAP7_75t_L   g15822(.A1(\a[47] ), .A2(new_n16078), .B(new_n16075), .C(new_n16071), .Y(new_n16079));
  OA21x2_ASAP7_75t_L        g15823(.A1(new_n16071), .A2(new_n16077), .B(new_n16079), .Y(new_n16080));
  A2O1A1O1Ixp25_ASAP7_75t_L g15824(.A1(new_n15730), .A2(new_n15729), .B(new_n15735), .C(new_n15736), .D(new_n15744), .Y(new_n16081));
  NAND2xp33_ASAP7_75t_L     g15825(.A(new_n16081), .B(new_n16080), .Y(new_n16082));
  O2A1O1Ixp33_ASAP7_75t_L   g15826(.A1(new_n16071), .A2(new_n16077), .B(new_n16079), .C(new_n16081), .Y(new_n16083));
  INVx1_ASAP7_75t_L         g15827(.A(new_n16083), .Y(new_n16084));
  NOR2xp33_ASAP7_75t_L      g15828(.A(new_n3456), .B(new_n6741), .Y(new_n16085));
  AOI221xp5_ASAP7_75t_L     g15829(.A1(\b[32] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[31] ), .C(new_n16085), .Y(new_n16086));
  O2A1O1Ixp33_ASAP7_75t_L   g15830(.A1(new_n6443), .A2(new_n3897), .B(new_n16086), .C(new_n6439), .Y(new_n16087));
  INVx1_ASAP7_75t_L         g15831(.A(new_n16087), .Y(new_n16088));
  O2A1O1Ixp33_ASAP7_75t_L   g15832(.A1(new_n6443), .A2(new_n3897), .B(new_n16086), .C(\a[44] ), .Y(new_n16089));
  AO221x2_ASAP7_75t_L       g15833(.A1(new_n16088), .A2(\a[44] ), .B1(new_n16082), .B2(new_n16084), .C(new_n16089), .Y(new_n16090));
  AND2x2_ASAP7_75t_L        g15834(.A(new_n16084), .B(new_n16082), .Y(new_n16091));
  A2O1A1Ixp33_ASAP7_75t_L   g15835(.A1(\a[44] ), .A2(new_n16088), .B(new_n16089), .C(new_n16091), .Y(new_n16092));
  NAND2xp33_ASAP7_75t_L     g15836(.A(new_n16090), .B(new_n16092), .Y(new_n16093));
  O2A1O1Ixp33_ASAP7_75t_L   g15837(.A1(new_n15748), .A2(new_n15750), .B(new_n15762), .C(new_n16093), .Y(new_n16094));
  AOI211xp5_ASAP7_75t_L     g15838(.A1(new_n16092), .A2(new_n16090), .B(new_n15752), .C(new_n15763), .Y(new_n16095));
  NOR2xp33_ASAP7_75t_L      g15839(.A(new_n16095), .B(new_n16094), .Y(new_n16096));
  NOR2xp33_ASAP7_75t_L      g15840(.A(new_n4581), .B(new_n5641), .Y(new_n16097));
  AOI221xp5_ASAP7_75t_L     g15841(.A1(\b[33] ), .A2(new_n5920), .B1(\b[34] ), .B2(new_n5623), .C(new_n16097), .Y(new_n16098));
  O2A1O1Ixp33_ASAP7_75t_L   g15842(.A1(new_n5630), .A2(new_n4589), .B(new_n16098), .C(new_n5626), .Y(new_n16099));
  INVx1_ASAP7_75t_L         g15843(.A(new_n16099), .Y(new_n16100));
  O2A1O1Ixp33_ASAP7_75t_L   g15844(.A1(new_n5630), .A2(new_n4589), .B(new_n16098), .C(\a[41] ), .Y(new_n16101));
  A2O1A1Ixp33_ASAP7_75t_L   g15845(.A1(\a[41] ), .A2(new_n16100), .B(new_n16101), .C(new_n16096), .Y(new_n16102));
  INVx1_ASAP7_75t_L         g15846(.A(new_n16101), .Y(new_n16103));
  O2A1O1Ixp33_ASAP7_75t_L   g15847(.A1(new_n16099), .A2(new_n5626), .B(new_n16103), .C(new_n16096), .Y(new_n16104));
  AOI21xp33_ASAP7_75t_L     g15848(.A1(new_n16102), .A2(new_n16096), .B(new_n16104), .Y(new_n16105));
  NAND3xp33_ASAP7_75t_L     g15849(.A(new_n16105), .B(new_n15766), .C(new_n15993), .Y(new_n16106));
  NAND2xp33_ASAP7_75t_L     g15850(.A(new_n15993), .B(new_n15766), .Y(new_n16107));
  A2O1A1Ixp33_ASAP7_75t_L   g15851(.A1(new_n16102), .A2(new_n16096), .B(new_n16104), .C(new_n16107), .Y(new_n16108));
  AND2x2_ASAP7_75t_L        g15852(.A(new_n16108), .B(new_n16106), .Y(new_n16109));
  NOR2xp33_ASAP7_75t_L      g15853(.A(new_n5311), .B(new_n4908), .Y(new_n16110));
  AOI221xp5_ASAP7_75t_L     g15854(.A1(\b[36] ), .A2(new_n5139), .B1(\b[37] ), .B2(new_n4916), .C(new_n16110), .Y(new_n16111));
  O2A1O1Ixp33_ASAP7_75t_L   g15855(.A1(new_n4911), .A2(new_n5318), .B(new_n16111), .C(new_n4906), .Y(new_n16112));
  INVx1_ASAP7_75t_L         g15856(.A(new_n16112), .Y(new_n16113));
  O2A1O1Ixp33_ASAP7_75t_L   g15857(.A1(new_n4911), .A2(new_n5318), .B(new_n16111), .C(\a[38] ), .Y(new_n16114));
  AOI21xp33_ASAP7_75t_L     g15858(.A1(new_n16113), .A2(\a[38] ), .B(new_n16114), .Y(new_n16115));
  XNOR2x2_ASAP7_75t_L       g15859(.A(new_n16115), .B(new_n16109), .Y(new_n16116));
  XNOR2x2_ASAP7_75t_L       g15860(.A(new_n15991), .B(new_n16116), .Y(new_n16117));
  INVx1_ASAP7_75t_L         g15861(.A(new_n16117), .Y(new_n16118));
  NOR2xp33_ASAP7_75t_L      g15862(.A(new_n6110), .B(new_n4147), .Y(new_n16119));
  AOI221xp5_ASAP7_75t_L     g15863(.A1(\b[39] ), .A2(new_n4402), .B1(\b[40] ), .B2(new_n4155), .C(new_n16119), .Y(new_n16120));
  O2A1O1Ixp33_ASAP7_75t_L   g15864(.A1(new_n4150), .A2(new_n6117), .B(new_n16120), .C(new_n4145), .Y(new_n16121));
  INVx1_ASAP7_75t_L         g15865(.A(new_n16121), .Y(new_n16122));
  O2A1O1Ixp33_ASAP7_75t_L   g15866(.A1(new_n4150), .A2(new_n6117), .B(new_n16120), .C(\a[35] ), .Y(new_n16123));
  A2O1A1Ixp33_ASAP7_75t_L   g15867(.A1(new_n16122), .A2(\a[35] ), .B(new_n16123), .C(new_n16117), .Y(new_n16124));
  INVx1_ASAP7_75t_L         g15868(.A(new_n16124), .Y(new_n16125));
  INVx1_ASAP7_75t_L         g15869(.A(new_n16123), .Y(new_n16126));
  O2A1O1Ixp33_ASAP7_75t_L   g15870(.A1(new_n4145), .A2(new_n16121), .B(new_n16126), .C(new_n16117), .Y(new_n16127));
  INVx1_ASAP7_75t_L         g15871(.A(new_n16127), .Y(new_n16128));
  O2A1O1Ixp33_ASAP7_75t_L   g15872(.A1(new_n16118), .A2(new_n16125), .B(new_n16128), .C(new_n15989), .Y(new_n16129));
  A2O1A1Ixp33_ASAP7_75t_L   g15873(.A1(new_n16117), .A2(new_n16124), .B(new_n16127), .C(new_n15989), .Y(new_n16130));
  OAI21xp33_ASAP7_75t_L     g15874(.A1(new_n15989), .A2(new_n16129), .B(new_n16130), .Y(new_n16131));
  NAND2xp33_ASAP7_75t_L     g15875(.A(new_n16131), .B(new_n15977), .Y(new_n16132));
  OA21x2_ASAP7_75t_L        g15876(.A1(new_n15989), .A2(new_n16129), .B(new_n16130), .Y(new_n16133));
  O2A1O1Ixp33_ASAP7_75t_L   g15877(.A1(new_n15975), .A2(new_n15976), .B(new_n16133), .C(new_n15968), .Y(new_n16134));
  OAI21xp33_ASAP7_75t_L     g15878(.A1(new_n15975), .A2(new_n15976), .B(new_n16133), .Y(new_n16135));
  NAND3xp33_ASAP7_75t_L     g15879(.A(new_n15968), .B(new_n16132), .C(new_n16135), .Y(new_n16136));
  A2O1A1Ixp33_ASAP7_75t_L   g15880(.A1(new_n16134), .A2(new_n16132), .B(new_n15968), .C(new_n16136), .Y(new_n16137));
  NOR2xp33_ASAP7_75t_L      g15881(.A(new_n9355), .B(new_n1962), .Y(new_n16138));
  AOI221xp5_ASAP7_75t_L     g15882(.A1(new_n1955), .A2(\b[53] ), .B1(new_n2093), .B2(\b[51] ), .C(new_n16138), .Y(new_n16139));
  INVx1_ASAP7_75t_L         g15883(.A(new_n16139), .Y(new_n16140));
  A2O1A1Ixp33_ASAP7_75t_L   g15884(.A1(new_n1951), .A2(new_n1953), .B(new_n1793), .C(new_n16139), .Y(new_n16141));
  A2O1A1O1Ixp25_ASAP7_75t_L g15885(.A1(new_n9689), .A2(new_n9686), .B(new_n16140), .C(new_n16141), .D(new_n1952), .Y(new_n16142));
  O2A1O1Ixp33_ASAP7_75t_L   g15886(.A1(new_n1956), .A2(new_n9691), .B(new_n16139), .C(\a[23] ), .Y(new_n16143));
  A2O1A1Ixp33_ASAP7_75t_L   g15887(.A1(new_n15824), .A2(\a[26] ), .B(new_n15825), .C(new_n15832), .Y(new_n16144));
  NOR2xp33_ASAP7_75t_L      g15888(.A(new_n16142), .B(new_n16143), .Y(new_n16145));
  A2O1A1O1Ixp25_ASAP7_75t_L g15889(.A1(new_n15830), .A2(new_n16144), .B(new_n15820), .C(new_n15834), .D(new_n16145), .Y(new_n16146));
  INVx1_ASAP7_75t_L         g15890(.A(new_n16146), .Y(new_n16147));
  INVx1_ASAP7_75t_L         g15891(.A(new_n16145), .Y(new_n16148));
  A2O1A1O1Ixp25_ASAP7_75t_L g15892(.A1(new_n15830), .A2(new_n15826), .B(new_n15820), .C(new_n15834), .D(new_n16148), .Y(new_n16149));
  O2A1O1Ixp33_ASAP7_75t_L   g15893(.A1(new_n16142), .A2(new_n16143), .B(new_n16147), .C(new_n16149), .Y(new_n16150));
  NAND2xp33_ASAP7_75t_L     g15894(.A(new_n16137), .B(new_n16150), .Y(new_n16151));
  NAND4xp25_ASAP7_75t_L     g15895(.A(new_n16135), .B(new_n16132), .C(new_n15965), .D(new_n15967), .Y(new_n16152));
  AOI21xp33_ASAP7_75t_L     g15896(.A1(new_n16135), .A2(new_n16132), .B(new_n15968), .Y(new_n16153));
  AOI31xp33_ASAP7_75t_L     g15897(.A1(new_n16135), .A2(new_n16132), .A3(new_n16152), .B(new_n16153), .Y(new_n16154));
  A2O1A1Ixp33_ASAP7_75t_L   g15898(.A1(new_n16148), .A2(new_n16147), .B(new_n16149), .C(new_n16154), .Y(new_n16155));
  NAND2xp33_ASAP7_75t_L     g15899(.A(new_n16155), .B(new_n16151), .Y(new_n16156));
  A2O1A1Ixp33_ASAP7_75t_L   g15900(.A1(new_n15397), .A2(new_n15396), .B(new_n15398), .C(new_n15568), .Y(new_n16157));
  A2O1A1Ixp33_ASAP7_75t_L   g15901(.A1(new_n16157), .A2(new_n15397), .B(new_n15827), .C(new_n16144), .Y(new_n16158));
  A2O1A1Ixp33_ASAP7_75t_L   g15902(.A1(new_n15818), .A2(new_n15845), .B(new_n15819), .C(new_n16158), .Y(new_n16159));
  A2O1A1Ixp33_ASAP7_75t_L   g15903(.A1(new_n15845), .A2(new_n15818), .B(new_n15819), .C(new_n16159), .Y(new_n16160));
  A2O1A1Ixp33_ASAP7_75t_L   g15904(.A1(new_n16160), .A2(new_n15837), .B(new_n15640), .C(new_n15639), .Y(new_n16161));
  O2A1O1Ixp33_ASAP7_75t_L   g15905(.A1(new_n15842), .A2(new_n15844), .B(new_n15843), .C(new_n16158), .Y(new_n16162));
  A2O1A1O1Ixp25_ASAP7_75t_L g15906(.A1(new_n15834), .A2(new_n15833), .B(new_n15836), .C(new_n16159), .D(new_n16162), .Y(new_n16163));
  NOR2xp33_ASAP7_75t_L      g15907(.A(new_n10332), .B(new_n1518), .Y(new_n16164));
  AOI221xp5_ASAP7_75t_L     g15908(.A1(\b[54] ), .A2(new_n1659), .B1(\b[55] ), .B2(new_n1507), .C(new_n16164), .Y(new_n16165));
  O2A1O1Ixp33_ASAP7_75t_L   g15909(.A1(new_n1521), .A2(new_n10339), .B(new_n16165), .C(new_n1501), .Y(new_n16166));
  O2A1O1Ixp33_ASAP7_75t_L   g15910(.A1(new_n1521), .A2(new_n10339), .B(new_n16165), .C(\a[20] ), .Y(new_n16167));
  INVx1_ASAP7_75t_L         g15911(.A(new_n16167), .Y(new_n16168));
  OAI21xp33_ASAP7_75t_L     g15912(.A1(new_n1501), .A2(new_n16166), .B(new_n16168), .Y(new_n16169));
  INVx1_ASAP7_75t_L         g15913(.A(new_n16169), .Y(new_n16170));
  O2A1O1Ixp33_ASAP7_75t_L   g15914(.A1(new_n15640), .A2(new_n16163), .B(new_n15639), .C(new_n16170), .Y(new_n16171));
  INVx1_ASAP7_75t_L         g15915(.A(new_n16171), .Y(new_n16172));
  O2A1O1Ixp33_ASAP7_75t_L   g15916(.A1(new_n1501), .A2(new_n16166), .B(new_n16168), .C(new_n16161), .Y(new_n16173));
  A2O1A1Ixp33_ASAP7_75t_L   g15917(.A1(new_n16172), .A2(new_n16161), .B(new_n16173), .C(new_n16156), .Y(new_n16174));
  O2A1O1Ixp33_ASAP7_75t_L   g15918(.A1(new_n15640), .A2(new_n16163), .B(new_n15639), .C(new_n16169), .Y(new_n16175));
  INVx1_ASAP7_75t_L         g15919(.A(new_n16175), .Y(new_n16176));
  O2A1O1Ixp33_ASAP7_75t_L   g15920(.A1(new_n16170), .A2(new_n16171), .B(new_n16176), .C(new_n16156), .Y(new_n16177));
  A2O1A1Ixp33_ASAP7_75t_L   g15921(.A1(new_n16156), .A2(new_n16174), .B(new_n16177), .C(new_n15957), .Y(new_n16178));
  INVx1_ASAP7_75t_L         g15922(.A(new_n16149), .Y(new_n16179));
  O2A1O1Ixp33_ASAP7_75t_L   g15923(.A1(new_n16145), .A2(new_n16146), .B(new_n16179), .C(new_n16154), .Y(new_n16180));
  A2O1A1O1Ixp25_ASAP7_75t_L g15924(.A1(new_n16132), .A2(new_n16134), .B(new_n15968), .C(new_n16136), .D(new_n16180), .Y(new_n16181));
  O2A1O1Ixp33_ASAP7_75t_L   g15925(.A1(new_n16145), .A2(new_n16146), .B(new_n16179), .C(new_n16137), .Y(new_n16182));
  O2A1O1Ixp33_ASAP7_75t_L   g15926(.A1(new_n16181), .A2(new_n16182), .B(new_n16174), .C(new_n16177), .Y(new_n16183));
  O2A1O1Ixp33_ASAP7_75t_L   g15927(.A1(new_n15955), .A2(new_n15956), .B(new_n16183), .C(new_n15945), .Y(new_n16184));
  INVx1_ASAP7_75t_L         g15928(.A(new_n15956), .Y(new_n16185));
  NAND2xp33_ASAP7_75t_L     g15929(.A(new_n15954), .B(new_n16185), .Y(new_n16186));
  NAND2xp33_ASAP7_75t_L     g15930(.A(new_n16183), .B(new_n16186), .Y(new_n16187));
  NAND3xp33_ASAP7_75t_L     g15931(.A(new_n15945), .B(new_n16178), .C(new_n16187), .Y(new_n16188));
  A2O1A1Ixp33_ASAP7_75t_L   g15932(.A1(new_n16184), .A2(new_n16178), .B(new_n15945), .C(new_n16188), .Y(new_n16189));
  O2A1O1Ixp33_ASAP7_75t_L   g15933(.A1(new_n15930), .A2(new_n15931), .B(new_n15933), .C(new_n16189), .Y(new_n16190));
  NAND2xp33_ASAP7_75t_L     g15934(.A(\a[11] ), .B(new_n15928), .Y(new_n16191));
  A2O1A1Ixp33_ASAP7_75t_L   g15935(.A1(new_n12986), .A2(new_n718), .B(new_n15927), .C(new_n637), .Y(new_n16192));
  A2O1A1Ixp33_ASAP7_75t_L   g15936(.A1(new_n16192), .A2(new_n16191), .B(new_n15931), .C(new_n15933), .Y(new_n16193));
  A2O1A1O1Ixp25_ASAP7_75t_L g15937(.A1(new_n16184), .A2(new_n16178), .B(new_n15945), .C(new_n16188), .D(new_n16193), .Y(new_n16194));
  NOR2xp33_ASAP7_75t_L      g15938(.A(new_n16190), .B(new_n16194), .Y(new_n16195));
  O2A1O1Ixp33_ASAP7_75t_L   g15939(.A1(new_n15913), .A2(new_n15914), .B(new_n15907), .C(new_n16195), .Y(new_n16196));
  AOI21xp33_ASAP7_75t_L     g15940(.A1(new_n16178), .A2(new_n16187), .B(new_n15945), .Y(new_n16197));
  INVx1_ASAP7_75t_L         g15941(.A(new_n16197), .Y(new_n16198));
  NAND3xp33_ASAP7_75t_L     g15942(.A(new_n16193), .B(new_n16188), .C(new_n16198), .Y(new_n16199));
  INVx1_ASAP7_75t_L         g15943(.A(new_n15931), .Y(new_n16200));
  A2O1A1Ixp33_ASAP7_75t_L   g15944(.A1(new_n15630), .A2(new_n15626), .B(new_n15880), .C(new_n15895), .Y(new_n16201));
  INVx1_ASAP7_75t_L         g15945(.A(new_n15928), .Y(new_n16202));
  O2A1O1Ixp33_ASAP7_75t_L   g15946(.A1(new_n16202), .A2(new_n637), .B(new_n16192), .C(new_n16201), .Y(new_n16203));
  O2A1O1Ixp33_ASAP7_75t_L   g15947(.A1(new_n15627), .A2(new_n15932), .B(new_n16200), .C(new_n16203), .Y(new_n16204));
  NAND2xp33_ASAP7_75t_L     g15948(.A(new_n16204), .B(new_n16189), .Y(new_n16205));
  OAI211xp5_ASAP7_75t_L     g15949(.A1(new_n15891), .A2(new_n15919), .B(new_n16205), .C(new_n16199), .Y(new_n16206));
  OAI21xp33_ASAP7_75t_L     g15950(.A1(new_n16190), .A2(new_n16194), .B(new_n15926), .Y(new_n16207));
  NAND2xp33_ASAP7_75t_L     g15951(.A(new_n16206), .B(new_n16207), .Y(new_n16208));
  A2O1A1Ixp33_ASAP7_75t_L   g15952(.A1(new_n15910), .A2(new_n15918), .B(new_n15922), .C(new_n16208), .Y(new_n16209));
  INVx1_ASAP7_75t_L         g15953(.A(new_n16209), .Y(new_n16210));
  OAI21xp33_ASAP7_75t_L     g15954(.A1(new_n15610), .A2(new_n15612), .B(new_n15341), .Y(new_n16211));
  INVx1_ASAP7_75t_L         g15955(.A(new_n15604), .Y(new_n16212));
  O2A1O1Ixp33_ASAP7_75t_L   g15956(.A1(new_n15344), .A2(new_n15346), .B(new_n15603), .C(new_n15601), .Y(new_n16213));
  A2O1A1Ixp33_ASAP7_75t_L   g15957(.A1(new_n15345), .A2(new_n16212), .B(new_n16213), .C(new_n15910), .Y(new_n16214));
  A2O1A1Ixp33_ASAP7_75t_L   g15958(.A1(new_n15911), .A2(new_n16211), .B(new_n15921), .C(new_n16214), .Y(new_n16215));
  O2A1O1Ixp33_ASAP7_75t_L   g15959(.A1(new_n16190), .A2(new_n16194), .B(new_n15926), .C(new_n16215), .Y(new_n16216));
  O2A1O1Ixp33_ASAP7_75t_L   g15960(.A1(new_n16196), .A2(new_n15926), .B(new_n16216), .C(new_n16210), .Y(\f[74] ));
  A2O1A1Ixp33_ASAP7_75t_L   g15961(.A1(new_n16188), .A2(new_n16198), .B(new_n16204), .C(new_n16200), .Y(new_n16218));
  INVx1_ASAP7_75t_L         g15962(.A(new_n15942), .Y(new_n16219));
  AOI31xp33_ASAP7_75t_L     g15963(.A1(new_n16178), .A2(new_n16187), .A3(new_n15944), .B(new_n16219), .Y(new_n16220));
  OAI22xp33_ASAP7_75t_L     g15964(.A1(new_n980), .A2(new_n12258), .B1(new_n12603), .B2(new_n864), .Y(new_n16221));
  AOI221xp5_ASAP7_75t_L     g15965(.A1(new_n886), .A2(\b[63] ), .B1(new_n873), .B2(new_n12961), .C(new_n16221), .Y(new_n16222));
  XNOR2x2_ASAP7_75t_L       g15966(.A(new_n867), .B(new_n16222), .Y(new_n16223));
  INVx1_ASAP7_75t_L         g15967(.A(new_n16223), .Y(new_n16224));
  NOR2xp33_ASAP7_75t_L      g15968(.A(new_n16224), .B(new_n16220), .Y(new_n16225));
  AND2x2_ASAP7_75t_L        g15969(.A(new_n16224), .B(new_n16220), .Y(new_n16226));
  OAI22xp33_ASAP7_75t_L     g15970(.A1(new_n1654), .A2(new_n10309), .B1(new_n10332), .B2(new_n1517), .Y(new_n16227));
  AOI221xp5_ASAP7_75t_L     g15971(.A1(new_n1511), .A2(\b[57] ), .B1(new_n1513), .B2(new_n10991), .C(new_n16227), .Y(new_n16228));
  XNOR2x2_ASAP7_75t_L       g15972(.A(new_n1501), .B(new_n16228), .Y(new_n16229));
  O2A1O1Ixp33_ASAP7_75t_L   g15973(.A1(new_n16173), .A2(new_n16175), .B(new_n16156), .C(new_n16171), .Y(new_n16230));
  NAND2xp33_ASAP7_75t_L     g15974(.A(new_n16229), .B(new_n16230), .Y(new_n16231));
  A2O1A1Ixp33_ASAP7_75t_L   g15975(.A1(new_n16148), .A2(new_n16147), .B(new_n16149), .C(new_n16137), .Y(new_n16232));
  AOI21xp33_ASAP7_75t_L     g15976(.A1(new_n16232), .A2(new_n16137), .B(new_n16182), .Y(new_n16233));
  A2O1A1O1Ixp25_ASAP7_75t_L g15977(.A1(new_n16176), .A2(new_n16170), .B(new_n16233), .C(new_n16172), .D(new_n16229), .Y(new_n16234));
  INVx1_ASAP7_75t_L         g15978(.A(new_n16234), .Y(new_n16235));
  NAND2xp33_ASAP7_75t_L     g15979(.A(new_n16231), .B(new_n16235), .Y(new_n16236));
  OAI22xp33_ASAP7_75t_L     g15980(.A1(new_n2572), .A2(new_n8427), .B1(new_n8755), .B2(new_n2410), .Y(new_n16237));
  AOI221xp5_ASAP7_75t_L     g15981(.A1(new_n2423), .A2(\b[51] ), .B1(new_n2417), .B2(new_n8790), .C(new_n16237), .Y(new_n16238));
  XNOR2x2_ASAP7_75t_L       g15982(.A(new_n2413), .B(new_n16238), .Y(new_n16239));
  NAND3xp33_ASAP7_75t_L     g15983(.A(new_n16152), .B(new_n15965), .C(new_n16239), .Y(new_n16240));
  INVx1_ASAP7_75t_L         g15984(.A(new_n16240), .Y(new_n16241));
  O2A1O1Ixp33_ASAP7_75t_L   g15985(.A1(new_n15966), .A2(new_n15963), .B(new_n16152), .C(new_n16239), .Y(new_n16242));
  NOR2xp33_ASAP7_75t_L      g15986(.A(new_n16242), .B(new_n16241), .Y(new_n16243));
  INVx1_ASAP7_75t_L         g15987(.A(new_n16243), .Y(new_n16244));
  INVx1_ASAP7_75t_L         g15988(.A(new_n16116), .Y(new_n16245));
  NOR2xp33_ASAP7_75t_L      g15989(.A(new_n15991), .B(new_n16245), .Y(new_n16246));
  A2O1A1O1Ixp25_ASAP7_75t_L g15990(.A1(new_n16122), .A2(\a[35] ), .B(new_n16123), .C(new_n16117), .D(new_n16246), .Y(new_n16247));
  INVx1_ASAP7_75t_L         g15991(.A(new_n16247), .Y(new_n16248));
  A2O1A1Ixp33_ASAP7_75t_L   g15992(.A1(\a[38] ), .A2(new_n16113), .B(new_n16114), .C(new_n16109), .Y(new_n16249));
  A2O1A1Ixp33_ASAP7_75t_L   g15993(.A1(new_n15766), .A2(new_n15993), .B(new_n16105), .C(new_n16249), .Y(new_n16250));
  A2O1A1Ixp33_ASAP7_75t_L   g15994(.A1(new_n15762), .A2(new_n15753), .B(new_n16093), .C(new_n16102), .Y(new_n16251));
  A2O1A1O1Ixp25_ASAP7_75t_L g15995(.A1(new_n16088), .A2(\a[44] ), .B(new_n16089), .C(new_n16082), .D(new_n16083), .Y(new_n16252));
  INVx1_ASAP7_75t_L         g15996(.A(new_n16252), .Y(new_n16253));
  NOR2xp33_ASAP7_75t_L      g15997(.A(new_n3891), .B(new_n7304), .Y(new_n16254));
  AOI221xp5_ASAP7_75t_L     g15998(.A1(\b[31] ), .A2(new_n6742), .B1(\b[33] ), .B2(new_n6442), .C(new_n16254), .Y(new_n16255));
  INVx1_ASAP7_75t_L         g15999(.A(new_n16255), .Y(new_n16256));
  A2O1A1Ixp33_ASAP7_75t_L   g16000(.A1(new_n4831), .A2(new_n6450), .B(new_n16256), .C(\a[44] ), .Y(new_n16257));
  O2A1O1Ixp33_ASAP7_75t_L   g16001(.A1(new_n6443), .A2(new_n4108), .B(new_n16255), .C(\a[44] ), .Y(new_n16258));
  NOR2xp33_ASAP7_75t_L      g16002(.A(new_n2703), .B(new_n10065), .Y(new_n16259));
  AOI221xp5_ASAP7_75t_L     g16003(.A1(new_n8175), .A2(\b[27] ), .B1(new_n8484), .B2(\b[25] ), .C(new_n16259), .Y(new_n16260));
  INVx1_ASAP7_75t_L         g16004(.A(new_n16260), .Y(new_n16261));
  A2O1A1Ixp33_ASAP7_75t_L   g16005(.A1(new_n2887), .A2(new_n8490), .B(new_n16261), .C(\a[50] ), .Y(new_n16262));
  O2A1O1Ixp33_ASAP7_75t_L   g16006(.A1(new_n8176), .A2(new_n2889), .B(new_n16260), .C(\a[50] ), .Y(new_n16263));
  NAND2xp33_ASAP7_75t_L     g16007(.A(new_n16008), .B(new_n16053), .Y(new_n16264));
  A2O1A1Ixp33_ASAP7_75t_L   g16008(.A1(new_n16054), .A2(new_n16009), .B(new_n16006), .C(new_n16264), .Y(new_n16265));
  NOR2xp33_ASAP7_75t_L      g16009(.A(new_n1150), .B(new_n11354), .Y(new_n16266));
  AOI221xp5_ASAP7_75t_L     g16010(.A1(\b[18] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[17] ), .C(new_n16266), .Y(new_n16267));
  INVx1_ASAP7_75t_L         g16011(.A(new_n16267), .Y(new_n16268));
  A2O1A1Ixp33_ASAP7_75t_L   g16012(.A1(new_n2329), .A2(new_n11351), .B(new_n16268), .C(\a[59] ), .Y(new_n16269));
  O2A1O1Ixp33_ASAP7_75t_L   g16013(.A1(new_n11053), .A2(new_n1464), .B(new_n16267), .C(\a[59] ), .Y(new_n16270));
  NOR2xp33_ASAP7_75t_L      g16014(.A(new_n748), .B(new_n13030), .Y(new_n16271));
  A2O1A1Ixp33_ASAP7_75t_L   g16015(.A1(new_n13028), .A2(\b[10] ), .B(new_n15655), .C(\a[11] ), .Y(new_n16272));
  NOR2xp33_ASAP7_75t_L      g16016(.A(\a[11] ), .B(new_n15657), .Y(new_n16273));
  INVx1_ASAP7_75t_L         g16017(.A(new_n16273), .Y(new_n16274));
  AND2x2_ASAP7_75t_L        g16018(.A(new_n16272), .B(new_n16274), .Y(new_n16275));
  INVx1_ASAP7_75t_L         g16019(.A(new_n16275), .Y(new_n16276));
  A2O1A1Ixp33_ASAP7_75t_L   g16020(.A1(new_n13028), .A2(\b[12] ), .B(new_n16271), .C(new_n16276), .Y(new_n16277));
  O2A1O1Ixp33_ASAP7_75t_L   g16021(.A1(new_n12669), .A2(new_n12671), .B(\b[12] ), .C(new_n16271), .Y(new_n16278));
  NAND2xp33_ASAP7_75t_L     g16022(.A(new_n16278), .B(new_n16275), .Y(new_n16279));
  AND2x2_ASAP7_75t_L        g16023(.A(new_n16279), .B(new_n16277), .Y(new_n16280));
  INVx1_ASAP7_75t_L         g16024(.A(new_n16280), .Y(new_n16281));
  NOR2xp33_ASAP7_75t_L      g16025(.A(new_n960), .B(new_n12318), .Y(new_n16282));
  AOI221xp5_ASAP7_75t_L     g16026(.A1(new_n11995), .A2(\b[15] ), .B1(new_n13314), .B2(\b[13] ), .C(new_n16282), .Y(new_n16283));
  INVx1_ASAP7_75t_L         g16027(.A(new_n16283), .Y(new_n16284));
  A2O1A1Ixp33_ASAP7_75t_L   g16028(.A1(new_n1052), .A2(new_n11997), .B(new_n16284), .C(\a[62] ), .Y(new_n16285));
  INVx1_ASAP7_75t_L         g16029(.A(new_n16285), .Y(new_n16286));
  A2O1A1Ixp33_ASAP7_75t_L   g16030(.A1(new_n1052), .A2(new_n11997), .B(new_n16284), .C(new_n11987), .Y(new_n16287));
  O2A1O1Ixp33_ASAP7_75t_L   g16031(.A1(new_n11987), .A2(new_n16286), .B(new_n16287), .C(new_n16281), .Y(new_n16288));
  O2A1O1Ixp33_ASAP7_75t_L   g16032(.A1(new_n11987), .A2(new_n16286), .B(new_n16287), .C(new_n16280), .Y(new_n16289));
  INVx1_ASAP7_75t_L         g16033(.A(new_n16289), .Y(new_n16290));
  OAI21xp33_ASAP7_75t_L     g16034(.A1(new_n16281), .A2(new_n16288), .B(new_n16290), .Y(new_n16291));
  O2A1O1Ixp33_ASAP7_75t_L   g16035(.A1(new_n12669), .A2(new_n12671), .B(\b[11] ), .C(new_n16015), .Y(new_n16292));
  INVx1_ASAP7_75t_L         g16036(.A(new_n16292), .Y(new_n16293));
  A2O1A1Ixp33_ASAP7_75t_L   g16037(.A1(new_n16293), .A2(new_n15656), .B(new_n16020), .C(new_n16291), .Y(new_n16294));
  INVx1_ASAP7_75t_L         g16038(.A(new_n16020), .Y(new_n16295));
  O2A1O1Ixp33_ASAP7_75t_L   g16039(.A1(new_n15657), .A2(new_n16292), .B(new_n16295), .C(new_n16291), .Y(new_n16296));
  AO21x2_ASAP7_75t_L        g16040(.A1(\a[59] ), .A2(new_n16269), .B(new_n16270), .Y(new_n16297));
  A2O1A1Ixp33_ASAP7_75t_L   g16041(.A1(new_n16294), .A2(new_n16291), .B(new_n16296), .C(new_n16297), .Y(new_n16298));
  O2A1O1Ixp33_ASAP7_75t_L   g16042(.A1(new_n15656), .A2(new_n16018), .B(new_n16021), .C(new_n16017), .Y(new_n16299));
  INVx1_ASAP7_75t_L         g16043(.A(new_n16294), .Y(new_n16300));
  INVx1_ASAP7_75t_L         g16044(.A(new_n16288), .Y(new_n16301));
  A2O1A1Ixp33_ASAP7_75t_L   g16045(.A1(new_n16301), .A2(new_n16280), .B(new_n16289), .C(new_n16299), .Y(new_n16302));
  O2A1O1Ixp33_ASAP7_75t_L   g16046(.A1(new_n16299), .A2(new_n16300), .B(new_n16302), .C(new_n16297), .Y(new_n16303));
  A2O1A1O1Ixp25_ASAP7_75t_L g16047(.A1(new_n16269), .A2(\a[59] ), .B(new_n16270), .C(new_n16298), .D(new_n16303), .Y(new_n16304));
  O2A1O1Ixp33_ASAP7_75t_L   g16048(.A1(new_n16013), .A2(new_n16026), .B(new_n16032), .C(new_n16024), .Y(new_n16305));
  NAND2xp33_ASAP7_75t_L     g16049(.A(new_n16305), .B(new_n16304), .Y(new_n16306));
  INVx1_ASAP7_75t_L         g16050(.A(new_n16305), .Y(new_n16307));
  A2O1A1Ixp33_ASAP7_75t_L   g16051(.A1(new_n16298), .A2(new_n16297), .B(new_n16303), .C(new_n16307), .Y(new_n16308));
  NAND2xp33_ASAP7_75t_L     g16052(.A(new_n16308), .B(new_n16306), .Y(new_n16309));
  INVx1_ASAP7_75t_L         g16053(.A(new_n16309), .Y(new_n16310));
  NOR2xp33_ASAP7_75t_L      g16054(.A(new_n1745), .B(new_n10388), .Y(new_n16311));
  AOI221xp5_ASAP7_75t_L     g16055(.A1(new_n10086), .A2(\b[21] ), .B1(new_n11361), .B2(\b[19] ), .C(new_n16311), .Y(new_n16312));
  O2A1O1Ixp33_ASAP7_75t_L   g16056(.A1(new_n10088), .A2(new_n1901), .B(new_n16312), .C(new_n10083), .Y(new_n16313));
  O2A1O1Ixp33_ASAP7_75t_L   g16057(.A1(new_n10088), .A2(new_n1901), .B(new_n16312), .C(\a[56] ), .Y(new_n16314));
  INVx1_ASAP7_75t_L         g16058(.A(new_n16314), .Y(new_n16315));
  O2A1O1Ixp33_ASAP7_75t_L   g16059(.A1(new_n16313), .A2(new_n10083), .B(new_n16315), .C(new_n16309), .Y(new_n16316));
  INVx1_ASAP7_75t_L         g16060(.A(new_n16316), .Y(new_n16317));
  INVx1_ASAP7_75t_L         g16061(.A(new_n16313), .Y(new_n16318));
  A2O1A1Ixp33_ASAP7_75t_L   g16062(.A1(\a[56] ), .A2(new_n16318), .B(new_n16314), .C(new_n16309), .Y(new_n16319));
  INVx1_ASAP7_75t_L         g16063(.A(new_n16319), .Y(new_n16320));
  O2A1O1Ixp33_ASAP7_75t_L   g16064(.A1(new_n16035), .A2(new_n16038), .B(new_n16040), .C(new_n16051), .Y(new_n16321));
  INVx1_ASAP7_75t_L         g16065(.A(new_n16321), .Y(new_n16322));
  A2O1A1Ixp33_ASAP7_75t_L   g16066(.A1(new_n16317), .A2(new_n16310), .B(new_n16320), .C(new_n16322), .Y(new_n16323));
  OAI211xp5_ASAP7_75t_L     g16067(.A1(new_n16309), .A2(new_n16316), .B(new_n16321), .C(new_n16319), .Y(new_n16324));
  NAND2xp33_ASAP7_75t_L     g16068(.A(new_n16324), .B(new_n16323), .Y(new_n16325));
  INVx1_ASAP7_75t_L         g16069(.A(new_n16325), .Y(new_n16326));
  NOR2xp33_ASAP7_75t_L      g16070(.A(new_n2188), .B(new_n10400), .Y(new_n16327));
  AOI221xp5_ASAP7_75t_L     g16071(.A1(new_n9102), .A2(\b[24] ), .B1(new_n10398), .B2(\b[22] ), .C(new_n16327), .Y(new_n16328));
  O2A1O1Ixp33_ASAP7_75t_L   g16072(.A1(new_n9104), .A2(new_n2853), .B(new_n16328), .C(new_n9099), .Y(new_n16329));
  O2A1O1Ixp33_ASAP7_75t_L   g16073(.A1(new_n9104), .A2(new_n2853), .B(new_n16328), .C(\a[53] ), .Y(new_n16330));
  INVx1_ASAP7_75t_L         g16074(.A(new_n16330), .Y(new_n16331));
  O2A1O1Ixp33_ASAP7_75t_L   g16075(.A1(new_n9099), .A2(new_n16329), .B(new_n16331), .C(new_n16325), .Y(new_n16332));
  INVx1_ASAP7_75t_L         g16076(.A(new_n16332), .Y(new_n16333));
  O2A1O1Ixp33_ASAP7_75t_L   g16077(.A1(new_n9099), .A2(new_n16329), .B(new_n16331), .C(new_n16326), .Y(new_n16334));
  A2O1A1Ixp33_ASAP7_75t_L   g16078(.A1(new_n16333), .A2(new_n16326), .B(new_n16334), .C(new_n16265), .Y(new_n16335));
  INVx1_ASAP7_75t_L         g16079(.A(new_n16334), .Y(new_n16336));
  O2A1O1Ixp33_ASAP7_75t_L   g16080(.A1(new_n16325), .A2(new_n16332), .B(new_n16336), .C(new_n16265), .Y(new_n16337));
  AO21x2_ASAP7_75t_L        g16081(.A1(\a[50] ), .A2(new_n16262), .B(new_n16263), .Y(new_n16338));
  A2O1A1Ixp33_ASAP7_75t_L   g16082(.A1(new_n16335), .A2(new_n16265), .B(new_n16337), .C(new_n16338), .Y(new_n16339));
  A2O1A1O1Ixp25_ASAP7_75t_L g16083(.A1(new_n16004), .A2(\a[53] ), .B(new_n16005), .C(new_n16062), .D(new_n16052), .Y(new_n16340));
  O2A1O1Ixp33_ASAP7_75t_L   g16084(.A1(new_n16325), .A2(new_n16332), .B(new_n16336), .C(new_n16340), .Y(new_n16341));
  A2O1A1Ixp33_ASAP7_75t_L   g16085(.A1(new_n16326), .A2(new_n16333), .B(new_n16334), .C(new_n16340), .Y(new_n16342));
  O2A1O1Ixp33_ASAP7_75t_L   g16086(.A1(new_n16340), .A2(new_n16341), .B(new_n16342), .C(new_n16338), .Y(new_n16343));
  A2O1A1O1Ixp25_ASAP7_75t_L g16087(.A1(new_n16262), .A2(\a[50] ), .B(new_n16263), .C(new_n16339), .D(new_n16343), .Y(new_n16344));
  A2O1A1O1Ixp25_ASAP7_75t_L g16088(.A1(new_n15998), .A2(\a[50] ), .B(new_n15999), .C(new_n16068), .D(new_n16059), .Y(new_n16345));
  NAND2xp33_ASAP7_75t_L     g16089(.A(new_n16345), .B(new_n16344), .Y(new_n16346));
  INVx1_ASAP7_75t_L         g16090(.A(new_n15706), .Y(new_n16347));
  A2O1A1Ixp33_ASAP7_75t_L   g16091(.A1(new_n16008), .A2(new_n16264), .B(new_n16056), .C(new_n16063), .Y(new_n16348));
  A2O1A1Ixp33_ASAP7_75t_L   g16092(.A1(new_n15713), .A2(new_n16347), .B(new_n16348), .C(new_n16066), .Y(new_n16349));
  A2O1A1Ixp33_ASAP7_75t_L   g16093(.A1(new_n16339), .A2(new_n16338), .B(new_n16343), .C(new_n16349), .Y(new_n16350));
  NOR2xp33_ASAP7_75t_L      g16094(.A(new_n3098), .B(new_n7312), .Y(new_n16351));
  AOI221xp5_ASAP7_75t_L     g16095(.A1(\b[28] ), .A2(new_n7609), .B1(\b[30] ), .B2(new_n7334), .C(new_n16351), .Y(new_n16352));
  OAI211xp5_ASAP7_75t_L     g16096(.A1(new_n7321), .A2(new_n3464), .B(\a[47] ), .C(new_n16352), .Y(new_n16353));
  INVx1_ASAP7_75t_L         g16097(.A(new_n16352), .Y(new_n16354));
  A2O1A1Ixp33_ASAP7_75t_L   g16098(.A1(new_n4813), .A2(new_n7322), .B(new_n16354), .C(new_n7316), .Y(new_n16355));
  NAND2xp33_ASAP7_75t_L     g16099(.A(new_n16353), .B(new_n16355), .Y(new_n16356));
  AOI21xp33_ASAP7_75t_L     g16100(.A1(new_n16350), .A2(new_n16346), .B(new_n16356), .Y(new_n16357));
  INVx1_ASAP7_75t_L         g16101(.A(new_n16357), .Y(new_n16358));
  O2A1O1Ixp33_ASAP7_75t_L   g16102(.A1(new_n15716), .A2(new_n15720), .B(new_n15730), .C(new_n16070), .Y(new_n16359));
  NOR2xp33_ASAP7_75t_L      g16103(.A(new_n16359), .B(new_n16077), .Y(new_n16360));
  NAND2xp33_ASAP7_75t_L     g16104(.A(new_n16346), .B(new_n16350), .Y(new_n16361));
  O2A1O1Ixp33_ASAP7_75t_L   g16105(.A1(new_n7321), .A2(new_n3464), .B(new_n16352), .C(new_n7316), .Y(new_n16362));
  O2A1O1Ixp33_ASAP7_75t_L   g16106(.A1(new_n16362), .A2(new_n7316), .B(new_n16355), .C(new_n16361), .Y(new_n16363));
  NOR3xp33_ASAP7_75t_L      g16107(.A(new_n16360), .B(new_n16363), .C(new_n16357), .Y(new_n16364));
  NOR2xp33_ASAP7_75t_L      g16108(.A(new_n16360), .B(new_n16364), .Y(new_n16365));
  INVx1_ASAP7_75t_L         g16109(.A(new_n16363), .Y(new_n16366));
  OAI21xp33_ASAP7_75t_L     g16110(.A1(new_n16357), .A2(new_n16360), .B(new_n16366), .Y(new_n16367));
  INVx1_ASAP7_75t_L         g16111(.A(new_n16367), .Y(new_n16368));
  AO21x2_ASAP7_75t_L        g16112(.A1(\a[44] ), .A2(new_n16257), .B(new_n16258), .Y(new_n16369));
  A2O1A1Ixp33_ASAP7_75t_L   g16113(.A1(new_n16368), .A2(new_n16358), .B(new_n16365), .C(new_n16369), .Y(new_n16370));
  A2O1A1Ixp33_ASAP7_75t_L   g16114(.A1(new_n16350), .A2(new_n16346), .B(new_n16356), .C(new_n16368), .Y(new_n16371));
  O2A1O1Ixp33_ASAP7_75t_L   g16115(.A1(new_n16360), .A2(new_n16364), .B(new_n16371), .C(new_n16369), .Y(new_n16372));
  A2O1A1O1Ixp25_ASAP7_75t_L g16116(.A1(new_n16257), .A2(\a[44] ), .B(new_n16258), .C(new_n16370), .D(new_n16372), .Y(new_n16373));
  NAND2xp33_ASAP7_75t_L     g16117(.A(new_n16253), .B(new_n16373), .Y(new_n16374));
  A2O1A1Ixp33_ASAP7_75t_L   g16118(.A1(new_n16369), .A2(new_n16370), .B(new_n16372), .C(new_n16252), .Y(new_n16375));
  AND2x2_ASAP7_75t_L        g16119(.A(new_n16375), .B(new_n16374), .Y(new_n16376));
  NOR2xp33_ASAP7_75t_L      g16120(.A(new_n4613), .B(new_n5641), .Y(new_n16377));
  AOI221xp5_ASAP7_75t_L     g16121(.A1(\b[34] ), .A2(new_n5920), .B1(\b[35] ), .B2(new_n5623), .C(new_n16377), .Y(new_n16378));
  O2A1O1Ixp33_ASAP7_75t_L   g16122(.A1(new_n5630), .A2(new_n4622), .B(new_n16378), .C(new_n5626), .Y(new_n16379));
  O2A1O1Ixp33_ASAP7_75t_L   g16123(.A1(new_n5630), .A2(new_n4622), .B(new_n16378), .C(\a[41] ), .Y(new_n16380));
  INVx1_ASAP7_75t_L         g16124(.A(new_n16380), .Y(new_n16381));
  O2A1O1Ixp33_ASAP7_75t_L   g16125(.A1(new_n16379), .A2(new_n5626), .B(new_n16381), .C(new_n16376), .Y(new_n16382));
  OA21x2_ASAP7_75t_L        g16126(.A1(new_n5626), .A2(new_n16379), .B(new_n16381), .Y(new_n16383));
  NAND2xp33_ASAP7_75t_L     g16127(.A(new_n16383), .B(new_n16376), .Y(new_n16384));
  INVx1_ASAP7_75t_L         g16128(.A(new_n16384), .Y(new_n16385));
  NOR2xp33_ASAP7_75t_L      g16129(.A(new_n16382), .B(new_n16385), .Y(new_n16386));
  XNOR2x2_ASAP7_75t_L       g16130(.A(new_n16251), .B(new_n16386), .Y(new_n16387));
  NOR2xp33_ASAP7_75t_L      g16131(.A(new_n5570), .B(new_n4908), .Y(new_n16388));
  AOI221xp5_ASAP7_75t_L     g16132(.A1(\b[37] ), .A2(new_n5139), .B1(\b[38] ), .B2(new_n4916), .C(new_n16388), .Y(new_n16389));
  O2A1O1Ixp33_ASAP7_75t_L   g16133(.A1(new_n4911), .A2(new_n5578), .B(new_n16389), .C(new_n4906), .Y(new_n16390));
  INVx1_ASAP7_75t_L         g16134(.A(new_n16390), .Y(new_n16391));
  O2A1O1Ixp33_ASAP7_75t_L   g16135(.A1(new_n4911), .A2(new_n5578), .B(new_n16389), .C(\a[38] ), .Y(new_n16392));
  AOI21xp33_ASAP7_75t_L     g16136(.A1(new_n16391), .A2(\a[38] ), .B(new_n16392), .Y(new_n16393));
  XNOR2x2_ASAP7_75t_L       g16137(.A(new_n16393), .B(new_n16387), .Y(new_n16394));
  NAND2xp33_ASAP7_75t_L     g16138(.A(new_n16250), .B(new_n16394), .Y(new_n16395));
  INVx1_ASAP7_75t_L         g16139(.A(new_n16392), .Y(new_n16396));
  O2A1O1Ixp33_ASAP7_75t_L   g16140(.A1(new_n16390), .A2(new_n4906), .B(new_n16396), .C(new_n16387), .Y(new_n16397));
  A2O1A1Ixp33_ASAP7_75t_L   g16141(.A1(\a[38] ), .A2(new_n16391), .B(new_n16392), .C(new_n16387), .Y(new_n16398));
  O2A1O1Ixp33_ASAP7_75t_L   g16142(.A1(new_n16387), .A2(new_n16397), .B(new_n16398), .C(new_n16250), .Y(new_n16399));
  INVx1_ASAP7_75t_L         g16143(.A(new_n16399), .Y(new_n16400));
  NAND2xp33_ASAP7_75t_L     g16144(.A(new_n16395), .B(new_n16400), .Y(new_n16401));
  NOR2xp33_ASAP7_75t_L      g16145(.A(new_n6378), .B(new_n4147), .Y(new_n16402));
  AOI221xp5_ASAP7_75t_L     g16146(.A1(\b[40] ), .A2(new_n4402), .B1(\b[41] ), .B2(new_n4155), .C(new_n16402), .Y(new_n16403));
  O2A1O1Ixp33_ASAP7_75t_L   g16147(.A1(new_n4150), .A2(new_n6386), .B(new_n16403), .C(new_n4145), .Y(new_n16404));
  INVx1_ASAP7_75t_L         g16148(.A(new_n16404), .Y(new_n16405));
  O2A1O1Ixp33_ASAP7_75t_L   g16149(.A1(new_n4150), .A2(new_n6386), .B(new_n16403), .C(\a[35] ), .Y(new_n16406));
  A2O1A1Ixp33_ASAP7_75t_L   g16150(.A1(\a[35] ), .A2(new_n16405), .B(new_n16406), .C(new_n16401), .Y(new_n16407));
  OAI21xp33_ASAP7_75t_L     g16151(.A1(new_n16387), .A2(new_n16397), .B(new_n16398), .Y(new_n16408));
  A2O1A1O1Ixp25_ASAP7_75t_L g16152(.A1(new_n15766), .A2(new_n15993), .B(new_n16105), .C(new_n16249), .D(new_n16408), .Y(new_n16409));
  NOR2xp33_ASAP7_75t_L      g16153(.A(new_n16399), .B(new_n16409), .Y(new_n16410));
  AOI21xp33_ASAP7_75t_L     g16154(.A1(new_n16405), .A2(\a[35] ), .B(new_n16406), .Y(new_n16411));
  NAND2xp33_ASAP7_75t_L     g16155(.A(new_n16411), .B(new_n16410), .Y(new_n16412));
  AOI21xp33_ASAP7_75t_L     g16156(.A1(new_n16412), .A2(new_n16407), .B(new_n16248), .Y(new_n16413));
  NOR2xp33_ASAP7_75t_L      g16157(.A(new_n16411), .B(new_n16410), .Y(new_n16414));
  INVx1_ASAP7_75t_L         g16158(.A(new_n16411), .Y(new_n16415));
  NOR2xp33_ASAP7_75t_L      g16159(.A(new_n16415), .B(new_n16401), .Y(new_n16416));
  NOR3xp33_ASAP7_75t_L      g16160(.A(new_n16414), .B(new_n16416), .C(new_n16247), .Y(new_n16417));
  OR2x4_ASAP7_75t_L         g16161(.A(new_n16413), .B(new_n16417), .Y(new_n16418));
  A2O1A1O1Ixp25_ASAP7_75t_L g16162(.A1(new_n16117), .A2(new_n16124), .B(new_n16127), .C(new_n15988), .D(new_n15985), .Y(new_n16419));
  NOR2xp33_ASAP7_75t_L      g16163(.A(new_n7249), .B(new_n3510), .Y(new_n16420));
  AOI221xp5_ASAP7_75t_L     g16164(.A1(\b[43] ), .A2(new_n3708), .B1(\b[44] ), .B2(new_n3499), .C(new_n16420), .Y(new_n16421));
  O2A1O1Ixp33_ASAP7_75t_L   g16165(.A1(new_n3513), .A2(new_n7255), .B(new_n16421), .C(new_n3493), .Y(new_n16422));
  O2A1O1Ixp33_ASAP7_75t_L   g16166(.A1(new_n3513), .A2(new_n7255), .B(new_n16421), .C(\a[32] ), .Y(new_n16423));
  INVx1_ASAP7_75t_L         g16167(.A(new_n16423), .Y(new_n16424));
  O2A1O1Ixp33_ASAP7_75t_L   g16168(.A1(new_n16422), .A2(new_n3493), .B(new_n16424), .C(new_n16419), .Y(new_n16425));
  INVx1_ASAP7_75t_L         g16169(.A(new_n16422), .Y(new_n16426));
  A2O1A1Ixp33_ASAP7_75t_L   g16170(.A1(\a[32] ), .A2(new_n16426), .B(new_n16423), .C(new_n16419), .Y(new_n16427));
  OAI21xp33_ASAP7_75t_L     g16171(.A1(new_n16419), .A2(new_n16425), .B(new_n16427), .Y(new_n16428));
  INVx1_ASAP7_75t_L         g16172(.A(new_n16428), .Y(new_n16429));
  NOR2xp33_ASAP7_75t_L      g16173(.A(new_n7860), .B(new_n2930), .Y(new_n16430));
  AOI221xp5_ASAP7_75t_L     g16174(.A1(\b[46] ), .A2(new_n3129), .B1(\b[47] ), .B2(new_n2936), .C(new_n16430), .Y(new_n16431));
  O2A1O1Ixp33_ASAP7_75t_L   g16175(.A1(new_n2940), .A2(new_n7868), .B(new_n16431), .C(new_n2928), .Y(new_n16432));
  INVx1_ASAP7_75t_L         g16176(.A(new_n16432), .Y(new_n16433));
  O2A1O1Ixp33_ASAP7_75t_L   g16177(.A1(new_n2940), .A2(new_n7868), .B(new_n16431), .C(\a[29] ), .Y(new_n16434));
  AOI21xp33_ASAP7_75t_L     g16178(.A1(new_n16433), .A2(\a[29] ), .B(new_n16434), .Y(new_n16435));
  A2O1A1Ixp33_ASAP7_75t_L   g16179(.A1(new_n15977), .A2(new_n16131), .B(new_n15976), .C(new_n16435), .Y(new_n16436));
  INVx1_ASAP7_75t_L         g16180(.A(new_n15976), .Y(new_n16437));
  INVx1_ASAP7_75t_L         g16181(.A(new_n16435), .Y(new_n16438));
  NAND3xp33_ASAP7_75t_L     g16182(.A(new_n16132), .B(new_n16437), .C(new_n16438), .Y(new_n16439));
  AOI21xp33_ASAP7_75t_L     g16183(.A1(new_n16426), .A2(\a[32] ), .B(new_n16423), .Y(new_n16440));
  INVx1_ASAP7_75t_L         g16184(.A(new_n15987), .Y(new_n16441));
  A2O1A1Ixp33_ASAP7_75t_L   g16185(.A1(new_n15983), .A2(new_n16441), .B(new_n16129), .C(new_n16440), .Y(new_n16442));
  O2A1O1Ixp33_ASAP7_75t_L   g16186(.A1(new_n16440), .A2(new_n16425), .B(new_n16442), .C(new_n16418), .Y(new_n16443));
  INVx1_ASAP7_75t_L         g16187(.A(new_n16443), .Y(new_n16444));
  NOR2xp33_ASAP7_75t_L      g16188(.A(new_n16413), .B(new_n16417), .Y(new_n16445));
  NOR2xp33_ASAP7_75t_L      g16189(.A(new_n16445), .B(new_n16428), .Y(new_n16446));
  INVx1_ASAP7_75t_L         g16190(.A(new_n16446), .Y(new_n16447));
  AOI22xp33_ASAP7_75t_L     g16191(.A1(new_n16439), .A2(new_n16436), .B1(new_n16447), .B2(new_n16444), .Y(new_n16448));
  A2O1A1Ixp33_ASAP7_75t_L   g16192(.A1(new_n16439), .A2(new_n16436), .B(new_n16443), .C(new_n16447), .Y(new_n16449));
  INVx1_ASAP7_75t_L         g16193(.A(new_n16449), .Y(new_n16450));
  O2A1O1Ixp33_ASAP7_75t_L   g16194(.A1(new_n16429), .A2(new_n16418), .B(new_n16450), .C(new_n16448), .Y(new_n16451));
  NAND2xp33_ASAP7_75t_L     g16195(.A(\b[54] ), .B(new_n1955), .Y(new_n16452));
  OAI221xp5_ASAP7_75t_L     g16196(.A1(new_n1962), .A2(new_n9683), .B1(new_n9355), .B2(new_n2089), .C(new_n16452), .Y(new_n16453));
  A2O1A1Ixp33_ASAP7_75t_L   g16197(.A1(new_n9717), .A2(new_n1964), .B(new_n16453), .C(\a[23] ), .Y(new_n16454));
  AOI21xp33_ASAP7_75t_L     g16198(.A1(new_n9717), .A2(new_n1964), .B(new_n16453), .Y(new_n16455));
  NOR2xp33_ASAP7_75t_L      g16199(.A(\a[23] ), .B(new_n16455), .Y(new_n16456));
  AOI21xp33_ASAP7_75t_L     g16200(.A1(new_n16454), .A2(\a[23] ), .B(new_n16456), .Y(new_n16457));
  A2O1A1O1Ixp25_ASAP7_75t_L g16201(.A1(new_n16179), .A2(new_n16145), .B(new_n16154), .C(new_n16147), .D(new_n16457), .Y(new_n16458));
  INVx1_ASAP7_75t_L         g16202(.A(new_n16458), .Y(new_n16459));
  A2O1A1Ixp33_ASAP7_75t_L   g16203(.A1(new_n16179), .A2(new_n16145), .B(new_n16154), .C(new_n16147), .Y(new_n16460));
  NOR2xp33_ASAP7_75t_L      g16204(.A(new_n16457), .B(new_n16460), .Y(new_n16461));
  O2A1O1Ixp33_ASAP7_75t_L   g16205(.A1(new_n16146), .A2(new_n16180), .B(new_n16459), .C(new_n16461), .Y(new_n16462));
  A2O1A1Ixp33_ASAP7_75t_L   g16206(.A1(new_n16450), .A2(new_n16444), .B(new_n16448), .C(new_n16243), .Y(new_n16463));
  NAND2xp33_ASAP7_75t_L     g16207(.A(new_n16436), .B(new_n16439), .Y(new_n16464));
  OAI21xp33_ASAP7_75t_L     g16208(.A1(new_n16443), .A2(new_n16446), .B(new_n16464), .Y(new_n16465));
  A2O1A1Ixp33_ASAP7_75t_L   g16209(.A1(new_n16445), .A2(new_n16428), .B(new_n16449), .C(new_n16465), .Y(new_n16466));
  NOR2xp33_ASAP7_75t_L      g16210(.A(new_n16243), .B(new_n16466), .Y(new_n16467));
  INVx1_ASAP7_75t_L         g16211(.A(new_n16467), .Y(new_n16468));
  AOI21xp33_ASAP7_75t_L     g16212(.A1(new_n16468), .A2(new_n16463), .B(new_n16462), .Y(new_n16469));
  A2O1A1O1Ixp25_ASAP7_75t_L g16213(.A1(new_n16460), .A2(new_n16459), .B(new_n16461), .C(new_n16463), .D(new_n16467), .Y(new_n16470));
  O2A1O1Ixp33_ASAP7_75t_L   g16214(.A1(new_n16451), .A2(new_n16244), .B(new_n16470), .C(new_n16469), .Y(new_n16471));
  O2A1O1Ixp33_ASAP7_75t_L   g16215(.A1(new_n16170), .A2(new_n16171), .B(new_n16176), .C(new_n16233), .Y(new_n16472));
  A2O1A1Ixp33_ASAP7_75t_L   g16216(.A1(new_n16172), .A2(new_n16161), .B(new_n16173), .C(new_n16233), .Y(new_n16473));
  A2O1A1Ixp33_ASAP7_75t_L   g16217(.A1(new_n16155), .A2(new_n16151), .B(new_n16472), .C(new_n16473), .Y(new_n16474));
  NOR2xp33_ASAP7_75t_L      g16218(.A(new_n11626), .B(new_n1284), .Y(new_n16475));
  AOI221xp5_ASAP7_75t_L     g16219(.A1(\b[58] ), .A2(new_n1290), .B1(\b[59] ), .B2(new_n1204), .C(new_n16475), .Y(new_n16476));
  O2A1O1Ixp33_ASAP7_75t_L   g16220(.A1(new_n1210), .A2(new_n11634), .B(new_n16476), .C(new_n1206), .Y(new_n16477));
  INVx1_ASAP7_75t_L         g16221(.A(new_n16477), .Y(new_n16478));
  O2A1O1Ixp33_ASAP7_75t_L   g16222(.A1(new_n1210), .A2(new_n11634), .B(new_n16476), .C(\a[17] ), .Y(new_n16479));
  AOI21xp33_ASAP7_75t_L     g16223(.A1(new_n16478), .A2(\a[17] ), .B(new_n16479), .Y(new_n16480));
  A2O1A1Ixp33_ASAP7_75t_L   g16224(.A1(new_n16474), .A2(new_n15954), .B(new_n15956), .C(new_n16480), .Y(new_n16481));
  A2O1A1O1Ixp25_ASAP7_75t_L g16225(.A1(new_n16174), .A2(new_n16156), .B(new_n16177), .C(new_n15954), .D(new_n15956), .Y(new_n16482));
  A2O1A1Ixp33_ASAP7_75t_L   g16226(.A1(\a[17] ), .A2(new_n16478), .B(new_n16479), .C(new_n16482), .Y(new_n16483));
  INVx1_ASAP7_75t_L         g16227(.A(new_n16229), .Y(new_n16484));
  A2O1A1Ixp33_ASAP7_75t_L   g16228(.A1(new_n16170), .A2(new_n16176), .B(new_n16233), .C(new_n16172), .Y(new_n16485));
  NOR2xp33_ASAP7_75t_L      g16229(.A(new_n16484), .B(new_n16485), .Y(new_n16486));
  NOR2xp33_ASAP7_75t_L      g16230(.A(new_n16234), .B(new_n16486), .Y(new_n16487));
  A2O1A1Ixp33_ASAP7_75t_L   g16231(.A1(new_n16470), .A2(new_n16463), .B(new_n16469), .C(new_n16487), .Y(new_n16488));
  NAND2xp33_ASAP7_75t_L     g16232(.A(new_n16471), .B(new_n16236), .Y(new_n16489));
  AOI22xp33_ASAP7_75t_L     g16233(.A1(new_n16483), .A2(new_n16481), .B1(new_n16489), .B2(new_n16488), .Y(new_n16490));
  INVx1_ASAP7_75t_L         g16234(.A(new_n16480), .Y(new_n16491));
  O2A1O1Ixp33_ASAP7_75t_L   g16235(.A1(new_n15955), .A2(new_n16183), .B(new_n16185), .C(new_n16491), .Y(new_n16492));
  AOI211xp5_ASAP7_75t_L     g16236(.A1(new_n16474), .A2(new_n15954), .B(new_n16480), .C(new_n15956), .Y(new_n16493));
  AO21x2_ASAP7_75t_L        g16237(.A1(new_n16470), .A2(new_n16463), .B(new_n16469), .Y(new_n16494));
  NOR2xp33_ASAP7_75t_L      g16238(.A(new_n16487), .B(new_n16494), .Y(new_n16495));
  O2A1O1Ixp33_ASAP7_75t_L   g16239(.A1(new_n16492), .A2(new_n16493), .B(new_n16488), .C(new_n16495), .Y(new_n16496));
  O2A1O1Ixp33_ASAP7_75t_L   g16240(.A1(new_n16471), .A2(new_n16236), .B(new_n16496), .C(new_n16490), .Y(new_n16497));
  OAI21xp33_ASAP7_75t_L     g16241(.A1(new_n16225), .A2(new_n16226), .B(new_n16497), .Y(new_n16498));
  A2O1A1Ixp33_ASAP7_75t_L   g16242(.A1(new_n16184), .A2(new_n16178), .B(new_n16219), .C(new_n16223), .Y(new_n16499));
  NAND2xp33_ASAP7_75t_L     g16243(.A(new_n16224), .B(new_n16220), .Y(new_n16500));
  NOR3xp33_ASAP7_75t_L      g16244(.A(new_n16464), .B(new_n16443), .C(new_n16446), .Y(new_n16501));
  A2O1A1Ixp33_ASAP7_75t_L   g16245(.A1(new_n16459), .A2(new_n16460), .B(new_n16461), .C(new_n16468), .Y(new_n16502));
  O2A1O1Ixp33_ASAP7_75t_L   g16246(.A1(new_n16448), .A2(new_n16501), .B(new_n16243), .C(new_n16502), .Y(new_n16503));
  A2O1A1Ixp33_ASAP7_75t_L   g16247(.A1(new_n16442), .A2(new_n16427), .B(new_n16418), .C(new_n16450), .Y(new_n16504));
  A2O1A1Ixp33_ASAP7_75t_L   g16248(.A1(new_n16465), .A2(new_n16504), .B(new_n16244), .C(new_n16470), .Y(new_n16505));
  O2A1O1Ixp33_ASAP7_75t_L   g16249(.A1(new_n16462), .A2(new_n16503), .B(new_n16505), .C(new_n16236), .Y(new_n16506));
  OAI22xp33_ASAP7_75t_L     g16250(.A1(new_n16495), .A2(new_n16506), .B1(new_n16493), .B2(new_n16492), .Y(new_n16507));
  A2O1A1Ixp33_ASAP7_75t_L   g16251(.A1(new_n16483), .A2(new_n16481), .B(new_n16506), .C(new_n16489), .Y(new_n16508));
  A2O1A1Ixp33_ASAP7_75t_L   g16252(.A1(new_n16487), .A2(new_n16494), .B(new_n16508), .C(new_n16507), .Y(new_n16509));
  NAND3xp33_ASAP7_75t_L     g16253(.A(new_n16509), .B(new_n16499), .C(new_n16500), .Y(new_n16510));
  NAND3xp33_ASAP7_75t_L     g16254(.A(new_n16510), .B(new_n16498), .C(new_n16218), .Y(new_n16511));
  O2A1O1Ixp33_ASAP7_75t_L   g16255(.A1(new_n16203), .A2(new_n16201), .B(new_n16189), .C(new_n15931), .Y(new_n16512));
  NOR2xp33_ASAP7_75t_L      g16256(.A(new_n16223), .B(new_n16220), .Y(new_n16513));
  O2A1O1Ixp33_ASAP7_75t_L   g16257(.A1(new_n16220), .A2(new_n16513), .B(new_n16500), .C(new_n16509), .Y(new_n16514));
  NOR3xp33_ASAP7_75t_L      g16258(.A(new_n16497), .B(new_n16226), .C(new_n16225), .Y(new_n16515));
  OAI21xp33_ASAP7_75t_L     g16259(.A1(new_n16514), .A2(new_n16515), .B(new_n16512), .Y(new_n16516));
  NAND2xp33_ASAP7_75t_L     g16260(.A(new_n16511), .B(new_n16516), .Y(new_n16517));
  A2O1A1O1Ixp25_ASAP7_75t_L g16261(.A1(new_n16184), .A2(new_n16178), .B(new_n15945), .C(new_n16188), .D(new_n16204), .Y(new_n16518));
  NAND2xp33_ASAP7_75t_L     g16262(.A(new_n16510), .B(new_n16498), .Y(new_n16519));
  A2O1A1Ixp33_ASAP7_75t_L   g16263(.A1(new_n16193), .A2(new_n16189), .B(new_n15931), .C(new_n16519), .Y(new_n16520));
  A2O1A1O1Ixp25_ASAP7_75t_L g16264(.A1(new_n15910), .A2(new_n15918), .B(new_n15922), .C(new_n16208), .D(new_n16196), .Y(new_n16521));
  A2O1A1Ixp33_ASAP7_75t_L   g16265(.A1(new_n16498), .A2(new_n16510), .B(new_n16218), .C(new_n16521), .Y(new_n16522));
  O2A1O1Ixp33_ASAP7_75t_L   g16266(.A1(new_n15931), .A2(new_n16518), .B(new_n16520), .C(new_n16522), .Y(new_n16523));
  O2A1O1Ixp33_ASAP7_75t_L   g16267(.A1(new_n16196), .A2(new_n16210), .B(new_n16517), .C(new_n16523), .Y(\f[75] ));
  O2A1O1Ixp33_ASAP7_75t_L   g16268(.A1(new_n16224), .A2(new_n16225), .B(new_n16509), .C(new_n16513), .Y(new_n16525));
  NOR2xp33_ASAP7_75t_L      g16269(.A(new_n9709), .B(new_n1962), .Y(new_n16526));
  AOI221xp5_ASAP7_75t_L     g16270(.A1(new_n1955), .A2(\b[55] ), .B1(new_n2093), .B2(\b[53] ), .C(new_n16526), .Y(new_n16527));
  INVx1_ASAP7_75t_L         g16271(.A(new_n16527), .Y(new_n16528));
  O2A1O1Ixp33_ASAP7_75t_L   g16272(.A1(new_n1956), .A2(new_n15849), .B(new_n16527), .C(new_n1952), .Y(new_n16529));
  INVx1_ASAP7_75t_L         g16273(.A(new_n16529), .Y(new_n16530));
  NOR2xp33_ASAP7_75t_L      g16274(.A(new_n1952), .B(new_n16529), .Y(new_n16531));
  A2O1A1O1Ixp25_ASAP7_75t_L g16275(.A1(new_n10320), .A2(new_n1964), .B(new_n16528), .C(new_n16530), .D(new_n16531), .Y(new_n16532));
  INVx1_ASAP7_75t_L         g16276(.A(new_n16532), .Y(new_n16533));
  A2O1A1Ixp33_ASAP7_75t_L   g16277(.A1(new_n16466), .A2(new_n16240), .B(new_n16242), .C(new_n16533), .Y(new_n16534));
  INVx1_ASAP7_75t_L         g16278(.A(new_n16242), .Y(new_n16535));
  O2A1O1Ixp33_ASAP7_75t_L   g16279(.A1(new_n16241), .A2(new_n16451), .B(new_n16535), .C(new_n16533), .Y(new_n16536));
  NOR2xp33_ASAP7_75t_L      g16280(.A(new_n8427), .B(new_n2930), .Y(new_n16537));
  AOI221xp5_ASAP7_75t_L     g16281(.A1(\b[47] ), .A2(new_n3129), .B1(\b[48] ), .B2(new_n2936), .C(new_n16537), .Y(new_n16538));
  O2A1O1Ixp33_ASAP7_75t_L   g16282(.A1(new_n2940), .A2(new_n14802), .B(new_n16538), .C(new_n2928), .Y(new_n16539));
  INVx1_ASAP7_75t_L         g16283(.A(new_n16539), .Y(new_n16540));
  O2A1O1Ixp33_ASAP7_75t_L   g16284(.A1(new_n2940), .A2(new_n14802), .B(new_n16538), .C(\a[29] ), .Y(new_n16541));
  AOI21xp33_ASAP7_75t_L     g16285(.A1(new_n16540), .A2(\a[29] ), .B(new_n16541), .Y(new_n16542));
  INVx1_ASAP7_75t_L         g16286(.A(new_n16542), .Y(new_n16543));
  A2O1A1Ixp33_ASAP7_75t_L   g16287(.A1(new_n16428), .A2(new_n16445), .B(new_n16425), .C(new_n16543), .Y(new_n16544));
  INVx1_ASAP7_75t_L         g16288(.A(new_n16425), .Y(new_n16545));
  A2O1A1O1Ixp25_ASAP7_75t_L g16289(.A1(new_n16427), .A2(new_n16419), .B(new_n16418), .C(new_n16545), .D(new_n16543), .Y(new_n16546));
  NAND2xp33_ASAP7_75t_L     g16290(.A(\b[39] ), .B(new_n4916), .Y(new_n16547));
  OAI221xp5_ASAP7_75t_L     g16291(.A1(new_n4908), .A2(new_n5855), .B1(new_n5311), .B2(new_n5144), .C(new_n16547), .Y(new_n16548));
  A2O1A1Ixp33_ASAP7_75t_L   g16292(.A1(new_n6651), .A2(new_n4912), .B(new_n16548), .C(\a[38] ), .Y(new_n16549));
  AOI211xp5_ASAP7_75t_L     g16293(.A1(new_n6651), .A2(new_n4912), .B(new_n16548), .C(new_n4906), .Y(new_n16550));
  A2O1A1O1Ixp25_ASAP7_75t_L g16294(.A1(new_n6651), .A2(new_n4912), .B(new_n16548), .C(new_n16549), .D(new_n16550), .Y(new_n16551));
  OAI21xp33_ASAP7_75t_L     g16295(.A1(new_n5626), .A2(new_n16099), .B(new_n16103), .Y(new_n16552));
  A2O1A1O1Ixp25_ASAP7_75t_L g16296(.A1(new_n16096), .A2(new_n16552), .B(new_n16094), .C(new_n16384), .D(new_n16382), .Y(new_n16553));
  NOR2xp33_ASAP7_75t_L      g16297(.A(new_n5074), .B(new_n5641), .Y(new_n16554));
  AOI221xp5_ASAP7_75t_L     g16298(.A1(\b[35] ), .A2(new_n5920), .B1(\b[36] ), .B2(new_n5623), .C(new_n16554), .Y(new_n16555));
  O2A1O1Ixp33_ASAP7_75t_L   g16299(.A1(new_n5630), .A2(new_n5083), .B(new_n16555), .C(new_n5626), .Y(new_n16556));
  NOR2xp33_ASAP7_75t_L      g16300(.A(new_n5626), .B(new_n16556), .Y(new_n16557));
  O2A1O1Ixp33_ASAP7_75t_L   g16301(.A1(new_n5630), .A2(new_n5083), .B(new_n16555), .C(\a[41] ), .Y(new_n16558));
  O2A1O1Ixp33_ASAP7_75t_L   g16302(.A1(new_n16080), .A2(new_n16081), .B(new_n16092), .C(new_n16373), .Y(new_n16559));
  INVx1_ASAP7_75t_L         g16303(.A(new_n16559), .Y(new_n16560));
  NOR2xp33_ASAP7_75t_L      g16304(.A(new_n3891), .B(new_n6741), .Y(new_n16561));
  AOI221xp5_ASAP7_75t_L     g16305(.A1(\b[34] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[33] ), .C(new_n16561), .Y(new_n16562));
  O2A1O1Ixp33_ASAP7_75t_L   g16306(.A1(new_n6443), .A2(new_n4352), .B(new_n16562), .C(new_n6439), .Y(new_n16563));
  INVx1_ASAP7_75t_L         g16307(.A(new_n16563), .Y(new_n16564));
  O2A1O1Ixp33_ASAP7_75t_L   g16308(.A1(new_n6443), .A2(new_n4352), .B(new_n16562), .C(\a[44] ), .Y(new_n16565));
  NOR2xp33_ASAP7_75t_L      g16309(.A(new_n3674), .B(new_n7318), .Y(new_n16566));
  AOI221xp5_ASAP7_75t_L     g16310(.A1(new_n7333), .A2(\b[30] ), .B1(new_n7609), .B2(\b[29] ), .C(new_n16566), .Y(new_n16567));
  O2A1O1Ixp33_ASAP7_75t_L   g16311(.A1(new_n7321), .A2(new_n3681), .B(new_n16567), .C(new_n7316), .Y(new_n16568));
  NOR2xp33_ASAP7_75t_L      g16312(.A(new_n7316), .B(new_n16568), .Y(new_n16569));
  O2A1O1Ixp33_ASAP7_75t_L   g16313(.A1(new_n7321), .A2(new_n3681), .B(new_n16567), .C(\a[47] ), .Y(new_n16570));
  NOR2xp33_ASAP7_75t_L      g16314(.A(new_n16570), .B(new_n16569), .Y(new_n16571));
  INVx1_ASAP7_75t_L         g16315(.A(new_n16571), .Y(new_n16572));
  O2A1O1Ixp33_ASAP7_75t_L   g16316(.A1(new_n16052), .A2(new_n16055), .B(new_n16335), .C(new_n16337), .Y(new_n16573));
  A2O1A1Ixp33_ASAP7_75t_L   g16317(.A1(\a[50] ), .A2(new_n16262), .B(new_n16263), .C(new_n16573), .Y(new_n16574));
  A2O1A1Ixp33_ASAP7_75t_L   g16318(.A1(new_n16574), .A2(new_n16573), .B(new_n16345), .C(new_n16339), .Y(new_n16575));
  NOR2xp33_ASAP7_75t_L      g16319(.A(new_n2205), .B(new_n10400), .Y(new_n16576));
  AOI221xp5_ASAP7_75t_L     g16320(.A1(new_n9102), .A2(\b[25] ), .B1(new_n10398), .B2(\b[23] ), .C(new_n16576), .Y(new_n16577));
  O2A1O1Ixp33_ASAP7_75t_L   g16321(.A1(new_n9104), .A2(new_n2385), .B(new_n16577), .C(new_n9099), .Y(new_n16578));
  INVx1_ASAP7_75t_L         g16322(.A(new_n16578), .Y(new_n16579));
  O2A1O1Ixp33_ASAP7_75t_L   g16323(.A1(new_n9104), .A2(new_n2385), .B(new_n16577), .C(\a[53] ), .Y(new_n16580));
  NOR2xp33_ASAP7_75t_L      g16324(.A(new_n1895), .B(new_n10388), .Y(new_n16581));
  AOI221xp5_ASAP7_75t_L     g16325(.A1(new_n10086), .A2(\b[22] ), .B1(new_n11361), .B2(\b[20] ), .C(new_n16581), .Y(new_n16582));
  O2A1O1Ixp33_ASAP7_75t_L   g16326(.A1(new_n10088), .A2(new_n2522), .B(new_n16582), .C(new_n10083), .Y(new_n16583));
  INVx1_ASAP7_75t_L         g16327(.A(new_n16583), .Y(new_n16584));
  O2A1O1Ixp33_ASAP7_75t_L   g16328(.A1(new_n10088), .A2(new_n2522), .B(new_n16582), .C(\a[56] ), .Y(new_n16585));
  A2O1A1Ixp33_ASAP7_75t_L   g16329(.A1(new_n13028), .A2(\b[10] ), .B(new_n15655), .C(new_n637), .Y(new_n16586));
  NOR2xp33_ASAP7_75t_L      g16330(.A(new_n833), .B(new_n13030), .Y(new_n16587));
  O2A1O1Ixp33_ASAP7_75t_L   g16331(.A1(new_n12669), .A2(new_n12671), .B(\b[13] ), .C(new_n16587), .Y(new_n16588));
  INVx1_ASAP7_75t_L         g16332(.A(new_n16588), .Y(new_n16589));
  A2O1A1O1Ixp25_ASAP7_75t_L g16333(.A1(new_n16272), .A2(new_n16274), .B(new_n16278), .C(new_n16586), .D(new_n16589), .Y(new_n16590));
  INVx1_ASAP7_75t_L         g16334(.A(new_n16590), .Y(new_n16591));
  NAND2xp33_ASAP7_75t_L     g16335(.A(new_n16588), .B(new_n16591), .Y(new_n16592));
  NOR2xp33_ASAP7_75t_L      g16336(.A(new_n1043), .B(new_n12318), .Y(new_n16593));
  AOI221xp5_ASAP7_75t_L     g16337(.A1(new_n11995), .A2(\b[16] ), .B1(new_n13314), .B2(\b[14] ), .C(new_n16593), .Y(new_n16594));
  O2A1O1Ixp33_ASAP7_75t_L   g16338(.A1(new_n11998), .A2(new_n1161), .B(new_n16594), .C(new_n11987), .Y(new_n16595));
  INVx1_ASAP7_75t_L         g16339(.A(new_n16594), .Y(new_n16596));
  A2O1A1Ixp33_ASAP7_75t_L   g16340(.A1(new_n1156), .A2(new_n11997), .B(new_n16596), .C(new_n11987), .Y(new_n16597));
  OAI21xp33_ASAP7_75t_L     g16341(.A1(new_n11987), .A2(new_n16595), .B(new_n16597), .Y(new_n16598));
  A2O1A1O1Ixp25_ASAP7_75t_L g16342(.A1(new_n16586), .A2(new_n16277), .B(new_n16590), .C(new_n16592), .D(new_n16598), .Y(new_n16599));
  A2O1A1Ixp33_ASAP7_75t_L   g16343(.A1(new_n16277), .A2(new_n16586), .B(new_n16590), .C(new_n16592), .Y(new_n16600));
  O2A1O1Ixp33_ASAP7_75t_L   g16344(.A1(new_n11987), .A2(new_n16595), .B(new_n16597), .C(new_n16600), .Y(new_n16601));
  NOR2xp33_ASAP7_75t_L      g16345(.A(new_n16601), .B(new_n16599), .Y(new_n16602));
  NAND3xp33_ASAP7_75t_L     g16346(.A(new_n16602), .B(new_n16294), .C(new_n16301), .Y(new_n16603));
  A2O1A1O1Ixp25_ASAP7_75t_L g16347(.A1(new_n16290), .A2(new_n16281), .B(new_n16299), .C(new_n16301), .D(new_n16602), .Y(new_n16604));
  INVx1_ASAP7_75t_L         g16348(.A(new_n16604), .Y(new_n16605));
  AND2x2_ASAP7_75t_L        g16349(.A(new_n16603), .B(new_n16605), .Y(new_n16606));
  NOR2xp33_ASAP7_75t_L      g16350(.A(new_n1349), .B(new_n11354), .Y(new_n16607));
  AOI221xp5_ASAP7_75t_L     g16351(.A1(\b[19] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[18] ), .C(new_n16607), .Y(new_n16608));
  O2A1O1Ixp33_ASAP7_75t_L   g16352(.A1(new_n11053), .A2(new_n1628), .B(new_n16608), .C(new_n11048), .Y(new_n16609));
  INVx1_ASAP7_75t_L         g16353(.A(new_n16609), .Y(new_n16610));
  O2A1O1Ixp33_ASAP7_75t_L   g16354(.A1(new_n11053), .A2(new_n1628), .B(new_n16608), .C(\a[59] ), .Y(new_n16611));
  A2O1A1Ixp33_ASAP7_75t_L   g16355(.A1(\a[59] ), .A2(new_n16610), .B(new_n16611), .C(new_n16606), .Y(new_n16612));
  INVx1_ASAP7_75t_L         g16356(.A(new_n16611), .Y(new_n16613));
  O2A1O1Ixp33_ASAP7_75t_L   g16357(.A1(new_n16609), .A2(new_n11048), .B(new_n16613), .C(new_n16606), .Y(new_n16614));
  AOI21xp33_ASAP7_75t_L     g16358(.A1(new_n16612), .A2(new_n16606), .B(new_n16614), .Y(new_n16615));
  A2O1A1O1Ixp25_ASAP7_75t_L g16359(.A1(new_n16301), .A2(new_n16280), .B(new_n16289), .C(new_n16294), .D(new_n16296), .Y(new_n16616));
  A2O1A1Ixp33_ASAP7_75t_L   g16360(.A1(\a[59] ), .A2(new_n16269), .B(new_n16270), .C(new_n16616), .Y(new_n16617));
  A2O1A1Ixp33_ASAP7_75t_L   g16361(.A1(new_n16617), .A2(new_n16616), .B(new_n16305), .C(new_n16298), .Y(new_n16618));
  INVx1_ASAP7_75t_L         g16362(.A(new_n16618), .Y(new_n16619));
  NAND2xp33_ASAP7_75t_L     g16363(.A(new_n16619), .B(new_n16615), .Y(new_n16620));
  O2A1O1Ixp33_ASAP7_75t_L   g16364(.A1(new_n16304), .A2(new_n16305), .B(new_n16298), .C(new_n16615), .Y(new_n16621));
  INVx1_ASAP7_75t_L         g16365(.A(new_n16621), .Y(new_n16622));
  AO21x2_ASAP7_75t_L        g16366(.A1(\a[56] ), .A2(new_n16584), .B(new_n16585), .Y(new_n16623));
  NAND3xp33_ASAP7_75t_L     g16367(.A(new_n16622), .B(new_n16620), .C(new_n16623), .Y(new_n16624));
  NAND2xp33_ASAP7_75t_L     g16368(.A(new_n16620), .B(new_n16622), .Y(new_n16625));
  NOR2xp33_ASAP7_75t_L      g16369(.A(new_n16623), .B(new_n16625), .Y(new_n16626));
  A2O1A1O1Ixp25_ASAP7_75t_L g16370(.A1(new_n16584), .A2(\a[56] ), .B(new_n16585), .C(new_n16624), .D(new_n16626), .Y(new_n16627));
  O2A1O1Ixp33_ASAP7_75t_L   g16371(.A1(new_n16310), .A2(new_n16320), .B(new_n16322), .C(new_n16316), .Y(new_n16628));
  NAND2xp33_ASAP7_75t_L     g16372(.A(new_n16628), .B(new_n16627), .Y(new_n16629));
  INVx1_ASAP7_75t_L         g16373(.A(new_n16628), .Y(new_n16630));
  A2O1A1Ixp33_ASAP7_75t_L   g16374(.A1(new_n16624), .A2(new_n16623), .B(new_n16626), .C(new_n16630), .Y(new_n16631));
  INVx1_ASAP7_75t_L         g16375(.A(new_n16580), .Y(new_n16632));
  OAI21xp33_ASAP7_75t_L     g16376(.A1(new_n9099), .A2(new_n16578), .B(new_n16632), .Y(new_n16633));
  NAND3xp33_ASAP7_75t_L     g16377(.A(new_n16629), .B(new_n16631), .C(new_n16633), .Y(new_n16634));
  NAND2xp33_ASAP7_75t_L     g16378(.A(new_n16631), .B(new_n16629), .Y(new_n16635));
  NOR2xp33_ASAP7_75t_L      g16379(.A(new_n16633), .B(new_n16635), .Y(new_n16636));
  A2O1A1O1Ixp25_ASAP7_75t_L g16380(.A1(new_n16579), .A2(\a[53] ), .B(new_n16580), .C(new_n16634), .D(new_n16636), .Y(new_n16637));
  O2A1O1Ixp33_ASAP7_75t_L   g16381(.A1(new_n16326), .A2(new_n16334), .B(new_n16265), .C(new_n16332), .Y(new_n16638));
  NAND2xp33_ASAP7_75t_L     g16382(.A(new_n16638), .B(new_n16637), .Y(new_n16639));
  INVx1_ASAP7_75t_L         g16383(.A(new_n16638), .Y(new_n16640));
  A2O1A1Ixp33_ASAP7_75t_L   g16384(.A1(new_n16634), .A2(new_n16633), .B(new_n16636), .C(new_n16640), .Y(new_n16641));
  AND2x2_ASAP7_75t_L        g16385(.A(new_n16641), .B(new_n16639), .Y(new_n16642));
  NOR2xp33_ASAP7_75t_L      g16386(.A(new_n2879), .B(new_n10065), .Y(new_n16643));
  AOI221xp5_ASAP7_75t_L     g16387(.A1(new_n8175), .A2(\b[28] ), .B1(new_n8484), .B2(\b[26] ), .C(new_n16643), .Y(new_n16644));
  O2A1O1Ixp33_ASAP7_75t_L   g16388(.A1(new_n8176), .A2(new_n3087), .B(new_n16644), .C(new_n8172), .Y(new_n16645));
  INVx1_ASAP7_75t_L         g16389(.A(new_n16645), .Y(new_n16646));
  O2A1O1Ixp33_ASAP7_75t_L   g16390(.A1(new_n8176), .A2(new_n3087), .B(new_n16644), .C(\a[50] ), .Y(new_n16647));
  AOI21xp33_ASAP7_75t_L     g16391(.A1(new_n16646), .A2(\a[50] ), .B(new_n16647), .Y(new_n16648));
  XNOR2x2_ASAP7_75t_L       g16392(.A(new_n16648), .B(new_n16642), .Y(new_n16649));
  INVx1_ASAP7_75t_L         g16393(.A(new_n16649), .Y(new_n16650));
  O2A1O1Ixp33_ASAP7_75t_L   g16394(.A1(new_n16344), .A2(new_n16345), .B(new_n16339), .C(new_n16650), .Y(new_n16651));
  INVx1_ASAP7_75t_L         g16395(.A(new_n16651), .Y(new_n16652));
  NOR2xp33_ASAP7_75t_L      g16396(.A(new_n16575), .B(new_n16650), .Y(new_n16653));
  A2O1A1Ixp33_ASAP7_75t_L   g16397(.A1(new_n16652), .A2(new_n16575), .B(new_n16653), .C(new_n16572), .Y(new_n16654));
  NOR2xp33_ASAP7_75t_L      g16398(.A(new_n16572), .B(new_n16653), .Y(new_n16655));
  A2O1A1Ixp33_ASAP7_75t_L   g16399(.A1(new_n16350), .A2(new_n16339), .B(new_n16649), .C(new_n16655), .Y(new_n16656));
  NAND3xp33_ASAP7_75t_L     g16400(.A(new_n16654), .B(new_n16367), .C(new_n16656), .Y(new_n16657));
  O2A1O1Ixp33_ASAP7_75t_L   g16401(.A1(new_n16344), .A2(new_n16345), .B(new_n16339), .C(new_n16649), .Y(new_n16658));
  INVx1_ASAP7_75t_L         g16402(.A(new_n16658), .Y(new_n16659));
  INVx1_ASAP7_75t_L         g16403(.A(new_n16654), .Y(new_n16660));
  A2O1A1Ixp33_ASAP7_75t_L   g16404(.A1(new_n16655), .A2(new_n16659), .B(new_n16660), .C(new_n16368), .Y(new_n16661));
  AND2x2_ASAP7_75t_L        g16405(.A(new_n16657), .B(new_n16661), .Y(new_n16662));
  A2O1A1Ixp33_ASAP7_75t_L   g16406(.A1(new_n16564), .A2(\a[44] ), .B(new_n16565), .C(new_n16662), .Y(new_n16663));
  NOR2xp33_ASAP7_75t_L      g16407(.A(new_n6439), .B(new_n16563), .Y(new_n16664));
  OR3x1_ASAP7_75t_L         g16408(.A(new_n16662), .B(new_n16664), .C(new_n16565), .Y(new_n16665));
  NAND2xp33_ASAP7_75t_L     g16409(.A(new_n16663), .B(new_n16665), .Y(new_n16666));
  O2A1O1Ixp33_ASAP7_75t_L   g16410(.A1(new_n16252), .A2(new_n16373), .B(new_n16370), .C(new_n16666), .Y(new_n16667));
  A2O1A1O1Ixp25_ASAP7_75t_L g16411(.A1(new_n16358), .A2(new_n16368), .B(new_n16365), .C(new_n16369), .D(new_n16559), .Y(new_n16668));
  NAND3xp33_ASAP7_75t_L     g16412(.A(new_n16668), .B(new_n16663), .C(new_n16665), .Y(new_n16669));
  A2O1A1Ixp33_ASAP7_75t_L   g16413(.A1(new_n16560), .A2(new_n16370), .B(new_n16667), .C(new_n16669), .Y(new_n16670));
  NOR2xp33_ASAP7_75t_L      g16414(.A(new_n16558), .B(new_n16557), .Y(new_n16671));
  NOR2xp33_ASAP7_75t_L      g16415(.A(new_n16357), .B(new_n16360), .Y(new_n16672));
  A2O1A1Ixp33_ASAP7_75t_L   g16416(.A1(new_n16366), .A2(new_n16672), .B(new_n16360), .C(new_n16371), .Y(new_n16673));
  A2O1A1Ixp33_ASAP7_75t_L   g16417(.A1(new_n16369), .A2(new_n16673), .B(new_n16559), .C(new_n16666), .Y(new_n16674));
  AND3x1_ASAP7_75t_L        g16418(.A(new_n16674), .B(new_n16669), .C(new_n16671), .Y(new_n16675));
  O2A1O1Ixp33_ASAP7_75t_L   g16419(.A1(new_n16557), .A2(new_n16558), .B(new_n16670), .C(new_n16675), .Y(new_n16676));
  A2O1A1Ixp33_ASAP7_75t_L   g16420(.A1(new_n16384), .A2(new_n16251), .B(new_n16382), .C(new_n16676), .Y(new_n16677));
  INVx1_ASAP7_75t_L         g16421(.A(new_n16677), .Y(new_n16678));
  NAND2xp33_ASAP7_75t_L     g16422(.A(new_n16553), .B(new_n16676), .Y(new_n16679));
  O2A1O1Ixp33_ASAP7_75t_L   g16423(.A1(new_n16553), .A2(new_n16678), .B(new_n16679), .C(new_n16551), .Y(new_n16680));
  A2O1A1Ixp33_ASAP7_75t_L   g16424(.A1(new_n16096), .A2(new_n16552), .B(new_n16094), .C(new_n16386), .Y(new_n16681));
  INVx1_ASAP7_75t_L         g16425(.A(new_n16681), .Y(new_n16682));
  NAND2xp33_ASAP7_75t_L     g16426(.A(new_n16551), .B(new_n16679), .Y(new_n16683));
  O2A1O1Ixp33_ASAP7_75t_L   g16427(.A1(new_n16382), .A2(new_n16682), .B(new_n16677), .C(new_n16683), .Y(new_n16684));
  NOR2xp33_ASAP7_75t_L      g16428(.A(new_n16684), .B(new_n16680), .Y(new_n16685));
  A2O1A1Ixp33_ASAP7_75t_L   g16429(.A1(new_n16408), .A2(new_n16250), .B(new_n16397), .C(new_n16685), .Y(new_n16686));
  INVx1_ASAP7_75t_L         g16430(.A(new_n16397), .Y(new_n16687));
  A2O1A1Ixp33_ASAP7_75t_L   g16431(.A1(new_n16108), .A2(new_n16249), .B(new_n16394), .C(new_n16687), .Y(new_n16688));
  INVx1_ASAP7_75t_L         g16432(.A(new_n16688), .Y(new_n16689));
  OAI21xp33_ASAP7_75t_L     g16433(.A1(new_n16680), .A2(new_n16684), .B(new_n16689), .Y(new_n16690));
  NOR2xp33_ASAP7_75t_L      g16434(.A(new_n6671), .B(new_n4147), .Y(new_n16691));
  AOI221xp5_ASAP7_75t_L     g16435(.A1(\b[41] ), .A2(new_n4402), .B1(\b[42] ), .B2(new_n4155), .C(new_n16691), .Y(new_n16692));
  O2A1O1Ixp33_ASAP7_75t_L   g16436(.A1(new_n4150), .A2(new_n6679), .B(new_n16692), .C(new_n4145), .Y(new_n16693));
  INVx1_ASAP7_75t_L         g16437(.A(new_n16693), .Y(new_n16694));
  O2A1O1Ixp33_ASAP7_75t_L   g16438(.A1(new_n4150), .A2(new_n6679), .B(new_n16692), .C(\a[35] ), .Y(new_n16695));
  AOI21xp33_ASAP7_75t_L     g16439(.A1(new_n16694), .A2(\a[35] ), .B(new_n16695), .Y(new_n16696));
  NAND3xp33_ASAP7_75t_L     g16440(.A(new_n16690), .B(new_n16686), .C(new_n16696), .Y(new_n16697));
  NAND2xp33_ASAP7_75t_L     g16441(.A(new_n16686), .B(new_n16690), .Y(new_n16698));
  A2O1A1Ixp33_ASAP7_75t_L   g16442(.A1(\a[35] ), .A2(new_n16694), .B(new_n16695), .C(new_n16698), .Y(new_n16699));
  NAND2xp33_ASAP7_75t_L     g16443(.A(new_n16697), .B(new_n16699), .Y(new_n16700));
  NAND2xp33_ASAP7_75t_L     g16444(.A(\b[45] ), .B(new_n3499), .Y(new_n16701));
  OAI221xp5_ASAP7_75t_L     g16445(.A1(new_n3510), .A2(new_n7270), .B1(new_n6944), .B2(new_n3703), .C(new_n16701), .Y(new_n16702));
  AOI21xp33_ASAP7_75t_L     g16446(.A1(new_n7278), .A2(new_n3505), .B(new_n16702), .Y(new_n16703));
  NAND2xp33_ASAP7_75t_L     g16447(.A(\a[32] ), .B(new_n16703), .Y(new_n16704));
  A2O1A1Ixp33_ASAP7_75t_L   g16448(.A1(new_n7278), .A2(new_n3505), .B(new_n16702), .C(new_n3493), .Y(new_n16705));
  NAND2xp33_ASAP7_75t_L     g16449(.A(new_n16705), .B(new_n16704), .Y(new_n16706));
  A2O1A1Ixp33_ASAP7_75t_L   g16450(.A1(new_n16412), .A2(new_n16248), .B(new_n16414), .C(new_n16706), .Y(new_n16707));
  O2A1O1Ixp33_ASAP7_75t_L   g16451(.A1(new_n16247), .A2(new_n16416), .B(new_n16407), .C(new_n16706), .Y(new_n16708));
  A2O1A1Ixp33_ASAP7_75t_L   g16452(.A1(new_n16706), .A2(new_n16707), .B(new_n16708), .C(new_n16700), .Y(new_n16709));
  AOI21xp33_ASAP7_75t_L     g16453(.A1(new_n16707), .A2(new_n16706), .B(new_n16708), .Y(new_n16710));
  NOR2xp33_ASAP7_75t_L      g16454(.A(new_n16710), .B(new_n16700), .Y(new_n16711));
  AOI21xp33_ASAP7_75t_L     g16455(.A1(new_n16709), .A2(new_n16700), .B(new_n16711), .Y(new_n16712));
  A2O1A1Ixp33_ASAP7_75t_L   g16456(.A1(new_n16544), .A2(new_n16543), .B(new_n16546), .C(new_n16712), .Y(new_n16713));
  INVx1_ASAP7_75t_L         g16457(.A(new_n16713), .Y(new_n16714));
  INVx1_ASAP7_75t_L         g16458(.A(new_n16544), .Y(new_n16715));
  INVx1_ASAP7_75t_L         g16459(.A(new_n16546), .Y(new_n16716));
  O2A1O1Ixp33_ASAP7_75t_L   g16460(.A1(new_n16542), .A2(new_n16715), .B(new_n16716), .C(new_n16712), .Y(new_n16717));
  NOR2xp33_ASAP7_75t_L      g16461(.A(new_n16712), .B(new_n16717), .Y(new_n16718));
  A2O1A1Ixp33_ASAP7_75t_L   g16462(.A1(new_n16540), .A2(\a[29] ), .B(new_n16541), .C(new_n16544), .Y(new_n16719));
  A2O1A1O1Ixp25_ASAP7_75t_L g16463(.A1(new_n16540), .A2(\a[29] ), .B(new_n16541), .C(new_n16544), .D(new_n16546), .Y(new_n16720));
  A2O1A1Ixp33_ASAP7_75t_L   g16464(.A1(new_n16700), .A2(new_n16709), .B(new_n16711), .C(new_n16720), .Y(new_n16721));
  A2O1A1Ixp33_ASAP7_75t_L   g16465(.A1(new_n16716), .A2(new_n16719), .B(new_n16717), .C(new_n16721), .Y(new_n16722));
  NAND2xp33_ASAP7_75t_L     g16466(.A(new_n16437), .B(new_n16132), .Y(new_n16723));
  AOI211xp5_ASAP7_75t_L     g16467(.A1(new_n16439), .A2(new_n16436), .B(new_n16443), .C(new_n16446), .Y(new_n16724));
  NAND2xp33_ASAP7_75t_L     g16468(.A(\b[51] ), .B(new_n2421), .Y(new_n16725));
  OAI221xp5_ASAP7_75t_L     g16469(.A1(new_n2415), .A2(new_n9355), .B1(new_n8755), .B2(new_n2572), .C(new_n16725), .Y(new_n16726));
  AOI21xp33_ASAP7_75t_L     g16470(.A1(new_n9367), .A2(new_n2417), .B(new_n16726), .Y(new_n16727));
  NAND2xp33_ASAP7_75t_L     g16471(.A(\a[26] ), .B(new_n16727), .Y(new_n16728));
  A2O1A1Ixp33_ASAP7_75t_L   g16472(.A1(new_n9367), .A2(new_n2417), .B(new_n16726), .C(new_n2413), .Y(new_n16729));
  NAND2xp33_ASAP7_75t_L     g16473(.A(new_n16729), .B(new_n16728), .Y(new_n16730));
  A2O1A1Ixp33_ASAP7_75t_L   g16474(.A1(new_n16438), .A2(new_n16723), .B(new_n16724), .C(new_n16730), .Y(new_n16731));
  O2A1O1Ixp33_ASAP7_75t_L   g16475(.A1(new_n15975), .A2(new_n16133), .B(new_n16437), .C(new_n16435), .Y(new_n16732));
  NOR3xp33_ASAP7_75t_L      g16476(.A(new_n16724), .B(new_n16732), .C(new_n16730), .Y(new_n16733));
  INVx1_ASAP7_75t_L         g16477(.A(new_n16733), .Y(new_n16734));
  NAND3xp33_ASAP7_75t_L     g16478(.A(new_n16722), .B(new_n16731), .C(new_n16734), .Y(new_n16735));
  INVx1_ASAP7_75t_L         g16479(.A(new_n16731), .Y(new_n16736));
  NOR3xp33_ASAP7_75t_L      g16480(.A(new_n16722), .B(new_n16736), .C(new_n16733), .Y(new_n16737));
  O2A1O1Ixp33_ASAP7_75t_L   g16481(.A1(new_n16714), .A2(new_n16718), .B(new_n16735), .C(new_n16737), .Y(new_n16738));
  A2O1A1Ixp33_ASAP7_75t_L   g16482(.A1(new_n16534), .A2(new_n16533), .B(new_n16536), .C(new_n16738), .Y(new_n16739));
  O2A1O1Ixp33_ASAP7_75t_L   g16483(.A1(new_n1956), .A2(new_n15849), .B(new_n16527), .C(\a[23] ), .Y(new_n16740));
  O2A1O1Ixp33_ASAP7_75t_L   g16484(.A1(new_n16531), .A2(new_n16740), .B(new_n16534), .C(new_n16536), .Y(new_n16741));
  A2O1A1Ixp33_ASAP7_75t_L   g16485(.A1(new_n16722), .A2(new_n16735), .B(new_n16737), .C(new_n16741), .Y(new_n16742));
  NAND2xp33_ASAP7_75t_L     g16486(.A(\b[57] ), .B(new_n1507), .Y(new_n16743));
  OAI221xp5_ASAP7_75t_L     g16487(.A1(new_n1518), .A2(new_n11303), .B1(new_n10332), .B2(new_n1654), .C(new_n16743), .Y(new_n16744));
  AOI21xp33_ASAP7_75t_L     g16488(.A1(new_n11314), .A2(new_n1513), .B(new_n16744), .Y(new_n16745));
  NAND2xp33_ASAP7_75t_L     g16489(.A(\a[20] ), .B(new_n16745), .Y(new_n16746));
  A2O1A1Ixp33_ASAP7_75t_L   g16490(.A1(new_n11314), .A2(new_n1513), .B(new_n16744), .C(new_n1501), .Y(new_n16747));
  NAND2xp33_ASAP7_75t_L     g16491(.A(new_n16747), .B(new_n16746), .Y(new_n16748));
  A2O1A1Ixp33_ASAP7_75t_L   g16492(.A1(new_n15826), .A2(new_n15830), .B(new_n15820), .C(new_n15834), .Y(new_n16749));
  A2O1A1Ixp33_ASAP7_75t_L   g16493(.A1(new_n16148), .A2(new_n16749), .B(new_n16180), .C(new_n16457), .Y(new_n16750));
  O2A1O1Ixp33_ASAP7_75t_L   g16494(.A1(new_n16457), .A2(new_n16458), .B(new_n16750), .C(new_n16467), .Y(new_n16751));
  A2O1A1Ixp33_ASAP7_75t_L   g16495(.A1(new_n16751), .A2(new_n16463), .B(new_n16458), .C(new_n16748), .Y(new_n16752));
  INVx1_ASAP7_75t_L         g16496(.A(new_n16460), .Y(new_n16753));
  O2A1O1Ixp33_ASAP7_75t_L   g16497(.A1(new_n16154), .A2(new_n16150), .B(new_n16147), .C(new_n16458), .Y(new_n16754));
  OAI211xp5_ASAP7_75t_L     g16498(.A1(new_n16754), .A2(new_n16461), .B(new_n16468), .C(new_n16463), .Y(new_n16755));
  O2A1O1Ixp33_ASAP7_75t_L   g16499(.A1(new_n16753), .A2(new_n16457), .B(new_n16755), .C(new_n16748), .Y(new_n16756));
  AO221x2_ASAP7_75t_L       g16500(.A1(new_n16752), .A2(new_n16748), .B1(new_n16742), .B2(new_n16739), .C(new_n16756), .Y(new_n16757));
  XNOR2x2_ASAP7_75t_L       g16501(.A(new_n16738), .B(new_n16741), .Y(new_n16758));
  A2O1A1Ixp33_ASAP7_75t_L   g16502(.A1(new_n16748), .A2(new_n16752), .B(new_n16756), .C(new_n16758), .Y(new_n16759));
  NAND2xp33_ASAP7_75t_L     g16503(.A(new_n16757), .B(new_n16759), .Y(new_n16760));
  NOR2xp33_ASAP7_75t_L      g16504(.A(new_n12258), .B(new_n1284), .Y(new_n16761));
  AOI221xp5_ASAP7_75t_L     g16505(.A1(\b[59] ), .A2(new_n1290), .B1(\b[60] ), .B2(new_n1204), .C(new_n16761), .Y(new_n16762));
  INVx1_ASAP7_75t_L         g16506(.A(new_n16762), .Y(new_n16763));
  O2A1O1Ixp33_ASAP7_75t_L   g16507(.A1(new_n1210), .A2(new_n14764), .B(new_n16762), .C(new_n1206), .Y(new_n16764));
  INVx1_ASAP7_75t_L         g16508(.A(new_n16764), .Y(new_n16765));
  NOR2xp33_ASAP7_75t_L      g16509(.A(new_n1206), .B(new_n16764), .Y(new_n16766));
  A2O1A1O1Ixp25_ASAP7_75t_L g16510(.A1(new_n12269), .A2(new_n1216), .B(new_n16763), .C(new_n16765), .D(new_n16766), .Y(new_n16767));
  INVx1_ASAP7_75t_L         g16511(.A(new_n16767), .Y(new_n16768));
  A2O1A1Ixp33_ASAP7_75t_L   g16512(.A1(new_n16459), .A2(new_n16460), .B(new_n16461), .C(new_n16755), .Y(new_n16769));
  A2O1A1O1Ixp25_ASAP7_75t_L g16513(.A1(new_n16505), .A2(new_n16769), .B(new_n16486), .C(new_n16235), .D(new_n16767), .Y(new_n16770));
  INVx1_ASAP7_75t_L         g16514(.A(new_n16770), .Y(new_n16771));
  A2O1A1O1Ixp25_ASAP7_75t_L g16515(.A1(new_n16505), .A2(new_n16769), .B(new_n16486), .C(new_n16235), .D(new_n16768), .Y(new_n16772));
  A2O1A1Ixp33_ASAP7_75t_L   g16516(.A1(new_n16771), .A2(new_n16768), .B(new_n16772), .C(new_n16760), .Y(new_n16773));
  A2O1A1O1Ixp25_ASAP7_75t_L g16517(.A1(new_n16470), .A2(new_n16463), .B(new_n16469), .C(new_n16231), .D(new_n16234), .Y(new_n16774));
  O2A1O1Ixp33_ASAP7_75t_L   g16518(.A1(new_n1210), .A2(new_n14764), .B(new_n16762), .C(\a[17] ), .Y(new_n16775));
  A2O1A1Ixp33_ASAP7_75t_L   g16519(.A1(new_n16765), .A2(\a[17] ), .B(new_n16775), .C(new_n16774), .Y(new_n16776));
  O2A1O1Ixp33_ASAP7_75t_L   g16520(.A1(new_n16774), .A2(new_n16770), .B(new_n16776), .C(new_n16760), .Y(new_n16777));
  OAI211xp5_ASAP7_75t_L     g16521(.A1(new_n16493), .A2(new_n16492), .B(new_n16488), .C(new_n16489), .Y(new_n16778));
  O2A1O1Ixp33_ASAP7_75t_L   g16522(.A1(new_n15955), .A2(new_n16183), .B(new_n16185), .C(new_n16480), .Y(new_n16779));
  INVx1_ASAP7_75t_L         g16523(.A(new_n16779), .Y(new_n16780));
  AOI22xp33_ASAP7_75t_L     g16524(.A1(new_n885), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n985), .Y(new_n16781));
  A2O1A1Ixp33_ASAP7_75t_L   g16525(.A1(new_n12990), .A2(new_n12988), .B(new_n872), .C(new_n16781), .Y(new_n16782));
  XNOR2x2_ASAP7_75t_L       g16526(.A(new_n867), .B(new_n16782), .Y(new_n16783));
  AO21x2_ASAP7_75t_L        g16527(.A1(new_n16780), .A2(new_n16778), .B(new_n16783), .Y(new_n16784));
  NAND3xp33_ASAP7_75t_L     g16528(.A(new_n16778), .B(new_n16780), .C(new_n16783), .Y(new_n16785));
  NAND2xp33_ASAP7_75t_L     g16529(.A(new_n16785), .B(new_n16784), .Y(new_n16786));
  A2O1A1Ixp33_ASAP7_75t_L   g16530(.A1(new_n16773), .A2(new_n16760), .B(new_n16777), .C(new_n16786), .Y(new_n16787));
  AOI21xp33_ASAP7_75t_L     g16531(.A1(new_n16773), .A2(new_n16760), .B(new_n16777), .Y(new_n16788));
  NAND3xp33_ASAP7_75t_L     g16532(.A(new_n16788), .B(new_n16784), .C(new_n16785), .Y(new_n16789));
  A2O1A1Ixp33_ASAP7_75t_L   g16533(.A1(new_n16215), .A2(new_n16208), .B(new_n16196), .C(new_n16517), .Y(new_n16790));
  INVx1_ASAP7_75t_L         g16534(.A(new_n16525), .Y(new_n16791));
  NAND3xp33_ASAP7_75t_L     g16535(.A(new_n16789), .B(new_n16787), .C(new_n16791), .Y(new_n16792));
  AOI21xp33_ASAP7_75t_L     g16536(.A1(new_n16789), .A2(new_n16787), .B(new_n16525), .Y(new_n16793));
  AOI31xp33_ASAP7_75t_L     g16537(.A1(new_n16792), .A2(new_n16787), .A3(new_n16789), .B(new_n16793), .Y(new_n16794));
  A2O1A1O1Ixp25_ASAP7_75t_L g16538(.A1(new_n16498), .A2(new_n16510), .B(new_n16512), .C(new_n16790), .D(new_n16794), .Y(new_n16795));
  A2O1A1Ixp33_ASAP7_75t_L   g16539(.A1(new_n16498), .A2(new_n16510), .B(new_n16512), .C(new_n16790), .Y(new_n16796));
  AOI31xp33_ASAP7_75t_L     g16540(.A1(new_n16792), .A2(new_n16789), .A3(new_n16787), .B(new_n16796), .Y(new_n16797));
  A2O1A1O1Ixp25_ASAP7_75t_L g16541(.A1(new_n16787), .A2(new_n16789), .B(new_n16525), .C(new_n16797), .D(new_n16795), .Y(\f[76] ));
  NOR2xp33_ASAP7_75t_L      g16542(.A(new_n16492), .B(new_n16493), .Y(new_n16799));
  O2A1O1Ixp33_ASAP7_75t_L   g16543(.A1(new_n16486), .A2(new_n16234), .B(new_n16471), .C(new_n16799), .Y(new_n16800));
  O2A1O1Ixp33_ASAP7_75t_L   g16544(.A1(new_n16236), .A2(new_n16471), .B(new_n16800), .C(new_n16779), .Y(new_n16801));
  A2O1A1Ixp33_ASAP7_75t_L   g16545(.A1(new_n16800), .A2(new_n16488), .B(new_n16779), .C(new_n16783), .Y(new_n16802));
  A2O1A1Ixp33_ASAP7_75t_L   g16546(.A1(new_n16785), .A2(new_n16801), .B(new_n16788), .C(new_n16802), .Y(new_n16803));
  INVx1_ASAP7_75t_L         g16547(.A(new_n16803), .Y(new_n16804));
  NOR2xp33_ASAP7_75t_L      g16548(.A(new_n12956), .B(new_n980), .Y(new_n16805));
  A2O1A1Ixp33_ASAP7_75t_L   g16549(.A1(new_n12986), .A2(new_n873), .B(new_n16805), .C(\a[14] ), .Y(new_n16806));
  A2O1A1O1Ixp25_ASAP7_75t_L g16550(.A1(new_n873), .A2(new_n14172), .B(new_n985), .C(\b[63] ), .D(new_n867), .Y(new_n16807));
  A2O1A1O1Ixp25_ASAP7_75t_L g16551(.A1(new_n12986), .A2(new_n873), .B(new_n16805), .C(new_n16806), .D(new_n16807), .Y(new_n16808));
  O2A1O1Ixp33_ASAP7_75t_L   g16552(.A1(new_n16766), .A2(new_n16775), .B(new_n16771), .C(new_n16772), .Y(new_n16809));
  A2O1A1O1Ixp25_ASAP7_75t_L g16553(.A1(new_n16759), .A2(new_n16757), .B(new_n16809), .C(new_n16771), .D(new_n16808), .Y(new_n16810));
  INVx1_ASAP7_75t_L         g16554(.A(new_n16808), .Y(new_n16811));
  A2O1A1O1Ixp25_ASAP7_75t_L g16555(.A1(new_n16759), .A2(new_n16757), .B(new_n16809), .C(new_n16771), .D(new_n16811), .Y(new_n16812));
  INVx1_ASAP7_75t_L         g16556(.A(new_n16812), .Y(new_n16813));
  NOR2xp33_ASAP7_75t_L      g16557(.A(new_n11591), .B(new_n1518), .Y(new_n16814));
  AOI221xp5_ASAP7_75t_L     g16558(.A1(\b[57] ), .A2(new_n1659), .B1(\b[58] ), .B2(new_n1507), .C(new_n16814), .Y(new_n16815));
  O2A1O1Ixp33_ASAP7_75t_L   g16559(.A1(new_n1521), .A2(new_n11597), .B(new_n16815), .C(new_n1501), .Y(new_n16816));
  INVx1_ASAP7_75t_L         g16560(.A(new_n16816), .Y(new_n16817));
  O2A1O1Ixp33_ASAP7_75t_L   g16561(.A1(new_n1521), .A2(new_n11597), .B(new_n16815), .C(\a[20] ), .Y(new_n16818));
  AOI21xp33_ASAP7_75t_L     g16562(.A1(new_n16817), .A2(\a[20] ), .B(new_n16818), .Y(new_n16819));
  INVx1_ASAP7_75t_L         g16563(.A(new_n16534), .Y(new_n16820));
  O2A1O1Ixp33_ASAP7_75t_L   g16564(.A1(new_n16448), .A2(new_n16501), .B(new_n16240), .C(new_n16242), .Y(new_n16821));
  A2O1A1Ixp33_ASAP7_75t_L   g16565(.A1(new_n16530), .A2(\a[23] ), .B(new_n16740), .C(new_n16821), .Y(new_n16822));
  A2O1A1Ixp33_ASAP7_75t_L   g16566(.A1(new_n16463), .A2(new_n16535), .B(new_n16820), .C(new_n16822), .Y(new_n16823));
  A2O1A1O1Ixp25_ASAP7_75t_L g16567(.A1(new_n16735), .A2(new_n16722), .B(new_n16737), .C(new_n16823), .D(new_n16820), .Y(new_n16824));
  NAND2xp33_ASAP7_75t_L     g16568(.A(new_n16819), .B(new_n16824), .Y(new_n16825));
  A2O1A1O1Ixp25_ASAP7_75t_L g16569(.A1(new_n16822), .A2(new_n16821), .B(new_n16738), .C(new_n16534), .D(new_n16819), .Y(new_n16826));
  INVx1_ASAP7_75t_L         g16570(.A(new_n16826), .Y(new_n16827));
  NOR2xp33_ASAP7_75t_L      g16571(.A(new_n10309), .B(new_n1962), .Y(new_n16828));
  AOI221xp5_ASAP7_75t_L     g16572(.A1(new_n1955), .A2(\b[56] ), .B1(new_n2093), .B2(\b[54] ), .C(new_n16828), .Y(new_n16829));
  O2A1O1Ixp33_ASAP7_75t_L   g16573(.A1(new_n1956), .A2(new_n10339), .B(new_n16829), .C(new_n1952), .Y(new_n16830));
  INVx1_ASAP7_75t_L         g16574(.A(new_n16830), .Y(new_n16831));
  O2A1O1Ixp33_ASAP7_75t_L   g16575(.A1(new_n1956), .A2(new_n10339), .B(new_n16829), .C(\a[23] ), .Y(new_n16832));
  AOI21xp33_ASAP7_75t_L     g16576(.A1(new_n16831), .A2(\a[23] ), .B(new_n16832), .Y(new_n16833));
  INVx1_ASAP7_75t_L         g16577(.A(new_n16833), .Y(new_n16834));
  A2O1A1Ixp33_ASAP7_75t_L   g16578(.A1(new_n16713), .A2(new_n16721), .B(new_n16733), .C(new_n16731), .Y(new_n16835));
  NOR2xp33_ASAP7_75t_L      g16579(.A(new_n16834), .B(new_n16835), .Y(new_n16836));
  A2O1A1O1Ixp25_ASAP7_75t_L g16580(.A1(new_n16713), .A2(new_n16721), .B(new_n16733), .C(new_n16731), .D(new_n16833), .Y(new_n16837));
  NOR2xp33_ASAP7_75t_L      g16581(.A(new_n16837), .B(new_n16836), .Y(new_n16838));
  NAND2xp33_ASAP7_75t_L     g16582(.A(\b[49] ), .B(new_n2936), .Y(new_n16839));
  OAI221xp5_ASAP7_75t_L     g16583(.A1(new_n2930), .A2(new_n8755), .B1(new_n7860), .B2(new_n3133), .C(new_n16839), .Y(new_n16840));
  AOI21xp33_ASAP7_75t_L     g16584(.A1(new_n8763), .A2(new_n2932), .B(new_n16840), .Y(new_n16841));
  NAND2xp33_ASAP7_75t_L     g16585(.A(\a[29] ), .B(new_n16841), .Y(new_n16842));
  A2O1A1Ixp33_ASAP7_75t_L   g16586(.A1(new_n8763), .A2(new_n2932), .B(new_n16840), .C(new_n2928), .Y(new_n16843));
  AND2x2_ASAP7_75t_L        g16587(.A(new_n16843), .B(new_n16842), .Y(new_n16844));
  A2O1A1O1Ixp25_ASAP7_75t_L g16588(.A1(new_n16699), .A2(new_n16697), .B(new_n16710), .C(new_n16707), .D(new_n16844), .Y(new_n16845));
  AND3x1_ASAP7_75t_L        g16589(.A(new_n16709), .B(new_n16844), .C(new_n16707), .Y(new_n16846));
  NOR2xp33_ASAP7_75t_L      g16590(.A(new_n16845), .B(new_n16846), .Y(new_n16847));
  INVx1_ASAP7_75t_L         g16591(.A(new_n16690), .Y(new_n16848));
  NAND2xp33_ASAP7_75t_L     g16592(.A(\b[46] ), .B(new_n3499), .Y(new_n16849));
  OAI221xp5_ASAP7_75t_L     g16593(.A1(new_n3510), .A2(new_n7552), .B1(new_n7249), .B2(new_n3703), .C(new_n16849), .Y(new_n16850));
  AOI21xp33_ASAP7_75t_L     g16594(.A1(new_n8726), .A2(new_n3505), .B(new_n16850), .Y(new_n16851));
  NAND2xp33_ASAP7_75t_L     g16595(.A(\a[32] ), .B(new_n16851), .Y(new_n16852));
  A2O1A1Ixp33_ASAP7_75t_L   g16596(.A1(new_n8726), .A2(new_n3505), .B(new_n16850), .C(new_n3493), .Y(new_n16853));
  NAND2xp33_ASAP7_75t_L     g16597(.A(new_n16853), .B(new_n16852), .Y(new_n16854));
  INVx1_ASAP7_75t_L         g16598(.A(new_n16854), .Y(new_n16855));
  O2A1O1Ixp33_ASAP7_75t_L   g16599(.A1(new_n16696), .A2(new_n16848), .B(new_n16686), .C(new_n16855), .Y(new_n16856));
  INVx1_ASAP7_75t_L         g16600(.A(new_n16856), .Y(new_n16857));
  OAI211xp5_ASAP7_75t_L     g16601(.A1(new_n16848), .A2(new_n16696), .B(new_n16686), .C(new_n16855), .Y(new_n16858));
  NAND2xp33_ASAP7_75t_L     g16602(.A(new_n16858), .B(new_n16857), .Y(new_n16859));
  O2A1O1Ixp33_ASAP7_75t_L   g16603(.A1(new_n16382), .A2(new_n16682), .B(new_n16676), .C(new_n16680), .Y(new_n16860));
  NOR2xp33_ASAP7_75t_L      g16604(.A(new_n6110), .B(new_n4908), .Y(new_n16861));
  AOI221xp5_ASAP7_75t_L     g16605(.A1(\b[39] ), .A2(new_n5139), .B1(\b[40] ), .B2(new_n4916), .C(new_n16861), .Y(new_n16862));
  O2A1O1Ixp33_ASAP7_75t_L   g16606(.A1(new_n4911), .A2(new_n6117), .B(new_n16862), .C(new_n4906), .Y(new_n16863));
  INVx1_ASAP7_75t_L         g16607(.A(new_n16863), .Y(new_n16864));
  O2A1O1Ixp33_ASAP7_75t_L   g16608(.A1(new_n4911), .A2(new_n6117), .B(new_n16862), .C(\a[38] ), .Y(new_n16865));
  O2A1O1Ixp33_ASAP7_75t_L   g16609(.A1(new_n16558), .A2(new_n16557), .B(new_n16670), .C(new_n16667), .Y(new_n16866));
  INVx1_ASAP7_75t_L         g16610(.A(new_n16866), .Y(new_n16867));
  O2A1O1Ixp33_ASAP7_75t_L   g16611(.A1(new_n16649), .A2(new_n16658), .B(new_n16572), .C(new_n16651), .Y(new_n16868));
  A2O1A1Ixp33_ASAP7_75t_L   g16612(.A1(new_n16323), .A2(new_n16317), .B(new_n16627), .C(new_n16634), .Y(new_n16869));
  NOR2xp33_ASAP7_75t_L      g16613(.A(new_n2377), .B(new_n10400), .Y(new_n16870));
  AOI221xp5_ASAP7_75t_L     g16614(.A1(new_n9102), .A2(\b[26] ), .B1(new_n10398), .B2(\b[24] ), .C(new_n16870), .Y(new_n16871));
  O2A1O1Ixp33_ASAP7_75t_L   g16615(.A1(new_n9104), .A2(new_n2708), .B(new_n16871), .C(new_n9099), .Y(new_n16872));
  INVx1_ASAP7_75t_L         g16616(.A(new_n16872), .Y(new_n16873));
  O2A1O1Ixp33_ASAP7_75t_L   g16617(.A1(new_n9104), .A2(new_n2708), .B(new_n16871), .C(\a[53] ), .Y(new_n16874));
  A2O1A1O1Ixp25_ASAP7_75t_L g16618(.A1(new_n16272), .A2(new_n16274), .B(new_n16278), .C(new_n16586), .D(new_n16588), .Y(new_n16875));
  A2O1A1Ixp33_ASAP7_75t_L   g16619(.A1(new_n16591), .A2(new_n16588), .B(new_n16875), .C(new_n16598), .Y(new_n16876));
  NOR2xp33_ASAP7_75t_L      g16620(.A(new_n936), .B(new_n13030), .Y(new_n16877));
  A2O1A1Ixp33_ASAP7_75t_L   g16621(.A1(\b[14] ), .A2(new_n13028), .B(new_n16877), .C(new_n16588), .Y(new_n16878));
  O2A1O1Ixp33_ASAP7_75t_L   g16622(.A1(new_n12669), .A2(new_n12671), .B(\b[14] ), .C(new_n16877), .Y(new_n16879));
  A2O1A1Ixp33_ASAP7_75t_L   g16623(.A1(new_n13028), .A2(\b[13] ), .B(new_n16587), .C(new_n16879), .Y(new_n16880));
  NAND2xp33_ASAP7_75t_L     g16624(.A(new_n16880), .B(new_n16878), .Y(new_n16881));
  NOR2xp33_ASAP7_75t_L      g16625(.A(new_n1150), .B(new_n12318), .Y(new_n16882));
  AOI221xp5_ASAP7_75t_L     g16626(.A1(new_n11995), .A2(\b[17] ), .B1(new_n13314), .B2(\b[15] ), .C(new_n16882), .Y(new_n16883));
  INVx1_ASAP7_75t_L         g16627(.A(new_n16883), .Y(new_n16884));
  A2O1A1Ixp33_ASAP7_75t_L   g16628(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n16883), .Y(new_n16885));
  A2O1A1Ixp33_ASAP7_75t_L   g16629(.A1(new_n1354), .A2(new_n1355), .B(new_n16884), .C(new_n16885), .Y(new_n16886));
  NAND2xp33_ASAP7_75t_L     g16630(.A(\a[62] ), .B(new_n16886), .Y(new_n16887));
  A2O1A1Ixp33_ASAP7_75t_L   g16631(.A1(new_n1633), .A2(new_n11997), .B(new_n16884), .C(new_n11987), .Y(new_n16888));
  AOI21xp33_ASAP7_75t_L     g16632(.A1(new_n16887), .A2(new_n16888), .B(new_n16881), .Y(new_n16889));
  INVx1_ASAP7_75t_L         g16633(.A(new_n16889), .Y(new_n16890));
  NAND3xp33_ASAP7_75t_L     g16634(.A(new_n16887), .B(new_n16888), .C(new_n16881), .Y(new_n16891));
  NAND2xp33_ASAP7_75t_L     g16635(.A(new_n16891), .B(new_n16890), .Y(new_n16892));
  A2O1A1O1Ixp25_ASAP7_75t_L g16636(.A1(new_n16277), .A2(new_n16586), .B(new_n16589), .C(new_n16876), .D(new_n16892), .Y(new_n16893));
  A2O1A1Ixp33_ASAP7_75t_L   g16637(.A1(new_n16586), .A2(new_n16277), .B(new_n16589), .C(new_n16876), .Y(new_n16894));
  AOI21xp33_ASAP7_75t_L     g16638(.A1(new_n16891), .A2(new_n16890), .B(new_n16894), .Y(new_n16895));
  NOR2xp33_ASAP7_75t_L      g16639(.A(new_n16895), .B(new_n16893), .Y(new_n16896));
  NOR2xp33_ASAP7_75t_L      g16640(.A(new_n1458), .B(new_n11354), .Y(new_n16897));
  AOI221xp5_ASAP7_75t_L     g16641(.A1(\b[20] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[19] ), .C(new_n16897), .Y(new_n16898));
  O2A1O1Ixp33_ASAP7_75t_L   g16642(.A1(new_n11053), .A2(new_n1754), .B(new_n16898), .C(new_n11048), .Y(new_n16899));
  INVx1_ASAP7_75t_L         g16643(.A(new_n16899), .Y(new_n16900));
  O2A1O1Ixp33_ASAP7_75t_L   g16644(.A1(new_n11053), .A2(new_n1754), .B(new_n16898), .C(\a[59] ), .Y(new_n16901));
  A2O1A1Ixp33_ASAP7_75t_L   g16645(.A1(\a[59] ), .A2(new_n16900), .B(new_n16901), .C(new_n16896), .Y(new_n16902));
  INVx1_ASAP7_75t_L         g16646(.A(new_n16901), .Y(new_n16903));
  O2A1O1Ixp33_ASAP7_75t_L   g16647(.A1(new_n16899), .A2(new_n11048), .B(new_n16903), .C(new_n16896), .Y(new_n16904));
  AOI21xp33_ASAP7_75t_L     g16648(.A1(new_n16902), .A2(new_n16896), .B(new_n16904), .Y(new_n16905));
  A2O1A1O1Ixp25_ASAP7_75t_L g16649(.A1(new_n16610), .A2(\a[59] ), .B(new_n16611), .C(new_n16603), .D(new_n16604), .Y(new_n16906));
  NAND2xp33_ASAP7_75t_L     g16650(.A(new_n16906), .B(new_n16905), .Y(new_n16907));
  INVx1_ASAP7_75t_L         g16651(.A(new_n16906), .Y(new_n16908));
  A2O1A1Ixp33_ASAP7_75t_L   g16652(.A1(new_n16902), .A2(new_n16896), .B(new_n16904), .C(new_n16908), .Y(new_n16909));
  AND2x2_ASAP7_75t_L        g16653(.A(new_n16909), .B(new_n16907), .Y(new_n16910));
  INVx1_ASAP7_75t_L         g16654(.A(new_n16910), .Y(new_n16911));
  NOR2xp33_ASAP7_75t_L      g16655(.A(new_n2045), .B(new_n10388), .Y(new_n16912));
  AOI221xp5_ASAP7_75t_L     g16656(.A1(new_n10086), .A2(\b[23] ), .B1(new_n11361), .B2(\b[21] ), .C(new_n16912), .Y(new_n16913));
  O2A1O1Ixp33_ASAP7_75t_L   g16657(.A1(new_n10088), .A2(new_n2194), .B(new_n16913), .C(new_n10083), .Y(new_n16914));
  O2A1O1Ixp33_ASAP7_75t_L   g16658(.A1(new_n10088), .A2(new_n2194), .B(new_n16913), .C(\a[56] ), .Y(new_n16915));
  INVx1_ASAP7_75t_L         g16659(.A(new_n16915), .Y(new_n16916));
  OAI211xp5_ASAP7_75t_L     g16660(.A1(new_n10083), .A2(new_n16914), .B(new_n16911), .C(new_n16916), .Y(new_n16917));
  INVx1_ASAP7_75t_L         g16661(.A(new_n16914), .Y(new_n16918));
  A2O1A1Ixp33_ASAP7_75t_L   g16662(.A1(\a[56] ), .A2(new_n16918), .B(new_n16915), .C(new_n16910), .Y(new_n16919));
  NAND2xp33_ASAP7_75t_L     g16663(.A(new_n16919), .B(new_n16917), .Y(new_n16920));
  O2A1O1Ixp33_ASAP7_75t_L   g16664(.A1(new_n16615), .A2(new_n16619), .B(new_n16624), .C(new_n16920), .Y(new_n16921));
  INVx1_ASAP7_75t_L         g16665(.A(new_n16921), .Y(new_n16922));
  A2O1A1O1Ixp25_ASAP7_75t_L g16666(.A1(new_n16584), .A2(\a[56] ), .B(new_n16585), .C(new_n16620), .D(new_n16621), .Y(new_n16923));
  NAND2xp33_ASAP7_75t_L     g16667(.A(new_n16923), .B(new_n16920), .Y(new_n16924));
  AND2x2_ASAP7_75t_L        g16668(.A(new_n16924), .B(new_n16922), .Y(new_n16925));
  A2O1A1Ixp33_ASAP7_75t_L   g16669(.A1(new_n16873), .A2(\a[53] ), .B(new_n16874), .C(new_n16925), .Y(new_n16926));
  AO221x2_ASAP7_75t_L       g16670(.A1(\a[53] ), .A2(new_n16873), .B1(new_n16922), .B2(new_n16924), .C(new_n16874), .Y(new_n16927));
  NAND3xp33_ASAP7_75t_L     g16671(.A(new_n16926), .B(new_n16869), .C(new_n16927), .Y(new_n16928));
  NAND2xp33_ASAP7_75t_L     g16672(.A(new_n16927), .B(new_n16926), .Y(new_n16929));
  NAND3xp33_ASAP7_75t_L     g16673(.A(new_n16929), .B(new_n16634), .C(new_n16631), .Y(new_n16930));
  AND2x2_ASAP7_75t_L        g16674(.A(new_n16928), .B(new_n16930), .Y(new_n16931));
  NOR2xp33_ASAP7_75t_L      g16675(.A(new_n3079), .B(new_n10065), .Y(new_n16932));
  AOI221xp5_ASAP7_75t_L     g16676(.A1(new_n8175), .A2(\b[29] ), .B1(new_n8484), .B2(\b[27] ), .C(new_n16932), .Y(new_n16933));
  O2A1O1Ixp33_ASAP7_75t_L   g16677(.A1(new_n8176), .A2(new_n3104), .B(new_n16933), .C(new_n8172), .Y(new_n16934));
  INVx1_ASAP7_75t_L         g16678(.A(new_n16934), .Y(new_n16935));
  O2A1O1Ixp33_ASAP7_75t_L   g16679(.A1(new_n8176), .A2(new_n3104), .B(new_n16933), .C(\a[50] ), .Y(new_n16936));
  A2O1A1Ixp33_ASAP7_75t_L   g16680(.A1(\a[50] ), .A2(new_n16935), .B(new_n16936), .C(new_n16931), .Y(new_n16937));
  INVx1_ASAP7_75t_L         g16681(.A(new_n16936), .Y(new_n16938));
  O2A1O1Ixp33_ASAP7_75t_L   g16682(.A1(new_n16934), .A2(new_n8172), .B(new_n16938), .C(new_n16931), .Y(new_n16939));
  AO21x2_ASAP7_75t_L        g16683(.A1(new_n16931), .A2(new_n16937), .B(new_n16939), .Y(new_n16940));
  A2O1A1Ixp33_ASAP7_75t_L   g16684(.A1(\a[50] ), .A2(new_n16646), .B(new_n16647), .C(new_n16642), .Y(new_n16941));
  A2O1A1Ixp33_ASAP7_75t_L   g16685(.A1(new_n16335), .A2(new_n16333), .B(new_n16637), .C(new_n16941), .Y(new_n16942));
  A2O1A1Ixp33_ASAP7_75t_L   g16686(.A1(new_n16937), .A2(new_n16931), .B(new_n16939), .C(new_n16942), .Y(new_n16943));
  O2A1O1Ixp33_ASAP7_75t_L   g16687(.A1(new_n16637), .A2(new_n16638), .B(new_n16941), .C(new_n16940), .Y(new_n16944));
  NOR2xp33_ASAP7_75t_L      g16688(.A(new_n3891), .B(new_n7318), .Y(new_n16945));
  AOI221xp5_ASAP7_75t_L     g16689(.A1(new_n7333), .A2(\b[31] ), .B1(new_n7609), .B2(\b[30] ), .C(new_n16945), .Y(new_n16946));
  O2A1O1Ixp33_ASAP7_75t_L   g16690(.A1(new_n7321), .A2(new_n3897), .B(new_n16946), .C(new_n7316), .Y(new_n16947));
  INVx1_ASAP7_75t_L         g16691(.A(new_n16947), .Y(new_n16948));
  O2A1O1Ixp33_ASAP7_75t_L   g16692(.A1(new_n7321), .A2(new_n3897), .B(new_n16946), .C(\a[47] ), .Y(new_n16949));
  AOI21xp33_ASAP7_75t_L     g16693(.A1(new_n16948), .A2(\a[47] ), .B(new_n16949), .Y(new_n16950));
  A2O1A1Ixp33_ASAP7_75t_L   g16694(.A1(new_n16943), .A2(new_n16940), .B(new_n16944), .C(new_n16950), .Y(new_n16951));
  A2O1A1O1Ixp25_ASAP7_75t_L g16695(.A1(new_n16937), .A2(new_n16931), .B(new_n16939), .C(new_n16943), .D(new_n16944), .Y(new_n16952));
  A2O1A1Ixp33_ASAP7_75t_L   g16696(.A1(\a[47] ), .A2(new_n16948), .B(new_n16949), .C(new_n16952), .Y(new_n16953));
  NAND2xp33_ASAP7_75t_L     g16697(.A(new_n16951), .B(new_n16953), .Y(new_n16954));
  INVx1_ASAP7_75t_L         g16698(.A(new_n16954), .Y(new_n16955));
  NAND2xp33_ASAP7_75t_L     g16699(.A(new_n16868), .B(new_n16955), .Y(new_n16956));
  A2O1A1Ixp33_ASAP7_75t_L   g16700(.A1(new_n16649), .A2(new_n16575), .B(new_n16660), .C(new_n16954), .Y(new_n16957));
  NAND2xp33_ASAP7_75t_L     g16701(.A(new_n16957), .B(new_n16956), .Y(new_n16958));
  NOR2xp33_ASAP7_75t_L      g16702(.A(new_n4101), .B(new_n6741), .Y(new_n16959));
  AOI221xp5_ASAP7_75t_L     g16703(.A1(\b[35] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[34] ), .C(new_n16959), .Y(new_n16960));
  O2A1O1Ixp33_ASAP7_75t_L   g16704(.A1(new_n6443), .A2(new_n4589), .B(new_n16960), .C(new_n6439), .Y(new_n16961));
  O2A1O1Ixp33_ASAP7_75t_L   g16705(.A1(new_n6443), .A2(new_n4589), .B(new_n16960), .C(\a[44] ), .Y(new_n16962));
  INVx1_ASAP7_75t_L         g16706(.A(new_n16962), .Y(new_n16963));
  O2A1O1Ixp33_ASAP7_75t_L   g16707(.A1(new_n16961), .A2(new_n6439), .B(new_n16963), .C(new_n16958), .Y(new_n16964));
  INVx1_ASAP7_75t_L         g16708(.A(new_n16961), .Y(new_n16965));
  A2O1A1Ixp33_ASAP7_75t_L   g16709(.A1(\a[44] ), .A2(new_n16965), .B(new_n16962), .C(new_n16958), .Y(new_n16966));
  OA21x2_ASAP7_75t_L        g16710(.A1(new_n16958), .A2(new_n16964), .B(new_n16966), .Y(new_n16967));
  INVx1_ASAP7_75t_L         g16711(.A(new_n16657), .Y(new_n16968));
  O2A1O1Ixp33_ASAP7_75t_L   g16712(.A1(new_n16565), .A2(new_n16664), .B(new_n16661), .C(new_n16968), .Y(new_n16969));
  NAND2xp33_ASAP7_75t_L     g16713(.A(new_n16969), .B(new_n16967), .Y(new_n16970));
  O2A1O1Ixp33_ASAP7_75t_L   g16714(.A1(new_n16958), .A2(new_n16964), .B(new_n16966), .C(new_n16969), .Y(new_n16971));
  INVx1_ASAP7_75t_L         g16715(.A(new_n16971), .Y(new_n16972));
  AND2x2_ASAP7_75t_L        g16716(.A(new_n16972), .B(new_n16970), .Y(new_n16973));
  NOR2xp33_ASAP7_75t_L      g16717(.A(new_n5311), .B(new_n5641), .Y(new_n16974));
  AOI221xp5_ASAP7_75t_L     g16718(.A1(\b[36] ), .A2(new_n5920), .B1(\b[37] ), .B2(new_n5623), .C(new_n16974), .Y(new_n16975));
  O2A1O1Ixp33_ASAP7_75t_L   g16719(.A1(new_n5630), .A2(new_n5318), .B(new_n16975), .C(new_n5626), .Y(new_n16976));
  O2A1O1Ixp33_ASAP7_75t_L   g16720(.A1(new_n5630), .A2(new_n5318), .B(new_n16975), .C(\a[41] ), .Y(new_n16977));
  INVx1_ASAP7_75t_L         g16721(.A(new_n16977), .Y(new_n16978));
  OAI21xp33_ASAP7_75t_L     g16722(.A1(new_n5626), .A2(new_n16976), .B(new_n16978), .Y(new_n16979));
  NOR2xp33_ASAP7_75t_L      g16723(.A(new_n16979), .B(new_n16973), .Y(new_n16980));
  NAND2xp33_ASAP7_75t_L     g16724(.A(new_n16972), .B(new_n16970), .Y(new_n16981));
  O2A1O1Ixp33_ASAP7_75t_L   g16725(.A1(new_n16976), .A2(new_n5626), .B(new_n16978), .C(new_n16981), .Y(new_n16982));
  NOR2xp33_ASAP7_75t_L      g16726(.A(new_n16982), .B(new_n16980), .Y(new_n16983));
  NAND2xp33_ASAP7_75t_L     g16727(.A(new_n16867), .B(new_n16983), .Y(new_n16984));
  OAI211xp5_ASAP7_75t_L     g16728(.A1(new_n5626), .A2(new_n16976), .B(new_n16981), .C(new_n16978), .Y(new_n16985));
  INVx1_ASAP7_75t_L         g16729(.A(new_n16976), .Y(new_n16986));
  A2O1A1Ixp33_ASAP7_75t_L   g16730(.A1(\a[41] ), .A2(new_n16986), .B(new_n16977), .C(new_n16973), .Y(new_n16987));
  NAND2xp33_ASAP7_75t_L     g16731(.A(new_n16985), .B(new_n16987), .Y(new_n16988));
  NAND2xp33_ASAP7_75t_L     g16732(.A(new_n16866), .B(new_n16988), .Y(new_n16989));
  AND2x2_ASAP7_75t_L        g16733(.A(new_n16984), .B(new_n16989), .Y(new_n16990));
  A2O1A1Ixp33_ASAP7_75t_L   g16734(.A1(new_n16864), .A2(\a[38] ), .B(new_n16865), .C(new_n16990), .Y(new_n16991));
  AOI21xp33_ASAP7_75t_L     g16735(.A1(new_n16864), .A2(\a[38] ), .B(new_n16865), .Y(new_n16992));
  NAND2xp33_ASAP7_75t_L     g16736(.A(new_n16984), .B(new_n16989), .Y(new_n16993));
  NAND2xp33_ASAP7_75t_L     g16737(.A(new_n16992), .B(new_n16993), .Y(new_n16994));
  NAND2xp33_ASAP7_75t_L     g16738(.A(new_n16994), .B(new_n16991), .Y(new_n16995));
  XOR2x2_ASAP7_75t_L        g16739(.A(new_n16860), .B(new_n16995), .Y(new_n16996));
  NOR2xp33_ASAP7_75t_L      g16740(.A(new_n6944), .B(new_n4147), .Y(new_n16997));
  AOI221xp5_ASAP7_75t_L     g16741(.A1(\b[42] ), .A2(new_n4402), .B1(\b[43] ), .B2(new_n4155), .C(new_n16997), .Y(new_n16998));
  O2A1O1Ixp33_ASAP7_75t_L   g16742(.A1(new_n4150), .A2(new_n6951), .B(new_n16998), .C(new_n4145), .Y(new_n16999));
  INVx1_ASAP7_75t_L         g16743(.A(new_n16999), .Y(new_n17000));
  O2A1O1Ixp33_ASAP7_75t_L   g16744(.A1(new_n4150), .A2(new_n6951), .B(new_n16998), .C(\a[35] ), .Y(new_n17001));
  A2O1A1Ixp33_ASAP7_75t_L   g16745(.A1(new_n17000), .A2(\a[35] ), .B(new_n17001), .C(new_n16996), .Y(new_n17002));
  INVx1_ASAP7_75t_L         g16746(.A(new_n17001), .Y(new_n17003));
  O2A1O1Ixp33_ASAP7_75t_L   g16747(.A1(new_n4145), .A2(new_n16999), .B(new_n17003), .C(new_n16996), .Y(new_n17004));
  AO21x2_ASAP7_75t_L        g16748(.A1(new_n16996), .A2(new_n17002), .B(new_n17004), .Y(new_n17005));
  AND3x1_ASAP7_75t_L        g16749(.A(new_n17005), .B(new_n16858), .C(new_n16857), .Y(new_n17006));
  A2O1A1Ixp33_ASAP7_75t_L   g16750(.A1(new_n16996), .A2(new_n17002), .B(new_n17004), .C(new_n16859), .Y(new_n17007));
  OAI21xp33_ASAP7_75t_L     g16751(.A1(new_n16859), .A2(new_n17006), .B(new_n17007), .Y(new_n17008));
  NAND2xp33_ASAP7_75t_L     g16752(.A(new_n16847), .B(new_n17008), .Y(new_n17009));
  O2A1O1Ixp33_ASAP7_75t_L   g16753(.A1(new_n16859), .A2(new_n17006), .B(new_n17007), .C(new_n16847), .Y(new_n17010));
  AO21x2_ASAP7_75t_L        g16754(.A1(new_n16847), .A2(new_n17009), .B(new_n17010), .Y(new_n17011));
  NAND2xp33_ASAP7_75t_L     g16755(.A(\b[52] ), .B(new_n2421), .Y(new_n17012));
  OAI221xp5_ASAP7_75t_L     g16756(.A1(new_n2415), .A2(new_n9683), .B1(new_n8779), .B2(new_n2572), .C(new_n17012), .Y(new_n17013));
  A2O1A1Ixp33_ASAP7_75t_L   g16757(.A1(new_n9690), .A2(new_n2417), .B(new_n17013), .C(\a[26] ), .Y(new_n17014));
  NAND2xp33_ASAP7_75t_L     g16758(.A(\a[26] ), .B(new_n17014), .Y(new_n17015));
  A2O1A1Ixp33_ASAP7_75t_L   g16759(.A1(new_n9690), .A2(new_n2417), .B(new_n17013), .C(new_n2413), .Y(new_n17016));
  NAND2xp33_ASAP7_75t_L     g16760(.A(new_n17016), .B(new_n17015), .Y(new_n17017));
  A2O1A1Ixp33_ASAP7_75t_L   g16761(.A1(new_n16716), .A2(new_n16542), .B(new_n16712), .C(new_n16544), .Y(new_n17018));
  NOR2xp33_ASAP7_75t_L      g16762(.A(new_n17017), .B(new_n17018), .Y(new_n17019));
  AOI211xp5_ASAP7_75t_L     g16763(.A1(new_n9690), .A2(new_n2417), .B(new_n17013), .C(new_n2413), .Y(new_n17020));
  A2O1A1O1Ixp25_ASAP7_75t_L g16764(.A1(new_n9690), .A2(new_n2417), .B(new_n17013), .C(new_n17014), .D(new_n17020), .Y(new_n17021));
  A2O1A1O1Ixp25_ASAP7_75t_L g16765(.A1(new_n16716), .A2(new_n16542), .B(new_n16712), .C(new_n16544), .D(new_n17021), .Y(new_n17022));
  NOR2xp33_ASAP7_75t_L      g16766(.A(new_n17022), .B(new_n17019), .Y(new_n17023));
  A2O1A1Ixp33_ASAP7_75t_L   g16767(.A1(new_n16847), .A2(new_n17009), .B(new_n17010), .C(new_n17023), .Y(new_n17024));
  NOR3xp33_ASAP7_75t_L      g16768(.A(new_n17011), .B(new_n17022), .C(new_n17019), .Y(new_n17025));
  A2O1A1Ixp33_ASAP7_75t_L   g16769(.A1(new_n17011), .A2(new_n17024), .B(new_n17025), .C(new_n16838), .Y(new_n17026));
  INVx1_ASAP7_75t_L         g16770(.A(new_n17026), .Y(new_n17027));
  AOI211xp5_ASAP7_75t_L     g16771(.A1(new_n17011), .A2(new_n17024), .B(new_n17025), .C(new_n16838), .Y(new_n17028));
  OAI211xp5_ASAP7_75t_L     g16772(.A1(new_n17027), .A2(new_n17028), .B(new_n16825), .C(new_n16827), .Y(new_n17029));
  INVx1_ASAP7_75t_L         g16773(.A(new_n16536), .Y(new_n17030));
  A2O1A1Ixp33_ASAP7_75t_L   g16774(.A1(new_n16532), .A2(new_n17030), .B(new_n16738), .C(new_n16534), .Y(new_n17031));
  AOI211xp5_ASAP7_75t_L     g16775(.A1(\a[20] ), .A2(new_n16817), .B(new_n16818), .C(new_n17031), .Y(new_n17032));
  INVx1_ASAP7_75t_L         g16776(.A(new_n17028), .Y(new_n17033));
  OAI211xp5_ASAP7_75t_L     g16777(.A1(new_n16826), .A2(new_n17032), .B(new_n17026), .C(new_n17033), .Y(new_n17034));
  NOR2xp33_ASAP7_75t_L      g16778(.A(new_n12258), .B(new_n2118), .Y(new_n17035));
  AOI221xp5_ASAP7_75t_L     g16779(.A1(\b[60] ), .A2(new_n1290), .B1(\b[62] ), .B2(new_n1209), .C(new_n17035), .Y(new_n17036));
  INVx1_ASAP7_75t_L         g16780(.A(new_n17036), .Y(new_n17037));
  A2O1A1Ixp33_ASAP7_75t_L   g16781(.A1(new_n1205), .A2(new_n1207), .B(new_n1076), .C(new_n17036), .Y(new_n17038));
  A2O1A1O1Ixp25_ASAP7_75t_L g16782(.A1(new_n12609), .A2(new_n12606), .B(new_n17037), .C(new_n17038), .D(new_n1206), .Y(new_n17039));
  O2A1O1Ixp33_ASAP7_75t_L   g16783(.A1(new_n1210), .A2(new_n12610), .B(new_n17036), .C(\a[17] ), .Y(new_n17040));
  O2A1O1Ixp33_ASAP7_75t_L   g16784(.A1(new_n16821), .A2(new_n16820), .B(new_n16822), .C(new_n16738), .Y(new_n17041));
  A2O1A1Ixp33_ASAP7_75t_L   g16785(.A1(new_n17030), .A2(new_n16822), .B(new_n17041), .C(new_n16742), .Y(new_n17042));
  INVx1_ASAP7_75t_L         g16786(.A(new_n16752), .Y(new_n17043));
  INVx1_ASAP7_75t_L         g16787(.A(new_n16748), .Y(new_n17044));
  A2O1A1Ixp33_ASAP7_75t_L   g16788(.A1(new_n16751), .A2(new_n16463), .B(new_n16458), .C(new_n17044), .Y(new_n17045));
  A2O1A1Ixp33_ASAP7_75t_L   g16789(.A1(new_n16747), .A2(new_n16746), .B(new_n17043), .C(new_n17045), .Y(new_n17046));
  NOR2xp33_ASAP7_75t_L      g16790(.A(new_n17039), .B(new_n17040), .Y(new_n17047));
  INVx1_ASAP7_75t_L         g16791(.A(new_n17047), .Y(new_n17048));
  A2O1A1Ixp33_ASAP7_75t_L   g16792(.A1(new_n17046), .A2(new_n17042), .B(new_n17043), .C(new_n17048), .Y(new_n17049));
  A2O1A1O1Ixp25_ASAP7_75t_L g16793(.A1(new_n17045), .A2(new_n17044), .B(new_n16758), .C(new_n16752), .D(new_n17048), .Y(new_n17050));
  O2A1O1Ixp33_ASAP7_75t_L   g16794(.A1(new_n17039), .A2(new_n17040), .B(new_n17049), .C(new_n17050), .Y(new_n17051));
  AND2x2_ASAP7_75t_L        g16795(.A(new_n17034), .B(new_n17029), .Y(new_n17052));
  INVx1_ASAP7_75t_L         g16796(.A(new_n17050), .Y(new_n17053));
  O2A1O1Ixp33_ASAP7_75t_L   g16797(.A1(new_n16756), .A2(new_n16748), .B(new_n17042), .C(new_n17043), .Y(new_n17054));
  NAND2xp33_ASAP7_75t_L     g16798(.A(new_n17048), .B(new_n17054), .Y(new_n17055));
  NAND3xp33_ASAP7_75t_L     g16799(.A(new_n17052), .B(new_n17055), .C(new_n17053), .Y(new_n17056));
  A2O1A1Ixp33_ASAP7_75t_L   g16800(.A1(new_n17034), .A2(new_n17029), .B(new_n17051), .C(new_n17056), .Y(new_n17057));
  O2A1O1Ixp33_ASAP7_75t_L   g16801(.A1(new_n16808), .A2(new_n16810), .B(new_n16813), .C(new_n17057), .Y(new_n17058));
  O2A1O1Ixp33_ASAP7_75t_L   g16802(.A1(new_n16772), .A2(new_n16768), .B(new_n16760), .C(new_n16770), .Y(new_n17059));
  A2O1A1O1Ixp25_ASAP7_75t_L g16803(.A1(new_n12603), .A2(new_n14444), .B(new_n872), .C(new_n980), .D(new_n12956), .Y(new_n17060));
  A2O1A1Ixp33_ASAP7_75t_L   g16804(.A1(new_n17060), .A2(new_n16806), .B(new_n16807), .C(new_n17059), .Y(new_n17061));
  A2O1A1Ixp33_ASAP7_75t_L   g16805(.A1(new_n16773), .A2(new_n16771), .B(new_n16810), .C(new_n17061), .Y(new_n17062));
  O2A1O1Ixp33_ASAP7_75t_L   g16806(.A1(new_n17052), .A2(new_n17051), .B(new_n17056), .C(new_n17062), .Y(new_n17063));
  NOR3xp33_ASAP7_75t_L      g16807(.A(new_n17063), .B(new_n17058), .C(new_n16804), .Y(new_n17064));
  INVx1_ASAP7_75t_L         g16808(.A(new_n16810), .Y(new_n17065));
  INVx1_ASAP7_75t_L         g16809(.A(new_n17049), .Y(new_n17066));
  O2A1O1Ixp33_ASAP7_75t_L   g16810(.A1(new_n17054), .A2(new_n17066), .B(new_n17055), .C(new_n17052), .Y(new_n17067));
  NAND2xp33_ASAP7_75t_L     g16811(.A(new_n17034), .B(new_n17029), .Y(new_n17068));
  O2A1O1Ixp33_ASAP7_75t_L   g16812(.A1(new_n17039), .A2(new_n17040), .B(new_n17049), .C(new_n17068), .Y(new_n17069));
  O2A1O1Ixp33_ASAP7_75t_L   g16813(.A1(new_n17066), .A2(new_n17054), .B(new_n17069), .C(new_n17067), .Y(new_n17070));
  A2O1A1Ixp33_ASAP7_75t_L   g16814(.A1(new_n17065), .A2(new_n16811), .B(new_n16812), .C(new_n17070), .Y(new_n17071));
  NAND3xp33_ASAP7_75t_L     g16815(.A(new_n17057), .B(new_n17061), .C(new_n16813), .Y(new_n17072));
  AOI21xp33_ASAP7_75t_L     g16816(.A1(new_n17071), .A2(new_n17072), .B(new_n16803), .Y(new_n17073));
  NOR2xp33_ASAP7_75t_L      g16817(.A(new_n17073), .B(new_n17064), .Y(new_n17074));
  INVx1_ASAP7_75t_L         g16818(.A(new_n17074), .Y(new_n17075));
  A2O1A1O1Ixp25_ASAP7_75t_L g16819(.A1(new_n16790), .A2(new_n16520), .B(new_n16794), .C(new_n16792), .D(new_n17075), .Y(new_n17076));
  A2O1A1Ixp33_ASAP7_75t_L   g16820(.A1(new_n16790), .A2(new_n16520), .B(new_n16794), .C(new_n16792), .Y(new_n17077));
  NOR2xp33_ASAP7_75t_L      g16821(.A(new_n17074), .B(new_n17077), .Y(new_n17078));
  NOR2xp33_ASAP7_75t_L      g16822(.A(new_n17078), .B(new_n17076), .Y(\f[77] ));
  OAI22xp33_ASAP7_75t_L     g16823(.A1(new_n1285), .A2(new_n12258), .B1(new_n12603), .B2(new_n2118), .Y(new_n17080));
  AOI221xp5_ASAP7_75t_L     g16824(.A1(new_n1209), .A2(\b[63] ), .B1(new_n1216), .B2(new_n12961), .C(new_n17080), .Y(new_n17081));
  XNOR2x2_ASAP7_75t_L       g16825(.A(new_n1206), .B(new_n17081), .Y(new_n17082));
  INVx1_ASAP7_75t_L         g16826(.A(new_n17082), .Y(new_n17083));
  A2O1A1O1Ixp25_ASAP7_75t_L g16827(.A1(new_n17034), .A2(new_n17029), .B(new_n17051), .C(new_n17049), .D(new_n17083), .Y(new_n17084));
  INVx1_ASAP7_75t_L         g16828(.A(new_n17084), .Y(new_n17085));
  O2A1O1Ixp33_ASAP7_75t_L   g16829(.A1(new_n17050), .A2(new_n17048), .B(new_n17068), .C(new_n17066), .Y(new_n17086));
  NAND2xp33_ASAP7_75t_L     g16830(.A(new_n17083), .B(new_n17086), .Y(new_n17087));
  OAI22xp33_ASAP7_75t_L     g16831(.A1(new_n1654), .A2(new_n11303), .B1(new_n11591), .B2(new_n1517), .Y(new_n17088));
  AOI221xp5_ASAP7_75t_L     g16832(.A1(new_n1511), .A2(\b[60] ), .B1(new_n1513), .B2(new_n13839), .C(new_n17088), .Y(new_n17089));
  XNOR2x2_ASAP7_75t_L       g16833(.A(new_n1501), .B(new_n17089), .Y(new_n17090));
  INVx1_ASAP7_75t_L         g16834(.A(new_n17090), .Y(new_n17091));
  AOI31xp33_ASAP7_75t_L     g16835(.A1(new_n16825), .A2(new_n17033), .A3(new_n17026), .B(new_n16826), .Y(new_n17092));
  XNOR2x2_ASAP7_75t_L       g16836(.A(new_n17091), .B(new_n17092), .Y(new_n17093));
  INVx1_ASAP7_75t_L         g16837(.A(new_n16837), .Y(new_n17094));
  A2O1A1O1Ixp25_ASAP7_75t_L g16838(.A1(new_n17009), .A2(new_n16847), .B(new_n17010), .C(new_n17024), .D(new_n17025), .Y(new_n17095));
  INVx1_ASAP7_75t_L         g16839(.A(new_n10991), .Y(new_n17096));
  NOR2xp33_ASAP7_75t_L      g16840(.A(new_n10332), .B(new_n1962), .Y(new_n17097));
  AOI221xp5_ASAP7_75t_L     g16841(.A1(new_n1955), .A2(\b[57] ), .B1(new_n2093), .B2(\b[55] ), .C(new_n17097), .Y(new_n17098));
  O2A1O1Ixp33_ASAP7_75t_L   g16842(.A1(new_n1956), .A2(new_n17096), .B(new_n17098), .C(new_n1952), .Y(new_n17099));
  INVx1_ASAP7_75t_L         g16843(.A(new_n17099), .Y(new_n17100));
  O2A1O1Ixp33_ASAP7_75t_L   g16844(.A1(new_n1956), .A2(new_n17096), .B(new_n17098), .C(\a[23] ), .Y(new_n17101));
  AOI21xp33_ASAP7_75t_L     g16845(.A1(new_n17100), .A2(\a[23] ), .B(new_n17101), .Y(new_n17102));
  INVx1_ASAP7_75t_L         g16846(.A(new_n17102), .Y(new_n17103));
  O2A1O1Ixp33_ASAP7_75t_L   g16847(.A1(new_n16836), .A2(new_n17095), .B(new_n17094), .C(new_n17103), .Y(new_n17104));
  INVx1_ASAP7_75t_L         g16848(.A(new_n17104), .Y(new_n17105));
  A2O1A1O1Ixp25_ASAP7_75t_L g16849(.A1(new_n17024), .A2(new_n17011), .B(new_n17025), .C(new_n16838), .D(new_n16837), .Y(new_n17106));
  A2O1A1Ixp33_ASAP7_75t_L   g16850(.A1(\a[23] ), .A2(new_n17100), .B(new_n17101), .C(new_n17106), .Y(new_n17107));
  NAND2xp33_ASAP7_75t_L     g16851(.A(new_n17107), .B(new_n17105), .Y(new_n17108));
  OAI22xp33_ASAP7_75t_L     g16852(.A1(new_n2572), .A2(new_n9355), .B1(new_n9683), .B2(new_n2410), .Y(new_n17109));
  AOI221xp5_ASAP7_75t_L     g16853(.A1(new_n2423), .A2(\b[54] ), .B1(new_n2417), .B2(new_n9717), .C(new_n17109), .Y(new_n17110));
  XNOR2x2_ASAP7_75t_L       g16854(.A(new_n2413), .B(new_n17110), .Y(new_n17111));
  A2O1A1O1Ixp25_ASAP7_75t_L g16855(.A1(new_n17009), .A2(new_n16847), .B(new_n17010), .C(new_n17023), .D(new_n17022), .Y(new_n17112));
  NAND2xp33_ASAP7_75t_L     g16856(.A(new_n17111), .B(new_n17112), .Y(new_n17113));
  INVx1_ASAP7_75t_L         g16857(.A(new_n17111), .Y(new_n17114));
  A2O1A1Ixp33_ASAP7_75t_L   g16858(.A1(new_n17011), .A2(new_n17023), .B(new_n17022), .C(new_n17114), .Y(new_n17115));
  OAI22xp33_ASAP7_75t_L     g16859(.A1(new_n3133), .A2(new_n8427), .B1(new_n8755), .B2(new_n2925), .Y(new_n17116));
  AOI221xp5_ASAP7_75t_L     g16860(.A1(new_n2938), .A2(\b[51] ), .B1(new_n2932), .B2(new_n8790), .C(new_n17116), .Y(new_n17117));
  XNOR2x2_ASAP7_75t_L       g16861(.A(new_n2928), .B(new_n17117), .Y(new_n17118));
  AOI21xp33_ASAP7_75t_L     g16862(.A1(new_n17008), .A2(new_n16847), .B(new_n16845), .Y(new_n17119));
  NAND2xp33_ASAP7_75t_L     g16863(.A(new_n17118), .B(new_n17119), .Y(new_n17120));
  OR2x4_ASAP7_75t_L         g16864(.A(new_n17118), .B(new_n17119), .Y(new_n17121));
  NOR2xp33_ASAP7_75t_L      g16865(.A(new_n16866), .B(new_n16988), .Y(new_n17122));
  A2O1A1O1Ixp25_ASAP7_75t_L g16866(.A1(new_n16864), .A2(\a[38] ), .B(new_n16865), .C(new_n16989), .D(new_n17122), .Y(new_n17123));
  A2O1A1O1Ixp25_ASAP7_75t_L g16867(.A1(new_n16659), .A2(new_n16650), .B(new_n16571), .C(new_n16652), .D(new_n16955), .Y(new_n17124));
  A2O1A1O1Ixp25_ASAP7_75t_L g16868(.A1(new_n16965), .A2(\a[44] ), .B(new_n16962), .C(new_n16956), .D(new_n17124), .Y(new_n17125));
  INVx1_ASAP7_75t_L         g16869(.A(new_n16942), .Y(new_n17126));
  A2O1A1Ixp33_ASAP7_75t_L   g16870(.A1(new_n16937), .A2(new_n16931), .B(new_n16939), .C(new_n17126), .Y(new_n17127));
  A2O1A1Ixp33_ASAP7_75t_L   g16871(.A1(new_n17127), .A2(new_n17126), .B(new_n16950), .C(new_n16943), .Y(new_n17128));
  NOR2xp33_ASAP7_75t_L      g16872(.A(new_n2703), .B(new_n10400), .Y(new_n17129));
  AOI221xp5_ASAP7_75t_L     g16873(.A1(new_n9102), .A2(\b[27] ), .B1(new_n10398), .B2(\b[25] ), .C(new_n17129), .Y(new_n17130));
  INVx1_ASAP7_75t_L         g16874(.A(new_n17130), .Y(new_n17131));
  A2O1A1Ixp33_ASAP7_75t_L   g16875(.A1(new_n2887), .A2(new_n9437), .B(new_n17131), .C(\a[53] ), .Y(new_n17132));
  O2A1O1Ixp33_ASAP7_75t_L   g16876(.A1(new_n9104), .A2(new_n2889), .B(new_n17130), .C(\a[53] ), .Y(new_n17133));
  NOR2xp33_ASAP7_75t_L      g16877(.A(new_n960), .B(new_n13030), .Y(new_n17134));
  INVx1_ASAP7_75t_L         g16878(.A(new_n17134), .Y(new_n17135));
  O2A1O1Ixp33_ASAP7_75t_L   g16879(.A1(new_n1043), .A2(new_n12672), .B(new_n17135), .C(\a[14] ), .Y(new_n17136));
  O2A1O1Ixp33_ASAP7_75t_L   g16880(.A1(new_n1043), .A2(new_n12672), .B(new_n17135), .C(new_n867), .Y(new_n17137));
  INVx1_ASAP7_75t_L         g16881(.A(new_n17137), .Y(new_n17138));
  O2A1O1Ixp33_ASAP7_75t_L   g16882(.A1(\a[14] ), .A2(new_n17136), .B(new_n17138), .C(new_n16588), .Y(new_n17139));
  INVx1_ASAP7_75t_L         g16883(.A(new_n17139), .Y(new_n17140));
  O2A1O1Ixp33_ASAP7_75t_L   g16884(.A1(\a[14] ), .A2(new_n17136), .B(new_n17138), .C(new_n16589), .Y(new_n17141));
  A2O1A1O1Ixp25_ASAP7_75t_L g16885(.A1(new_n13028), .A2(\b[13] ), .B(new_n16587), .C(new_n17140), .D(new_n17141), .Y(new_n17142));
  NOR2xp33_ASAP7_75t_L      g16886(.A(new_n1349), .B(new_n12318), .Y(new_n17143));
  AOI221xp5_ASAP7_75t_L     g16887(.A1(new_n11995), .A2(\b[18] ), .B1(new_n13314), .B2(\b[16] ), .C(new_n17143), .Y(new_n17144));
  O2A1O1Ixp33_ASAP7_75t_L   g16888(.A1(new_n11998), .A2(new_n1464), .B(new_n17144), .C(new_n11987), .Y(new_n17145));
  O2A1O1Ixp33_ASAP7_75t_L   g16889(.A1(new_n11998), .A2(new_n1464), .B(new_n17144), .C(\a[62] ), .Y(new_n17146));
  INVx1_ASAP7_75t_L         g16890(.A(new_n17146), .Y(new_n17147));
  O2A1O1Ixp33_ASAP7_75t_L   g16891(.A1(new_n17145), .A2(new_n11987), .B(new_n17147), .C(new_n17142), .Y(new_n17148));
  INVx1_ASAP7_75t_L         g16892(.A(new_n17148), .Y(new_n17149));
  INVx1_ASAP7_75t_L         g16893(.A(new_n17142), .Y(new_n17150));
  O2A1O1Ixp33_ASAP7_75t_L   g16894(.A1(new_n17145), .A2(new_n11987), .B(new_n17147), .C(new_n17150), .Y(new_n17151));
  A2O1A1O1Ixp25_ASAP7_75t_L g16895(.A1(new_n17140), .A2(new_n16589), .B(new_n17141), .C(new_n17149), .D(new_n17151), .Y(new_n17152));
  A2O1A1O1Ixp25_ASAP7_75t_L g16896(.A1(new_n13028), .A2(\b[14] ), .B(new_n16877), .C(new_n16588), .D(new_n16889), .Y(new_n17153));
  NAND2xp33_ASAP7_75t_L     g16897(.A(new_n17153), .B(new_n17152), .Y(new_n17154));
  INVx1_ASAP7_75t_L         g16898(.A(new_n17153), .Y(new_n17155));
  A2O1A1Ixp33_ASAP7_75t_L   g16899(.A1(new_n17149), .A2(new_n17150), .B(new_n17151), .C(new_n17155), .Y(new_n17156));
  NAND2xp33_ASAP7_75t_L     g16900(.A(new_n17156), .B(new_n17154), .Y(new_n17157));
  NOR2xp33_ASAP7_75t_L      g16901(.A(new_n1599), .B(new_n11354), .Y(new_n17158));
  AOI221xp5_ASAP7_75t_L     g16902(.A1(\b[21] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[20] ), .C(new_n17158), .Y(new_n17159));
  INVx1_ASAP7_75t_L         g16903(.A(new_n17159), .Y(new_n17160));
  A2O1A1Ixp33_ASAP7_75t_L   g16904(.A1(new_n2836), .A2(new_n11351), .B(new_n17160), .C(\a[59] ), .Y(new_n17161));
  A2O1A1Ixp33_ASAP7_75t_L   g16905(.A1(new_n2836), .A2(new_n11351), .B(new_n17160), .C(new_n11048), .Y(new_n17162));
  INVx1_ASAP7_75t_L         g16906(.A(new_n17162), .Y(new_n17163));
  AO21x2_ASAP7_75t_L        g16907(.A1(\a[59] ), .A2(new_n17161), .B(new_n17163), .Y(new_n17164));
  NAND3xp33_ASAP7_75t_L     g16908(.A(new_n17164), .B(new_n17156), .C(new_n17154), .Y(new_n17165));
  INVx1_ASAP7_75t_L         g16909(.A(new_n17165), .Y(new_n17166));
  A2O1A1Ixp33_ASAP7_75t_L   g16910(.A1(\a[59] ), .A2(new_n17161), .B(new_n17163), .C(new_n17157), .Y(new_n17167));
  OAI21xp33_ASAP7_75t_L     g16911(.A1(new_n17157), .A2(new_n17166), .B(new_n17167), .Y(new_n17168));
  NAND3xp33_ASAP7_75t_L     g16912(.A(new_n16892), .B(new_n16876), .C(new_n16591), .Y(new_n17169));
  A2O1A1O1Ixp25_ASAP7_75t_L g16913(.A1(\a[59] ), .A2(new_n16900), .B(new_n16901), .C(new_n17169), .D(new_n16893), .Y(new_n17170));
  XOR2x2_ASAP7_75t_L        g16914(.A(new_n17170), .B(new_n17168), .Y(new_n17171));
  NOR2xp33_ASAP7_75t_L      g16915(.A(new_n2188), .B(new_n10388), .Y(new_n17172));
  AOI221xp5_ASAP7_75t_L     g16916(.A1(new_n10086), .A2(\b[24] ), .B1(new_n11361), .B2(\b[22] ), .C(new_n17172), .Y(new_n17173));
  O2A1O1Ixp33_ASAP7_75t_L   g16917(.A1(new_n10088), .A2(new_n2853), .B(new_n17173), .C(new_n10083), .Y(new_n17174));
  O2A1O1Ixp33_ASAP7_75t_L   g16918(.A1(new_n10088), .A2(new_n2853), .B(new_n17173), .C(\a[56] ), .Y(new_n17175));
  INVx1_ASAP7_75t_L         g16919(.A(new_n17175), .Y(new_n17176));
  OAI211xp5_ASAP7_75t_L     g16920(.A1(new_n10083), .A2(new_n17174), .B(new_n17171), .C(new_n17176), .Y(new_n17177));
  INVx1_ASAP7_75t_L         g16921(.A(new_n16909), .Y(new_n17178));
  A2O1A1O1Ixp25_ASAP7_75t_L g16922(.A1(new_n16918), .A2(\a[56] ), .B(new_n16915), .C(new_n16907), .D(new_n17178), .Y(new_n17179));
  O2A1O1Ixp33_ASAP7_75t_L   g16923(.A1(new_n17174), .A2(new_n10083), .B(new_n17176), .C(new_n17171), .Y(new_n17180));
  INVx1_ASAP7_75t_L         g16924(.A(new_n17180), .Y(new_n17181));
  AOI21xp33_ASAP7_75t_L     g16925(.A1(new_n17181), .A2(new_n17177), .B(new_n17179), .Y(new_n17182));
  INVx1_ASAP7_75t_L         g16926(.A(new_n16919), .Y(new_n17183));
  O2A1O1Ixp33_ASAP7_75t_L   g16927(.A1(new_n17183), .A2(new_n17178), .B(new_n17177), .C(new_n17180), .Y(new_n17184));
  AO21x2_ASAP7_75t_L        g16928(.A1(\a[53] ), .A2(new_n17132), .B(new_n17133), .Y(new_n17185));
  A2O1A1Ixp33_ASAP7_75t_L   g16929(.A1(new_n17184), .A2(new_n17177), .B(new_n17182), .C(new_n17185), .Y(new_n17186));
  A2O1A1Ixp33_ASAP7_75t_L   g16930(.A1(new_n17184), .A2(new_n17177), .B(new_n17182), .C(new_n17186), .Y(new_n17187));
  INVx1_ASAP7_75t_L         g16931(.A(new_n17187), .Y(new_n17188));
  A2O1A1O1Ixp25_ASAP7_75t_L g16932(.A1(new_n17132), .A2(\a[53] ), .B(new_n17133), .C(new_n17186), .D(new_n17188), .Y(new_n17189));
  A2O1A1O1Ixp25_ASAP7_75t_L g16933(.A1(new_n16873), .A2(\a[53] ), .B(new_n16874), .C(new_n16924), .D(new_n16921), .Y(new_n17190));
  NAND2xp33_ASAP7_75t_L     g16934(.A(new_n17190), .B(new_n17189), .Y(new_n17191));
  INVx1_ASAP7_75t_L         g16935(.A(new_n17190), .Y(new_n17192));
  A2O1A1Ixp33_ASAP7_75t_L   g16936(.A1(new_n17186), .A2(new_n17185), .B(new_n17188), .C(new_n17192), .Y(new_n17193));
  NAND2xp33_ASAP7_75t_L     g16937(.A(new_n17193), .B(new_n17191), .Y(new_n17194));
  INVx1_ASAP7_75t_L         g16938(.A(new_n17194), .Y(new_n17195));
  NOR2xp33_ASAP7_75t_L      g16939(.A(new_n3098), .B(new_n10065), .Y(new_n17196));
  AOI221xp5_ASAP7_75t_L     g16940(.A1(new_n8175), .A2(\b[30] ), .B1(new_n8484), .B2(\b[28] ), .C(new_n17196), .Y(new_n17197));
  O2A1O1Ixp33_ASAP7_75t_L   g16941(.A1(new_n8176), .A2(new_n3464), .B(new_n17197), .C(new_n8172), .Y(new_n17198));
  O2A1O1Ixp33_ASAP7_75t_L   g16942(.A1(new_n8176), .A2(new_n3464), .B(new_n17197), .C(\a[50] ), .Y(new_n17199));
  INVx1_ASAP7_75t_L         g16943(.A(new_n17199), .Y(new_n17200));
  O2A1O1Ixp33_ASAP7_75t_L   g16944(.A1(new_n17198), .A2(new_n8172), .B(new_n17200), .C(new_n17194), .Y(new_n17201));
  INVx1_ASAP7_75t_L         g16945(.A(new_n17201), .Y(new_n17202));
  INVx1_ASAP7_75t_L         g16946(.A(new_n17198), .Y(new_n17203));
  A2O1A1Ixp33_ASAP7_75t_L   g16947(.A1(\a[50] ), .A2(new_n17203), .B(new_n17199), .C(new_n17194), .Y(new_n17204));
  INVx1_ASAP7_75t_L         g16948(.A(new_n17204), .Y(new_n17205));
  A2O1A1Ixp33_ASAP7_75t_L   g16949(.A1(new_n16634), .A2(new_n16631), .B(new_n16929), .C(new_n16937), .Y(new_n17206));
  AOI211xp5_ASAP7_75t_L     g16950(.A1(new_n17202), .A2(new_n17195), .B(new_n17205), .C(new_n17206), .Y(new_n17207));
  INVx1_ASAP7_75t_L         g16951(.A(new_n17206), .Y(new_n17208));
  O2A1O1Ixp33_ASAP7_75t_L   g16952(.A1(new_n17194), .A2(new_n17201), .B(new_n17204), .C(new_n17208), .Y(new_n17209));
  NOR2xp33_ASAP7_75t_L      g16953(.A(new_n17207), .B(new_n17209), .Y(new_n17210));
  NOR2xp33_ASAP7_75t_L      g16954(.A(new_n3891), .B(new_n7312), .Y(new_n17211));
  AOI221xp5_ASAP7_75t_L     g16955(.A1(\b[31] ), .A2(new_n7609), .B1(\b[33] ), .B2(new_n7334), .C(new_n17211), .Y(new_n17212));
  O2A1O1Ixp33_ASAP7_75t_L   g16956(.A1(new_n7321), .A2(new_n4108), .B(new_n17212), .C(new_n7316), .Y(new_n17213));
  INVx1_ASAP7_75t_L         g16957(.A(new_n17213), .Y(new_n17214));
  O2A1O1Ixp33_ASAP7_75t_L   g16958(.A1(new_n7321), .A2(new_n4108), .B(new_n17212), .C(\a[47] ), .Y(new_n17215));
  A2O1A1Ixp33_ASAP7_75t_L   g16959(.A1(\a[47] ), .A2(new_n17214), .B(new_n17215), .C(new_n17210), .Y(new_n17216));
  INVx1_ASAP7_75t_L         g16960(.A(new_n17215), .Y(new_n17217));
  O2A1O1Ixp33_ASAP7_75t_L   g16961(.A1(new_n17213), .A2(new_n7316), .B(new_n17217), .C(new_n17210), .Y(new_n17218));
  AOI21xp33_ASAP7_75t_L     g16962(.A1(new_n17216), .A2(new_n17210), .B(new_n17218), .Y(new_n17219));
  XOR2x2_ASAP7_75t_L        g16963(.A(new_n17128), .B(new_n17219), .Y(new_n17220));
  NOR2xp33_ASAP7_75t_L      g16964(.A(new_n4344), .B(new_n6741), .Y(new_n17221));
  AOI221xp5_ASAP7_75t_L     g16965(.A1(\b[36] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[35] ), .C(new_n17221), .Y(new_n17222));
  O2A1O1Ixp33_ASAP7_75t_L   g16966(.A1(new_n6443), .A2(new_n4622), .B(new_n17222), .C(new_n6439), .Y(new_n17223));
  O2A1O1Ixp33_ASAP7_75t_L   g16967(.A1(new_n6443), .A2(new_n4622), .B(new_n17222), .C(\a[44] ), .Y(new_n17224));
  INVx1_ASAP7_75t_L         g16968(.A(new_n17224), .Y(new_n17225));
  OAI21xp33_ASAP7_75t_L     g16969(.A1(new_n6439), .A2(new_n17223), .B(new_n17225), .Y(new_n17226));
  XOR2x2_ASAP7_75t_L        g16970(.A(new_n17226), .B(new_n17220), .Y(new_n17227));
  XNOR2x2_ASAP7_75t_L       g16971(.A(new_n17125), .B(new_n17227), .Y(new_n17228));
  INVx1_ASAP7_75t_L         g16972(.A(new_n17228), .Y(new_n17229));
  NOR2xp33_ASAP7_75t_L      g16973(.A(new_n5570), .B(new_n5641), .Y(new_n17230));
  AOI221xp5_ASAP7_75t_L     g16974(.A1(\b[37] ), .A2(new_n5920), .B1(\b[38] ), .B2(new_n5623), .C(new_n17230), .Y(new_n17231));
  O2A1O1Ixp33_ASAP7_75t_L   g16975(.A1(new_n5630), .A2(new_n5578), .B(new_n17231), .C(new_n5626), .Y(new_n17232));
  O2A1O1Ixp33_ASAP7_75t_L   g16976(.A1(new_n5630), .A2(new_n5578), .B(new_n17231), .C(\a[41] ), .Y(new_n17233));
  INVx1_ASAP7_75t_L         g16977(.A(new_n17233), .Y(new_n17234));
  O2A1O1Ixp33_ASAP7_75t_L   g16978(.A1(new_n17232), .A2(new_n5626), .B(new_n17234), .C(new_n17228), .Y(new_n17235));
  INVx1_ASAP7_75t_L         g16979(.A(new_n17235), .Y(new_n17236));
  O2A1O1Ixp33_ASAP7_75t_L   g16980(.A1(new_n17232), .A2(new_n5626), .B(new_n17234), .C(new_n17229), .Y(new_n17237));
  AOI21xp33_ASAP7_75t_L     g16981(.A1(new_n17236), .A2(new_n17229), .B(new_n17237), .Y(new_n17238));
  A2O1A1Ixp33_ASAP7_75t_L   g16982(.A1(new_n16979), .A2(new_n16970), .B(new_n16971), .C(new_n17238), .Y(new_n17239));
  A2O1A1O1Ixp25_ASAP7_75t_L g16983(.A1(new_n16986), .A2(\a[41] ), .B(new_n16977), .C(new_n16970), .D(new_n16971), .Y(new_n17240));
  A2O1A1Ixp33_ASAP7_75t_L   g16984(.A1(new_n17236), .A2(new_n17229), .B(new_n17237), .C(new_n17240), .Y(new_n17241));
  NAND2xp33_ASAP7_75t_L     g16985(.A(new_n17241), .B(new_n17239), .Y(new_n17242));
  NOR2xp33_ASAP7_75t_L      g16986(.A(new_n6378), .B(new_n4908), .Y(new_n17243));
  AOI221xp5_ASAP7_75t_L     g16987(.A1(\b[40] ), .A2(new_n5139), .B1(\b[41] ), .B2(new_n4916), .C(new_n17243), .Y(new_n17244));
  O2A1O1Ixp33_ASAP7_75t_L   g16988(.A1(new_n4911), .A2(new_n6386), .B(new_n17244), .C(new_n4906), .Y(new_n17245));
  INVx1_ASAP7_75t_L         g16989(.A(new_n17245), .Y(new_n17246));
  O2A1O1Ixp33_ASAP7_75t_L   g16990(.A1(new_n4911), .A2(new_n6386), .B(new_n17244), .C(\a[38] ), .Y(new_n17247));
  A2O1A1Ixp33_ASAP7_75t_L   g16991(.A1(\a[38] ), .A2(new_n17246), .B(new_n17247), .C(new_n17242), .Y(new_n17248));
  INVx1_ASAP7_75t_L         g16992(.A(new_n17242), .Y(new_n17249));
  AOI21xp33_ASAP7_75t_L     g16993(.A1(new_n17246), .A2(\a[38] ), .B(new_n17247), .Y(new_n17250));
  NAND2xp33_ASAP7_75t_L     g16994(.A(new_n17250), .B(new_n17249), .Y(new_n17251));
  NAND2xp33_ASAP7_75t_L     g16995(.A(new_n17248), .B(new_n17251), .Y(new_n17252));
  NAND2xp33_ASAP7_75t_L     g16996(.A(new_n17123), .B(new_n17252), .Y(new_n17253));
  INVx1_ASAP7_75t_L         g16997(.A(new_n16991), .Y(new_n17254));
  XNOR2x2_ASAP7_75t_L       g16998(.A(new_n17250), .B(new_n17242), .Y(new_n17255));
  A2O1A1Ixp33_ASAP7_75t_L   g16999(.A1(new_n16983), .A2(new_n16867), .B(new_n17254), .C(new_n17255), .Y(new_n17256));
  NAND2xp33_ASAP7_75t_L     g17000(.A(new_n17256), .B(new_n17253), .Y(new_n17257));
  NOR2xp33_ASAP7_75t_L      g17001(.A(new_n7249), .B(new_n4147), .Y(new_n17258));
  AOI221xp5_ASAP7_75t_L     g17002(.A1(\b[43] ), .A2(new_n4402), .B1(\b[44] ), .B2(new_n4155), .C(new_n17258), .Y(new_n17259));
  O2A1O1Ixp33_ASAP7_75t_L   g17003(.A1(new_n4150), .A2(new_n7255), .B(new_n17259), .C(new_n4145), .Y(new_n17260));
  O2A1O1Ixp33_ASAP7_75t_L   g17004(.A1(new_n4150), .A2(new_n7255), .B(new_n17259), .C(\a[35] ), .Y(new_n17261));
  INVx1_ASAP7_75t_L         g17005(.A(new_n17261), .Y(new_n17262));
  O2A1O1Ixp33_ASAP7_75t_L   g17006(.A1(new_n17260), .A2(new_n4145), .B(new_n17262), .C(new_n17257), .Y(new_n17263));
  INVx1_ASAP7_75t_L         g17007(.A(new_n17260), .Y(new_n17264));
  A2O1A1Ixp33_ASAP7_75t_L   g17008(.A1(\a[35] ), .A2(new_n17264), .B(new_n17261), .C(new_n17257), .Y(new_n17265));
  A2O1A1O1Ixp25_ASAP7_75t_L g17009(.A1(new_n16679), .A2(new_n16553), .B(new_n16551), .C(new_n16677), .D(new_n16995), .Y(new_n17266));
  A2O1A1O1Ixp25_ASAP7_75t_L g17010(.A1(new_n17000), .A2(\a[35] ), .B(new_n17001), .C(new_n16996), .D(new_n17266), .Y(new_n17267));
  OAI211xp5_ASAP7_75t_L     g17011(.A1(new_n17257), .A2(new_n17263), .B(new_n17267), .C(new_n17265), .Y(new_n17268));
  O2A1O1Ixp33_ASAP7_75t_L   g17012(.A1(new_n17257), .A2(new_n17263), .B(new_n17265), .C(new_n17267), .Y(new_n17269));
  INVx1_ASAP7_75t_L         g17013(.A(new_n17269), .Y(new_n17270));
  NAND2xp33_ASAP7_75t_L     g17014(.A(new_n17268), .B(new_n17270), .Y(new_n17271));
  A2O1A1O1Ixp25_ASAP7_75t_L g17015(.A1(new_n16996), .A2(new_n17002), .B(new_n17004), .C(new_n16858), .D(new_n16856), .Y(new_n17272));
  NOR2xp33_ASAP7_75t_L      g17016(.A(new_n7860), .B(new_n3510), .Y(new_n17273));
  AOI221xp5_ASAP7_75t_L     g17017(.A1(\b[46] ), .A2(new_n3708), .B1(\b[47] ), .B2(new_n3499), .C(new_n17273), .Y(new_n17274));
  O2A1O1Ixp33_ASAP7_75t_L   g17018(.A1(new_n3513), .A2(new_n7868), .B(new_n17274), .C(new_n3493), .Y(new_n17275));
  O2A1O1Ixp33_ASAP7_75t_L   g17019(.A1(new_n3513), .A2(new_n7868), .B(new_n17274), .C(\a[32] ), .Y(new_n17276));
  INVx1_ASAP7_75t_L         g17020(.A(new_n17276), .Y(new_n17277));
  O2A1O1Ixp33_ASAP7_75t_L   g17021(.A1(new_n17275), .A2(new_n3493), .B(new_n17277), .C(new_n17272), .Y(new_n17278));
  INVx1_ASAP7_75t_L         g17022(.A(new_n17275), .Y(new_n17279));
  A2O1A1Ixp33_ASAP7_75t_L   g17023(.A1(\a[32] ), .A2(new_n17279), .B(new_n17276), .C(new_n17272), .Y(new_n17280));
  O2A1O1Ixp33_ASAP7_75t_L   g17024(.A1(new_n17272), .A2(new_n17278), .B(new_n17280), .C(new_n17271), .Y(new_n17281));
  AOI21xp33_ASAP7_75t_L     g17025(.A1(new_n17279), .A2(\a[32] ), .B(new_n17276), .Y(new_n17282));
  A2O1A1Ixp33_ASAP7_75t_L   g17026(.A1(new_n17005), .A2(new_n16858), .B(new_n16856), .C(new_n17282), .Y(new_n17283));
  NAND3xp33_ASAP7_75t_L     g17027(.A(new_n17271), .B(new_n17283), .C(new_n17280), .Y(new_n17284));
  INVx1_ASAP7_75t_L         g17028(.A(new_n17284), .Y(new_n17285));
  OA211x2_ASAP7_75t_L       g17029(.A1(new_n17281), .A2(new_n17285), .B(new_n17121), .C(new_n17120), .Y(new_n17286));
  AOI211xp5_ASAP7_75t_L     g17030(.A1(new_n17121), .A2(new_n17120), .B(new_n17281), .C(new_n17285), .Y(new_n17287));
  OR2x4_ASAP7_75t_L         g17031(.A(new_n17287), .B(new_n17286), .Y(new_n17288));
  NAND3xp33_ASAP7_75t_L     g17032(.A(new_n17288), .B(new_n17115), .C(new_n17113), .Y(new_n17289));
  AOI21xp33_ASAP7_75t_L     g17033(.A1(new_n17113), .A2(new_n17115), .B(new_n17288), .Y(new_n17290));
  INVx1_ASAP7_75t_L         g17034(.A(new_n17290), .Y(new_n17291));
  NAND3xp33_ASAP7_75t_L     g17035(.A(new_n17108), .B(new_n17291), .C(new_n17289), .Y(new_n17292));
  AND3x1_ASAP7_75t_L        g17036(.A(new_n17288), .B(new_n17115), .C(new_n17113), .Y(new_n17293));
  NOR3xp33_ASAP7_75t_L      g17037(.A(new_n17108), .B(new_n17293), .C(new_n17290), .Y(new_n17294));
  A2O1A1Ixp33_ASAP7_75t_L   g17038(.A1(new_n17108), .A2(new_n17292), .B(new_n17294), .C(new_n17093), .Y(new_n17295));
  XNOR2x2_ASAP7_75t_L       g17039(.A(new_n17090), .B(new_n17092), .Y(new_n17296));
  A2O1A1Ixp33_ASAP7_75t_L   g17040(.A1(new_n17113), .A2(new_n17115), .B(new_n17288), .C(new_n17108), .Y(new_n17297));
  O2A1O1Ixp33_ASAP7_75t_L   g17041(.A1(new_n17293), .A2(new_n17297), .B(new_n17108), .C(new_n17294), .Y(new_n17298));
  NAND2xp33_ASAP7_75t_L     g17042(.A(new_n17296), .B(new_n17298), .Y(new_n17299));
  AOI22xp33_ASAP7_75t_L     g17043(.A1(new_n17085), .A2(new_n17087), .B1(new_n17295), .B2(new_n17299), .Y(new_n17300));
  A2O1A1Ixp33_ASAP7_75t_L   g17044(.A1(new_n17029), .A2(new_n17034), .B(new_n17051), .C(new_n17049), .Y(new_n17301));
  NOR2xp33_ASAP7_75t_L      g17045(.A(new_n17082), .B(new_n17301), .Y(new_n17302));
  AOI211xp5_ASAP7_75t_L     g17046(.A1(new_n17107), .A2(new_n17105), .B(new_n17290), .C(new_n17293), .Y(new_n17303));
  NAND4xp25_ASAP7_75t_L     g17047(.A(new_n17291), .B(new_n17105), .C(new_n17107), .D(new_n17289), .Y(new_n17304));
  A2O1A1O1Ixp25_ASAP7_75t_L g17048(.A1(new_n17107), .A2(new_n17105), .B(new_n17303), .C(new_n17304), .D(new_n17296), .Y(new_n17305));
  A2O1A1Ixp33_ASAP7_75t_L   g17049(.A1(new_n17107), .A2(new_n17105), .B(new_n17303), .C(new_n17304), .Y(new_n17306));
  NOR2xp33_ASAP7_75t_L      g17050(.A(new_n17093), .B(new_n17306), .Y(new_n17307));
  NOR4xp25_ASAP7_75t_L      g17051(.A(new_n17302), .B(new_n17305), .C(new_n17307), .D(new_n17084), .Y(new_n17308));
  A2O1A1Ixp33_ASAP7_75t_L   g17052(.A1(new_n16808), .A2(new_n16813), .B(new_n17057), .C(new_n17065), .Y(new_n17309));
  NOR3xp33_ASAP7_75t_L      g17053(.A(new_n17300), .B(new_n17308), .C(new_n17309), .Y(new_n17310));
  A2O1A1O1Ixp25_ASAP7_75t_L g17054(.A1(new_n17034), .A2(new_n17029), .B(new_n17051), .C(new_n17049), .D(new_n17082), .Y(new_n17311));
  INVx1_ASAP7_75t_L         g17055(.A(new_n17311), .Y(new_n17312));
  O2A1O1Ixp33_ASAP7_75t_L   g17056(.A1(new_n17066), .A2(new_n17067), .B(new_n17312), .C(new_n17302), .Y(new_n17313));
  O2A1O1Ixp33_ASAP7_75t_L   g17057(.A1(new_n17086), .A2(new_n17311), .B(new_n17087), .C(new_n17307), .Y(new_n17314));
  NAND4xp25_ASAP7_75t_L     g17058(.A(new_n17299), .B(new_n17085), .C(new_n17087), .D(new_n17295), .Y(new_n17315));
  O2A1O1Ixp33_ASAP7_75t_L   g17059(.A1(new_n16812), .A2(new_n16811), .B(new_n17070), .C(new_n16810), .Y(new_n17316));
  A2O1A1O1Ixp25_ASAP7_75t_L g17060(.A1(new_n17295), .A2(new_n17314), .B(new_n17313), .C(new_n17315), .D(new_n17316), .Y(new_n17317));
  NOR2xp33_ASAP7_75t_L      g17061(.A(new_n17310), .B(new_n17317), .Y(new_n17318));
  A2O1A1Ixp33_ASAP7_75t_L   g17062(.A1(new_n17077), .A2(new_n17074), .B(new_n17064), .C(new_n17318), .Y(new_n17319));
  INVx1_ASAP7_75t_L         g17063(.A(new_n17319), .Y(new_n17320));
  NOR3xp33_ASAP7_75t_L      g17064(.A(new_n17076), .B(new_n17318), .C(new_n17064), .Y(new_n17321));
  NOR2xp33_ASAP7_75t_L      g17065(.A(new_n17320), .B(new_n17321), .Y(\f[78] ));
  O2A1O1Ixp33_ASAP7_75t_L   g17066(.A1(new_n17084), .A2(new_n17302), .B(new_n17295), .C(new_n17307), .Y(new_n17323));
  O2A1O1Ixp33_ASAP7_75t_L   g17067(.A1(new_n17298), .A2(new_n17296), .B(new_n17323), .C(new_n17300), .Y(new_n17324));
  NAND2xp33_ASAP7_75t_L     g17068(.A(new_n16827), .B(new_n16825), .Y(new_n17325));
  O2A1O1Ixp33_ASAP7_75t_L   g17069(.A1(new_n16836), .A2(new_n16837), .B(new_n17095), .C(new_n17325), .Y(new_n17326));
  A2O1A1Ixp33_ASAP7_75t_L   g17070(.A1(new_n17326), .A2(new_n17026), .B(new_n16826), .C(new_n17091), .Y(new_n17327));
  NAND2xp33_ASAP7_75t_L     g17071(.A(new_n17108), .B(new_n17292), .Y(new_n17328));
  INVx1_ASAP7_75t_L         g17072(.A(new_n12993), .Y(new_n17329));
  AOI22xp33_ASAP7_75t_L     g17073(.A1(new_n1204), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1290), .Y(new_n17330));
  INVx1_ASAP7_75t_L         g17074(.A(new_n17330), .Y(new_n17331));
  A2O1A1Ixp33_ASAP7_75t_L   g17075(.A1(new_n1205), .A2(new_n1207), .B(new_n1076), .C(new_n17330), .Y(new_n17332));
  O2A1O1Ixp33_ASAP7_75t_L   g17076(.A1(new_n17331), .A2(new_n17329), .B(new_n17332), .C(new_n1206), .Y(new_n17333));
  O2A1O1Ixp33_ASAP7_75t_L   g17077(.A1(new_n1210), .A2(new_n12993), .B(new_n17330), .C(\a[17] ), .Y(new_n17334));
  NOR2xp33_ASAP7_75t_L      g17078(.A(new_n17334), .B(new_n17333), .Y(new_n17335));
  A2O1A1O1Ixp25_ASAP7_75t_L g17079(.A1(new_n17304), .A2(new_n17328), .B(new_n17296), .C(new_n17327), .D(new_n17335), .Y(new_n17336));
  A2O1A1Ixp33_ASAP7_75t_L   g17080(.A1(new_n17328), .A2(new_n17304), .B(new_n17296), .C(new_n17327), .Y(new_n17337));
  NOR3xp33_ASAP7_75t_L      g17081(.A(new_n17337), .B(new_n17333), .C(new_n17334), .Y(new_n17338));
  NOR2xp33_ASAP7_75t_L      g17082(.A(new_n12258), .B(new_n1518), .Y(new_n17339));
  AOI221xp5_ASAP7_75t_L     g17083(.A1(\b[59] ), .A2(new_n1659), .B1(\b[60] ), .B2(new_n1507), .C(new_n17339), .Y(new_n17340));
  O2A1O1Ixp33_ASAP7_75t_L   g17084(.A1(new_n1521), .A2(new_n14764), .B(new_n17340), .C(new_n1501), .Y(new_n17341));
  INVx1_ASAP7_75t_L         g17085(.A(new_n17341), .Y(new_n17342));
  O2A1O1Ixp33_ASAP7_75t_L   g17086(.A1(new_n1521), .A2(new_n14764), .B(new_n17340), .C(\a[20] ), .Y(new_n17343));
  AOI21xp33_ASAP7_75t_L     g17087(.A1(new_n17342), .A2(\a[20] ), .B(new_n17343), .Y(new_n17344));
  O2A1O1Ixp33_ASAP7_75t_L   g17088(.A1(new_n16837), .A2(new_n17027), .B(new_n17103), .C(new_n17303), .Y(new_n17345));
  NAND2xp33_ASAP7_75t_L     g17089(.A(new_n17344), .B(new_n17345), .Y(new_n17346));
  O2A1O1Ixp33_ASAP7_75t_L   g17090(.A1(new_n17106), .A2(new_n17102), .B(new_n17292), .C(new_n17344), .Y(new_n17347));
  INVx1_ASAP7_75t_L         g17091(.A(new_n17347), .Y(new_n17348));
  NAND2xp33_ASAP7_75t_L     g17092(.A(new_n17120), .B(new_n17121), .Y(new_n17349));
  NOR2xp33_ASAP7_75t_L      g17093(.A(new_n10309), .B(new_n2415), .Y(new_n17350));
  AOI221xp5_ASAP7_75t_L     g17094(.A1(\b[53] ), .A2(new_n2577), .B1(\b[54] ), .B2(new_n2421), .C(new_n17350), .Y(new_n17351));
  O2A1O1Ixp33_ASAP7_75t_L   g17095(.A1(new_n2425), .A2(new_n15849), .B(new_n17351), .C(new_n2413), .Y(new_n17352));
  INVx1_ASAP7_75t_L         g17096(.A(new_n17352), .Y(new_n17353));
  O2A1O1Ixp33_ASAP7_75t_L   g17097(.A1(new_n2425), .A2(new_n15849), .B(new_n17351), .C(\a[26] ), .Y(new_n17354));
  AOI21xp33_ASAP7_75t_L     g17098(.A1(new_n17353), .A2(\a[26] ), .B(new_n17354), .Y(new_n17355));
  OAI311xp33_ASAP7_75t_L    g17099(.A1(new_n17349), .A2(new_n17285), .A3(new_n17281), .B1(new_n17355), .C1(new_n17121), .Y(new_n17356));
  A2O1A1O1Ixp25_ASAP7_75t_L g17100(.A1(new_n16709), .A2(new_n16707), .B(new_n16844), .C(new_n17009), .D(new_n17118), .Y(new_n17357));
  INVx1_ASAP7_75t_L         g17101(.A(new_n17281), .Y(new_n17358));
  NOR2xp33_ASAP7_75t_L      g17102(.A(new_n17285), .B(new_n17349), .Y(new_n17359));
  INVx1_ASAP7_75t_L         g17103(.A(new_n17355), .Y(new_n17360));
  A2O1A1Ixp33_ASAP7_75t_L   g17104(.A1(new_n17359), .A2(new_n17358), .B(new_n17357), .C(new_n17360), .Y(new_n17361));
  NAND2xp33_ASAP7_75t_L     g17105(.A(new_n17356), .B(new_n17361), .Y(new_n17362));
  INVx1_ASAP7_75t_L         g17106(.A(new_n9367), .Y(new_n17363));
  NOR2xp33_ASAP7_75t_L      g17107(.A(new_n9355), .B(new_n2930), .Y(new_n17364));
  AOI221xp5_ASAP7_75t_L     g17108(.A1(\b[50] ), .A2(new_n3129), .B1(\b[51] ), .B2(new_n2936), .C(new_n17364), .Y(new_n17365));
  O2A1O1Ixp33_ASAP7_75t_L   g17109(.A1(new_n2940), .A2(new_n17363), .B(new_n17365), .C(new_n2928), .Y(new_n17366));
  O2A1O1Ixp33_ASAP7_75t_L   g17110(.A1(new_n2940), .A2(new_n17363), .B(new_n17365), .C(\a[29] ), .Y(new_n17367));
  INVx1_ASAP7_75t_L         g17111(.A(new_n17367), .Y(new_n17368));
  OAI21xp33_ASAP7_75t_L     g17112(.A1(new_n2928), .A2(new_n17366), .B(new_n17368), .Y(new_n17369));
  INVx1_ASAP7_75t_L         g17113(.A(new_n17366), .Y(new_n17370));
  INVx1_ASAP7_75t_L         g17114(.A(new_n17278), .Y(new_n17371));
  A2O1A1Ixp33_ASAP7_75t_L   g17115(.A1(new_n17283), .A2(new_n17282), .B(new_n17271), .C(new_n17371), .Y(new_n17372));
  A2O1A1Ixp33_ASAP7_75t_L   g17116(.A1(new_n17370), .A2(\a[29] ), .B(new_n17367), .C(new_n17372), .Y(new_n17373));
  A2O1A1O1Ixp25_ASAP7_75t_L g17117(.A1(new_n17283), .A2(new_n17282), .B(new_n17271), .C(new_n17371), .D(new_n17369), .Y(new_n17374));
  AO21x2_ASAP7_75t_L        g17118(.A1(new_n17369), .A2(new_n17373), .B(new_n17374), .Y(new_n17375));
  NOR2xp33_ASAP7_75t_L      g17119(.A(new_n8427), .B(new_n3510), .Y(new_n17376));
  AOI221xp5_ASAP7_75t_L     g17120(.A1(\b[47] ), .A2(new_n3708), .B1(\b[48] ), .B2(new_n3499), .C(new_n17376), .Y(new_n17377));
  O2A1O1Ixp33_ASAP7_75t_L   g17121(.A1(new_n3513), .A2(new_n14802), .B(new_n17377), .C(new_n3493), .Y(new_n17378));
  O2A1O1Ixp33_ASAP7_75t_L   g17122(.A1(new_n3513), .A2(new_n14802), .B(new_n17377), .C(\a[32] ), .Y(new_n17379));
  INVx1_ASAP7_75t_L         g17123(.A(new_n17379), .Y(new_n17380));
  OAI21xp33_ASAP7_75t_L     g17124(.A1(new_n3493), .A2(new_n17378), .B(new_n17380), .Y(new_n17381));
  OR3x1_ASAP7_75t_L         g17125(.A(new_n17269), .B(new_n17263), .C(new_n17381), .Y(new_n17382));
  NOR2xp33_ASAP7_75t_L      g17126(.A(new_n17263), .B(new_n17269), .Y(new_n17383));
  O2A1O1Ixp33_ASAP7_75t_L   g17127(.A1(new_n3493), .A2(new_n17378), .B(new_n17380), .C(new_n17383), .Y(new_n17384));
  INVx1_ASAP7_75t_L         g17128(.A(new_n17384), .Y(new_n17385));
  NAND2xp33_ASAP7_75t_L     g17129(.A(new_n17382), .B(new_n17385), .Y(new_n17386));
  A2O1A1Ixp33_ASAP7_75t_L   g17130(.A1(new_n16972), .A2(new_n16987), .B(new_n17238), .C(new_n17236), .Y(new_n17387));
  NOR2xp33_ASAP7_75t_L      g17131(.A(new_n5855), .B(new_n5641), .Y(new_n17388));
  AOI221xp5_ASAP7_75t_L     g17132(.A1(\b[38] ), .A2(new_n5920), .B1(\b[39] ), .B2(new_n5623), .C(new_n17388), .Y(new_n17389));
  O2A1O1Ixp33_ASAP7_75t_L   g17133(.A1(new_n5630), .A2(new_n5862), .B(new_n17389), .C(new_n5626), .Y(new_n17390));
  NOR2xp33_ASAP7_75t_L      g17134(.A(new_n5626), .B(new_n17390), .Y(new_n17391));
  O2A1O1Ixp33_ASAP7_75t_L   g17135(.A1(new_n5630), .A2(new_n5862), .B(new_n17389), .C(\a[41] ), .Y(new_n17392));
  NOR2xp33_ASAP7_75t_L      g17136(.A(new_n17392), .B(new_n17391), .Y(new_n17393));
  O2A1O1Ixp33_ASAP7_75t_L   g17137(.A1(new_n17223), .A2(new_n6439), .B(new_n17225), .C(new_n17220), .Y(new_n17394));
  NOR2xp33_ASAP7_75t_L      g17138(.A(new_n17125), .B(new_n17227), .Y(new_n17395));
  NAND2xp33_ASAP7_75t_L     g17139(.A(\b[37] ), .B(new_n6442), .Y(new_n17396));
  OAI221xp5_ASAP7_75t_L     g17140(.A1(new_n7304), .A2(new_n4613), .B1(new_n4581), .B2(new_n6741), .C(new_n17396), .Y(new_n17397));
  A2O1A1Ixp33_ASAP7_75t_L   g17141(.A1(new_n10229), .A2(new_n6450), .B(new_n17397), .C(\a[44] ), .Y(new_n17398));
  AOI211xp5_ASAP7_75t_L     g17142(.A1(new_n10229), .A2(new_n6450), .B(new_n17397), .C(new_n6439), .Y(new_n17399));
  A2O1A1O1Ixp25_ASAP7_75t_L g17143(.A1(new_n6450), .A2(new_n10229), .B(new_n17397), .C(new_n17398), .D(new_n17399), .Y(new_n17400));
  INVx1_ASAP7_75t_L         g17144(.A(new_n17179), .Y(new_n17401));
  NOR2xp33_ASAP7_75t_L      g17145(.A(new_n1043), .B(new_n13030), .Y(new_n17402));
  O2A1O1Ixp33_ASAP7_75t_L   g17146(.A1(new_n867), .A2(new_n17137), .B(new_n16589), .C(new_n17136), .Y(new_n17403));
  A2O1A1Ixp33_ASAP7_75t_L   g17147(.A1(new_n13028), .A2(\b[16] ), .B(new_n17402), .C(new_n17403), .Y(new_n17404));
  O2A1O1Ixp33_ASAP7_75t_L   g17148(.A1(new_n12669), .A2(new_n12671), .B(\b[15] ), .C(new_n17134), .Y(new_n17405));
  O2A1O1Ixp33_ASAP7_75t_L   g17149(.A1(new_n12669), .A2(new_n12671), .B(\b[16] ), .C(new_n17402), .Y(new_n17406));
  INVx1_ASAP7_75t_L         g17150(.A(new_n17406), .Y(new_n17407));
  O2A1O1Ixp33_ASAP7_75t_L   g17151(.A1(\a[14] ), .A2(new_n17405), .B(new_n17140), .C(new_n17407), .Y(new_n17408));
  INVx1_ASAP7_75t_L         g17152(.A(new_n17408), .Y(new_n17409));
  AND2x2_ASAP7_75t_L        g17153(.A(new_n17404), .B(new_n17409), .Y(new_n17410));
  NAND2xp33_ASAP7_75t_L     g17154(.A(\b[19] ), .B(new_n11995), .Y(new_n17411));
  OAI221xp5_ASAP7_75t_L     g17155(.A1(new_n12318), .A2(new_n1458), .B1(new_n1349), .B2(new_n12320), .C(new_n17411), .Y(new_n17412));
  AOI21xp33_ASAP7_75t_L     g17156(.A1(new_n1607), .A2(new_n11997), .B(new_n17412), .Y(new_n17413));
  NAND2xp33_ASAP7_75t_L     g17157(.A(\a[62] ), .B(new_n17413), .Y(new_n17414));
  A2O1A1Ixp33_ASAP7_75t_L   g17158(.A1(new_n1607), .A2(new_n11997), .B(new_n17412), .C(new_n11987), .Y(new_n17415));
  NAND2xp33_ASAP7_75t_L     g17159(.A(new_n17415), .B(new_n17414), .Y(new_n17416));
  XNOR2x2_ASAP7_75t_L       g17160(.A(new_n17410), .B(new_n17416), .Y(new_n17417));
  O2A1O1Ixp33_ASAP7_75t_L   g17161(.A1(new_n17153), .A2(new_n17152), .B(new_n17149), .C(new_n17417), .Y(new_n17418));
  INVx1_ASAP7_75t_L         g17162(.A(new_n17418), .Y(new_n17419));
  NAND3xp33_ASAP7_75t_L     g17163(.A(new_n17417), .B(new_n17156), .C(new_n17149), .Y(new_n17420));
  AND2x2_ASAP7_75t_L        g17164(.A(new_n17420), .B(new_n17419), .Y(new_n17421));
  NOR2xp33_ASAP7_75t_L      g17165(.A(new_n1745), .B(new_n11354), .Y(new_n17422));
  AOI221xp5_ASAP7_75t_L     g17166(.A1(\b[22] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[21] ), .C(new_n17422), .Y(new_n17423));
  O2A1O1Ixp33_ASAP7_75t_L   g17167(.A1(new_n11053), .A2(new_n2522), .B(new_n17423), .C(new_n11048), .Y(new_n17424));
  INVx1_ASAP7_75t_L         g17168(.A(new_n17424), .Y(new_n17425));
  O2A1O1Ixp33_ASAP7_75t_L   g17169(.A1(new_n11053), .A2(new_n2522), .B(new_n17423), .C(\a[59] ), .Y(new_n17426));
  A2O1A1Ixp33_ASAP7_75t_L   g17170(.A1(\a[59] ), .A2(new_n17425), .B(new_n17426), .C(new_n17421), .Y(new_n17427));
  INVx1_ASAP7_75t_L         g17171(.A(new_n17426), .Y(new_n17428));
  O2A1O1Ixp33_ASAP7_75t_L   g17172(.A1(new_n17424), .A2(new_n11048), .B(new_n17428), .C(new_n17421), .Y(new_n17429));
  A2O1A1Ixp33_ASAP7_75t_L   g17173(.A1(new_n17167), .A2(new_n17157), .B(new_n17170), .C(new_n17165), .Y(new_n17430));
  AOI211xp5_ASAP7_75t_L     g17174(.A1(new_n17427), .A2(new_n17421), .B(new_n17429), .C(new_n17430), .Y(new_n17431));
  A2O1A1Ixp33_ASAP7_75t_L   g17175(.A1(new_n17427), .A2(new_n17421), .B(new_n17429), .C(new_n17430), .Y(new_n17432));
  INVx1_ASAP7_75t_L         g17176(.A(new_n17432), .Y(new_n17433));
  NOR2xp33_ASAP7_75t_L      g17177(.A(new_n17431), .B(new_n17433), .Y(new_n17434));
  NOR2xp33_ASAP7_75t_L      g17178(.A(new_n2205), .B(new_n10388), .Y(new_n17435));
  AOI221xp5_ASAP7_75t_L     g17179(.A1(new_n10086), .A2(\b[25] ), .B1(new_n11361), .B2(\b[23] ), .C(new_n17435), .Y(new_n17436));
  O2A1O1Ixp33_ASAP7_75t_L   g17180(.A1(new_n10088), .A2(new_n2385), .B(new_n17436), .C(new_n10083), .Y(new_n17437));
  INVx1_ASAP7_75t_L         g17181(.A(new_n17437), .Y(new_n17438));
  O2A1O1Ixp33_ASAP7_75t_L   g17182(.A1(new_n10088), .A2(new_n2385), .B(new_n17436), .C(\a[56] ), .Y(new_n17439));
  A2O1A1Ixp33_ASAP7_75t_L   g17183(.A1(\a[56] ), .A2(new_n17438), .B(new_n17439), .C(new_n17434), .Y(new_n17440));
  INVx1_ASAP7_75t_L         g17184(.A(new_n17439), .Y(new_n17441));
  O2A1O1Ixp33_ASAP7_75t_L   g17185(.A1(new_n17437), .A2(new_n10083), .B(new_n17441), .C(new_n17434), .Y(new_n17442));
  AOI21xp33_ASAP7_75t_L     g17186(.A1(new_n17440), .A2(new_n17434), .B(new_n17442), .Y(new_n17443));
  A2O1A1Ixp33_ASAP7_75t_L   g17187(.A1(new_n17177), .A2(new_n17401), .B(new_n17180), .C(new_n17443), .Y(new_n17444));
  A2O1A1Ixp33_ASAP7_75t_L   g17188(.A1(new_n17440), .A2(new_n17434), .B(new_n17442), .C(new_n17184), .Y(new_n17445));
  NAND2xp33_ASAP7_75t_L     g17189(.A(new_n17445), .B(new_n17444), .Y(new_n17446));
  NOR2xp33_ASAP7_75t_L      g17190(.A(new_n2879), .B(new_n10400), .Y(new_n17447));
  AOI221xp5_ASAP7_75t_L     g17191(.A1(new_n9102), .A2(\b[28] ), .B1(new_n10398), .B2(\b[26] ), .C(new_n17447), .Y(new_n17448));
  O2A1O1Ixp33_ASAP7_75t_L   g17192(.A1(new_n9104), .A2(new_n3087), .B(new_n17448), .C(new_n9099), .Y(new_n17449));
  NOR2xp33_ASAP7_75t_L      g17193(.A(new_n9099), .B(new_n17449), .Y(new_n17450));
  O2A1O1Ixp33_ASAP7_75t_L   g17194(.A1(new_n9104), .A2(new_n3087), .B(new_n17448), .C(\a[53] ), .Y(new_n17451));
  NOR2xp33_ASAP7_75t_L      g17195(.A(new_n17451), .B(new_n17450), .Y(new_n17452));
  XOR2x2_ASAP7_75t_L        g17196(.A(new_n17452), .B(new_n17446), .Y(new_n17453));
  O2A1O1Ixp33_ASAP7_75t_L   g17197(.A1(new_n17189), .A2(new_n17190), .B(new_n17186), .C(new_n17453), .Y(new_n17454));
  AND3x1_ASAP7_75t_L        g17198(.A(new_n17453), .B(new_n17193), .C(new_n17186), .Y(new_n17455));
  NOR2xp33_ASAP7_75t_L      g17199(.A(new_n17454), .B(new_n17455), .Y(new_n17456));
  NOR2xp33_ASAP7_75t_L      g17200(.A(new_n3456), .B(new_n10065), .Y(new_n17457));
  AOI221xp5_ASAP7_75t_L     g17201(.A1(new_n8175), .A2(\b[31] ), .B1(new_n8484), .B2(\b[29] ), .C(new_n17457), .Y(new_n17458));
  O2A1O1Ixp33_ASAP7_75t_L   g17202(.A1(new_n8176), .A2(new_n3681), .B(new_n17458), .C(new_n8172), .Y(new_n17459));
  INVx1_ASAP7_75t_L         g17203(.A(new_n17459), .Y(new_n17460));
  O2A1O1Ixp33_ASAP7_75t_L   g17204(.A1(new_n8176), .A2(new_n3681), .B(new_n17458), .C(\a[50] ), .Y(new_n17461));
  A2O1A1Ixp33_ASAP7_75t_L   g17205(.A1(\a[50] ), .A2(new_n17460), .B(new_n17461), .C(new_n17456), .Y(new_n17462));
  INVx1_ASAP7_75t_L         g17206(.A(new_n17461), .Y(new_n17463));
  O2A1O1Ixp33_ASAP7_75t_L   g17207(.A1(new_n17459), .A2(new_n8172), .B(new_n17463), .C(new_n17456), .Y(new_n17464));
  AOI21xp33_ASAP7_75t_L     g17208(.A1(new_n17462), .A2(new_n17456), .B(new_n17464), .Y(new_n17465));
  O2A1O1Ixp33_ASAP7_75t_L   g17209(.A1(new_n17195), .A2(new_n17205), .B(new_n17206), .C(new_n17201), .Y(new_n17466));
  NAND2xp33_ASAP7_75t_L     g17210(.A(new_n17466), .B(new_n17465), .Y(new_n17467));
  A2O1A1O1Ixp25_ASAP7_75t_L g17211(.A1(new_n17204), .A2(new_n17194), .B(new_n17208), .C(new_n17202), .D(new_n17465), .Y(new_n17468));
  INVx1_ASAP7_75t_L         g17212(.A(new_n17468), .Y(new_n17469));
  NAND2xp33_ASAP7_75t_L     g17213(.A(new_n17467), .B(new_n17469), .Y(new_n17470));
  INVx1_ASAP7_75t_L         g17214(.A(new_n17470), .Y(new_n17471));
  NOR2xp33_ASAP7_75t_L      g17215(.A(new_n4344), .B(new_n7318), .Y(new_n17472));
  AOI221xp5_ASAP7_75t_L     g17216(.A1(new_n7333), .A2(\b[33] ), .B1(new_n7609), .B2(\b[32] ), .C(new_n17472), .Y(new_n17473));
  O2A1O1Ixp33_ASAP7_75t_L   g17217(.A1(new_n7321), .A2(new_n4352), .B(new_n17473), .C(new_n7316), .Y(new_n17474));
  INVx1_ASAP7_75t_L         g17218(.A(new_n17474), .Y(new_n17475));
  O2A1O1Ixp33_ASAP7_75t_L   g17219(.A1(new_n7321), .A2(new_n4352), .B(new_n17473), .C(\a[47] ), .Y(new_n17476));
  AOI211xp5_ASAP7_75t_L     g17220(.A1(new_n17475), .A2(\a[47] ), .B(new_n17476), .C(new_n17471), .Y(new_n17477));
  A2O1A1Ixp33_ASAP7_75t_L   g17221(.A1(\a[47] ), .A2(new_n17475), .B(new_n17476), .C(new_n17471), .Y(new_n17478));
  INVx1_ASAP7_75t_L         g17222(.A(new_n17478), .Y(new_n17479));
  NOR2xp33_ASAP7_75t_L      g17223(.A(new_n17477), .B(new_n17479), .Y(new_n17480));
  INVx1_ASAP7_75t_L         g17224(.A(new_n17480), .Y(new_n17481));
  INVx1_ASAP7_75t_L         g17225(.A(new_n16950), .Y(new_n17482));
  A2O1A1Ixp33_ASAP7_75t_L   g17226(.A1(new_n16943), .A2(new_n16940), .B(new_n16944), .C(new_n17482), .Y(new_n17483));
  A2O1A1Ixp33_ASAP7_75t_L   g17227(.A1(new_n16943), .A2(new_n17483), .B(new_n17219), .C(new_n17216), .Y(new_n17484));
  NAND2xp33_ASAP7_75t_L     g17228(.A(new_n17484), .B(new_n17480), .Y(new_n17485));
  INVx1_ASAP7_75t_L         g17229(.A(new_n17485), .Y(new_n17486));
  NAND2xp33_ASAP7_75t_L     g17230(.A(new_n17484), .B(new_n17481), .Y(new_n17487));
  O2A1O1Ixp33_ASAP7_75t_L   g17231(.A1(new_n17481), .A2(new_n17486), .B(new_n17487), .C(new_n17400), .Y(new_n17488));
  O2A1O1Ixp33_ASAP7_75t_L   g17232(.A1(new_n16952), .A2(new_n16950), .B(new_n16943), .C(new_n17219), .Y(new_n17489));
  A2O1A1O1Ixp25_ASAP7_75t_L g17233(.A1(new_n17214), .A2(\a[47] ), .B(new_n17215), .C(new_n17210), .D(new_n17489), .Y(new_n17490));
  NAND2xp33_ASAP7_75t_L     g17234(.A(new_n17490), .B(new_n17480), .Y(new_n17491));
  NAND2xp33_ASAP7_75t_L     g17235(.A(new_n17400), .B(new_n17491), .Y(new_n17492));
  O2A1O1Ixp33_ASAP7_75t_L   g17236(.A1(new_n17477), .A2(new_n17479), .B(new_n17484), .C(new_n17492), .Y(new_n17493));
  OAI22xp33_ASAP7_75t_L     g17237(.A1(new_n17488), .A2(new_n17493), .B1(new_n17394), .B2(new_n17395), .Y(new_n17494));
  NOR2xp33_ASAP7_75t_L      g17238(.A(new_n17394), .B(new_n17395), .Y(new_n17495));
  NOR2xp33_ASAP7_75t_L      g17239(.A(new_n17493), .B(new_n17488), .Y(new_n17496));
  NAND2xp33_ASAP7_75t_L     g17240(.A(new_n17495), .B(new_n17496), .Y(new_n17497));
  AOI21xp33_ASAP7_75t_L     g17241(.A1(new_n17497), .A2(new_n17494), .B(new_n17393), .Y(new_n17498));
  AND3x1_ASAP7_75t_L        g17242(.A(new_n17497), .B(new_n17494), .C(new_n17393), .Y(new_n17499));
  NOR2xp33_ASAP7_75t_L      g17243(.A(new_n17498), .B(new_n17499), .Y(new_n17500));
  NAND2xp33_ASAP7_75t_L     g17244(.A(new_n17387), .B(new_n17500), .Y(new_n17501));
  INVx1_ASAP7_75t_L         g17245(.A(new_n17501), .Y(new_n17502));
  NOR2xp33_ASAP7_75t_L      g17246(.A(new_n17387), .B(new_n17500), .Y(new_n17503));
  NOR2xp33_ASAP7_75t_L      g17247(.A(new_n17503), .B(new_n17502), .Y(new_n17504));
  NOR2xp33_ASAP7_75t_L      g17248(.A(new_n6671), .B(new_n4908), .Y(new_n17505));
  AOI221xp5_ASAP7_75t_L     g17249(.A1(\b[41] ), .A2(new_n5139), .B1(\b[42] ), .B2(new_n4916), .C(new_n17505), .Y(new_n17506));
  O2A1O1Ixp33_ASAP7_75t_L   g17250(.A1(new_n4911), .A2(new_n6679), .B(new_n17506), .C(new_n4906), .Y(new_n17507));
  INVx1_ASAP7_75t_L         g17251(.A(new_n17507), .Y(new_n17508));
  O2A1O1Ixp33_ASAP7_75t_L   g17252(.A1(new_n4911), .A2(new_n6679), .B(new_n17506), .C(\a[38] ), .Y(new_n17509));
  A2O1A1Ixp33_ASAP7_75t_L   g17253(.A1(\a[38] ), .A2(new_n17508), .B(new_n17509), .C(new_n17504), .Y(new_n17510));
  INVx1_ASAP7_75t_L         g17254(.A(new_n17509), .Y(new_n17511));
  O2A1O1Ixp33_ASAP7_75t_L   g17255(.A1(new_n17507), .A2(new_n4906), .B(new_n17511), .C(new_n17504), .Y(new_n17512));
  AOI21xp33_ASAP7_75t_L     g17256(.A1(new_n17510), .A2(new_n17504), .B(new_n17512), .Y(new_n17513));
  A2O1A1Ixp33_ASAP7_75t_L   g17257(.A1(new_n16984), .A2(new_n16991), .B(new_n17252), .C(new_n17248), .Y(new_n17514));
  XNOR2x2_ASAP7_75t_L       g17258(.A(new_n17514), .B(new_n17513), .Y(new_n17515));
  NOR2xp33_ASAP7_75t_L      g17259(.A(new_n7249), .B(new_n4142), .Y(new_n17516));
  AOI221xp5_ASAP7_75t_L     g17260(.A1(\b[44] ), .A2(new_n4402), .B1(\b[46] ), .B2(new_n4156), .C(new_n17516), .Y(new_n17517));
  INVx1_ASAP7_75t_L         g17261(.A(new_n17517), .Y(new_n17518));
  A2O1A1Ixp33_ASAP7_75t_L   g17262(.A1(new_n7278), .A2(new_n4151), .B(new_n17518), .C(\a[35] ), .Y(new_n17519));
  O2A1O1Ixp33_ASAP7_75t_L   g17263(.A1(new_n4150), .A2(new_n7279), .B(new_n17517), .C(\a[35] ), .Y(new_n17520));
  A2O1A1Ixp33_ASAP7_75t_L   g17264(.A1(\a[35] ), .A2(new_n17519), .B(new_n17520), .C(new_n17515), .Y(new_n17521));
  NAND2xp33_ASAP7_75t_L     g17265(.A(new_n17515), .B(new_n17521), .Y(new_n17522));
  A2O1A1Ixp33_ASAP7_75t_L   g17266(.A1(new_n17519), .A2(\a[35] ), .B(new_n17520), .C(new_n17521), .Y(new_n17523));
  AND2x2_ASAP7_75t_L        g17267(.A(new_n17522), .B(new_n17523), .Y(new_n17524));
  NOR2xp33_ASAP7_75t_L      g17268(.A(new_n17524), .B(new_n17386), .Y(new_n17525));
  NAND2xp33_ASAP7_75t_L     g17269(.A(new_n17524), .B(new_n17386), .Y(new_n17526));
  A2O1A1Ixp33_ASAP7_75t_L   g17270(.A1(new_n17373), .A2(new_n17369), .B(new_n17374), .C(new_n17526), .Y(new_n17527));
  INVx1_ASAP7_75t_L         g17271(.A(new_n17525), .Y(new_n17528));
  AND3x1_ASAP7_75t_L        g17272(.A(new_n17527), .B(new_n17526), .C(new_n17528), .Y(new_n17529));
  O2A1O1Ixp33_ASAP7_75t_L   g17273(.A1(new_n17525), .A2(new_n17527), .B(new_n17375), .C(new_n17529), .Y(new_n17530));
  NOR2xp33_ASAP7_75t_L      g17274(.A(new_n17530), .B(new_n17362), .Y(new_n17531));
  INVx1_ASAP7_75t_L         g17275(.A(new_n17531), .Y(new_n17532));
  INVx1_ASAP7_75t_L         g17276(.A(new_n17115), .Y(new_n17533));
  NAND2xp33_ASAP7_75t_L     g17277(.A(\b[58] ), .B(new_n1955), .Y(new_n17534));
  OAI221xp5_ASAP7_75t_L     g17278(.A1(new_n1962), .A2(new_n10978), .B1(new_n10332), .B2(new_n2089), .C(new_n17534), .Y(new_n17535));
  AOI21xp33_ASAP7_75t_L     g17279(.A1(new_n11314), .A2(new_n1964), .B(new_n17535), .Y(new_n17536));
  NAND2xp33_ASAP7_75t_L     g17280(.A(\a[23] ), .B(new_n17536), .Y(new_n17537));
  A2O1A1Ixp33_ASAP7_75t_L   g17281(.A1(new_n11314), .A2(new_n1964), .B(new_n17535), .C(new_n1952), .Y(new_n17538));
  AND2x2_ASAP7_75t_L        g17282(.A(new_n17538), .B(new_n17537), .Y(new_n17539));
  INVx1_ASAP7_75t_L         g17283(.A(new_n17539), .Y(new_n17540));
  A2O1A1Ixp33_ASAP7_75t_L   g17284(.A1(new_n17288), .A2(new_n17113), .B(new_n17533), .C(new_n17540), .Y(new_n17541));
  O2A1O1Ixp33_ASAP7_75t_L   g17285(.A1(new_n17287), .A2(new_n17286), .B(new_n17113), .C(new_n17533), .Y(new_n17542));
  NAND2xp33_ASAP7_75t_L     g17286(.A(new_n17539), .B(new_n17542), .Y(new_n17543));
  NAND2xp33_ASAP7_75t_L     g17287(.A(new_n17543), .B(new_n17541), .Y(new_n17544));
  NAND2xp33_ASAP7_75t_L     g17288(.A(new_n17530), .B(new_n17362), .Y(new_n17545));
  AOI21xp33_ASAP7_75t_L     g17289(.A1(new_n17532), .A2(new_n17545), .B(new_n17544), .Y(new_n17546));
  AND2x2_ASAP7_75t_L        g17290(.A(new_n17356), .B(new_n17361), .Y(new_n17547));
  INVx1_ASAP7_75t_L         g17291(.A(new_n17530), .Y(new_n17548));
  NOR2xp33_ASAP7_75t_L      g17292(.A(new_n17548), .B(new_n17547), .Y(new_n17549));
  AOI31xp33_ASAP7_75t_L     g17293(.A1(new_n17532), .A2(new_n17541), .A3(new_n17543), .B(new_n17549), .Y(new_n17550));
  AO21x2_ASAP7_75t_L        g17294(.A1(new_n17532), .A2(new_n17550), .B(new_n17546), .Y(new_n17551));
  NAND3xp33_ASAP7_75t_L     g17295(.A(new_n17551), .B(new_n17348), .C(new_n17346), .Y(new_n17552));
  INVx1_ASAP7_75t_L         g17296(.A(new_n17344), .Y(new_n17553));
  A2O1A1Ixp33_ASAP7_75t_L   g17297(.A1(new_n17026), .A2(new_n17094), .B(new_n17102), .C(new_n17292), .Y(new_n17554));
  NOR2xp33_ASAP7_75t_L      g17298(.A(new_n17553), .B(new_n17554), .Y(new_n17555));
  O2A1O1Ixp33_ASAP7_75t_L   g17299(.A1(new_n17530), .A2(new_n17362), .B(new_n17550), .C(new_n17546), .Y(new_n17556));
  OAI21xp33_ASAP7_75t_L     g17300(.A1(new_n17347), .A2(new_n17555), .B(new_n17556), .Y(new_n17557));
  AO211x2_ASAP7_75t_L       g17301(.A1(new_n17552), .A2(new_n17557), .B(new_n17336), .C(new_n17338), .Y(new_n17558));
  OAI211xp5_ASAP7_75t_L     g17302(.A1(new_n17336), .A2(new_n17338), .B(new_n17557), .C(new_n17552), .Y(new_n17559));
  NAND2xp33_ASAP7_75t_L     g17303(.A(new_n17559), .B(new_n17558), .Y(new_n17560));
  INVx1_ASAP7_75t_L         g17304(.A(new_n17314), .Y(new_n17561));
  A2O1A1Ixp33_ASAP7_75t_L   g17305(.A1(new_n17093), .A2(new_n17306), .B(new_n17561), .C(new_n17312), .Y(new_n17562));
  NOR2xp33_ASAP7_75t_L      g17306(.A(new_n17562), .B(new_n17560), .Y(new_n17563));
  A2O1A1O1Ixp25_ASAP7_75t_L g17307(.A1(new_n17292), .A2(new_n17108), .B(new_n17294), .C(new_n17093), .D(new_n17561), .Y(new_n17564));
  A2O1A1Ixp33_ASAP7_75t_L   g17308(.A1(new_n17083), .A2(new_n17301), .B(new_n17564), .C(new_n17560), .Y(new_n17565));
  INVx1_ASAP7_75t_L         g17309(.A(new_n17565), .Y(new_n17566));
  NOR2xp33_ASAP7_75t_L      g17310(.A(new_n17563), .B(new_n17566), .Y(new_n17567));
  INVx1_ASAP7_75t_L         g17311(.A(new_n17567), .Y(new_n17568));
  O2A1O1Ixp33_ASAP7_75t_L   g17312(.A1(new_n17324), .A2(new_n17316), .B(new_n17319), .C(new_n17568), .Y(new_n17569));
  A2O1A1Ixp33_ASAP7_75t_L   g17313(.A1(new_n17071), .A2(new_n17065), .B(new_n17324), .C(new_n17319), .Y(new_n17570));
  NOR2xp33_ASAP7_75t_L      g17314(.A(new_n17570), .B(new_n17567), .Y(new_n17571));
  NOR2xp33_ASAP7_75t_L      g17315(.A(new_n17571), .B(new_n17569), .Y(\f[79] ));
  INVx1_ASAP7_75t_L         g17316(.A(new_n17336), .Y(new_n17573));
  INVx1_ASAP7_75t_L         g17317(.A(new_n17337), .Y(new_n17574));
  NAND2xp33_ASAP7_75t_L     g17318(.A(new_n17335), .B(new_n17574), .Y(new_n17575));
  NAND4xp25_ASAP7_75t_L     g17319(.A(new_n17575), .B(new_n17552), .C(new_n17557), .D(new_n17573), .Y(new_n17576));
  A2O1A1Ixp33_ASAP7_75t_L   g17320(.A1(new_n17295), .A2(new_n17327), .B(new_n17335), .C(new_n17576), .Y(new_n17577));
  NOR2xp33_ASAP7_75t_L      g17321(.A(new_n12956), .B(new_n1285), .Y(new_n17578));
  A2O1A1Ixp33_ASAP7_75t_L   g17322(.A1(new_n12986), .A2(new_n1216), .B(new_n17578), .C(\a[17] ), .Y(new_n17579));
  A2O1A1O1Ixp25_ASAP7_75t_L g17323(.A1(new_n1216), .A2(new_n14172), .B(new_n1290), .C(\b[63] ), .D(new_n1206), .Y(new_n17580));
  A2O1A1O1Ixp25_ASAP7_75t_L g17324(.A1(new_n12986), .A2(new_n1216), .B(new_n17578), .C(new_n17579), .D(new_n17580), .Y(new_n17581));
  O2A1O1Ixp33_ASAP7_75t_L   g17325(.A1(new_n17556), .A2(new_n17555), .B(new_n17348), .C(new_n17581), .Y(new_n17582));
  A2O1A1Ixp33_ASAP7_75t_L   g17326(.A1(new_n17551), .A2(new_n17346), .B(new_n17347), .C(new_n17581), .Y(new_n17583));
  NOR2xp33_ASAP7_75t_L      g17327(.A(new_n12603), .B(new_n1518), .Y(new_n17584));
  AOI221xp5_ASAP7_75t_L     g17328(.A1(\b[60] ), .A2(new_n1659), .B1(\b[61] ), .B2(new_n1507), .C(new_n17584), .Y(new_n17585));
  O2A1O1Ixp33_ASAP7_75t_L   g17329(.A1(new_n1521), .A2(new_n12610), .B(new_n17585), .C(new_n1501), .Y(new_n17586));
  INVx1_ASAP7_75t_L         g17330(.A(new_n17586), .Y(new_n17587));
  O2A1O1Ixp33_ASAP7_75t_L   g17331(.A1(new_n1521), .A2(new_n12610), .B(new_n17585), .C(\a[20] ), .Y(new_n17588));
  OAI31xp33_ASAP7_75t_L     g17332(.A1(new_n17544), .A2(new_n17549), .A3(new_n17531), .B(new_n17541), .Y(new_n17589));
  AOI211xp5_ASAP7_75t_L     g17333(.A1(\a[20] ), .A2(new_n17587), .B(new_n17588), .C(new_n17589), .Y(new_n17590));
  NAND3xp33_ASAP7_75t_L     g17334(.A(new_n17545), .B(new_n17543), .C(new_n17541), .Y(new_n17591));
  AOI21xp33_ASAP7_75t_L     g17335(.A1(new_n17587), .A2(\a[20] ), .B(new_n17588), .Y(new_n17592));
  O2A1O1Ixp33_ASAP7_75t_L   g17336(.A1(new_n17531), .A2(new_n17591), .B(new_n17541), .C(new_n17592), .Y(new_n17593));
  NOR2xp33_ASAP7_75t_L      g17337(.A(new_n17593), .B(new_n17590), .Y(new_n17594));
  NOR2xp33_ASAP7_75t_L      g17338(.A(new_n11303), .B(new_n1962), .Y(new_n17595));
  AOI221xp5_ASAP7_75t_L     g17339(.A1(new_n1955), .A2(\b[59] ), .B1(new_n2093), .B2(\b[57] ), .C(new_n17595), .Y(new_n17596));
  O2A1O1Ixp33_ASAP7_75t_L   g17340(.A1(new_n1956), .A2(new_n11597), .B(new_n17596), .C(new_n1952), .Y(new_n17597));
  INVx1_ASAP7_75t_L         g17341(.A(new_n17597), .Y(new_n17598));
  O2A1O1Ixp33_ASAP7_75t_L   g17342(.A1(new_n1956), .A2(new_n11597), .B(new_n17596), .C(\a[23] ), .Y(new_n17599));
  AOI21xp33_ASAP7_75t_L     g17343(.A1(new_n17598), .A2(\a[23] ), .B(new_n17599), .Y(new_n17600));
  INVx1_ASAP7_75t_L         g17344(.A(new_n17356), .Y(new_n17601));
  O2A1O1Ixp33_ASAP7_75t_L   g17345(.A1(new_n17601), .A2(new_n17530), .B(new_n17361), .C(new_n17600), .Y(new_n17602));
  INVx1_ASAP7_75t_L         g17346(.A(new_n17361), .Y(new_n17603));
  A2O1A1Ixp33_ASAP7_75t_L   g17347(.A1(new_n17548), .A2(new_n17356), .B(new_n17603), .C(new_n17600), .Y(new_n17604));
  OAI21xp33_ASAP7_75t_L     g17348(.A1(new_n17600), .A2(new_n17602), .B(new_n17604), .Y(new_n17605));
  NAND3xp33_ASAP7_75t_L     g17349(.A(new_n17375), .B(new_n17528), .C(new_n17526), .Y(new_n17606));
  NOR2xp33_ASAP7_75t_L      g17350(.A(new_n10332), .B(new_n2415), .Y(new_n17607));
  AOI221xp5_ASAP7_75t_L     g17351(.A1(\b[54] ), .A2(new_n2577), .B1(\b[55] ), .B2(new_n2421), .C(new_n17607), .Y(new_n17608));
  O2A1O1Ixp33_ASAP7_75t_L   g17352(.A1(new_n2425), .A2(new_n10339), .B(new_n17608), .C(new_n2413), .Y(new_n17609));
  INVx1_ASAP7_75t_L         g17353(.A(new_n17609), .Y(new_n17610));
  O2A1O1Ixp33_ASAP7_75t_L   g17354(.A1(new_n2425), .A2(new_n10339), .B(new_n17608), .C(\a[26] ), .Y(new_n17611));
  AOI21xp33_ASAP7_75t_L     g17355(.A1(new_n17610), .A2(\a[26] ), .B(new_n17611), .Y(new_n17612));
  AND3x1_ASAP7_75t_L        g17356(.A(new_n17606), .B(new_n17612), .C(new_n17373), .Y(new_n17613));
  O2A1O1Ixp33_ASAP7_75t_L   g17357(.A1(new_n17525), .A2(new_n17527), .B(new_n17373), .C(new_n17612), .Y(new_n17614));
  NOR2xp33_ASAP7_75t_L      g17358(.A(new_n17614), .B(new_n17613), .Y(new_n17615));
  INVx1_ASAP7_75t_L         g17359(.A(new_n17383), .Y(new_n17616));
  NOR2xp33_ASAP7_75t_L      g17360(.A(new_n9683), .B(new_n2930), .Y(new_n17617));
  AOI221xp5_ASAP7_75t_L     g17361(.A1(\b[51] ), .A2(new_n3129), .B1(\b[52] ), .B2(new_n2936), .C(new_n17617), .Y(new_n17618));
  O2A1O1Ixp33_ASAP7_75t_L   g17362(.A1(new_n2940), .A2(new_n9691), .B(new_n17618), .C(new_n2928), .Y(new_n17619));
  O2A1O1Ixp33_ASAP7_75t_L   g17363(.A1(new_n2940), .A2(new_n9691), .B(new_n17618), .C(\a[29] ), .Y(new_n17620));
  INVx1_ASAP7_75t_L         g17364(.A(new_n17620), .Y(new_n17621));
  OAI21xp33_ASAP7_75t_L     g17365(.A1(new_n2928), .A2(new_n17619), .B(new_n17621), .Y(new_n17622));
  A2O1A1Ixp33_ASAP7_75t_L   g17366(.A1(new_n17616), .A2(new_n17381), .B(new_n17525), .C(new_n17622), .Y(new_n17623));
  INVx1_ASAP7_75t_L         g17367(.A(new_n17623), .Y(new_n17624));
  A2O1A1Ixp33_ASAP7_75t_L   g17368(.A1(new_n17522), .A2(new_n17523), .B(new_n17386), .C(new_n17385), .Y(new_n17625));
  O2A1O1Ixp33_ASAP7_75t_L   g17369(.A1(new_n2928), .A2(new_n17619), .B(new_n17621), .C(new_n17625), .Y(new_n17626));
  INVx1_ASAP7_75t_L         g17370(.A(new_n17626), .Y(new_n17627));
  A2O1A1Ixp33_ASAP7_75t_L   g17371(.A1(new_n17528), .A2(new_n17385), .B(new_n17624), .C(new_n17627), .Y(new_n17628));
  O2A1O1Ixp33_ASAP7_75t_L   g17372(.A1(new_n17524), .A2(new_n17386), .B(new_n17385), .C(new_n17622), .Y(new_n17629));
  NOR2xp33_ASAP7_75t_L      g17373(.A(new_n8427), .B(new_n3509), .Y(new_n17630));
  AOI221xp5_ASAP7_75t_L     g17374(.A1(\b[48] ), .A2(new_n3708), .B1(\b[50] ), .B2(new_n3503), .C(new_n17630), .Y(new_n17631));
  INVx1_ASAP7_75t_L         g17375(.A(new_n17631), .Y(new_n17632));
  O2A1O1Ixp33_ASAP7_75t_L   g17376(.A1(new_n3513), .A2(new_n8764), .B(new_n17631), .C(new_n3493), .Y(new_n17633));
  INVx1_ASAP7_75t_L         g17377(.A(new_n17633), .Y(new_n17634));
  NOR2xp33_ASAP7_75t_L      g17378(.A(new_n3493), .B(new_n17633), .Y(new_n17635));
  A2O1A1O1Ixp25_ASAP7_75t_L g17379(.A1(new_n8763), .A2(new_n3505), .B(new_n17632), .C(new_n17634), .D(new_n17635), .Y(new_n17636));
  O2A1O1Ixp33_ASAP7_75t_L   g17380(.A1(new_n17249), .A2(new_n17250), .B(new_n17256), .C(new_n17513), .Y(new_n17637));
  A2O1A1O1Ixp25_ASAP7_75t_L g17381(.A1(new_n17519), .A2(\a[35] ), .B(new_n17520), .C(new_n17515), .D(new_n17637), .Y(new_n17638));
  XOR2x2_ASAP7_75t_L        g17382(.A(new_n17636), .B(new_n17638), .Y(new_n17639));
  NOR2xp33_ASAP7_75t_L      g17383(.A(new_n6944), .B(new_n4908), .Y(new_n17640));
  AOI221xp5_ASAP7_75t_L     g17384(.A1(\b[42] ), .A2(new_n5139), .B1(\b[43] ), .B2(new_n4916), .C(new_n17640), .Y(new_n17641));
  O2A1O1Ixp33_ASAP7_75t_L   g17385(.A1(new_n4911), .A2(new_n6951), .B(new_n17641), .C(new_n4906), .Y(new_n17642));
  INVx1_ASAP7_75t_L         g17386(.A(new_n17642), .Y(new_n17643));
  O2A1O1Ixp33_ASAP7_75t_L   g17387(.A1(new_n4911), .A2(new_n6951), .B(new_n17641), .C(\a[38] ), .Y(new_n17644));
  AOI21xp33_ASAP7_75t_L     g17388(.A1(new_n17643), .A2(\a[38] ), .B(new_n17644), .Y(new_n17645));
  O2A1O1Ixp33_ASAP7_75t_L   g17389(.A1(new_n17394), .A2(new_n17395), .B(new_n17496), .C(new_n17498), .Y(new_n17646));
  NOR2xp33_ASAP7_75t_L      g17390(.A(new_n5855), .B(new_n5640), .Y(new_n17647));
  AOI221xp5_ASAP7_75t_L     g17391(.A1(\b[39] ), .A2(new_n5920), .B1(\b[41] ), .B2(new_n5629), .C(new_n17647), .Y(new_n17648));
  O2A1O1Ixp33_ASAP7_75t_L   g17392(.A1(new_n5630), .A2(new_n6117), .B(new_n17648), .C(new_n5626), .Y(new_n17649));
  INVx1_ASAP7_75t_L         g17393(.A(new_n17649), .Y(new_n17650));
  O2A1O1Ixp33_ASAP7_75t_L   g17394(.A1(new_n5630), .A2(new_n6117), .B(new_n17648), .C(\a[41] ), .Y(new_n17651));
  AOI21xp33_ASAP7_75t_L     g17395(.A1(new_n17650), .A2(\a[41] ), .B(new_n17651), .Y(new_n17652));
  A2O1A1Ixp33_ASAP7_75t_L   g17396(.A1(new_n17491), .A2(new_n17490), .B(new_n17400), .C(new_n17485), .Y(new_n17653));
  INVx1_ASAP7_75t_L         g17397(.A(new_n17653), .Y(new_n17654));
  A2O1A1O1Ixp25_ASAP7_75t_L g17398(.A1(new_n17475), .A2(\a[47] ), .B(new_n17476), .C(new_n17467), .D(new_n17468), .Y(new_n17655));
  INVx1_ASAP7_75t_L         g17399(.A(new_n17655), .Y(new_n17656));
  MAJIxp5_ASAP7_75t_L       g17400(.A(new_n17443), .B(new_n17452), .C(new_n17184), .Y(new_n17657));
  NAND2xp33_ASAP7_75t_L     g17401(.A(\a[56] ), .B(new_n17438), .Y(new_n17658));
  A2O1A1Ixp33_ASAP7_75t_L   g17402(.A1(new_n17658), .A2(new_n17441), .B(new_n17431), .C(new_n17432), .Y(new_n17659));
  NOR2xp33_ASAP7_75t_L      g17403(.A(new_n2377), .B(new_n10388), .Y(new_n17660));
  AOI221xp5_ASAP7_75t_L     g17404(.A1(new_n10086), .A2(\b[26] ), .B1(new_n11361), .B2(\b[24] ), .C(new_n17660), .Y(new_n17661));
  O2A1O1Ixp33_ASAP7_75t_L   g17405(.A1(new_n10088), .A2(new_n2708), .B(new_n17661), .C(new_n10083), .Y(new_n17662));
  INVx1_ASAP7_75t_L         g17406(.A(new_n17662), .Y(new_n17663));
  O2A1O1Ixp33_ASAP7_75t_L   g17407(.A1(new_n10088), .A2(new_n2708), .B(new_n17661), .C(\a[56] ), .Y(new_n17664));
  AO21x2_ASAP7_75t_L        g17408(.A1(\a[56] ), .A2(new_n17663), .B(new_n17664), .Y(new_n17665));
  A2O1A1O1Ixp25_ASAP7_75t_L g17409(.A1(new_n17425), .A2(\a[59] ), .B(new_n17426), .C(new_n17420), .D(new_n17418), .Y(new_n17666));
  NOR2xp33_ASAP7_75t_L      g17410(.A(new_n1150), .B(new_n13030), .Y(new_n17667));
  O2A1O1Ixp33_ASAP7_75t_L   g17411(.A1(new_n12669), .A2(new_n12671), .B(\b[17] ), .C(new_n17667), .Y(new_n17668));
  NOR2xp33_ASAP7_75t_L      g17412(.A(new_n1599), .B(new_n12318), .Y(new_n17669));
  AOI221xp5_ASAP7_75t_L     g17413(.A1(new_n11995), .A2(\b[20] ), .B1(new_n13314), .B2(\b[18] ), .C(new_n17669), .Y(new_n17670));
  O2A1O1Ixp33_ASAP7_75t_L   g17414(.A1(new_n11998), .A2(new_n1754), .B(new_n17670), .C(new_n11987), .Y(new_n17671));
  INVx1_ASAP7_75t_L         g17415(.A(new_n17670), .Y(new_n17672));
  A2O1A1Ixp33_ASAP7_75t_L   g17416(.A1(new_n1752), .A2(new_n11997), .B(new_n17672), .C(new_n11987), .Y(new_n17673));
  INVx1_ASAP7_75t_L         g17417(.A(new_n17671), .Y(new_n17674));
  INVx1_ASAP7_75t_L         g17418(.A(new_n17673), .Y(new_n17675));
  A2O1A1Ixp33_ASAP7_75t_L   g17419(.A1(new_n13028), .A2(\b[16] ), .B(new_n17402), .C(new_n17668), .Y(new_n17676));
  A2O1A1Ixp33_ASAP7_75t_L   g17420(.A1(new_n17674), .A2(\a[62] ), .B(new_n17675), .C(new_n17676), .Y(new_n17677));
  A2O1A1O1Ixp25_ASAP7_75t_L g17421(.A1(new_n13028), .A2(\b[17] ), .B(new_n17667), .C(new_n17406), .D(new_n17677), .Y(new_n17678));
  O2A1O1Ixp33_ASAP7_75t_L   g17422(.A1(new_n11987), .A2(new_n17671), .B(new_n17673), .C(new_n17678), .Y(new_n17679));
  NAND2xp33_ASAP7_75t_L     g17423(.A(\a[62] ), .B(new_n17674), .Y(new_n17680));
  INVx1_ASAP7_75t_L         g17424(.A(new_n17667), .Y(new_n17681));
  O2A1O1Ixp33_ASAP7_75t_L   g17425(.A1(new_n12672), .A2(new_n1349), .B(new_n17681), .C(new_n17407), .Y(new_n17682));
  A2O1A1Ixp33_ASAP7_75t_L   g17426(.A1(new_n17680), .A2(new_n17673), .B(new_n17682), .C(new_n17676), .Y(new_n17683));
  INVx1_ASAP7_75t_L         g17427(.A(new_n17683), .Y(new_n17684));
  O2A1O1Ixp33_ASAP7_75t_L   g17428(.A1(new_n17668), .A2(new_n17407), .B(new_n17684), .C(new_n17679), .Y(new_n17685));
  INVx1_ASAP7_75t_L         g17429(.A(new_n17410), .Y(new_n17686));
  A2O1A1Ixp33_ASAP7_75t_L   g17430(.A1(new_n17414), .A2(new_n17415), .B(new_n17686), .C(new_n17409), .Y(new_n17687));
  XOR2x2_ASAP7_75t_L        g17431(.A(new_n17687), .B(new_n17685), .Y(new_n17688));
  NOR2xp33_ASAP7_75t_L      g17432(.A(new_n1895), .B(new_n11354), .Y(new_n17689));
  AOI221xp5_ASAP7_75t_L     g17433(.A1(\b[23] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[22] ), .C(new_n17689), .Y(new_n17690));
  INVx1_ASAP7_75t_L         g17434(.A(new_n17690), .Y(new_n17691));
  A2O1A1Ixp33_ASAP7_75t_L   g17435(.A1(new_n2679), .A2(new_n11351), .B(new_n17691), .C(\a[59] ), .Y(new_n17692));
  O2A1O1Ixp33_ASAP7_75t_L   g17436(.A1(new_n11053), .A2(new_n2194), .B(new_n17690), .C(new_n11048), .Y(new_n17693));
  NOR2xp33_ASAP7_75t_L      g17437(.A(new_n11048), .B(new_n17693), .Y(new_n17694));
  A2O1A1O1Ixp25_ASAP7_75t_L g17438(.A1(new_n11351), .A2(new_n2679), .B(new_n17691), .C(new_n17692), .D(new_n17694), .Y(new_n17695));
  XNOR2x2_ASAP7_75t_L       g17439(.A(new_n17695), .B(new_n17688), .Y(new_n17696));
  XOR2x2_ASAP7_75t_L        g17440(.A(new_n17666), .B(new_n17696), .Y(new_n17697));
  XNOR2x2_ASAP7_75t_L       g17441(.A(new_n17665), .B(new_n17697), .Y(new_n17698));
  XOR2x2_ASAP7_75t_L        g17442(.A(new_n17659), .B(new_n17698), .Y(new_n17699));
  NOR2xp33_ASAP7_75t_L      g17443(.A(new_n3079), .B(new_n10400), .Y(new_n17700));
  AOI221xp5_ASAP7_75t_L     g17444(.A1(new_n9102), .A2(\b[29] ), .B1(new_n10398), .B2(\b[27] ), .C(new_n17700), .Y(new_n17701));
  O2A1O1Ixp33_ASAP7_75t_L   g17445(.A1(new_n9104), .A2(new_n3104), .B(new_n17701), .C(new_n9099), .Y(new_n17702));
  O2A1O1Ixp33_ASAP7_75t_L   g17446(.A1(new_n9104), .A2(new_n3104), .B(new_n17701), .C(\a[53] ), .Y(new_n17703));
  INVx1_ASAP7_75t_L         g17447(.A(new_n17703), .Y(new_n17704));
  OAI21xp33_ASAP7_75t_L     g17448(.A1(new_n9099), .A2(new_n17702), .B(new_n17704), .Y(new_n17705));
  XNOR2x2_ASAP7_75t_L       g17449(.A(new_n17705), .B(new_n17699), .Y(new_n17706));
  NAND2xp33_ASAP7_75t_L     g17450(.A(new_n17657), .B(new_n17706), .Y(new_n17707));
  O2A1O1Ixp33_ASAP7_75t_L   g17451(.A1(new_n17702), .A2(new_n9099), .B(new_n17704), .C(new_n17699), .Y(new_n17708));
  INVx1_ASAP7_75t_L         g17452(.A(new_n17702), .Y(new_n17709));
  A2O1A1Ixp33_ASAP7_75t_L   g17453(.A1(\a[53] ), .A2(new_n17709), .B(new_n17703), .C(new_n17699), .Y(new_n17710));
  O2A1O1Ixp33_ASAP7_75t_L   g17454(.A1(new_n17699), .A2(new_n17708), .B(new_n17710), .C(new_n17657), .Y(new_n17711));
  AOI21xp33_ASAP7_75t_L     g17455(.A1(new_n17707), .A2(new_n17657), .B(new_n17711), .Y(new_n17712));
  NOR2xp33_ASAP7_75t_L      g17456(.A(new_n3674), .B(new_n10065), .Y(new_n17713));
  AOI221xp5_ASAP7_75t_L     g17457(.A1(new_n8175), .A2(\b[32] ), .B1(new_n8484), .B2(\b[30] ), .C(new_n17713), .Y(new_n17714));
  O2A1O1Ixp33_ASAP7_75t_L   g17458(.A1(new_n8176), .A2(new_n3897), .B(new_n17714), .C(new_n8172), .Y(new_n17715));
  NOR2xp33_ASAP7_75t_L      g17459(.A(new_n8172), .B(new_n17715), .Y(new_n17716));
  O2A1O1Ixp33_ASAP7_75t_L   g17460(.A1(new_n8176), .A2(new_n3897), .B(new_n17714), .C(\a[50] ), .Y(new_n17717));
  NOR2xp33_ASAP7_75t_L      g17461(.A(new_n17717), .B(new_n17716), .Y(new_n17718));
  XNOR2x2_ASAP7_75t_L       g17462(.A(new_n17718), .B(new_n17712), .Y(new_n17719));
  A2O1A1O1Ixp25_ASAP7_75t_L g17463(.A1(new_n17460), .A2(\a[50] ), .B(new_n17461), .C(new_n17456), .D(new_n17454), .Y(new_n17720));
  NAND2xp33_ASAP7_75t_L     g17464(.A(new_n17720), .B(new_n17719), .Y(new_n17721));
  A2O1A1O1Ixp25_ASAP7_75t_L g17465(.A1(new_n17193), .A2(new_n17186), .B(new_n17453), .C(new_n17462), .D(new_n17719), .Y(new_n17722));
  INVx1_ASAP7_75t_L         g17466(.A(new_n17722), .Y(new_n17723));
  NAND2xp33_ASAP7_75t_L     g17467(.A(new_n17721), .B(new_n17723), .Y(new_n17724));
  NOR2xp33_ASAP7_75t_L      g17468(.A(new_n4581), .B(new_n7318), .Y(new_n17725));
  AOI221xp5_ASAP7_75t_L     g17469(.A1(new_n7333), .A2(\b[34] ), .B1(new_n7609), .B2(\b[33] ), .C(new_n17725), .Y(new_n17726));
  O2A1O1Ixp33_ASAP7_75t_L   g17470(.A1(new_n7321), .A2(new_n4589), .B(new_n17726), .C(new_n7316), .Y(new_n17727));
  O2A1O1Ixp33_ASAP7_75t_L   g17471(.A1(new_n7321), .A2(new_n4589), .B(new_n17726), .C(\a[47] ), .Y(new_n17728));
  INVx1_ASAP7_75t_L         g17472(.A(new_n17728), .Y(new_n17729));
  O2A1O1Ixp33_ASAP7_75t_L   g17473(.A1(new_n17727), .A2(new_n7316), .B(new_n17729), .C(new_n17724), .Y(new_n17730));
  INVx1_ASAP7_75t_L         g17474(.A(new_n17727), .Y(new_n17731));
  A2O1A1Ixp33_ASAP7_75t_L   g17475(.A1(\a[47] ), .A2(new_n17731), .B(new_n17728), .C(new_n17724), .Y(new_n17732));
  O2A1O1Ixp33_ASAP7_75t_L   g17476(.A1(new_n17724), .A2(new_n17730), .B(new_n17732), .C(new_n17655), .Y(new_n17733));
  INVx1_ASAP7_75t_L         g17477(.A(new_n17733), .Y(new_n17734));
  O2A1O1Ixp33_ASAP7_75t_L   g17478(.A1(new_n17724), .A2(new_n17730), .B(new_n17732), .C(new_n17656), .Y(new_n17735));
  NOR2xp33_ASAP7_75t_L      g17479(.A(new_n4613), .B(new_n6741), .Y(new_n17736));
  AOI221xp5_ASAP7_75t_L     g17480(.A1(\b[38] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[37] ), .C(new_n17736), .Y(new_n17737));
  O2A1O1Ixp33_ASAP7_75t_L   g17481(.A1(new_n6443), .A2(new_n5318), .B(new_n17737), .C(new_n6439), .Y(new_n17738));
  INVx1_ASAP7_75t_L         g17482(.A(new_n17738), .Y(new_n17739));
  O2A1O1Ixp33_ASAP7_75t_L   g17483(.A1(new_n6443), .A2(new_n5318), .B(new_n17737), .C(\a[44] ), .Y(new_n17740));
  AOI21xp33_ASAP7_75t_L     g17484(.A1(new_n17739), .A2(\a[44] ), .B(new_n17740), .Y(new_n17741));
  A2O1A1Ixp33_ASAP7_75t_L   g17485(.A1(new_n17734), .A2(new_n17656), .B(new_n17735), .C(new_n17741), .Y(new_n17742));
  O2A1O1Ixp33_ASAP7_75t_L   g17486(.A1(new_n17468), .A2(new_n17479), .B(new_n17734), .C(new_n17735), .Y(new_n17743));
  A2O1A1Ixp33_ASAP7_75t_L   g17487(.A1(\a[44] ), .A2(new_n17739), .B(new_n17740), .C(new_n17743), .Y(new_n17744));
  AND2x2_ASAP7_75t_L        g17488(.A(new_n17742), .B(new_n17744), .Y(new_n17745));
  XNOR2x2_ASAP7_75t_L       g17489(.A(new_n17654), .B(new_n17745), .Y(new_n17746));
  OR2x4_ASAP7_75t_L         g17490(.A(new_n17652), .B(new_n17746), .Y(new_n17747));
  NAND2xp33_ASAP7_75t_L     g17491(.A(new_n17652), .B(new_n17746), .Y(new_n17748));
  NAND2xp33_ASAP7_75t_L     g17492(.A(new_n17748), .B(new_n17747), .Y(new_n17749));
  NOR2xp33_ASAP7_75t_L      g17493(.A(new_n17646), .B(new_n17749), .Y(new_n17750));
  INVx1_ASAP7_75t_L         g17494(.A(new_n17750), .Y(new_n17751));
  NAND2xp33_ASAP7_75t_L     g17495(.A(new_n17646), .B(new_n17749), .Y(new_n17752));
  NAND2xp33_ASAP7_75t_L     g17496(.A(new_n17752), .B(new_n17751), .Y(new_n17753));
  XNOR2x2_ASAP7_75t_L       g17497(.A(new_n17645), .B(new_n17753), .Y(new_n17754));
  AO21x2_ASAP7_75t_L        g17498(.A1(new_n17501), .A2(new_n17510), .B(new_n17754), .Y(new_n17755));
  NAND3xp33_ASAP7_75t_L     g17499(.A(new_n17754), .B(new_n17510), .C(new_n17501), .Y(new_n17756));
  NAND2xp33_ASAP7_75t_L     g17500(.A(new_n17756), .B(new_n17755), .Y(new_n17757));
  NOR2xp33_ASAP7_75t_L      g17501(.A(new_n7552), .B(new_n4147), .Y(new_n17758));
  AOI221xp5_ASAP7_75t_L     g17502(.A1(\b[45] ), .A2(new_n4402), .B1(\b[46] ), .B2(new_n4155), .C(new_n17758), .Y(new_n17759));
  O2A1O1Ixp33_ASAP7_75t_L   g17503(.A1(new_n4150), .A2(new_n7560), .B(new_n17759), .C(new_n4145), .Y(new_n17760));
  INVx1_ASAP7_75t_L         g17504(.A(new_n17760), .Y(new_n17761));
  O2A1O1Ixp33_ASAP7_75t_L   g17505(.A1(new_n4150), .A2(new_n7560), .B(new_n17759), .C(\a[35] ), .Y(new_n17762));
  AO21x2_ASAP7_75t_L        g17506(.A1(\a[35] ), .A2(new_n17761), .B(new_n17762), .Y(new_n17763));
  NAND3xp33_ASAP7_75t_L     g17507(.A(new_n17755), .B(new_n17756), .C(new_n17763), .Y(new_n17764));
  INVx1_ASAP7_75t_L         g17508(.A(new_n17764), .Y(new_n17765));
  A2O1A1Ixp33_ASAP7_75t_L   g17509(.A1(\a[35] ), .A2(new_n17761), .B(new_n17762), .C(new_n17757), .Y(new_n17766));
  OAI21xp33_ASAP7_75t_L     g17510(.A1(new_n17757), .A2(new_n17765), .B(new_n17766), .Y(new_n17767));
  NAND2xp33_ASAP7_75t_L     g17511(.A(new_n17767), .B(new_n17639), .Y(new_n17768));
  NOR2xp33_ASAP7_75t_L      g17512(.A(new_n17767), .B(new_n17639), .Y(new_n17769));
  INVx1_ASAP7_75t_L         g17513(.A(new_n17769), .Y(new_n17770));
  OAI211xp5_ASAP7_75t_L     g17514(.A1(new_n17629), .A2(new_n17626), .B(new_n17768), .C(new_n17770), .Y(new_n17771));
  INVx1_ASAP7_75t_L         g17515(.A(new_n17768), .Y(new_n17772));
  INVx1_ASAP7_75t_L         g17516(.A(new_n17629), .Y(new_n17773));
  A2O1A1Ixp33_ASAP7_75t_L   g17517(.A1(new_n17627), .A2(new_n17773), .B(new_n17772), .C(new_n17770), .Y(new_n17774));
  NOR2xp33_ASAP7_75t_L      g17518(.A(new_n17772), .B(new_n17774), .Y(new_n17775));
  A2O1A1Ixp33_ASAP7_75t_L   g17519(.A1(new_n17628), .A2(new_n17771), .B(new_n17775), .C(new_n17615), .Y(new_n17776));
  INVx1_ASAP7_75t_L         g17520(.A(new_n17776), .Y(new_n17777));
  A2O1A1Ixp33_ASAP7_75t_L   g17521(.A1(new_n17623), .A2(new_n17622), .B(new_n17629), .C(new_n17771), .Y(new_n17778));
  A2O1A1Ixp33_ASAP7_75t_L   g17522(.A1(new_n17639), .A2(new_n17767), .B(new_n17774), .C(new_n17778), .Y(new_n17779));
  NOR2xp33_ASAP7_75t_L      g17523(.A(new_n17615), .B(new_n17779), .Y(new_n17780));
  O2A1O1Ixp33_ASAP7_75t_L   g17524(.A1(new_n17600), .A2(new_n17602), .B(new_n17604), .C(new_n17780), .Y(new_n17781));
  INVx1_ASAP7_75t_L         g17525(.A(new_n17781), .Y(new_n17782));
  NOR3xp33_ASAP7_75t_L      g17526(.A(new_n17605), .B(new_n17777), .C(new_n17780), .Y(new_n17783));
  O2A1O1Ixp33_ASAP7_75t_L   g17527(.A1(new_n17777), .A2(new_n17782), .B(new_n17605), .C(new_n17783), .Y(new_n17784));
  XOR2x2_ASAP7_75t_L        g17528(.A(new_n17784), .B(new_n17594), .Y(new_n17785));
  O2A1O1Ixp33_ASAP7_75t_L   g17529(.A1(new_n17581), .A2(new_n17582), .B(new_n17583), .C(new_n17785), .Y(new_n17786));
  INVx1_ASAP7_75t_L         g17530(.A(new_n17580), .Y(new_n17787));
  A2O1A1Ixp33_ASAP7_75t_L   g17531(.A1(new_n12986), .A2(new_n1216), .B(new_n17578), .C(new_n1206), .Y(new_n17788));
  A2O1A1Ixp33_ASAP7_75t_L   g17532(.A1(new_n17788), .A2(new_n17787), .B(new_n17582), .C(new_n17583), .Y(new_n17789));
  XNOR2x2_ASAP7_75t_L       g17533(.A(new_n17784), .B(new_n17594), .Y(new_n17790));
  NOR2xp33_ASAP7_75t_L      g17534(.A(new_n17789), .B(new_n17790), .Y(new_n17791));
  OAI21xp33_ASAP7_75t_L     g17535(.A1(new_n17791), .A2(new_n17786), .B(new_n17577), .Y(new_n17792));
  INVx1_ASAP7_75t_L         g17536(.A(new_n17581), .Y(new_n17793));
  A2O1A1Ixp33_ASAP7_75t_L   g17537(.A1(new_n17551), .A2(new_n17346), .B(new_n17347), .C(new_n17793), .Y(new_n17794));
  O2A1O1Ixp33_ASAP7_75t_L   g17538(.A1(new_n17556), .A2(new_n17555), .B(new_n17348), .C(new_n17793), .Y(new_n17795));
  A2O1A1Ixp33_ASAP7_75t_L   g17539(.A1(new_n17794), .A2(new_n17793), .B(new_n17795), .C(new_n17790), .Y(new_n17796));
  A2O1A1O1Ixp25_ASAP7_75t_L g17540(.A1(new_n12603), .A2(new_n14444), .B(new_n1210), .C(new_n1285), .D(new_n12956), .Y(new_n17797));
  A2O1A1O1Ixp25_ASAP7_75t_L g17541(.A1(new_n17579), .A2(new_n17797), .B(new_n17580), .C(new_n17794), .D(new_n17795), .Y(new_n17798));
  NAND2xp33_ASAP7_75t_L     g17542(.A(new_n17798), .B(new_n17785), .Y(new_n17799));
  NAND4xp25_ASAP7_75t_L     g17543(.A(new_n17796), .B(new_n17799), .C(new_n17573), .D(new_n17576), .Y(new_n17800));
  NAND2xp33_ASAP7_75t_L     g17544(.A(new_n17800), .B(new_n17792), .Y(new_n17801));
  A2O1A1Ixp33_ASAP7_75t_L   g17545(.A1(new_n17314), .A2(new_n17295), .B(new_n17313), .C(new_n17315), .Y(new_n17802));
  A2O1A1Ixp33_ASAP7_75t_L   g17546(.A1(new_n17309), .A2(new_n17802), .B(new_n17320), .C(new_n17567), .Y(new_n17803));
  NAND3xp33_ASAP7_75t_L     g17547(.A(new_n17803), .B(new_n17565), .C(new_n17800), .Y(new_n17804));
  O2A1O1Ixp33_ASAP7_75t_L   g17548(.A1(new_n17786), .A2(new_n17791), .B(new_n17577), .C(new_n17804), .Y(new_n17805));
  O2A1O1Ixp33_ASAP7_75t_L   g17549(.A1(new_n17566), .A2(new_n17569), .B(new_n17801), .C(new_n17805), .Y(\f[80] ));
  INVx1_ASAP7_75t_L         g17550(.A(new_n17317), .Y(new_n17807));
  A2O1A1Ixp33_ASAP7_75t_L   g17551(.A1(new_n17319), .A2(new_n17807), .B(new_n17563), .C(new_n17565), .Y(new_n17808));
  NAND2xp33_ASAP7_75t_L     g17552(.A(new_n17799), .B(new_n17796), .Y(new_n17809));
  O2A1O1Ixp33_ASAP7_75t_L   g17553(.A1(new_n17574), .A2(new_n17335), .B(new_n17576), .C(new_n17809), .Y(new_n17810));
  A2O1A1O1Ixp25_ASAP7_75t_L g17554(.A1(new_n17550), .A2(new_n17532), .B(new_n17546), .C(new_n17346), .D(new_n17347), .Y(new_n17811));
  A2O1A1Ixp33_ASAP7_75t_L   g17555(.A1(new_n17797), .A2(new_n17579), .B(new_n17580), .C(new_n17811), .Y(new_n17812));
  A2O1A1Ixp33_ASAP7_75t_L   g17556(.A1(new_n17811), .A2(new_n17812), .B(new_n17785), .C(new_n17794), .Y(new_n17813));
  INVx1_ASAP7_75t_L         g17557(.A(new_n17593), .Y(new_n17814));
  INVx1_ASAP7_75t_L         g17558(.A(new_n12961), .Y(new_n17815));
  NOR2xp33_ASAP7_75t_L      g17559(.A(new_n12956), .B(new_n1518), .Y(new_n17816));
  AOI221xp5_ASAP7_75t_L     g17560(.A1(\b[61] ), .A2(new_n1659), .B1(\b[62] ), .B2(new_n1507), .C(new_n17816), .Y(new_n17817));
  O2A1O1Ixp33_ASAP7_75t_L   g17561(.A1(new_n1521), .A2(new_n17815), .B(new_n17817), .C(new_n1501), .Y(new_n17818));
  INVx1_ASAP7_75t_L         g17562(.A(new_n17818), .Y(new_n17819));
  O2A1O1Ixp33_ASAP7_75t_L   g17563(.A1(new_n1521), .A2(new_n17815), .B(new_n17817), .C(\a[20] ), .Y(new_n17820));
  AOI21xp33_ASAP7_75t_L     g17564(.A1(new_n17819), .A2(\a[20] ), .B(new_n17820), .Y(new_n17821));
  INVx1_ASAP7_75t_L         g17565(.A(new_n17821), .Y(new_n17822));
  O2A1O1Ixp33_ASAP7_75t_L   g17566(.A1(new_n17590), .A2(new_n17784), .B(new_n17814), .C(new_n17822), .Y(new_n17823));
  OAI21xp33_ASAP7_75t_L     g17567(.A1(new_n17590), .A2(new_n17784), .B(new_n17814), .Y(new_n17824));
  INVx1_ASAP7_75t_L         g17568(.A(new_n17820), .Y(new_n17825));
  O2A1O1Ixp33_ASAP7_75t_L   g17569(.A1(new_n17818), .A2(new_n1501), .B(new_n17825), .C(new_n17824), .Y(new_n17826));
  OAI22xp33_ASAP7_75t_L     g17570(.A1(new_n2089), .A2(new_n11303), .B1(new_n11591), .B2(new_n1962), .Y(new_n17827));
  AOI221xp5_ASAP7_75t_L     g17571(.A1(new_n1955), .A2(\b[60] ), .B1(new_n1964), .B2(new_n13839), .C(new_n17827), .Y(new_n17828));
  XNOR2x2_ASAP7_75t_L       g17572(.A(new_n1952), .B(new_n17828), .Y(new_n17829));
  INVx1_ASAP7_75t_L         g17573(.A(new_n17829), .Y(new_n17830));
  AOI211xp5_ASAP7_75t_L     g17574(.A1(new_n17781), .A2(new_n17776), .B(new_n17830), .C(new_n17602), .Y(new_n17831));
  A2O1A1Ixp33_ASAP7_75t_L   g17575(.A1(new_n17781), .A2(new_n17776), .B(new_n17602), .C(new_n17830), .Y(new_n17832));
  INVx1_ASAP7_75t_L         g17576(.A(new_n17832), .Y(new_n17833));
  OAI22xp33_ASAP7_75t_L     g17577(.A1(new_n3133), .A2(new_n9355), .B1(new_n9683), .B2(new_n2925), .Y(new_n17834));
  AOI221xp5_ASAP7_75t_L     g17578(.A1(new_n2938), .A2(\b[54] ), .B1(new_n2932), .B2(new_n9717), .C(new_n17834), .Y(new_n17835));
  XNOR2x2_ASAP7_75t_L       g17579(.A(new_n2928), .B(new_n17835), .Y(new_n17836));
  AND3x1_ASAP7_75t_L        g17580(.A(new_n17771), .B(new_n17836), .C(new_n17623), .Y(new_n17837));
  A2O1A1Ixp33_ASAP7_75t_L   g17581(.A1(new_n17623), .A2(new_n17622), .B(new_n17629), .C(new_n17770), .Y(new_n17838));
  O2A1O1Ixp33_ASAP7_75t_L   g17582(.A1(new_n17772), .A2(new_n17838), .B(new_n17623), .C(new_n17836), .Y(new_n17839));
  A2O1A1Ixp33_ASAP7_75t_L   g17583(.A1(new_n17742), .A2(new_n17744), .B(new_n17654), .C(new_n17747), .Y(new_n17840));
  INVx1_ASAP7_75t_L         g17584(.A(new_n17743), .Y(new_n17841));
  INVx1_ASAP7_75t_L         g17585(.A(new_n17741), .Y(new_n17842));
  A2O1A1O1Ixp25_ASAP7_75t_L g17586(.A1(new_n17731), .A2(\a[47] ), .B(new_n17728), .C(new_n17721), .D(new_n17722), .Y(new_n17843));
  INVx1_ASAP7_75t_L         g17587(.A(new_n17843), .Y(new_n17844));
  OAI21xp33_ASAP7_75t_L     g17588(.A1(new_n17407), .A2(new_n17668), .B(new_n17684), .Y(new_n17845));
  A2O1A1Ixp33_ASAP7_75t_L   g17589(.A1(new_n17673), .A2(new_n17680), .B(new_n17678), .C(new_n17845), .Y(new_n17846));
  A2O1A1Ixp33_ASAP7_75t_L   g17590(.A1(new_n2679), .A2(new_n11351), .B(new_n17691), .C(new_n11048), .Y(new_n17847));
  O2A1O1Ixp33_ASAP7_75t_L   g17591(.A1(new_n17693), .A2(new_n11048), .B(new_n17847), .C(new_n17688), .Y(new_n17848));
  NOR2xp33_ASAP7_75t_L      g17592(.A(new_n1349), .B(new_n13030), .Y(new_n17849));
  A2O1A1Ixp33_ASAP7_75t_L   g17593(.A1(new_n13028), .A2(\b[18] ), .B(new_n17849), .C(new_n1206), .Y(new_n17850));
  O2A1O1Ixp33_ASAP7_75t_L   g17594(.A1(new_n12669), .A2(new_n12671), .B(\b[18] ), .C(new_n17849), .Y(new_n17851));
  NAND2xp33_ASAP7_75t_L     g17595(.A(\a[17] ), .B(new_n17851), .Y(new_n17852));
  NAND2xp33_ASAP7_75t_L     g17596(.A(new_n17850), .B(new_n17852), .Y(new_n17853));
  O2A1O1Ixp33_ASAP7_75t_L   g17597(.A1(new_n1349), .A2(new_n12672), .B(new_n17681), .C(new_n17853), .Y(new_n17854));
  INVx1_ASAP7_75t_L         g17598(.A(new_n17854), .Y(new_n17855));
  NAND2xp33_ASAP7_75t_L     g17599(.A(new_n17668), .B(new_n17853), .Y(new_n17856));
  AND2x2_ASAP7_75t_L        g17600(.A(new_n17856), .B(new_n17855), .Y(new_n17857));
  INVx1_ASAP7_75t_L         g17601(.A(new_n17857), .Y(new_n17858));
  NOR2xp33_ASAP7_75t_L      g17602(.A(new_n1745), .B(new_n12318), .Y(new_n17859));
  AOI221xp5_ASAP7_75t_L     g17603(.A1(new_n11995), .A2(\b[21] ), .B1(new_n13314), .B2(\b[19] ), .C(new_n17859), .Y(new_n17860));
  INVx1_ASAP7_75t_L         g17604(.A(new_n17860), .Y(new_n17861));
  A2O1A1Ixp33_ASAP7_75t_L   g17605(.A1(new_n2836), .A2(new_n11997), .B(new_n17861), .C(\a[62] ), .Y(new_n17862));
  INVx1_ASAP7_75t_L         g17606(.A(new_n17862), .Y(new_n17863));
  O2A1O1Ixp33_ASAP7_75t_L   g17607(.A1(new_n11998), .A2(new_n1901), .B(new_n17860), .C(\a[62] ), .Y(new_n17864));
  INVx1_ASAP7_75t_L         g17608(.A(new_n17864), .Y(new_n17865));
  O2A1O1Ixp33_ASAP7_75t_L   g17609(.A1(new_n11987), .A2(new_n17863), .B(new_n17865), .C(new_n17858), .Y(new_n17866));
  O2A1O1Ixp33_ASAP7_75t_L   g17610(.A1(new_n11987), .A2(new_n17863), .B(new_n17865), .C(new_n17857), .Y(new_n17867));
  INVx1_ASAP7_75t_L         g17611(.A(new_n17867), .Y(new_n17868));
  O2A1O1Ixp33_ASAP7_75t_L   g17612(.A1(new_n17858), .A2(new_n17866), .B(new_n17868), .C(new_n17684), .Y(new_n17869));
  O2A1O1Ixp33_ASAP7_75t_L   g17613(.A1(new_n17682), .A2(new_n17677), .B(new_n17676), .C(new_n17869), .Y(new_n17870));
  O2A1O1Ixp33_ASAP7_75t_L   g17614(.A1(new_n17858), .A2(new_n17866), .B(new_n17868), .C(new_n17683), .Y(new_n17871));
  NOR2xp33_ASAP7_75t_L      g17615(.A(new_n2045), .B(new_n11354), .Y(new_n17872));
  AOI221xp5_ASAP7_75t_L     g17616(.A1(\b[24] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[23] ), .C(new_n17872), .Y(new_n17873));
  O2A1O1Ixp33_ASAP7_75t_L   g17617(.A1(new_n11053), .A2(new_n2853), .B(new_n17873), .C(new_n11048), .Y(new_n17874));
  O2A1O1Ixp33_ASAP7_75t_L   g17618(.A1(new_n11053), .A2(new_n2853), .B(new_n17873), .C(\a[59] ), .Y(new_n17875));
  INVx1_ASAP7_75t_L         g17619(.A(new_n17875), .Y(new_n17876));
  OAI21xp33_ASAP7_75t_L     g17620(.A1(new_n11048), .A2(new_n17874), .B(new_n17876), .Y(new_n17877));
  OR3x1_ASAP7_75t_L         g17621(.A(new_n17870), .B(new_n17871), .C(new_n17877), .Y(new_n17878));
  INVx1_ASAP7_75t_L         g17622(.A(new_n17869), .Y(new_n17879));
  A2O1A1Ixp33_ASAP7_75t_L   g17623(.A1(new_n17879), .A2(new_n17683), .B(new_n17871), .C(new_n17877), .Y(new_n17880));
  AND2x2_ASAP7_75t_L        g17624(.A(new_n17880), .B(new_n17878), .Y(new_n17881));
  A2O1A1Ixp33_ASAP7_75t_L   g17625(.A1(new_n17687), .A2(new_n17846), .B(new_n17848), .C(new_n17881), .Y(new_n17882));
  A2O1A1O1Ixp25_ASAP7_75t_L g17626(.A1(new_n17404), .A2(new_n17416), .B(new_n17408), .C(new_n17846), .D(new_n17848), .Y(new_n17883));
  INVx1_ASAP7_75t_L         g17627(.A(new_n17881), .Y(new_n17884));
  NAND2xp33_ASAP7_75t_L     g17628(.A(new_n17884), .B(new_n17883), .Y(new_n17885));
  NAND2xp33_ASAP7_75t_L     g17629(.A(new_n17882), .B(new_n17885), .Y(new_n17886));
  NOR2xp33_ASAP7_75t_L      g17630(.A(new_n2703), .B(new_n10388), .Y(new_n17887));
  AOI221xp5_ASAP7_75t_L     g17631(.A1(new_n10086), .A2(\b[27] ), .B1(new_n11361), .B2(\b[25] ), .C(new_n17887), .Y(new_n17888));
  O2A1O1Ixp33_ASAP7_75t_L   g17632(.A1(new_n10088), .A2(new_n2889), .B(new_n17888), .C(new_n10083), .Y(new_n17889));
  O2A1O1Ixp33_ASAP7_75t_L   g17633(.A1(new_n10088), .A2(new_n2889), .B(new_n17888), .C(\a[56] ), .Y(new_n17890));
  INVx1_ASAP7_75t_L         g17634(.A(new_n17890), .Y(new_n17891));
  O2A1O1Ixp33_ASAP7_75t_L   g17635(.A1(new_n17889), .A2(new_n10083), .B(new_n17891), .C(new_n17886), .Y(new_n17892));
  INVx1_ASAP7_75t_L         g17636(.A(new_n17886), .Y(new_n17893));
  O2A1O1Ixp33_ASAP7_75t_L   g17637(.A1(new_n17889), .A2(new_n10083), .B(new_n17891), .C(new_n17893), .Y(new_n17894));
  INVx1_ASAP7_75t_L         g17638(.A(new_n17894), .Y(new_n17895));
  A2O1A1O1Ixp25_ASAP7_75t_L g17639(.A1(new_n17156), .A2(new_n17149), .B(new_n17417), .C(new_n17427), .D(new_n17696), .Y(new_n17896));
  A2O1A1O1Ixp25_ASAP7_75t_L g17640(.A1(new_n17663), .A2(\a[56] ), .B(new_n17664), .C(new_n17697), .D(new_n17896), .Y(new_n17897));
  OAI211xp5_ASAP7_75t_L     g17641(.A1(new_n17892), .A2(new_n17886), .B(new_n17895), .C(new_n17897), .Y(new_n17898));
  INVx1_ASAP7_75t_L         g17642(.A(new_n17892), .Y(new_n17899));
  AO21x2_ASAP7_75t_L        g17643(.A1(new_n17893), .A2(new_n17899), .B(new_n17894), .Y(new_n17900));
  A2O1A1Ixp33_ASAP7_75t_L   g17644(.A1(new_n17697), .A2(new_n17665), .B(new_n17896), .C(new_n17900), .Y(new_n17901));
  NAND2xp33_ASAP7_75t_L     g17645(.A(new_n17898), .B(new_n17901), .Y(new_n17902));
  NOR2xp33_ASAP7_75t_L      g17646(.A(new_n3098), .B(new_n10400), .Y(new_n17903));
  AOI221xp5_ASAP7_75t_L     g17647(.A1(new_n9102), .A2(\b[30] ), .B1(new_n10398), .B2(\b[28] ), .C(new_n17903), .Y(new_n17904));
  O2A1O1Ixp33_ASAP7_75t_L   g17648(.A1(new_n9104), .A2(new_n3464), .B(new_n17904), .C(new_n9099), .Y(new_n17905));
  O2A1O1Ixp33_ASAP7_75t_L   g17649(.A1(new_n9104), .A2(new_n3464), .B(new_n17904), .C(\a[53] ), .Y(new_n17906));
  INVx1_ASAP7_75t_L         g17650(.A(new_n17906), .Y(new_n17907));
  O2A1O1Ixp33_ASAP7_75t_L   g17651(.A1(new_n17905), .A2(new_n9099), .B(new_n17907), .C(new_n17902), .Y(new_n17908));
  INVx1_ASAP7_75t_L         g17652(.A(new_n17902), .Y(new_n17909));
  O2A1O1Ixp33_ASAP7_75t_L   g17653(.A1(new_n17905), .A2(new_n9099), .B(new_n17907), .C(new_n17909), .Y(new_n17910));
  INVx1_ASAP7_75t_L         g17654(.A(new_n17910), .Y(new_n17911));
  A2O1A1O1Ixp25_ASAP7_75t_L g17655(.A1(new_n17658), .A2(new_n17441), .B(new_n17431), .C(new_n17432), .D(new_n17698), .Y(new_n17912));
  INVx1_ASAP7_75t_L         g17656(.A(new_n17699), .Y(new_n17913));
  A2O1A1O1Ixp25_ASAP7_75t_L g17657(.A1(new_n17709), .A2(\a[53] ), .B(new_n17703), .C(new_n17913), .D(new_n17912), .Y(new_n17914));
  OAI211xp5_ASAP7_75t_L     g17658(.A1(new_n17908), .A2(new_n17902), .B(new_n17911), .C(new_n17914), .Y(new_n17915));
  INVx1_ASAP7_75t_L         g17659(.A(new_n17908), .Y(new_n17916));
  INVx1_ASAP7_75t_L         g17660(.A(new_n17914), .Y(new_n17917));
  A2O1A1Ixp33_ASAP7_75t_L   g17661(.A1(new_n17916), .A2(new_n17909), .B(new_n17910), .C(new_n17917), .Y(new_n17918));
  NAND2xp33_ASAP7_75t_L     g17662(.A(new_n17918), .B(new_n17915), .Y(new_n17919));
  NOR2xp33_ASAP7_75t_L      g17663(.A(new_n3891), .B(new_n10065), .Y(new_n17920));
  AOI221xp5_ASAP7_75t_L     g17664(.A1(new_n8175), .A2(\b[33] ), .B1(new_n8484), .B2(\b[31] ), .C(new_n17920), .Y(new_n17921));
  O2A1O1Ixp33_ASAP7_75t_L   g17665(.A1(new_n8176), .A2(new_n4108), .B(new_n17921), .C(new_n8172), .Y(new_n17922));
  NOR2xp33_ASAP7_75t_L      g17666(.A(new_n8172), .B(new_n17922), .Y(new_n17923));
  O2A1O1Ixp33_ASAP7_75t_L   g17667(.A1(new_n8176), .A2(new_n4108), .B(new_n17921), .C(\a[50] ), .Y(new_n17924));
  NOR2xp33_ASAP7_75t_L      g17668(.A(new_n17924), .B(new_n17923), .Y(new_n17925));
  INVx1_ASAP7_75t_L         g17669(.A(new_n17707), .Y(new_n17926));
  INVx1_ASAP7_75t_L         g17670(.A(new_n17718), .Y(new_n17927));
  O2A1O1Ixp33_ASAP7_75t_L   g17671(.A1(new_n17711), .A2(new_n17657), .B(new_n17927), .C(new_n17926), .Y(new_n17928));
  XNOR2x2_ASAP7_75t_L       g17672(.A(new_n17925), .B(new_n17928), .Y(new_n17929));
  XOR2x2_ASAP7_75t_L        g17673(.A(new_n17919), .B(new_n17929), .Y(new_n17930));
  NOR2xp33_ASAP7_75t_L      g17674(.A(new_n4613), .B(new_n7318), .Y(new_n17931));
  AOI221xp5_ASAP7_75t_L     g17675(.A1(new_n7333), .A2(\b[35] ), .B1(new_n7609), .B2(\b[34] ), .C(new_n17931), .Y(new_n17932));
  O2A1O1Ixp33_ASAP7_75t_L   g17676(.A1(new_n7321), .A2(new_n4622), .B(new_n17932), .C(new_n7316), .Y(new_n17933));
  INVx1_ASAP7_75t_L         g17677(.A(new_n17933), .Y(new_n17934));
  O2A1O1Ixp33_ASAP7_75t_L   g17678(.A1(new_n7321), .A2(new_n4622), .B(new_n17932), .C(\a[47] ), .Y(new_n17935));
  A2O1A1Ixp33_ASAP7_75t_L   g17679(.A1(\a[47] ), .A2(new_n17934), .B(new_n17935), .C(new_n17930), .Y(new_n17936));
  INVx1_ASAP7_75t_L         g17680(.A(new_n17936), .Y(new_n17937));
  AOI211xp5_ASAP7_75t_L     g17681(.A1(new_n17934), .A2(\a[47] ), .B(new_n17935), .C(new_n17930), .Y(new_n17938));
  NOR2xp33_ASAP7_75t_L      g17682(.A(new_n17938), .B(new_n17937), .Y(new_n17939));
  NOR2xp33_ASAP7_75t_L      g17683(.A(new_n17844), .B(new_n17939), .Y(new_n17940));
  NOR3xp33_ASAP7_75t_L      g17684(.A(new_n17937), .B(new_n17938), .C(new_n17843), .Y(new_n17941));
  NOR2xp33_ASAP7_75t_L      g17685(.A(new_n17941), .B(new_n17940), .Y(new_n17942));
  NOR2xp33_ASAP7_75t_L      g17686(.A(new_n5311), .B(new_n7304), .Y(new_n17943));
  AOI221xp5_ASAP7_75t_L     g17687(.A1(\b[37] ), .A2(new_n6742), .B1(\b[39] ), .B2(new_n6442), .C(new_n17943), .Y(new_n17944));
  O2A1O1Ixp33_ASAP7_75t_L   g17688(.A1(new_n6443), .A2(new_n5578), .B(new_n17944), .C(new_n6439), .Y(new_n17945));
  INVx1_ASAP7_75t_L         g17689(.A(new_n17945), .Y(new_n17946));
  O2A1O1Ixp33_ASAP7_75t_L   g17690(.A1(new_n6443), .A2(new_n5578), .B(new_n17944), .C(\a[44] ), .Y(new_n17947));
  A2O1A1Ixp33_ASAP7_75t_L   g17691(.A1(\a[44] ), .A2(new_n17946), .B(new_n17947), .C(new_n17942), .Y(new_n17948));
  INVx1_ASAP7_75t_L         g17692(.A(new_n17947), .Y(new_n17949));
  O2A1O1Ixp33_ASAP7_75t_L   g17693(.A1(new_n17945), .A2(new_n6439), .B(new_n17949), .C(new_n17942), .Y(new_n17950));
  AOI21xp33_ASAP7_75t_L     g17694(.A1(new_n17948), .A2(new_n17942), .B(new_n17950), .Y(new_n17951));
  A2O1A1Ixp33_ASAP7_75t_L   g17695(.A1(new_n17841), .A2(new_n17842), .B(new_n17733), .C(new_n17951), .Y(new_n17952));
  INVx1_ASAP7_75t_L         g17696(.A(new_n17735), .Y(new_n17953));
  A2O1A1Ixp33_ASAP7_75t_L   g17697(.A1(new_n17953), .A2(new_n17655), .B(new_n17741), .C(new_n17734), .Y(new_n17954));
  INVx1_ASAP7_75t_L         g17698(.A(new_n17954), .Y(new_n17955));
  A2O1A1Ixp33_ASAP7_75t_L   g17699(.A1(new_n17948), .A2(new_n17942), .B(new_n17950), .C(new_n17955), .Y(new_n17956));
  AND2x2_ASAP7_75t_L        g17700(.A(new_n17956), .B(new_n17952), .Y(new_n17957));
  NOR2xp33_ASAP7_75t_L      g17701(.A(new_n6378), .B(new_n5641), .Y(new_n17958));
  AOI221xp5_ASAP7_75t_L     g17702(.A1(\b[40] ), .A2(new_n5920), .B1(\b[41] ), .B2(new_n5623), .C(new_n17958), .Y(new_n17959));
  O2A1O1Ixp33_ASAP7_75t_L   g17703(.A1(new_n5630), .A2(new_n6386), .B(new_n17959), .C(new_n5626), .Y(new_n17960));
  O2A1O1Ixp33_ASAP7_75t_L   g17704(.A1(new_n5630), .A2(new_n6386), .B(new_n17959), .C(\a[41] ), .Y(new_n17961));
  INVx1_ASAP7_75t_L         g17705(.A(new_n17961), .Y(new_n17962));
  OAI21xp33_ASAP7_75t_L     g17706(.A1(new_n5626), .A2(new_n17960), .B(new_n17962), .Y(new_n17963));
  XNOR2x2_ASAP7_75t_L       g17707(.A(new_n17963), .B(new_n17957), .Y(new_n17964));
  XNOR2x2_ASAP7_75t_L       g17708(.A(new_n17964), .B(new_n17840), .Y(new_n17965));
  NOR2xp33_ASAP7_75t_L      g17709(.A(new_n7249), .B(new_n4908), .Y(new_n17966));
  AOI221xp5_ASAP7_75t_L     g17710(.A1(\b[43] ), .A2(new_n5139), .B1(\b[44] ), .B2(new_n4916), .C(new_n17966), .Y(new_n17967));
  O2A1O1Ixp33_ASAP7_75t_L   g17711(.A1(new_n4911), .A2(new_n7255), .B(new_n17967), .C(new_n4906), .Y(new_n17968));
  O2A1O1Ixp33_ASAP7_75t_L   g17712(.A1(new_n4911), .A2(new_n7255), .B(new_n17967), .C(\a[38] ), .Y(new_n17969));
  INVx1_ASAP7_75t_L         g17713(.A(new_n17969), .Y(new_n17970));
  O2A1O1Ixp33_ASAP7_75t_L   g17714(.A1(new_n17968), .A2(new_n4906), .B(new_n17970), .C(new_n17965), .Y(new_n17971));
  INVx1_ASAP7_75t_L         g17715(.A(new_n17968), .Y(new_n17972));
  A2O1A1Ixp33_ASAP7_75t_L   g17716(.A1(\a[38] ), .A2(new_n17972), .B(new_n17969), .C(new_n17965), .Y(new_n17973));
  OAI21xp33_ASAP7_75t_L     g17717(.A1(new_n17965), .A2(new_n17971), .B(new_n17973), .Y(new_n17974));
  A2O1A1O1Ixp25_ASAP7_75t_L g17718(.A1(new_n17643), .A2(\a[38] ), .B(new_n17644), .C(new_n17752), .D(new_n17750), .Y(new_n17975));
  INVx1_ASAP7_75t_L         g17719(.A(new_n17975), .Y(new_n17976));
  NOR2xp33_ASAP7_75t_L      g17720(.A(new_n17976), .B(new_n17974), .Y(new_n17977));
  O2A1O1Ixp33_ASAP7_75t_L   g17721(.A1(new_n17965), .A2(new_n17971), .B(new_n17973), .C(new_n17975), .Y(new_n17978));
  NOR2xp33_ASAP7_75t_L      g17722(.A(new_n17978), .B(new_n17977), .Y(new_n17979));
  NOR2xp33_ASAP7_75t_L      g17723(.A(new_n7860), .B(new_n4147), .Y(new_n17980));
  AOI221xp5_ASAP7_75t_L     g17724(.A1(\b[46] ), .A2(new_n4402), .B1(\b[47] ), .B2(new_n4155), .C(new_n17980), .Y(new_n17981));
  O2A1O1Ixp33_ASAP7_75t_L   g17725(.A1(new_n4150), .A2(new_n7868), .B(new_n17981), .C(new_n4145), .Y(new_n17982));
  INVx1_ASAP7_75t_L         g17726(.A(new_n17982), .Y(new_n17983));
  O2A1O1Ixp33_ASAP7_75t_L   g17727(.A1(new_n4150), .A2(new_n7868), .B(new_n17981), .C(\a[35] ), .Y(new_n17984));
  A2O1A1Ixp33_ASAP7_75t_L   g17728(.A1(\a[35] ), .A2(new_n17983), .B(new_n17984), .C(new_n17979), .Y(new_n17985));
  INVx1_ASAP7_75t_L         g17729(.A(new_n17985), .Y(new_n17986));
  A2O1A1Ixp33_ASAP7_75t_L   g17730(.A1(new_n17983), .A2(\a[35] ), .B(new_n17984), .C(new_n17985), .Y(new_n17987));
  OAI31xp33_ASAP7_75t_L     g17731(.A1(new_n17977), .A2(new_n17986), .A3(new_n17978), .B(new_n17987), .Y(new_n17988));
  A2O1A1Ixp33_ASAP7_75t_L   g17732(.A1(new_n17510), .A2(new_n17501), .B(new_n17754), .C(new_n17764), .Y(new_n17989));
  NOR2xp33_ASAP7_75t_L      g17733(.A(new_n17989), .B(new_n17988), .Y(new_n17990));
  INVx1_ASAP7_75t_L         g17734(.A(new_n17984), .Y(new_n17991));
  O2A1O1Ixp33_ASAP7_75t_L   g17735(.A1(new_n17982), .A2(new_n4145), .B(new_n17991), .C(new_n17979), .Y(new_n17992));
  A2O1A1Ixp33_ASAP7_75t_L   g17736(.A1(new_n17985), .A2(new_n17979), .B(new_n17992), .C(new_n17989), .Y(new_n17993));
  INVx1_ASAP7_75t_L         g17737(.A(new_n17993), .Y(new_n17994));
  NOR2xp33_ASAP7_75t_L      g17738(.A(new_n17994), .B(new_n17990), .Y(new_n17995));
  OAI22xp33_ASAP7_75t_L     g17739(.A1(new_n3703), .A2(new_n8427), .B1(new_n8755), .B2(new_n3509), .Y(new_n17996));
  AOI221xp5_ASAP7_75t_L     g17740(.A1(new_n3503), .A2(\b[51] ), .B1(new_n3505), .B2(new_n8790), .C(new_n17996), .Y(new_n17997));
  XNOR2x2_ASAP7_75t_L       g17741(.A(new_n3493), .B(new_n17997), .Y(new_n17998));
  O2A1O1Ixp33_ASAP7_75t_L   g17742(.A1(new_n17636), .A2(new_n17638), .B(new_n17768), .C(new_n17998), .Y(new_n17999));
  INVx1_ASAP7_75t_L         g17743(.A(new_n17998), .Y(new_n18000));
  INVx1_ASAP7_75t_L         g17744(.A(new_n17637), .Y(new_n18001));
  A2O1A1Ixp33_ASAP7_75t_L   g17745(.A1(new_n17521), .A2(new_n18001), .B(new_n17636), .C(new_n17768), .Y(new_n18002));
  NOR2xp33_ASAP7_75t_L      g17746(.A(new_n18000), .B(new_n18002), .Y(new_n18003));
  NOR2xp33_ASAP7_75t_L      g17747(.A(new_n17999), .B(new_n18003), .Y(new_n18004));
  XOR2x2_ASAP7_75t_L        g17748(.A(new_n17995), .B(new_n18004), .Y(new_n18005));
  OR3x1_ASAP7_75t_L         g17749(.A(new_n17837), .B(new_n18005), .C(new_n17839), .Y(new_n18006));
  OAI21xp33_ASAP7_75t_L     g17750(.A1(new_n17839), .A2(new_n17837), .B(new_n18005), .Y(new_n18007));
  NAND2xp33_ASAP7_75t_L     g17751(.A(new_n18007), .B(new_n18006), .Y(new_n18008));
  INVx1_ASAP7_75t_L         g17752(.A(new_n18008), .Y(new_n18009));
  OAI22xp33_ASAP7_75t_L     g17753(.A1(new_n2572), .A2(new_n10309), .B1(new_n10332), .B2(new_n2410), .Y(new_n18010));
  AOI221xp5_ASAP7_75t_L     g17754(.A1(new_n2423), .A2(\b[57] ), .B1(new_n2417), .B2(new_n10991), .C(new_n18010), .Y(new_n18011));
  XNOR2x2_ASAP7_75t_L       g17755(.A(new_n2413), .B(new_n18011), .Y(new_n18012));
  INVx1_ASAP7_75t_L         g17756(.A(new_n18012), .Y(new_n18013));
  A2O1A1Ixp33_ASAP7_75t_L   g17757(.A1(new_n17779), .A2(new_n17615), .B(new_n17614), .C(new_n18013), .Y(new_n18014));
  INVx1_ASAP7_75t_L         g17758(.A(new_n18014), .Y(new_n18015));
  NOR3xp33_ASAP7_75t_L      g17759(.A(new_n17777), .B(new_n18013), .C(new_n17614), .Y(new_n18016));
  NOR3xp33_ASAP7_75t_L      g17760(.A(new_n18016), .B(new_n18015), .C(new_n18009), .Y(new_n18017));
  A2O1A1O1Ixp25_ASAP7_75t_L g17761(.A1(new_n17771), .A2(new_n17628), .B(new_n17775), .C(new_n17615), .D(new_n17614), .Y(new_n18018));
  NAND2xp33_ASAP7_75t_L     g17762(.A(new_n18012), .B(new_n18018), .Y(new_n18019));
  NAND3xp33_ASAP7_75t_L     g17763(.A(new_n18009), .B(new_n18014), .C(new_n18019), .Y(new_n18020));
  A2O1A1Ixp33_ASAP7_75t_L   g17764(.A1(new_n18007), .A2(new_n18006), .B(new_n18017), .C(new_n18020), .Y(new_n18021));
  NOR3xp33_ASAP7_75t_L      g17765(.A(new_n18021), .B(new_n17833), .C(new_n17831), .Y(new_n18022));
  INVx1_ASAP7_75t_L         g17766(.A(new_n17831), .Y(new_n18023));
  OAI21xp33_ASAP7_75t_L     g17767(.A1(new_n18015), .A2(new_n18016), .B(new_n18008), .Y(new_n18024));
  AND2x2_ASAP7_75t_L        g17768(.A(new_n18020), .B(new_n18024), .Y(new_n18025));
  AOI21xp33_ASAP7_75t_L     g17769(.A1(new_n18023), .A2(new_n17832), .B(new_n18025), .Y(new_n18026));
  NOR2xp33_ASAP7_75t_L      g17770(.A(new_n18026), .B(new_n18022), .Y(new_n18027));
  OAI21xp33_ASAP7_75t_L     g17771(.A1(new_n17823), .A2(new_n17826), .B(new_n18027), .Y(new_n18028));
  O2A1O1Ixp33_ASAP7_75t_L   g17772(.A1(new_n17590), .A2(new_n17784), .B(new_n17814), .C(new_n17821), .Y(new_n18029));
  INVx1_ASAP7_75t_L         g17773(.A(new_n17823), .Y(new_n18030));
  NAND3xp33_ASAP7_75t_L     g17774(.A(new_n18025), .B(new_n17832), .C(new_n18023), .Y(new_n18031));
  OAI21xp33_ASAP7_75t_L     g17775(.A1(new_n17831), .A2(new_n17833), .B(new_n18021), .Y(new_n18032));
  NAND2xp33_ASAP7_75t_L     g17776(.A(new_n18032), .B(new_n18031), .Y(new_n18033));
  OAI211xp5_ASAP7_75t_L     g17777(.A1(new_n17821), .A2(new_n18029), .B(new_n18033), .C(new_n18030), .Y(new_n18034));
  NAND3xp33_ASAP7_75t_L     g17778(.A(new_n18034), .B(new_n18028), .C(new_n17813), .Y(new_n18035));
  O2A1O1Ixp33_ASAP7_75t_L   g17779(.A1(new_n17795), .A2(new_n17793), .B(new_n17790), .C(new_n17582), .Y(new_n18036));
  O2A1O1Ixp33_ASAP7_75t_L   g17780(.A1(new_n17821), .A2(new_n18029), .B(new_n18030), .C(new_n18033), .Y(new_n18037));
  NOR3xp33_ASAP7_75t_L      g17781(.A(new_n18027), .B(new_n17826), .C(new_n17823), .Y(new_n18038));
  OAI21xp33_ASAP7_75t_L     g17782(.A1(new_n18037), .A2(new_n18038), .B(new_n18036), .Y(new_n18039));
  NAND2xp33_ASAP7_75t_L     g17783(.A(new_n18035), .B(new_n18039), .Y(new_n18040));
  NAND2xp33_ASAP7_75t_L     g17784(.A(new_n18028), .B(new_n18034), .Y(new_n18041));
  A2O1A1Ixp33_ASAP7_75t_L   g17785(.A1(new_n17789), .A2(new_n17790), .B(new_n17582), .C(new_n18041), .Y(new_n18042));
  A2O1A1O1Ixp25_ASAP7_75t_L g17786(.A1(new_n17570), .A2(new_n17567), .B(new_n17566), .C(new_n17801), .D(new_n17810), .Y(new_n18043));
  A2O1A1Ixp33_ASAP7_75t_L   g17787(.A1(new_n18028), .A2(new_n18034), .B(new_n17813), .C(new_n18043), .Y(new_n18044));
  O2A1O1Ixp33_ASAP7_75t_L   g17788(.A1(new_n17582), .A2(new_n17786), .B(new_n18042), .C(new_n18044), .Y(new_n18045));
  A2O1A1O1Ixp25_ASAP7_75t_L g17789(.A1(new_n17808), .A2(new_n17801), .B(new_n17810), .C(new_n18040), .D(new_n18045), .Y(\f[81] ));
  O2A1O1Ixp33_ASAP7_75t_L   g17790(.A1(new_n17823), .A2(new_n17822), .B(new_n18033), .C(new_n18029), .Y(new_n18047));
  A2O1A1Ixp33_ASAP7_75t_L   g17791(.A1(new_n18024), .A2(new_n18020), .B(new_n17831), .C(new_n17832), .Y(new_n18048));
  INVx1_ASAP7_75t_L         g17792(.A(new_n18048), .Y(new_n18049));
  NOR2xp33_ASAP7_75t_L      g17793(.A(new_n12956), .B(new_n1517), .Y(new_n18050));
  AOI21xp33_ASAP7_75t_L     g17794(.A1(new_n1659), .A2(\b[62] ), .B(new_n18050), .Y(new_n18051));
  INVx1_ASAP7_75t_L         g17795(.A(new_n18051), .Y(new_n18052));
  A2O1A1Ixp33_ASAP7_75t_L   g17796(.A1(new_n1508), .A2(new_n1509), .B(new_n1389), .C(new_n18051), .Y(new_n18053));
  O2A1O1Ixp33_ASAP7_75t_L   g17797(.A1(new_n18052), .A2(new_n17329), .B(new_n18053), .C(new_n1501), .Y(new_n18054));
  O2A1O1Ixp33_ASAP7_75t_L   g17798(.A1(new_n1521), .A2(new_n12993), .B(new_n18051), .C(\a[20] ), .Y(new_n18055));
  NOR2xp33_ASAP7_75t_L      g17799(.A(new_n18055), .B(new_n18054), .Y(new_n18056));
  INVx1_ASAP7_75t_L         g17800(.A(new_n18056), .Y(new_n18057));
  NOR2xp33_ASAP7_75t_L      g17801(.A(new_n11626), .B(new_n1962), .Y(new_n18058));
  AOI221xp5_ASAP7_75t_L     g17802(.A1(new_n1955), .A2(\b[61] ), .B1(new_n2093), .B2(\b[59] ), .C(new_n18058), .Y(new_n18059));
  O2A1O1Ixp33_ASAP7_75t_L   g17803(.A1(new_n1956), .A2(new_n14764), .B(new_n18059), .C(new_n1952), .Y(new_n18060));
  INVx1_ASAP7_75t_L         g17804(.A(new_n18060), .Y(new_n18061));
  O2A1O1Ixp33_ASAP7_75t_L   g17805(.A1(new_n1956), .A2(new_n14764), .B(new_n18059), .C(\a[23] ), .Y(new_n18062));
  AOI21xp33_ASAP7_75t_L     g17806(.A1(new_n18061), .A2(\a[23] ), .B(new_n18062), .Y(new_n18063));
  AOI21xp33_ASAP7_75t_L     g17807(.A1(new_n18019), .A2(new_n18008), .B(new_n18015), .Y(new_n18064));
  AND2x2_ASAP7_75t_L        g17808(.A(new_n18063), .B(new_n18064), .Y(new_n18065));
  O2A1O1Ixp33_ASAP7_75t_L   g17809(.A1(new_n18009), .A2(new_n18016), .B(new_n18014), .C(new_n18063), .Y(new_n18066));
  NOR2xp33_ASAP7_75t_L      g17810(.A(new_n18066), .B(new_n18065), .Y(new_n18067));
  NAND2xp33_ASAP7_75t_L     g17811(.A(\b[57] ), .B(new_n2421), .Y(new_n18068));
  OAI221xp5_ASAP7_75t_L     g17812(.A1(new_n2415), .A2(new_n11303), .B1(new_n10332), .B2(new_n2572), .C(new_n18068), .Y(new_n18069));
  A2O1A1Ixp33_ASAP7_75t_L   g17813(.A1(new_n11314), .A2(new_n2417), .B(new_n18069), .C(\a[26] ), .Y(new_n18070));
  NAND2xp33_ASAP7_75t_L     g17814(.A(\a[26] ), .B(new_n18070), .Y(new_n18071));
  A2O1A1Ixp33_ASAP7_75t_L   g17815(.A1(new_n11314), .A2(new_n2417), .B(new_n18069), .C(new_n2413), .Y(new_n18072));
  NAND2xp33_ASAP7_75t_L     g17816(.A(new_n18072), .B(new_n18071), .Y(new_n18073));
  NOR2xp33_ASAP7_75t_L      g17817(.A(new_n17839), .B(new_n17837), .Y(new_n18074));
  AO21x2_ASAP7_75t_L        g17818(.A1(new_n18005), .A2(new_n18074), .B(new_n17839), .Y(new_n18075));
  XNOR2x2_ASAP7_75t_L       g17819(.A(new_n18073), .B(new_n18075), .Y(new_n18076));
  NOR2xp33_ASAP7_75t_L      g17820(.A(new_n10309), .B(new_n2930), .Y(new_n18077));
  AOI221xp5_ASAP7_75t_L     g17821(.A1(\b[53] ), .A2(new_n3129), .B1(\b[54] ), .B2(new_n2936), .C(new_n18077), .Y(new_n18078));
  O2A1O1Ixp33_ASAP7_75t_L   g17822(.A1(new_n2940), .A2(new_n15849), .B(new_n18078), .C(new_n2928), .Y(new_n18079));
  INVx1_ASAP7_75t_L         g17823(.A(new_n18079), .Y(new_n18080));
  O2A1O1Ixp33_ASAP7_75t_L   g17824(.A1(new_n2940), .A2(new_n15849), .B(new_n18078), .C(\a[29] ), .Y(new_n18081));
  AOI21xp33_ASAP7_75t_L     g17825(.A1(new_n18080), .A2(\a[29] ), .B(new_n18081), .Y(new_n18082));
  INVx1_ASAP7_75t_L         g17826(.A(new_n18082), .Y(new_n18083));
  AOI211xp5_ASAP7_75t_L     g17827(.A1(new_n18004), .A2(new_n17995), .B(new_n18083), .C(new_n17999), .Y(new_n18084));
  A2O1A1Ixp33_ASAP7_75t_L   g17828(.A1(new_n18004), .A2(new_n17995), .B(new_n17999), .C(new_n18083), .Y(new_n18085));
  INVx1_ASAP7_75t_L         g17829(.A(new_n18085), .Y(new_n18086));
  NOR2xp33_ASAP7_75t_L      g17830(.A(new_n18084), .B(new_n18086), .Y(new_n18087));
  NOR2xp33_ASAP7_75t_L      g17831(.A(new_n9355), .B(new_n3510), .Y(new_n18088));
  AOI221xp5_ASAP7_75t_L     g17832(.A1(\b[50] ), .A2(new_n3708), .B1(\b[51] ), .B2(new_n3499), .C(new_n18088), .Y(new_n18089));
  O2A1O1Ixp33_ASAP7_75t_L   g17833(.A1(new_n3513), .A2(new_n17363), .B(new_n18089), .C(new_n3493), .Y(new_n18090));
  O2A1O1Ixp33_ASAP7_75t_L   g17834(.A1(new_n3513), .A2(new_n17363), .B(new_n18089), .C(\a[32] ), .Y(new_n18091));
  INVx1_ASAP7_75t_L         g17835(.A(new_n18091), .Y(new_n18092));
  OAI21xp33_ASAP7_75t_L     g17836(.A1(new_n3493), .A2(new_n18090), .B(new_n18092), .Y(new_n18093));
  NOR3xp33_ASAP7_75t_L      g17837(.A(new_n17994), .B(new_n18093), .C(new_n17986), .Y(new_n18094));
  A2O1A1Ixp33_ASAP7_75t_L   g17838(.A1(new_n17988), .A2(new_n17989), .B(new_n17986), .C(new_n18093), .Y(new_n18095));
  INVx1_ASAP7_75t_L         g17839(.A(new_n18095), .Y(new_n18096));
  NOR2xp33_ASAP7_75t_L      g17840(.A(new_n18094), .B(new_n18096), .Y(new_n18097));
  A2O1A1Ixp33_ASAP7_75t_L   g17841(.A1(new_n17734), .A2(new_n17656), .B(new_n17735), .C(new_n17842), .Y(new_n18098));
  A2O1A1Ixp33_ASAP7_75t_L   g17842(.A1(new_n17734), .A2(new_n18098), .B(new_n17951), .C(new_n17948), .Y(new_n18099));
  NAND2xp33_ASAP7_75t_L     g17843(.A(\b[40] ), .B(new_n6442), .Y(new_n18100));
  OAI221xp5_ASAP7_75t_L     g17844(.A1(new_n7304), .A2(new_n5570), .B1(new_n5311), .B2(new_n6741), .C(new_n18100), .Y(new_n18101));
  A2O1A1Ixp33_ASAP7_75t_L   g17845(.A1(new_n6651), .A2(new_n6450), .B(new_n18101), .C(\a[44] ), .Y(new_n18102));
  AOI211xp5_ASAP7_75t_L     g17846(.A1(new_n6651), .A2(new_n6450), .B(new_n18101), .C(new_n6439), .Y(new_n18103));
  A2O1A1O1Ixp25_ASAP7_75t_L g17847(.A1(new_n6450), .A2(new_n6651), .B(new_n18101), .C(new_n18102), .D(new_n18103), .Y(new_n18104));
  INVx1_ASAP7_75t_L         g17848(.A(new_n17866), .Y(new_n18105));
  NOR2xp33_ASAP7_75t_L      g17849(.A(new_n1458), .B(new_n13030), .Y(new_n18106));
  INVx1_ASAP7_75t_L         g17850(.A(new_n17850), .Y(new_n18107));
  A2O1A1O1Ixp25_ASAP7_75t_L g17851(.A1(new_n13028), .A2(\b[17] ), .B(new_n17667), .C(new_n17852), .D(new_n18107), .Y(new_n18108));
  A2O1A1Ixp33_ASAP7_75t_L   g17852(.A1(new_n13028), .A2(\b[19] ), .B(new_n18106), .C(new_n18108), .Y(new_n18109));
  O2A1O1Ixp33_ASAP7_75t_L   g17853(.A1(new_n12669), .A2(new_n12671), .B(\b[19] ), .C(new_n18106), .Y(new_n18110));
  INVx1_ASAP7_75t_L         g17854(.A(new_n18110), .Y(new_n18111));
  O2A1O1Ixp33_ASAP7_75t_L   g17855(.A1(new_n17668), .A2(new_n17853), .B(new_n17850), .C(new_n18111), .Y(new_n18112));
  INVx1_ASAP7_75t_L         g17856(.A(new_n18112), .Y(new_n18113));
  NAND2xp33_ASAP7_75t_L     g17857(.A(new_n18109), .B(new_n18113), .Y(new_n18114));
  NOR2xp33_ASAP7_75t_L      g17858(.A(new_n1895), .B(new_n12318), .Y(new_n18115));
  AOI221xp5_ASAP7_75t_L     g17859(.A1(new_n11995), .A2(\b[22] ), .B1(new_n13314), .B2(\b[20] ), .C(new_n18115), .Y(new_n18116));
  O2A1O1Ixp33_ASAP7_75t_L   g17860(.A1(new_n11998), .A2(new_n2522), .B(new_n18116), .C(new_n11987), .Y(new_n18117));
  O2A1O1Ixp33_ASAP7_75t_L   g17861(.A1(new_n11998), .A2(new_n2522), .B(new_n18116), .C(\a[62] ), .Y(new_n18118));
  INVx1_ASAP7_75t_L         g17862(.A(new_n18118), .Y(new_n18119));
  OAI211xp5_ASAP7_75t_L     g17863(.A1(new_n11987), .A2(new_n18117), .B(new_n18119), .C(new_n18114), .Y(new_n18120));
  O2A1O1Ixp33_ASAP7_75t_L   g17864(.A1(new_n11987), .A2(new_n18117), .B(new_n18119), .C(new_n18114), .Y(new_n18121));
  INVx1_ASAP7_75t_L         g17865(.A(new_n18121), .Y(new_n18122));
  AND2x2_ASAP7_75t_L        g17866(.A(new_n18120), .B(new_n18122), .Y(new_n18123));
  INVx1_ASAP7_75t_L         g17867(.A(new_n18123), .Y(new_n18124));
  A2O1A1O1Ixp25_ASAP7_75t_L g17868(.A1(new_n17868), .A2(new_n17858), .B(new_n17684), .C(new_n18105), .D(new_n18124), .Y(new_n18125));
  INVx1_ASAP7_75t_L         g17869(.A(new_n18125), .Y(new_n18126));
  O2A1O1Ixp33_ASAP7_75t_L   g17870(.A1(new_n17857), .A2(new_n17867), .B(new_n17683), .C(new_n17866), .Y(new_n18127));
  NAND2xp33_ASAP7_75t_L     g17871(.A(new_n18127), .B(new_n18124), .Y(new_n18128));
  NAND2xp33_ASAP7_75t_L     g17872(.A(new_n18128), .B(new_n18126), .Y(new_n18129));
  NOR2xp33_ASAP7_75t_L      g17873(.A(new_n2188), .B(new_n11354), .Y(new_n18130));
  AOI221xp5_ASAP7_75t_L     g17874(.A1(\b[25] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[24] ), .C(new_n18130), .Y(new_n18131));
  O2A1O1Ixp33_ASAP7_75t_L   g17875(.A1(new_n11053), .A2(new_n2385), .B(new_n18131), .C(new_n11048), .Y(new_n18132));
  O2A1O1Ixp33_ASAP7_75t_L   g17876(.A1(new_n11053), .A2(new_n2385), .B(new_n18131), .C(\a[59] ), .Y(new_n18133));
  INVx1_ASAP7_75t_L         g17877(.A(new_n18133), .Y(new_n18134));
  O2A1O1Ixp33_ASAP7_75t_L   g17878(.A1(new_n18132), .A2(new_n11048), .B(new_n18134), .C(new_n18129), .Y(new_n18135));
  INVx1_ASAP7_75t_L         g17879(.A(new_n18132), .Y(new_n18136));
  A2O1A1Ixp33_ASAP7_75t_L   g17880(.A1(\a[59] ), .A2(new_n18136), .B(new_n18133), .C(new_n18129), .Y(new_n18137));
  OAI21xp33_ASAP7_75t_L     g17881(.A1(new_n18129), .A2(new_n18135), .B(new_n18137), .Y(new_n18138));
  O2A1O1Ixp33_ASAP7_75t_L   g17882(.A1(new_n17883), .A2(new_n17884), .B(new_n17880), .C(new_n18138), .Y(new_n18139));
  NAND2xp33_ASAP7_75t_L     g17883(.A(new_n17880), .B(new_n17882), .Y(new_n18140));
  O2A1O1Ixp33_ASAP7_75t_L   g17884(.A1(new_n18129), .A2(new_n18135), .B(new_n18137), .C(new_n18140), .Y(new_n18141));
  NOR2xp33_ASAP7_75t_L      g17885(.A(new_n18141), .B(new_n18139), .Y(new_n18142));
  NOR2xp33_ASAP7_75t_L      g17886(.A(new_n2879), .B(new_n10388), .Y(new_n18143));
  AOI221xp5_ASAP7_75t_L     g17887(.A1(new_n10086), .A2(\b[28] ), .B1(new_n11361), .B2(\b[26] ), .C(new_n18143), .Y(new_n18144));
  O2A1O1Ixp33_ASAP7_75t_L   g17888(.A1(new_n10088), .A2(new_n3087), .B(new_n18144), .C(new_n10083), .Y(new_n18145));
  NOR2xp33_ASAP7_75t_L      g17889(.A(new_n10083), .B(new_n18145), .Y(new_n18146));
  O2A1O1Ixp33_ASAP7_75t_L   g17890(.A1(new_n10088), .A2(new_n3087), .B(new_n18144), .C(\a[56] ), .Y(new_n18147));
  NOR2xp33_ASAP7_75t_L      g17891(.A(new_n18147), .B(new_n18146), .Y(new_n18148));
  XNOR2x2_ASAP7_75t_L       g17892(.A(new_n18148), .B(new_n18142), .Y(new_n18149));
  A2O1A1O1Ixp25_ASAP7_75t_L g17893(.A1(new_n17895), .A2(new_n17886), .B(new_n17897), .C(new_n17899), .D(new_n18149), .Y(new_n18150));
  INVx1_ASAP7_75t_L         g17894(.A(new_n18150), .Y(new_n18151));
  NAND3xp33_ASAP7_75t_L     g17895(.A(new_n17901), .B(new_n17899), .C(new_n18149), .Y(new_n18152));
  NAND2xp33_ASAP7_75t_L     g17896(.A(new_n18152), .B(new_n18151), .Y(new_n18153));
  NOR2xp33_ASAP7_75t_L      g17897(.A(new_n3456), .B(new_n10400), .Y(new_n18154));
  AOI221xp5_ASAP7_75t_L     g17898(.A1(new_n9102), .A2(\b[31] ), .B1(new_n10398), .B2(\b[29] ), .C(new_n18154), .Y(new_n18155));
  O2A1O1Ixp33_ASAP7_75t_L   g17899(.A1(new_n9104), .A2(new_n3681), .B(new_n18155), .C(new_n9099), .Y(new_n18156));
  O2A1O1Ixp33_ASAP7_75t_L   g17900(.A1(new_n9104), .A2(new_n3681), .B(new_n18155), .C(\a[53] ), .Y(new_n18157));
  INVx1_ASAP7_75t_L         g17901(.A(new_n18157), .Y(new_n18158));
  O2A1O1Ixp33_ASAP7_75t_L   g17902(.A1(new_n18156), .A2(new_n9099), .B(new_n18158), .C(new_n18153), .Y(new_n18159));
  INVx1_ASAP7_75t_L         g17903(.A(new_n18156), .Y(new_n18160));
  A2O1A1Ixp33_ASAP7_75t_L   g17904(.A1(\a[53] ), .A2(new_n18160), .B(new_n18157), .C(new_n18153), .Y(new_n18161));
  OA21x2_ASAP7_75t_L        g17905(.A1(new_n18153), .A2(new_n18159), .B(new_n18161), .Y(new_n18162));
  INVx1_ASAP7_75t_L         g17906(.A(new_n18162), .Y(new_n18163));
  A2O1A1Ixp33_ASAP7_75t_L   g17907(.A1(new_n17911), .A2(new_n17902), .B(new_n17914), .C(new_n17916), .Y(new_n18164));
  NOR2xp33_ASAP7_75t_L      g17908(.A(new_n18164), .B(new_n18163), .Y(new_n18165));
  A2O1A1O1Ixp25_ASAP7_75t_L g17909(.A1(new_n17911), .A2(new_n17902), .B(new_n17914), .C(new_n17916), .D(new_n18162), .Y(new_n18166));
  NOR2xp33_ASAP7_75t_L      g17910(.A(new_n18166), .B(new_n18165), .Y(new_n18167));
  NOR2xp33_ASAP7_75t_L      g17911(.A(new_n4101), .B(new_n10065), .Y(new_n18168));
  AOI221xp5_ASAP7_75t_L     g17912(.A1(new_n8175), .A2(\b[34] ), .B1(new_n8484), .B2(\b[32] ), .C(new_n18168), .Y(new_n18169));
  O2A1O1Ixp33_ASAP7_75t_L   g17913(.A1(new_n8176), .A2(new_n4352), .B(new_n18169), .C(new_n8172), .Y(new_n18170));
  INVx1_ASAP7_75t_L         g17914(.A(new_n18170), .Y(new_n18171));
  O2A1O1Ixp33_ASAP7_75t_L   g17915(.A1(new_n8176), .A2(new_n4352), .B(new_n18169), .C(\a[50] ), .Y(new_n18172));
  A2O1A1Ixp33_ASAP7_75t_L   g17916(.A1(\a[50] ), .A2(new_n18171), .B(new_n18172), .C(new_n18167), .Y(new_n18173));
  INVx1_ASAP7_75t_L         g17917(.A(new_n18172), .Y(new_n18174));
  O2A1O1Ixp33_ASAP7_75t_L   g17918(.A1(new_n18170), .A2(new_n8172), .B(new_n18174), .C(new_n18167), .Y(new_n18175));
  AOI21xp33_ASAP7_75t_L     g17919(.A1(new_n18173), .A2(new_n18167), .B(new_n18175), .Y(new_n18176));
  OR2x4_ASAP7_75t_L         g17920(.A(new_n17919), .B(new_n17929), .Y(new_n18177));
  OA21x2_ASAP7_75t_L        g17921(.A1(new_n17925), .A2(new_n17928), .B(new_n18177), .Y(new_n18178));
  XNOR2x2_ASAP7_75t_L       g17922(.A(new_n18178), .B(new_n18176), .Y(new_n18179));
  NOR2xp33_ASAP7_75t_L      g17923(.A(new_n5074), .B(new_n7318), .Y(new_n18180));
  AOI221xp5_ASAP7_75t_L     g17924(.A1(new_n7333), .A2(\b[36] ), .B1(new_n7609), .B2(\b[35] ), .C(new_n18180), .Y(new_n18181));
  O2A1O1Ixp33_ASAP7_75t_L   g17925(.A1(new_n7321), .A2(new_n5083), .B(new_n18181), .C(new_n7316), .Y(new_n18182));
  O2A1O1Ixp33_ASAP7_75t_L   g17926(.A1(new_n7321), .A2(new_n5083), .B(new_n18181), .C(\a[47] ), .Y(new_n18183));
  INVx1_ASAP7_75t_L         g17927(.A(new_n18183), .Y(new_n18184));
  OAI21xp33_ASAP7_75t_L     g17928(.A1(new_n7316), .A2(new_n18182), .B(new_n18184), .Y(new_n18185));
  XNOR2x2_ASAP7_75t_L       g17929(.A(new_n18185), .B(new_n18179), .Y(new_n18186));
  INVx1_ASAP7_75t_L         g17930(.A(new_n18186), .Y(new_n18187));
  A2O1A1Ixp33_ASAP7_75t_L   g17931(.A1(new_n17939), .A2(new_n17844), .B(new_n17937), .C(new_n18187), .Y(new_n18188));
  A2O1A1Ixp33_ASAP7_75t_L   g17932(.A1(new_n17939), .A2(new_n17844), .B(new_n17937), .C(new_n18186), .Y(new_n18189));
  NAND2xp33_ASAP7_75t_L     g17933(.A(new_n18186), .B(new_n18189), .Y(new_n18190));
  AO21x2_ASAP7_75t_L        g17934(.A1(new_n18188), .A2(new_n18190), .B(new_n18104), .Y(new_n18191));
  NAND3xp33_ASAP7_75t_L     g17935(.A(new_n18190), .B(new_n18188), .C(new_n18104), .Y(new_n18192));
  NAND3xp33_ASAP7_75t_L     g17936(.A(new_n18191), .B(new_n18099), .C(new_n18192), .Y(new_n18193));
  AO21x2_ASAP7_75t_L        g17937(.A1(new_n18192), .A2(new_n18191), .B(new_n18099), .Y(new_n18194));
  NAND2xp33_ASAP7_75t_L     g17938(.A(new_n18193), .B(new_n18194), .Y(new_n18195));
  NOR2xp33_ASAP7_75t_L      g17939(.A(new_n6378), .B(new_n5640), .Y(new_n18196));
  AOI221xp5_ASAP7_75t_L     g17940(.A1(\b[41] ), .A2(new_n5920), .B1(\b[43] ), .B2(new_n5629), .C(new_n18196), .Y(new_n18197));
  O2A1O1Ixp33_ASAP7_75t_L   g17941(.A1(new_n5630), .A2(new_n6679), .B(new_n18197), .C(new_n5626), .Y(new_n18198));
  O2A1O1Ixp33_ASAP7_75t_L   g17942(.A1(new_n5630), .A2(new_n6679), .B(new_n18197), .C(\a[41] ), .Y(new_n18199));
  INVx1_ASAP7_75t_L         g17943(.A(new_n18199), .Y(new_n18200));
  O2A1O1Ixp33_ASAP7_75t_L   g17944(.A1(new_n18198), .A2(new_n5626), .B(new_n18200), .C(new_n18195), .Y(new_n18201));
  INVx1_ASAP7_75t_L         g17945(.A(new_n18198), .Y(new_n18202));
  A2O1A1Ixp33_ASAP7_75t_L   g17946(.A1(\a[41] ), .A2(new_n18202), .B(new_n18199), .C(new_n18195), .Y(new_n18203));
  A2O1A1O1Ixp25_ASAP7_75t_L g17947(.A1(new_n17487), .A2(new_n17481), .B(new_n17400), .C(new_n17485), .D(new_n17745), .Y(new_n18204));
  INVx1_ASAP7_75t_L         g17948(.A(new_n17747), .Y(new_n18205));
  O2A1O1Ixp33_ASAP7_75t_L   g17949(.A1(new_n17960), .A2(new_n5626), .B(new_n17962), .C(new_n17957), .Y(new_n18206));
  O2A1O1Ixp33_ASAP7_75t_L   g17950(.A1(new_n18204), .A2(new_n18205), .B(new_n17964), .C(new_n18206), .Y(new_n18207));
  OA211x2_ASAP7_75t_L       g17951(.A1(new_n18195), .A2(new_n18201), .B(new_n18203), .C(new_n18207), .Y(new_n18208));
  O2A1O1Ixp33_ASAP7_75t_L   g17952(.A1(new_n18195), .A2(new_n18201), .B(new_n18203), .C(new_n18207), .Y(new_n18209));
  NOR2xp33_ASAP7_75t_L      g17953(.A(new_n18209), .B(new_n18208), .Y(new_n18210));
  INVx1_ASAP7_75t_L         g17954(.A(new_n18210), .Y(new_n18211));
  NOR2xp33_ASAP7_75t_L      g17955(.A(new_n7249), .B(new_n4903), .Y(new_n18212));
  AOI221xp5_ASAP7_75t_L     g17956(.A1(\b[44] ), .A2(new_n5139), .B1(\b[46] ), .B2(new_n4917), .C(new_n18212), .Y(new_n18213));
  O2A1O1Ixp33_ASAP7_75t_L   g17957(.A1(new_n4911), .A2(new_n7279), .B(new_n18213), .C(new_n4906), .Y(new_n18214));
  O2A1O1Ixp33_ASAP7_75t_L   g17958(.A1(new_n4911), .A2(new_n7279), .B(new_n18213), .C(\a[38] ), .Y(new_n18215));
  INVx1_ASAP7_75t_L         g17959(.A(new_n18215), .Y(new_n18216));
  O2A1O1Ixp33_ASAP7_75t_L   g17960(.A1(new_n18214), .A2(new_n4906), .B(new_n18216), .C(new_n18211), .Y(new_n18217));
  O2A1O1Ixp33_ASAP7_75t_L   g17961(.A1(new_n18214), .A2(new_n4906), .B(new_n18216), .C(new_n18210), .Y(new_n18218));
  INVx1_ASAP7_75t_L         g17962(.A(new_n18218), .Y(new_n18219));
  INVx1_ASAP7_75t_L         g17963(.A(new_n17644), .Y(new_n18220));
  O2A1O1Ixp33_ASAP7_75t_L   g17964(.A1(new_n4906), .A2(new_n17642), .B(new_n18220), .C(new_n17753), .Y(new_n18221));
  O2A1O1Ixp33_ASAP7_75t_L   g17965(.A1(new_n18221), .A2(new_n17750), .B(new_n17974), .C(new_n17971), .Y(new_n18222));
  OAI211xp5_ASAP7_75t_L     g17966(.A1(new_n18211), .A2(new_n18217), .B(new_n18219), .C(new_n18222), .Y(new_n18223));
  O2A1O1Ixp33_ASAP7_75t_L   g17967(.A1(new_n18211), .A2(new_n18217), .B(new_n18219), .C(new_n18222), .Y(new_n18224));
  INVx1_ASAP7_75t_L         g17968(.A(new_n18224), .Y(new_n18225));
  AND2x2_ASAP7_75t_L        g17969(.A(new_n18223), .B(new_n18225), .Y(new_n18226));
  NOR2xp33_ASAP7_75t_L      g17970(.A(new_n7860), .B(new_n4142), .Y(new_n18227));
  AOI221xp5_ASAP7_75t_L     g17971(.A1(\b[47] ), .A2(new_n4402), .B1(\b[49] ), .B2(new_n4156), .C(new_n18227), .Y(new_n18228));
  INVx1_ASAP7_75t_L         g17972(.A(new_n18228), .Y(new_n18229));
  A2O1A1Ixp33_ASAP7_75t_L   g17973(.A1(new_n8438), .A2(new_n4151), .B(new_n18229), .C(\a[35] ), .Y(new_n18230));
  O2A1O1Ixp33_ASAP7_75t_L   g17974(.A1(new_n4150), .A2(new_n14802), .B(new_n18228), .C(\a[35] ), .Y(new_n18231));
  A2O1A1Ixp33_ASAP7_75t_L   g17975(.A1(\a[35] ), .A2(new_n18230), .B(new_n18231), .C(new_n18226), .Y(new_n18232));
  O2A1O1Ixp33_ASAP7_75t_L   g17976(.A1(new_n4150), .A2(new_n14802), .B(new_n18228), .C(new_n4145), .Y(new_n18233));
  INVx1_ASAP7_75t_L         g17977(.A(new_n18231), .Y(new_n18234));
  O2A1O1Ixp33_ASAP7_75t_L   g17978(.A1(new_n18233), .A2(new_n4145), .B(new_n18234), .C(new_n18226), .Y(new_n18235));
  A2O1A1Ixp33_ASAP7_75t_L   g17979(.A1(new_n18226), .A2(new_n18232), .B(new_n18235), .C(new_n18097), .Y(new_n18236));
  INVx1_ASAP7_75t_L         g17980(.A(new_n18236), .Y(new_n18237));
  NAND2xp33_ASAP7_75t_L     g17981(.A(new_n18226), .B(new_n18232), .Y(new_n18238));
  A2O1A1Ixp33_ASAP7_75t_L   g17982(.A1(new_n18230), .A2(\a[35] ), .B(new_n18231), .C(new_n18232), .Y(new_n18239));
  NAND2xp33_ASAP7_75t_L     g17983(.A(new_n18238), .B(new_n18239), .Y(new_n18240));
  NOR2xp33_ASAP7_75t_L      g17984(.A(new_n18240), .B(new_n18097), .Y(new_n18241));
  INVx1_ASAP7_75t_L         g17985(.A(new_n18241), .Y(new_n18242));
  NAND2xp33_ASAP7_75t_L     g17986(.A(new_n18242), .B(new_n18087), .Y(new_n18243));
  NOR3xp33_ASAP7_75t_L      g17987(.A(new_n18087), .B(new_n18237), .C(new_n18241), .Y(new_n18244));
  O2A1O1Ixp33_ASAP7_75t_L   g17988(.A1(new_n18237), .A2(new_n18243), .B(new_n18087), .C(new_n18244), .Y(new_n18245));
  NOR2xp33_ASAP7_75t_L      g17989(.A(new_n18245), .B(new_n18076), .Y(new_n18246));
  NAND2xp33_ASAP7_75t_L     g17990(.A(new_n18245), .B(new_n18076), .Y(new_n18247));
  NAND2xp33_ASAP7_75t_L     g17991(.A(new_n18247), .B(new_n18067), .Y(new_n18248));
  INVx1_ASAP7_75t_L         g17992(.A(new_n18247), .Y(new_n18249));
  NOR3xp33_ASAP7_75t_L      g17993(.A(new_n18067), .B(new_n18246), .C(new_n18249), .Y(new_n18250));
  O2A1O1Ixp33_ASAP7_75t_L   g17994(.A1(new_n18246), .A2(new_n18248), .B(new_n18067), .C(new_n18250), .Y(new_n18251));
  A2O1A1O1Ixp25_ASAP7_75t_L g17995(.A1(new_n18020), .A2(new_n18024), .B(new_n17831), .C(new_n17832), .D(new_n18056), .Y(new_n18252));
  A2O1A1Ixp33_ASAP7_75t_L   g17996(.A1(new_n18021), .A2(new_n18023), .B(new_n17833), .C(new_n18056), .Y(new_n18253));
  O2A1O1Ixp33_ASAP7_75t_L   g17997(.A1(new_n18056), .A2(new_n18252), .B(new_n18253), .C(new_n18251), .Y(new_n18254));
  NOR2xp33_ASAP7_75t_L      g17998(.A(new_n18073), .B(new_n18075), .Y(new_n18255));
  A2O1A1Ixp33_ASAP7_75t_L   g17999(.A1(new_n18074), .A2(new_n18005), .B(new_n17839), .C(new_n18073), .Y(new_n18256));
  INVx1_ASAP7_75t_L         g18000(.A(new_n18256), .Y(new_n18257));
  NOR2xp33_ASAP7_75t_L      g18001(.A(new_n18257), .B(new_n18255), .Y(new_n18258));
  NAND3xp33_ASAP7_75t_L     g18002(.A(new_n18087), .B(new_n18236), .C(new_n18242), .Y(new_n18259));
  A2O1A1Ixp33_ASAP7_75t_L   g18003(.A1(new_n18087), .A2(new_n18259), .B(new_n18244), .C(new_n18258), .Y(new_n18260));
  NAND3xp33_ASAP7_75t_L     g18004(.A(new_n18067), .B(new_n18260), .C(new_n18247), .Y(new_n18261));
  AO21x2_ASAP7_75t_L        g18005(.A1(new_n18067), .A2(new_n18261), .B(new_n18250), .Y(new_n18262));
  INVx1_ASAP7_75t_L         g18006(.A(new_n18252), .Y(new_n18263));
  O2A1O1Ixp33_ASAP7_75t_L   g18007(.A1(new_n18054), .A2(new_n18055), .B(new_n18263), .C(new_n18262), .Y(new_n18264));
  O2A1O1Ixp33_ASAP7_75t_L   g18008(.A1(new_n18057), .A2(new_n18049), .B(new_n18264), .C(new_n18254), .Y(new_n18265));
  A2O1A1Ixp33_ASAP7_75t_L   g18009(.A1(new_n17808), .A2(new_n17801), .B(new_n17810), .C(new_n18040), .Y(new_n18266));
  A2O1A1O1Ixp25_ASAP7_75t_L g18010(.A1(new_n18020), .A2(new_n18024), .B(new_n17831), .C(new_n17832), .D(new_n18057), .Y(new_n18267));
  O2A1O1Ixp33_ASAP7_75t_L   g18011(.A1(new_n18054), .A2(new_n18055), .B(new_n18263), .C(new_n18267), .Y(new_n18268));
  OAI211xp5_ASAP7_75t_L     g18012(.A1(new_n18056), .A2(new_n18252), .B(new_n18251), .C(new_n18253), .Y(new_n18269));
  O2A1O1Ixp33_ASAP7_75t_L   g18013(.A1(new_n18251), .A2(new_n18268), .B(new_n18269), .C(new_n18047), .Y(new_n18270));
  A2O1A1Ixp33_ASAP7_75t_L   g18014(.A1(new_n18057), .A2(new_n18263), .B(new_n18267), .C(new_n18262), .Y(new_n18271));
  AND3x1_ASAP7_75t_L        g18015(.A(new_n18271), .B(new_n18269), .C(new_n18047), .Y(new_n18272));
  NOR2xp33_ASAP7_75t_L      g18016(.A(new_n18270), .B(new_n18272), .Y(new_n18273));
  A2O1A1O1Ixp25_ASAP7_75t_L g18017(.A1(new_n18028), .A2(new_n18034), .B(new_n18036), .C(new_n18266), .D(new_n18273), .Y(new_n18274));
  A2O1A1Ixp33_ASAP7_75t_L   g18018(.A1(new_n18028), .A2(new_n18034), .B(new_n18036), .C(new_n18266), .Y(new_n18275));
  NOR2xp33_ASAP7_75t_L      g18019(.A(new_n18272), .B(new_n18275), .Y(new_n18276));
  O2A1O1Ixp33_ASAP7_75t_L   g18020(.A1(new_n18265), .A2(new_n18047), .B(new_n18276), .C(new_n18274), .Y(\f[82] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18021(.A1(new_n17821), .A2(new_n18029), .B(new_n18030), .C(new_n18027), .Y(new_n18278));
  A2O1A1Ixp33_ASAP7_75t_L   g18022(.A1(new_n17822), .A2(new_n17824), .B(new_n18278), .C(new_n18265), .Y(new_n18279));
  NOR2xp33_ASAP7_75t_L      g18023(.A(new_n12956), .B(new_n1654), .Y(new_n18280));
  A2O1A1Ixp33_ASAP7_75t_L   g18024(.A1(new_n12986), .A2(new_n1513), .B(new_n18280), .C(\a[20] ), .Y(new_n18281));
  A2O1A1O1Ixp25_ASAP7_75t_L g18025(.A1(new_n1513), .A2(new_n14172), .B(new_n1659), .C(\b[63] ), .D(new_n1501), .Y(new_n18282));
  A2O1A1O1Ixp25_ASAP7_75t_L g18026(.A1(new_n12986), .A2(new_n1513), .B(new_n18280), .C(new_n18281), .D(new_n18282), .Y(new_n18283));
  INVx1_ASAP7_75t_L         g18027(.A(new_n18283), .Y(new_n18284));
  NAND2xp33_ASAP7_75t_L     g18028(.A(new_n18063), .B(new_n18064), .Y(new_n18285));
  INVx1_ASAP7_75t_L         g18029(.A(new_n18066), .Y(new_n18286));
  NAND2xp33_ASAP7_75t_L     g18030(.A(new_n18285), .B(new_n18286), .Y(new_n18287));
  O2A1O1Ixp33_ASAP7_75t_L   g18031(.A1(new_n18255), .A2(new_n18257), .B(new_n18245), .C(new_n18287), .Y(new_n18288));
  A2O1A1Ixp33_ASAP7_75t_L   g18032(.A1(new_n18288), .A2(new_n18260), .B(new_n18066), .C(new_n18284), .Y(new_n18289));
  O2A1O1Ixp33_ASAP7_75t_L   g18033(.A1(new_n18063), .A2(new_n18064), .B(new_n18261), .C(new_n18284), .Y(new_n18290));
  NOR2xp33_ASAP7_75t_L      g18034(.A(new_n12258), .B(new_n1962), .Y(new_n18291));
  AOI221xp5_ASAP7_75t_L     g18035(.A1(new_n1955), .A2(\b[62] ), .B1(new_n2093), .B2(\b[60] ), .C(new_n18291), .Y(new_n18292));
  O2A1O1Ixp33_ASAP7_75t_L   g18036(.A1(new_n1956), .A2(new_n12610), .B(new_n18292), .C(new_n1952), .Y(new_n18293));
  INVx1_ASAP7_75t_L         g18037(.A(new_n18293), .Y(new_n18294));
  O2A1O1Ixp33_ASAP7_75t_L   g18038(.A1(new_n1956), .A2(new_n12610), .B(new_n18292), .C(\a[23] ), .Y(new_n18295));
  AOI21xp33_ASAP7_75t_L     g18039(.A1(new_n18294), .A2(\a[23] ), .B(new_n18295), .Y(new_n18296));
  INVx1_ASAP7_75t_L         g18040(.A(new_n18296), .Y(new_n18297));
  O2A1O1Ixp33_ASAP7_75t_L   g18041(.A1(new_n18255), .A2(new_n18245), .B(new_n18256), .C(new_n18296), .Y(new_n18298));
  INVx1_ASAP7_75t_L         g18042(.A(new_n18298), .Y(new_n18299));
  O2A1O1Ixp33_ASAP7_75t_L   g18043(.A1(new_n18255), .A2(new_n18245), .B(new_n18256), .C(new_n18297), .Y(new_n18300));
  NOR2xp33_ASAP7_75t_L      g18044(.A(new_n10332), .B(new_n2930), .Y(new_n18301));
  AOI221xp5_ASAP7_75t_L     g18045(.A1(\b[54] ), .A2(new_n3129), .B1(\b[55] ), .B2(new_n2936), .C(new_n18301), .Y(new_n18302));
  O2A1O1Ixp33_ASAP7_75t_L   g18046(.A1(new_n2940), .A2(new_n10339), .B(new_n18302), .C(new_n2928), .Y(new_n18303));
  INVx1_ASAP7_75t_L         g18047(.A(new_n18303), .Y(new_n18304));
  O2A1O1Ixp33_ASAP7_75t_L   g18048(.A1(new_n2940), .A2(new_n10339), .B(new_n18302), .C(\a[29] ), .Y(new_n18305));
  A2O1A1Ixp33_ASAP7_75t_L   g18049(.A1(new_n18239), .A2(new_n18238), .B(new_n18094), .C(new_n18095), .Y(new_n18306));
  A2O1A1Ixp33_ASAP7_75t_L   g18050(.A1(new_n18304), .A2(\a[29] ), .B(new_n18305), .C(new_n18306), .Y(new_n18307));
  INVx1_ASAP7_75t_L         g18051(.A(new_n18307), .Y(new_n18308));
  A2O1A1Ixp33_ASAP7_75t_L   g18052(.A1(new_n18304), .A2(\a[29] ), .B(new_n18305), .C(new_n18307), .Y(new_n18309));
  A2O1A1Ixp33_ASAP7_75t_L   g18053(.A1(new_n18236), .A2(new_n18095), .B(new_n18308), .C(new_n18309), .Y(new_n18310));
  INVx1_ASAP7_75t_L         g18054(.A(new_n18193), .Y(new_n18311));
  A2O1A1O1Ixp25_ASAP7_75t_L g18055(.A1(new_n18202), .A2(\a[41] ), .B(new_n18199), .C(new_n18194), .D(new_n18311), .Y(new_n18312));
  NOR2xp33_ASAP7_75t_L      g18056(.A(new_n6944), .B(new_n5641), .Y(new_n18313));
  AOI221xp5_ASAP7_75t_L     g18057(.A1(\b[42] ), .A2(new_n5920), .B1(\b[43] ), .B2(new_n5623), .C(new_n18313), .Y(new_n18314));
  O2A1O1Ixp33_ASAP7_75t_L   g18058(.A1(new_n5630), .A2(new_n6951), .B(new_n18314), .C(new_n5626), .Y(new_n18315));
  O2A1O1Ixp33_ASAP7_75t_L   g18059(.A1(new_n5630), .A2(new_n6951), .B(new_n18314), .C(\a[41] ), .Y(new_n18316));
  INVx1_ASAP7_75t_L         g18060(.A(new_n18316), .Y(new_n18317));
  OA21x2_ASAP7_75t_L        g18061(.A1(new_n5626), .A2(new_n18315), .B(new_n18317), .Y(new_n18318));
  INVx1_ASAP7_75t_L         g18062(.A(new_n18189), .Y(new_n18319));
  O2A1O1Ixp33_ASAP7_75t_L   g18063(.A1(new_n18187), .A2(new_n18319), .B(new_n18188), .C(new_n18104), .Y(new_n18320));
  O2A1O1Ixp33_ASAP7_75t_L   g18064(.A1(new_n17937), .A2(new_n17941), .B(new_n18186), .C(new_n18320), .Y(new_n18321));
  NOR2xp33_ASAP7_75t_L      g18065(.A(new_n5570), .B(new_n6741), .Y(new_n18322));
  AOI221xp5_ASAP7_75t_L     g18066(.A1(\b[41] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[40] ), .C(new_n18322), .Y(new_n18323));
  O2A1O1Ixp33_ASAP7_75t_L   g18067(.A1(new_n6443), .A2(new_n6117), .B(new_n18323), .C(new_n6439), .Y(new_n18324));
  INVx1_ASAP7_75t_L         g18068(.A(new_n18324), .Y(new_n18325));
  O2A1O1Ixp33_ASAP7_75t_L   g18069(.A1(new_n6443), .A2(new_n6117), .B(new_n18323), .C(\a[44] ), .Y(new_n18326));
  AOI21xp33_ASAP7_75t_L     g18070(.A1(new_n18325), .A2(\a[44] ), .B(new_n18326), .Y(new_n18327));
  INVx1_ASAP7_75t_L         g18071(.A(new_n18178), .Y(new_n18328));
  O2A1O1Ixp33_ASAP7_75t_L   g18072(.A1(new_n18182), .A2(new_n7316), .B(new_n18184), .C(new_n18179), .Y(new_n18329));
  A2O1A1O1Ixp25_ASAP7_75t_L g18073(.A1(new_n18173), .A2(new_n18167), .B(new_n18175), .C(new_n18328), .D(new_n18329), .Y(new_n18330));
  NOR2xp33_ASAP7_75t_L      g18074(.A(new_n5311), .B(new_n7318), .Y(new_n18331));
  AOI221xp5_ASAP7_75t_L     g18075(.A1(new_n7333), .A2(\b[37] ), .B1(new_n7609), .B2(\b[36] ), .C(new_n18331), .Y(new_n18332));
  O2A1O1Ixp33_ASAP7_75t_L   g18076(.A1(new_n7321), .A2(new_n5318), .B(new_n18332), .C(new_n7316), .Y(new_n18333));
  O2A1O1Ixp33_ASAP7_75t_L   g18077(.A1(new_n7321), .A2(new_n5318), .B(new_n18332), .C(\a[47] ), .Y(new_n18334));
  INVx1_ASAP7_75t_L         g18078(.A(new_n18334), .Y(new_n18335));
  A2O1A1O1Ixp25_ASAP7_75t_L g18079(.A1(new_n18171), .A2(\a[50] ), .B(new_n18172), .C(new_n18167), .D(new_n18166), .Y(new_n18336));
  INVx1_ASAP7_75t_L         g18080(.A(new_n18336), .Y(new_n18337));
  NOR2xp33_ASAP7_75t_L      g18081(.A(new_n4344), .B(new_n10065), .Y(new_n18338));
  AOI221xp5_ASAP7_75t_L     g18082(.A1(new_n8175), .A2(\b[35] ), .B1(new_n8484), .B2(\b[33] ), .C(new_n18338), .Y(new_n18339));
  O2A1O1Ixp33_ASAP7_75t_L   g18083(.A1(new_n8176), .A2(new_n4589), .B(new_n18339), .C(new_n8172), .Y(new_n18340));
  INVx1_ASAP7_75t_L         g18084(.A(new_n18340), .Y(new_n18341));
  O2A1O1Ixp33_ASAP7_75t_L   g18085(.A1(new_n8176), .A2(new_n4589), .B(new_n18339), .C(\a[50] ), .Y(new_n18342));
  INVx1_ASAP7_75t_L         g18086(.A(new_n18149), .Y(new_n18343));
  A2O1A1Ixp33_ASAP7_75t_L   g18087(.A1(new_n17895), .A2(new_n17886), .B(new_n17897), .C(new_n17899), .Y(new_n18344));
  A2O1A1O1Ixp25_ASAP7_75t_L g18088(.A1(new_n17668), .A2(new_n17407), .B(new_n17678), .C(new_n17879), .D(new_n17871), .Y(new_n18345));
  INVx1_ASAP7_75t_L         g18089(.A(new_n18345), .Y(new_n18346));
  A2O1A1Ixp33_ASAP7_75t_L   g18090(.A1(new_n17410), .A2(new_n17416), .B(new_n17408), .C(new_n17846), .Y(new_n18347));
  O2A1O1Ixp33_ASAP7_75t_L   g18091(.A1(new_n17688), .A2(new_n17695), .B(new_n18347), .C(new_n17884), .Y(new_n18348));
  A2O1A1Ixp33_ASAP7_75t_L   g18092(.A1(new_n17877), .A2(new_n18346), .B(new_n18348), .C(new_n18138), .Y(new_n18349));
  OAI21xp33_ASAP7_75t_L     g18093(.A1(new_n18148), .A2(new_n18142), .B(new_n18349), .Y(new_n18350));
  A2O1A1O1Ixp25_ASAP7_75t_L g18094(.A1(new_n18136), .A2(\a[59] ), .B(new_n18133), .C(new_n18128), .D(new_n18125), .Y(new_n18351));
  NOR2xp33_ASAP7_75t_L      g18095(.A(new_n2205), .B(new_n11354), .Y(new_n18352));
  AOI221xp5_ASAP7_75t_L     g18096(.A1(\b[26] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[25] ), .C(new_n18352), .Y(new_n18353));
  O2A1O1Ixp33_ASAP7_75t_L   g18097(.A1(new_n11053), .A2(new_n2708), .B(new_n18353), .C(new_n11048), .Y(new_n18354));
  O2A1O1Ixp33_ASAP7_75t_L   g18098(.A1(new_n11053), .A2(new_n2708), .B(new_n18353), .C(\a[59] ), .Y(new_n18355));
  INVx1_ASAP7_75t_L         g18099(.A(new_n18355), .Y(new_n18356));
  OAI21xp33_ASAP7_75t_L     g18100(.A1(new_n11048), .A2(new_n18354), .B(new_n18356), .Y(new_n18357));
  NOR2xp33_ASAP7_75t_L      g18101(.A(new_n1599), .B(new_n13030), .Y(new_n18358));
  O2A1O1Ixp33_ASAP7_75t_L   g18102(.A1(new_n12669), .A2(new_n12671), .B(\b[20] ), .C(new_n18358), .Y(new_n18359));
  A2O1A1Ixp33_ASAP7_75t_L   g18103(.A1(new_n13028), .A2(\b[19] ), .B(new_n18106), .C(new_n18359), .Y(new_n18360));
  A2O1A1Ixp33_ASAP7_75t_L   g18104(.A1(\b[20] ), .A2(new_n13028), .B(new_n18358), .C(new_n18110), .Y(new_n18361));
  NAND2xp33_ASAP7_75t_L     g18105(.A(new_n18361), .B(new_n18360), .Y(new_n18362));
  NOR2xp33_ASAP7_75t_L      g18106(.A(new_n2045), .B(new_n12318), .Y(new_n18363));
  AOI221xp5_ASAP7_75t_L     g18107(.A1(new_n11995), .A2(\b[23] ), .B1(new_n13314), .B2(\b[21] ), .C(new_n18363), .Y(new_n18364));
  INVx1_ASAP7_75t_L         g18108(.A(new_n18364), .Y(new_n18365));
  A2O1A1Ixp33_ASAP7_75t_L   g18109(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n18364), .Y(new_n18366));
  A2O1A1O1Ixp25_ASAP7_75t_L g18110(.A1(new_n2191), .A2(new_n2193), .B(new_n18365), .C(new_n18366), .D(new_n11987), .Y(new_n18367));
  O2A1O1Ixp33_ASAP7_75t_L   g18111(.A1(new_n11998), .A2(new_n2194), .B(new_n18364), .C(\a[62] ), .Y(new_n18368));
  NOR2xp33_ASAP7_75t_L      g18112(.A(new_n18367), .B(new_n18368), .Y(new_n18369));
  NOR2xp33_ASAP7_75t_L      g18113(.A(new_n18362), .B(new_n18369), .Y(new_n18370));
  INVx1_ASAP7_75t_L         g18114(.A(new_n18370), .Y(new_n18371));
  NAND2xp33_ASAP7_75t_L     g18115(.A(new_n18362), .B(new_n18369), .Y(new_n18372));
  AND2x2_ASAP7_75t_L        g18116(.A(new_n18372), .B(new_n18371), .Y(new_n18373));
  INVx1_ASAP7_75t_L         g18117(.A(new_n18373), .Y(new_n18374));
  O2A1O1Ixp33_ASAP7_75t_L   g18118(.A1(new_n18111), .A2(new_n18108), .B(new_n18122), .C(new_n18374), .Y(new_n18375));
  INVx1_ASAP7_75t_L         g18119(.A(new_n18375), .Y(new_n18376));
  O2A1O1Ixp33_ASAP7_75t_L   g18120(.A1(new_n18107), .A2(new_n17854), .B(new_n18110), .C(new_n18121), .Y(new_n18377));
  NAND2xp33_ASAP7_75t_L     g18121(.A(new_n18377), .B(new_n18374), .Y(new_n18378));
  NAND2xp33_ASAP7_75t_L     g18122(.A(new_n18378), .B(new_n18376), .Y(new_n18379));
  XOR2x2_ASAP7_75t_L        g18123(.A(new_n18357), .B(new_n18379), .Y(new_n18380));
  XNOR2x2_ASAP7_75t_L       g18124(.A(new_n18351), .B(new_n18380), .Y(new_n18381));
  INVx1_ASAP7_75t_L         g18125(.A(new_n18381), .Y(new_n18382));
  NOR2xp33_ASAP7_75t_L      g18126(.A(new_n3079), .B(new_n10388), .Y(new_n18383));
  AOI221xp5_ASAP7_75t_L     g18127(.A1(new_n10086), .A2(\b[29] ), .B1(new_n11361), .B2(\b[27] ), .C(new_n18383), .Y(new_n18384));
  O2A1O1Ixp33_ASAP7_75t_L   g18128(.A1(new_n10088), .A2(new_n3104), .B(new_n18384), .C(new_n10083), .Y(new_n18385));
  O2A1O1Ixp33_ASAP7_75t_L   g18129(.A1(new_n10088), .A2(new_n3104), .B(new_n18384), .C(\a[56] ), .Y(new_n18386));
  INVx1_ASAP7_75t_L         g18130(.A(new_n18386), .Y(new_n18387));
  O2A1O1Ixp33_ASAP7_75t_L   g18131(.A1(new_n18385), .A2(new_n10083), .B(new_n18387), .C(new_n18381), .Y(new_n18388));
  INVx1_ASAP7_75t_L         g18132(.A(new_n18388), .Y(new_n18389));
  O2A1O1Ixp33_ASAP7_75t_L   g18133(.A1(new_n18385), .A2(new_n10083), .B(new_n18387), .C(new_n18382), .Y(new_n18390));
  A2O1A1Ixp33_ASAP7_75t_L   g18134(.A1(new_n18389), .A2(new_n18382), .B(new_n18390), .C(new_n18350), .Y(new_n18391));
  INVx1_ASAP7_75t_L         g18135(.A(new_n18390), .Y(new_n18392));
  O2A1O1Ixp33_ASAP7_75t_L   g18136(.A1(new_n18381), .A2(new_n18388), .B(new_n18392), .C(new_n18350), .Y(new_n18393));
  NOR2xp33_ASAP7_75t_L      g18137(.A(new_n3674), .B(new_n10400), .Y(new_n18394));
  AOI221xp5_ASAP7_75t_L     g18138(.A1(new_n9102), .A2(\b[32] ), .B1(new_n10398), .B2(\b[30] ), .C(new_n18394), .Y(new_n18395));
  INVx1_ASAP7_75t_L         g18139(.A(new_n18395), .Y(new_n18396));
  O2A1O1Ixp33_ASAP7_75t_L   g18140(.A1(new_n9104), .A2(new_n3897), .B(new_n18395), .C(new_n9099), .Y(new_n18397));
  INVx1_ASAP7_75t_L         g18141(.A(new_n18397), .Y(new_n18398));
  NOR2xp33_ASAP7_75t_L      g18142(.A(new_n9099), .B(new_n18397), .Y(new_n18399));
  A2O1A1O1Ixp25_ASAP7_75t_L g18143(.A1(new_n9437), .A2(new_n3900), .B(new_n18396), .C(new_n18398), .D(new_n18399), .Y(new_n18400));
  A2O1A1Ixp33_ASAP7_75t_L   g18144(.A1(new_n18391), .A2(new_n18350), .B(new_n18393), .C(new_n18400), .Y(new_n18401));
  INVx1_ASAP7_75t_L         g18145(.A(new_n18391), .Y(new_n18402));
  O2A1O1Ixp33_ASAP7_75t_L   g18146(.A1(new_n18142), .A2(new_n18148), .B(new_n18349), .C(new_n18402), .Y(new_n18403));
  A2O1A1O1Ixp25_ASAP7_75t_L g18147(.A1(new_n18389), .A2(new_n18382), .B(new_n18390), .C(new_n18391), .D(new_n18403), .Y(new_n18404));
  O2A1O1Ixp33_ASAP7_75t_L   g18148(.A1(new_n9104), .A2(new_n3897), .B(new_n18395), .C(\a[53] ), .Y(new_n18405));
  A2O1A1Ixp33_ASAP7_75t_L   g18149(.A1(\a[53] ), .A2(new_n18398), .B(new_n18405), .C(new_n18404), .Y(new_n18406));
  NAND2xp33_ASAP7_75t_L     g18150(.A(new_n18401), .B(new_n18406), .Y(new_n18407));
  A2O1A1Ixp33_ASAP7_75t_L   g18151(.A1(new_n18344), .A2(new_n18343), .B(new_n18159), .C(new_n18407), .Y(new_n18408));
  A2O1A1O1Ixp25_ASAP7_75t_L g18152(.A1(new_n18160), .A2(\a[53] ), .B(new_n18157), .C(new_n18152), .D(new_n18150), .Y(new_n18409));
  NAND3xp33_ASAP7_75t_L     g18153(.A(new_n18406), .B(new_n18401), .C(new_n18409), .Y(new_n18410));
  AND2x2_ASAP7_75t_L        g18154(.A(new_n18410), .B(new_n18408), .Y(new_n18411));
  A2O1A1Ixp33_ASAP7_75t_L   g18155(.A1(new_n18341), .A2(\a[50] ), .B(new_n18342), .C(new_n18411), .Y(new_n18412));
  AO221x2_ASAP7_75t_L       g18156(.A1(\a[50] ), .A2(new_n18341), .B1(new_n18408), .B2(new_n18410), .C(new_n18342), .Y(new_n18413));
  AND2x2_ASAP7_75t_L        g18157(.A(new_n18413), .B(new_n18412), .Y(new_n18414));
  NAND2xp33_ASAP7_75t_L     g18158(.A(new_n18337), .B(new_n18414), .Y(new_n18415));
  NAND2xp33_ASAP7_75t_L     g18159(.A(new_n18413), .B(new_n18412), .Y(new_n18416));
  NAND2xp33_ASAP7_75t_L     g18160(.A(new_n18336), .B(new_n18416), .Y(new_n18417));
  NAND2xp33_ASAP7_75t_L     g18161(.A(new_n18417), .B(new_n18415), .Y(new_n18418));
  O2A1O1Ixp33_ASAP7_75t_L   g18162(.A1(new_n7316), .A2(new_n18333), .B(new_n18335), .C(new_n18418), .Y(new_n18419));
  INVx1_ASAP7_75t_L         g18163(.A(new_n18333), .Y(new_n18420));
  AOI221xp5_ASAP7_75t_L     g18164(.A1(\a[47] ), .A2(new_n18420), .B1(new_n18417), .B2(new_n18415), .C(new_n18334), .Y(new_n18421));
  NOR2xp33_ASAP7_75t_L      g18165(.A(new_n18421), .B(new_n18419), .Y(new_n18422));
  XNOR2x2_ASAP7_75t_L       g18166(.A(new_n18330), .B(new_n18422), .Y(new_n18423));
  XNOR2x2_ASAP7_75t_L       g18167(.A(new_n18327), .B(new_n18423), .Y(new_n18424));
  XOR2x2_ASAP7_75t_L        g18168(.A(new_n18321), .B(new_n18424), .Y(new_n18425));
  XOR2x2_ASAP7_75t_L        g18169(.A(new_n18318), .B(new_n18425), .Y(new_n18426));
  XOR2x2_ASAP7_75t_L        g18170(.A(new_n18312), .B(new_n18426), .Y(new_n18427));
  NOR2xp33_ASAP7_75t_L      g18171(.A(new_n7552), .B(new_n4908), .Y(new_n18428));
  AOI221xp5_ASAP7_75t_L     g18172(.A1(\b[45] ), .A2(new_n5139), .B1(\b[46] ), .B2(new_n4916), .C(new_n18428), .Y(new_n18429));
  O2A1O1Ixp33_ASAP7_75t_L   g18173(.A1(new_n4911), .A2(new_n7560), .B(new_n18429), .C(new_n4906), .Y(new_n18430));
  O2A1O1Ixp33_ASAP7_75t_L   g18174(.A1(new_n4911), .A2(new_n7560), .B(new_n18429), .C(\a[38] ), .Y(new_n18431));
  INVx1_ASAP7_75t_L         g18175(.A(new_n18431), .Y(new_n18432));
  O2A1O1Ixp33_ASAP7_75t_L   g18176(.A1(new_n18430), .A2(new_n4906), .B(new_n18432), .C(new_n18427), .Y(new_n18433));
  INVx1_ASAP7_75t_L         g18177(.A(new_n18430), .Y(new_n18434));
  A2O1A1Ixp33_ASAP7_75t_L   g18178(.A1(\a[38] ), .A2(new_n18434), .B(new_n18431), .C(new_n18427), .Y(new_n18435));
  INVx1_ASAP7_75t_L         g18179(.A(new_n18214), .Y(new_n18436));
  A2O1A1O1Ixp25_ASAP7_75t_L g18180(.A1(new_n18436), .A2(\a[38] ), .B(new_n18215), .C(new_n18210), .D(new_n18209), .Y(new_n18437));
  OAI211xp5_ASAP7_75t_L     g18181(.A1(new_n18427), .A2(new_n18433), .B(new_n18435), .C(new_n18437), .Y(new_n18438));
  OAI21xp33_ASAP7_75t_L     g18182(.A1(new_n18427), .A2(new_n18433), .B(new_n18435), .Y(new_n18439));
  INVx1_ASAP7_75t_L         g18183(.A(new_n18437), .Y(new_n18440));
  NAND2xp33_ASAP7_75t_L     g18184(.A(new_n18440), .B(new_n18439), .Y(new_n18441));
  NAND2xp33_ASAP7_75t_L     g18185(.A(new_n18438), .B(new_n18441), .Y(new_n18442));
  NOR2xp33_ASAP7_75t_L      g18186(.A(new_n8755), .B(new_n4147), .Y(new_n18443));
  AOI221xp5_ASAP7_75t_L     g18187(.A1(\b[48] ), .A2(new_n4402), .B1(\b[49] ), .B2(new_n4155), .C(new_n18443), .Y(new_n18444));
  O2A1O1Ixp33_ASAP7_75t_L   g18188(.A1(new_n4150), .A2(new_n8764), .B(new_n18444), .C(new_n4145), .Y(new_n18445));
  O2A1O1Ixp33_ASAP7_75t_L   g18189(.A1(new_n4150), .A2(new_n8764), .B(new_n18444), .C(\a[35] ), .Y(new_n18446));
  INVx1_ASAP7_75t_L         g18190(.A(new_n18446), .Y(new_n18447));
  OA21x2_ASAP7_75t_L        g18191(.A1(new_n4145), .A2(new_n18445), .B(new_n18447), .Y(new_n18448));
  NOR2xp33_ASAP7_75t_L      g18192(.A(new_n9683), .B(new_n3510), .Y(new_n18449));
  AOI221xp5_ASAP7_75t_L     g18193(.A1(\b[51] ), .A2(new_n3708), .B1(\b[52] ), .B2(new_n3499), .C(new_n18449), .Y(new_n18450));
  O2A1O1Ixp33_ASAP7_75t_L   g18194(.A1(new_n3513), .A2(new_n9691), .B(new_n18450), .C(new_n3493), .Y(new_n18451));
  O2A1O1Ixp33_ASAP7_75t_L   g18195(.A1(new_n3513), .A2(new_n9691), .B(new_n18450), .C(\a[32] ), .Y(new_n18452));
  INVx1_ASAP7_75t_L         g18196(.A(new_n18452), .Y(new_n18453));
  A2O1A1O1Ixp25_ASAP7_75t_L g18197(.A1(new_n18230), .A2(\a[35] ), .B(new_n18231), .C(new_n18223), .D(new_n18224), .Y(new_n18454));
  OAI211xp5_ASAP7_75t_L     g18198(.A1(new_n3493), .A2(new_n18451), .B(new_n18454), .C(new_n18453), .Y(new_n18455));
  O2A1O1Ixp33_ASAP7_75t_L   g18199(.A1(new_n3493), .A2(new_n18451), .B(new_n18453), .C(new_n18454), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18456), .Y(new_n18457));
  NAND2xp33_ASAP7_75t_L     g18201(.A(new_n18448), .B(new_n18442), .Y(new_n18458));
  AND3x1_ASAP7_75t_L        g18202(.A(new_n18458), .B(new_n18457), .C(new_n18455), .Y(new_n18459));
  OAI21xp33_ASAP7_75t_L     g18203(.A1(new_n18442), .A2(new_n18448), .B(new_n18459), .Y(new_n18460));
  AND3x1_ASAP7_75t_L        g18204(.A(new_n18460), .B(new_n18457), .C(new_n18455), .Y(new_n18461));
  AND2x2_ASAP7_75t_L        g18205(.A(new_n18458), .B(new_n18460), .Y(new_n18462));
  O2A1O1Ixp33_ASAP7_75t_L   g18206(.A1(new_n18448), .A2(new_n18442), .B(new_n18462), .C(new_n18461), .Y(new_n18463));
  XNOR2x2_ASAP7_75t_L       g18207(.A(new_n18463), .B(new_n18310), .Y(new_n18464));
  NAND2xp33_ASAP7_75t_L     g18208(.A(\b[58] ), .B(new_n2421), .Y(new_n18465));
  OAI221xp5_ASAP7_75t_L     g18209(.A1(new_n2415), .A2(new_n11591), .B1(new_n10978), .B2(new_n2572), .C(new_n18465), .Y(new_n18466));
  A2O1A1Ixp33_ASAP7_75t_L   g18210(.A1(new_n12577), .A2(new_n2417), .B(new_n18466), .C(\a[26] ), .Y(new_n18467));
  NAND2xp33_ASAP7_75t_L     g18211(.A(\a[26] ), .B(new_n18467), .Y(new_n18468));
  A2O1A1Ixp33_ASAP7_75t_L   g18212(.A1(new_n12577), .A2(new_n2417), .B(new_n18466), .C(new_n2413), .Y(new_n18469));
  NAND2xp33_ASAP7_75t_L     g18213(.A(new_n18469), .B(new_n18468), .Y(new_n18470));
  OAI31xp33_ASAP7_75t_L     g18214(.A1(new_n18084), .A2(new_n18237), .A3(new_n18241), .B(new_n18085), .Y(new_n18471));
  NOR2xp33_ASAP7_75t_L      g18215(.A(new_n18470), .B(new_n18471), .Y(new_n18472));
  INVx1_ASAP7_75t_L         g18216(.A(new_n18471), .Y(new_n18473));
  AOI21xp33_ASAP7_75t_L     g18217(.A1(new_n18469), .A2(new_n18468), .B(new_n18473), .Y(new_n18474));
  NOR2xp33_ASAP7_75t_L      g18218(.A(new_n18472), .B(new_n18474), .Y(new_n18475));
  NAND2xp33_ASAP7_75t_L     g18219(.A(new_n18464), .B(new_n18475), .Y(new_n18476));
  NOR3xp33_ASAP7_75t_L      g18220(.A(new_n18464), .B(new_n18474), .C(new_n18472), .Y(new_n18477));
  AOI21xp33_ASAP7_75t_L     g18221(.A1(new_n18476), .A2(new_n18464), .B(new_n18477), .Y(new_n18478));
  A2O1A1Ixp33_ASAP7_75t_L   g18222(.A1(new_n18299), .A2(new_n18297), .B(new_n18300), .C(new_n18478), .Y(new_n18479));
  A2O1A1O1Ixp25_ASAP7_75t_L g18223(.A1(new_n18294), .A2(\a[23] ), .B(new_n18295), .C(new_n18299), .D(new_n18300), .Y(new_n18480));
  A2O1A1Ixp33_ASAP7_75t_L   g18224(.A1(new_n18464), .A2(new_n18476), .B(new_n18477), .C(new_n18480), .Y(new_n18481));
  NAND2xp33_ASAP7_75t_L     g18225(.A(new_n18479), .B(new_n18481), .Y(new_n18482));
  A2O1A1Ixp33_ASAP7_75t_L   g18226(.A1(new_n18289), .A2(new_n18284), .B(new_n18290), .C(new_n18482), .Y(new_n18483));
  A2O1A1Ixp33_ASAP7_75t_L   g18227(.A1(new_n18288), .A2(new_n18260), .B(new_n18066), .C(new_n18283), .Y(new_n18484));
  AOI31xp33_ASAP7_75t_L     g18228(.A1(new_n18260), .A2(new_n18247), .A3(new_n18285), .B(new_n18066), .Y(new_n18485));
  A2O1A1O1Ixp25_ASAP7_75t_L g18229(.A1(new_n12603), .A2(new_n14444), .B(new_n1521), .C(new_n1654), .D(new_n12956), .Y(new_n18486));
  A2O1A1Ixp33_ASAP7_75t_L   g18230(.A1(new_n18486), .A2(new_n18281), .B(new_n18282), .C(new_n18485), .Y(new_n18487));
  NAND4xp25_ASAP7_75t_L     g18231(.A(new_n18484), .B(new_n18481), .C(new_n18479), .D(new_n18487), .Y(new_n18488));
  NAND2xp33_ASAP7_75t_L     g18232(.A(new_n18488), .B(new_n18483), .Y(new_n18489));
  O2A1O1Ixp33_ASAP7_75t_L   g18233(.A1(new_n18049), .A2(new_n18056), .B(new_n18271), .C(new_n18489), .Y(new_n18490));
  A2O1A1Ixp33_ASAP7_75t_L   g18234(.A1(new_n18253), .A2(new_n18056), .B(new_n18251), .C(new_n18263), .Y(new_n18491));
  AOI21xp33_ASAP7_75t_L     g18235(.A1(new_n18483), .A2(new_n18488), .B(new_n18491), .Y(new_n18492));
  NOR2xp33_ASAP7_75t_L      g18236(.A(new_n18492), .B(new_n18490), .Y(new_n18493));
  INVx1_ASAP7_75t_L         g18237(.A(new_n18493), .Y(new_n18494));
  A2O1A1O1Ixp25_ASAP7_75t_L g18238(.A1(new_n18266), .A2(new_n18042), .B(new_n18273), .C(new_n18279), .D(new_n18494), .Y(new_n18495));
  A2O1A1Ixp33_ASAP7_75t_L   g18239(.A1(new_n18266), .A2(new_n18042), .B(new_n18273), .C(new_n18279), .Y(new_n18496));
  NOR2xp33_ASAP7_75t_L      g18240(.A(new_n18493), .B(new_n18496), .Y(new_n18497));
  NOR2xp33_ASAP7_75t_L      g18241(.A(new_n18497), .B(new_n18495), .Y(\f[83] ));
  INVx1_ASAP7_75t_L         g18242(.A(new_n18300), .Y(new_n18499));
  O2A1O1Ixp33_ASAP7_75t_L   g18243(.A1(new_n18296), .A2(new_n18298), .B(new_n18499), .C(new_n18478), .Y(new_n18500));
  OAI22xp33_ASAP7_75t_L     g18244(.A1(new_n2089), .A2(new_n12258), .B1(new_n12603), .B2(new_n1962), .Y(new_n18501));
  AOI221xp5_ASAP7_75t_L     g18245(.A1(new_n1955), .A2(\b[63] ), .B1(new_n1964), .B2(new_n12961), .C(new_n18501), .Y(new_n18502));
  XNOR2x2_ASAP7_75t_L       g18246(.A(new_n1952), .B(new_n18502), .Y(new_n18503));
  A2O1A1O1Ixp25_ASAP7_75t_L g18247(.A1(new_n18296), .A2(new_n18499), .B(new_n18478), .C(new_n18299), .D(new_n18503), .Y(new_n18504));
  INVx1_ASAP7_75t_L         g18248(.A(new_n18504), .Y(new_n18505));
  NOR2xp33_ASAP7_75t_L      g18249(.A(new_n18503), .B(new_n18504), .Y(new_n18506));
  O2A1O1Ixp33_ASAP7_75t_L   g18250(.A1(new_n18298), .A2(new_n18500), .B(new_n18505), .C(new_n18506), .Y(new_n18507));
  INVx1_ASAP7_75t_L         g18251(.A(new_n18507), .Y(new_n18508));
  OAI22xp33_ASAP7_75t_L     g18252(.A1(new_n2572), .A2(new_n11303), .B1(new_n11591), .B2(new_n2410), .Y(new_n18509));
  AOI221xp5_ASAP7_75t_L     g18253(.A1(new_n2423), .A2(\b[60] ), .B1(new_n2417), .B2(new_n13839), .C(new_n18509), .Y(new_n18510));
  XNOR2x2_ASAP7_75t_L       g18254(.A(new_n2413), .B(new_n18510), .Y(new_n18511));
  INVx1_ASAP7_75t_L         g18255(.A(new_n18511), .Y(new_n18512));
  A2O1A1Ixp33_ASAP7_75t_L   g18256(.A1(new_n18469), .A2(new_n18468), .B(new_n18473), .C(new_n18476), .Y(new_n18513));
  NOR2xp33_ASAP7_75t_L      g18257(.A(new_n18512), .B(new_n18513), .Y(new_n18514));
  A2O1A1Ixp33_ASAP7_75t_L   g18258(.A1(new_n18475), .A2(new_n18464), .B(new_n18474), .C(new_n18512), .Y(new_n18515));
  INVx1_ASAP7_75t_L         g18259(.A(new_n18515), .Y(new_n18516));
  NOR2xp33_ASAP7_75t_L      g18260(.A(new_n18516), .B(new_n18514), .Y(new_n18517));
  A2O1A1Ixp33_ASAP7_75t_L   g18261(.A1(new_n18097), .A2(new_n18240), .B(new_n18096), .C(new_n18307), .Y(new_n18518));
  A2O1A1Ixp33_ASAP7_75t_L   g18262(.A1(new_n18309), .A2(new_n18518), .B(new_n18463), .C(new_n18307), .Y(new_n18519));
  OAI22xp33_ASAP7_75t_L     g18263(.A1(new_n3133), .A2(new_n10309), .B1(new_n10332), .B2(new_n2925), .Y(new_n18520));
  AOI221xp5_ASAP7_75t_L     g18264(.A1(new_n2938), .A2(\b[57] ), .B1(new_n2932), .B2(new_n10991), .C(new_n18520), .Y(new_n18521));
  XNOR2x2_ASAP7_75t_L       g18265(.A(new_n2928), .B(new_n18521), .Y(new_n18522));
  XNOR2x2_ASAP7_75t_L       g18266(.A(new_n18522), .B(new_n18519), .Y(new_n18523));
  OAI22xp33_ASAP7_75t_L     g18267(.A1(new_n3703), .A2(new_n9355), .B1(new_n9683), .B2(new_n3509), .Y(new_n18524));
  AOI221xp5_ASAP7_75t_L     g18268(.A1(new_n3503), .A2(\b[54] ), .B1(new_n3505), .B2(new_n9717), .C(new_n18524), .Y(new_n18525));
  XNOR2x2_ASAP7_75t_L       g18269(.A(new_n3493), .B(new_n18525), .Y(new_n18526));
  O2A1O1Ixp33_ASAP7_75t_L   g18270(.A1(new_n18442), .A2(new_n18448), .B(new_n18459), .C(new_n18456), .Y(new_n18527));
  NAND2xp33_ASAP7_75t_L     g18271(.A(new_n18526), .B(new_n18527), .Y(new_n18528));
  AO21x2_ASAP7_75t_L        g18272(.A1(new_n18457), .A2(new_n18460), .B(new_n18526), .Y(new_n18529));
  AND2x2_ASAP7_75t_L        g18273(.A(new_n18528), .B(new_n18529), .Y(new_n18530));
  INVx1_ASAP7_75t_L         g18274(.A(new_n18412), .Y(new_n18531));
  O2A1O1Ixp33_ASAP7_75t_L   g18275(.A1(new_n18150), .A2(new_n18159), .B(new_n18407), .C(new_n18531), .Y(new_n18532));
  NOR2xp33_ASAP7_75t_L      g18276(.A(new_n1745), .B(new_n13030), .Y(new_n18533));
  A2O1A1Ixp33_ASAP7_75t_L   g18277(.A1(new_n13028), .A2(\b[21] ), .B(new_n18533), .C(new_n1501), .Y(new_n18534));
  INVx1_ASAP7_75t_L         g18278(.A(new_n18534), .Y(new_n18535));
  O2A1O1Ixp33_ASAP7_75t_L   g18279(.A1(new_n12669), .A2(new_n12671), .B(\b[21] ), .C(new_n18533), .Y(new_n18536));
  NAND2xp33_ASAP7_75t_L     g18280(.A(\a[20] ), .B(new_n18536), .Y(new_n18537));
  INVx1_ASAP7_75t_L         g18281(.A(new_n18537), .Y(new_n18538));
  NOR2xp33_ASAP7_75t_L      g18282(.A(new_n18535), .B(new_n18538), .Y(new_n18539));
  A2O1A1Ixp33_ASAP7_75t_L   g18283(.A1(new_n13028), .A2(\b[20] ), .B(new_n18358), .C(new_n18539), .Y(new_n18540));
  OAI21xp33_ASAP7_75t_L     g18284(.A1(new_n18535), .A2(new_n18538), .B(new_n18359), .Y(new_n18541));
  AND2x2_ASAP7_75t_L        g18285(.A(new_n18541), .B(new_n18540), .Y(new_n18542));
  INVx1_ASAP7_75t_L         g18286(.A(new_n18542), .Y(new_n18543));
  NOR2xp33_ASAP7_75t_L      g18287(.A(new_n2188), .B(new_n12318), .Y(new_n18544));
  AOI221xp5_ASAP7_75t_L     g18288(.A1(new_n11995), .A2(\b[24] ), .B1(new_n13314), .B2(\b[22] ), .C(new_n18544), .Y(new_n18545));
  O2A1O1Ixp33_ASAP7_75t_L   g18289(.A1(new_n11998), .A2(new_n2853), .B(new_n18545), .C(new_n11987), .Y(new_n18546));
  O2A1O1Ixp33_ASAP7_75t_L   g18290(.A1(new_n11998), .A2(new_n2853), .B(new_n18545), .C(\a[62] ), .Y(new_n18547));
  INVx1_ASAP7_75t_L         g18291(.A(new_n18547), .Y(new_n18548));
  O2A1O1Ixp33_ASAP7_75t_L   g18292(.A1(new_n11987), .A2(new_n18546), .B(new_n18548), .C(new_n18543), .Y(new_n18549));
  INVx1_ASAP7_75t_L         g18293(.A(new_n18549), .Y(new_n18550));
  O2A1O1Ixp33_ASAP7_75t_L   g18294(.A1(new_n11987), .A2(new_n18546), .B(new_n18548), .C(new_n18542), .Y(new_n18551));
  AOI21xp33_ASAP7_75t_L     g18295(.A1(new_n18550), .A2(new_n18542), .B(new_n18551), .Y(new_n18552));
  INVx1_ASAP7_75t_L         g18296(.A(new_n18552), .Y(new_n18553));
  INVx1_ASAP7_75t_L         g18297(.A(new_n18359), .Y(new_n18554));
  O2A1O1Ixp33_ASAP7_75t_L   g18298(.A1(new_n18110), .A2(new_n18554), .B(new_n18371), .C(new_n18552), .Y(new_n18555));
  INVx1_ASAP7_75t_L         g18299(.A(new_n18555), .Y(new_n18556));
  O2A1O1Ixp33_ASAP7_75t_L   g18300(.A1(new_n18110), .A2(new_n18554), .B(new_n18371), .C(new_n18553), .Y(new_n18557));
  A2O1A1O1Ixp25_ASAP7_75t_L g18301(.A1(new_n13028), .A2(\b[19] ), .B(new_n18106), .C(new_n18359), .D(new_n18370), .Y(new_n18558));
  A2O1A1Ixp33_ASAP7_75t_L   g18302(.A1(new_n18550), .A2(new_n18542), .B(new_n18551), .C(new_n18558), .Y(new_n18559));
  A2O1A1Ixp33_ASAP7_75t_L   g18303(.A1(new_n18371), .A2(new_n18360), .B(new_n18555), .C(new_n18559), .Y(new_n18560));
  NOR2xp33_ASAP7_75t_L      g18304(.A(new_n2377), .B(new_n11354), .Y(new_n18561));
  AOI221xp5_ASAP7_75t_L     g18305(.A1(\b[27] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[26] ), .C(new_n18561), .Y(new_n18562));
  O2A1O1Ixp33_ASAP7_75t_L   g18306(.A1(new_n11053), .A2(new_n2889), .B(new_n18562), .C(new_n11048), .Y(new_n18563));
  INVx1_ASAP7_75t_L         g18307(.A(new_n18563), .Y(new_n18564));
  O2A1O1Ixp33_ASAP7_75t_L   g18308(.A1(new_n11053), .A2(new_n2889), .B(new_n18562), .C(\a[59] ), .Y(new_n18565));
  A2O1A1Ixp33_ASAP7_75t_L   g18309(.A1(\a[59] ), .A2(new_n18564), .B(new_n18565), .C(new_n18560), .Y(new_n18566));
  INVx1_ASAP7_75t_L         g18310(.A(new_n18565), .Y(new_n18567));
  O2A1O1Ixp33_ASAP7_75t_L   g18311(.A1(new_n18563), .A2(new_n11048), .B(new_n18567), .C(new_n18560), .Y(new_n18568));
  A2O1A1O1Ixp25_ASAP7_75t_L g18312(.A1(new_n18556), .A2(new_n18553), .B(new_n18557), .C(new_n18566), .D(new_n18568), .Y(new_n18569));
  O2A1O1Ixp33_ASAP7_75t_L   g18313(.A1(new_n11048), .A2(new_n18354), .B(new_n18356), .C(new_n18379), .Y(new_n18570));
  O2A1O1Ixp33_ASAP7_75t_L   g18314(.A1(new_n18112), .A2(new_n18121), .B(new_n18373), .C(new_n18570), .Y(new_n18571));
  NAND2xp33_ASAP7_75t_L     g18315(.A(new_n18569), .B(new_n18571), .Y(new_n18572));
  INVx1_ASAP7_75t_L         g18316(.A(new_n18570), .Y(new_n18573));
  O2A1O1Ixp33_ASAP7_75t_L   g18317(.A1(new_n18377), .A2(new_n18374), .B(new_n18573), .C(new_n18569), .Y(new_n18574));
  INVx1_ASAP7_75t_L         g18318(.A(new_n18574), .Y(new_n18575));
  NAND2xp33_ASAP7_75t_L     g18319(.A(new_n18572), .B(new_n18575), .Y(new_n18576));
  INVx1_ASAP7_75t_L         g18320(.A(new_n18576), .Y(new_n18577));
  NOR2xp33_ASAP7_75t_L      g18321(.A(new_n3098), .B(new_n10388), .Y(new_n18578));
  AOI221xp5_ASAP7_75t_L     g18322(.A1(new_n10086), .A2(\b[30] ), .B1(new_n11361), .B2(\b[28] ), .C(new_n18578), .Y(new_n18579));
  O2A1O1Ixp33_ASAP7_75t_L   g18323(.A1(new_n10088), .A2(new_n3464), .B(new_n18579), .C(new_n10083), .Y(new_n18580));
  O2A1O1Ixp33_ASAP7_75t_L   g18324(.A1(new_n10088), .A2(new_n3464), .B(new_n18579), .C(\a[56] ), .Y(new_n18581));
  INVx1_ASAP7_75t_L         g18325(.A(new_n18581), .Y(new_n18582));
  O2A1O1Ixp33_ASAP7_75t_L   g18326(.A1(new_n18580), .A2(new_n10083), .B(new_n18582), .C(new_n18576), .Y(new_n18583));
  INVx1_ASAP7_75t_L         g18327(.A(new_n18583), .Y(new_n18584));
  O2A1O1Ixp33_ASAP7_75t_L   g18328(.A1(new_n18580), .A2(new_n10083), .B(new_n18582), .C(new_n18577), .Y(new_n18585));
  INVx1_ASAP7_75t_L         g18329(.A(new_n18135), .Y(new_n18586));
  O2A1O1Ixp33_ASAP7_75t_L   g18330(.A1(new_n18124), .A2(new_n18127), .B(new_n18586), .C(new_n18380), .Y(new_n18587));
  INVx1_ASAP7_75t_L         g18331(.A(new_n18385), .Y(new_n18588));
  A2O1A1O1Ixp25_ASAP7_75t_L g18332(.A1(new_n18588), .A2(\a[56] ), .B(new_n18386), .C(new_n18382), .D(new_n18587), .Y(new_n18589));
  INVx1_ASAP7_75t_L         g18333(.A(new_n18589), .Y(new_n18590));
  AOI211xp5_ASAP7_75t_L     g18334(.A1(new_n18584), .A2(new_n18577), .B(new_n18585), .C(new_n18590), .Y(new_n18591));
  INVx1_ASAP7_75t_L         g18335(.A(new_n18585), .Y(new_n18592));
  O2A1O1Ixp33_ASAP7_75t_L   g18336(.A1(new_n18576), .A2(new_n18583), .B(new_n18592), .C(new_n18589), .Y(new_n18593));
  NOR2xp33_ASAP7_75t_L      g18337(.A(new_n18591), .B(new_n18593), .Y(new_n18594));
  NOR2xp33_ASAP7_75t_L      g18338(.A(new_n3891), .B(new_n10400), .Y(new_n18595));
  AOI221xp5_ASAP7_75t_L     g18339(.A1(new_n9102), .A2(\b[33] ), .B1(new_n10398), .B2(\b[31] ), .C(new_n18595), .Y(new_n18596));
  O2A1O1Ixp33_ASAP7_75t_L   g18340(.A1(new_n9104), .A2(new_n4108), .B(new_n18596), .C(new_n9099), .Y(new_n18597));
  NOR2xp33_ASAP7_75t_L      g18341(.A(new_n9099), .B(new_n18597), .Y(new_n18598));
  O2A1O1Ixp33_ASAP7_75t_L   g18342(.A1(new_n9104), .A2(new_n4108), .B(new_n18596), .C(\a[53] ), .Y(new_n18599));
  NOR2xp33_ASAP7_75t_L      g18343(.A(new_n18599), .B(new_n18598), .Y(new_n18600));
  INVx1_ASAP7_75t_L         g18344(.A(new_n18400), .Y(new_n18601));
  O2A1O1Ixp33_ASAP7_75t_L   g18345(.A1(new_n18350), .A2(new_n18393), .B(new_n18601), .C(new_n18402), .Y(new_n18602));
  XNOR2x2_ASAP7_75t_L       g18346(.A(new_n18600), .B(new_n18602), .Y(new_n18603));
  XNOR2x2_ASAP7_75t_L       g18347(.A(new_n18594), .B(new_n18603), .Y(new_n18604));
  NOR2xp33_ASAP7_75t_L      g18348(.A(new_n4581), .B(new_n10065), .Y(new_n18605));
  AOI221xp5_ASAP7_75t_L     g18349(.A1(new_n8175), .A2(\b[36] ), .B1(new_n8484), .B2(\b[34] ), .C(new_n18605), .Y(new_n18606));
  O2A1O1Ixp33_ASAP7_75t_L   g18350(.A1(new_n8176), .A2(new_n4622), .B(new_n18606), .C(new_n8172), .Y(new_n18607));
  INVx1_ASAP7_75t_L         g18351(.A(new_n18607), .Y(new_n18608));
  O2A1O1Ixp33_ASAP7_75t_L   g18352(.A1(new_n8176), .A2(new_n4622), .B(new_n18606), .C(\a[50] ), .Y(new_n18609));
  A2O1A1Ixp33_ASAP7_75t_L   g18353(.A1(\a[50] ), .A2(new_n18608), .B(new_n18609), .C(new_n18604), .Y(new_n18610));
  NOR2xp33_ASAP7_75t_L      g18354(.A(new_n8172), .B(new_n18607), .Y(new_n18611));
  OR3x1_ASAP7_75t_L         g18355(.A(new_n18604), .B(new_n18611), .C(new_n18609), .Y(new_n18612));
  NAND2xp33_ASAP7_75t_L     g18356(.A(new_n18610), .B(new_n18612), .Y(new_n18613));
  NAND2xp33_ASAP7_75t_L     g18357(.A(new_n18613), .B(new_n18532), .Y(new_n18614));
  A2O1A1O1Ixp25_ASAP7_75t_L g18358(.A1(new_n18401), .A2(new_n18406), .B(new_n18409), .C(new_n18412), .D(new_n18613), .Y(new_n18615));
  INVx1_ASAP7_75t_L         g18359(.A(new_n18615), .Y(new_n18616));
  NAND2xp33_ASAP7_75t_L     g18360(.A(new_n18616), .B(new_n18614), .Y(new_n18617));
  NOR2xp33_ASAP7_75t_L      g18361(.A(new_n5570), .B(new_n7318), .Y(new_n18618));
  AOI221xp5_ASAP7_75t_L     g18362(.A1(new_n7333), .A2(\b[38] ), .B1(new_n7609), .B2(\b[37] ), .C(new_n18618), .Y(new_n18619));
  O2A1O1Ixp33_ASAP7_75t_L   g18363(.A1(new_n7321), .A2(new_n5578), .B(new_n18619), .C(new_n7316), .Y(new_n18620));
  O2A1O1Ixp33_ASAP7_75t_L   g18364(.A1(new_n7321), .A2(new_n5578), .B(new_n18619), .C(\a[47] ), .Y(new_n18621));
  INVx1_ASAP7_75t_L         g18365(.A(new_n18621), .Y(new_n18622));
  O2A1O1Ixp33_ASAP7_75t_L   g18366(.A1(new_n18620), .A2(new_n7316), .B(new_n18622), .C(new_n18617), .Y(new_n18623));
  INVx1_ASAP7_75t_L         g18367(.A(new_n18620), .Y(new_n18624));
  A2O1A1Ixp33_ASAP7_75t_L   g18368(.A1(\a[47] ), .A2(new_n18624), .B(new_n18621), .C(new_n18617), .Y(new_n18625));
  A2O1A1O1Ixp25_ASAP7_75t_L g18369(.A1(new_n17918), .A2(new_n17916), .B(new_n18162), .C(new_n18173), .D(new_n18416), .Y(new_n18626));
  A2O1A1O1Ixp25_ASAP7_75t_L g18370(.A1(new_n18420), .A2(\a[47] ), .B(new_n18334), .C(new_n18417), .D(new_n18626), .Y(new_n18627));
  OAI211xp5_ASAP7_75t_L     g18371(.A1(new_n18617), .A2(new_n18623), .B(new_n18625), .C(new_n18627), .Y(new_n18628));
  OAI21xp33_ASAP7_75t_L     g18372(.A1(new_n18617), .A2(new_n18623), .B(new_n18625), .Y(new_n18629));
  A2O1A1Ixp33_ASAP7_75t_L   g18373(.A1(new_n18414), .A2(new_n18337), .B(new_n18419), .C(new_n18629), .Y(new_n18630));
  NAND2xp33_ASAP7_75t_L     g18374(.A(new_n18628), .B(new_n18630), .Y(new_n18631));
  NOR2xp33_ASAP7_75t_L      g18375(.A(new_n5855), .B(new_n6741), .Y(new_n18632));
  AOI221xp5_ASAP7_75t_L     g18376(.A1(\b[42] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[41] ), .C(new_n18632), .Y(new_n18633));
  O2A1O1Ixp33_ASAP7_75t_L   g18377(.A1(new_n6443), .A2(new_n6386), .B(new_n18633), .C(new_n6439), .Y(new_n18634));
  O2A1O1Ixp33_ASAP7_75t_L   g18378(.A1(new_n6443), .A2(new_n6386), .B(new_n18633), .C(\a[44] ), .Y(new_n18635));
  INVx1_ASAP7_75t_L         g18379(.A(new_n18635), .Y(new_n18636));
  O2A1O1Ixp33_ASAP7_75t_L   g18380(.A1(new_n18634), .A2(new_n6439), .B(new_n18636), .C(new_n18631), .Y(new_n18637));
  INVx1_ASAP7_75t_L         g18381(.A(new_n18634), .Y(new_n18638));
  A2O1A1Ixp33_ASAP7_75t_L   g18382(.A1(\a[44] ), .A2(new_n18638), .B(new_n18635), .C(new_n18631), .Y(new_n18639));
  OAI21xp33_ASAP7_75t_L     g18383(.A1(new_n18631), .A2(new_n18637), .B(new_n18639), .Y(new_n18640));
  INVx1_ASAP7_75t_L         g18384(.A(new_n18329), .Y(new_n18641));
  INVx1_ASAP7_75t_L         g18385(.A(new_n18422), .Y(new_n18642));
  O2A1O1Ixp33_ASAP7_75t_L   g18386(.A1(new_n18176), .A2(new_n18178), .B(new_n18641), .C(new_n18642), .Y(new_n18643));
  A2O1A1O1Ixp25_ASAP7_75t_L g18387(.A1(new_n18325), .A2(\a[44] ), .B(new_n18326), .C(new_n18423), .D(new_n18643), .Y(new_n18644));
  XOR2x2_ASAP7_75t_L        g18388(.A(new_n18644), .B(new_n18640), .Y(new_n18645));
  NOR2xp33_ASAP7_75t_L      g18389(.A(new_n7249), .B(new_n5641), .Y(new_n18646));
  AOI221xp5_ASAP7_75t_L     g18390(.A1(\b[43] ), .A2(new_n5920), .B1(\b[44] ), .B2(new_n5623), .C(new_n18646), .Y(new_n18647));
  O2A1O1Ixp33_ASAP7_75t_L   g18391(.A1(new_n5630), .A2(new_n7255), .B(new_n18647), .C(new_n5626), .Y(new_n18648));
  O2A1O1Ixp33_ASAP7_75t_L   g18392(.A1(new_n5630), .A2(new_n7255), .B(new_n18647), .C(\a[41] ), .Y(new_n18649));
  INVx1_ASAP7_75t_L         g18393(.A(new_n18649), .Y(new_n18650));
  OAI21xp33_ASAP7_75t_L     g18394(.A1(new_n5626), .A2(new_n18648), .B(new_n18650), .Y(new_n18651));
  XOR2x2_ASAP7_75t_L        g18395(.A(new_n18651), .B(new_n18645), .Y(new_n18652));
  O2A1O1Ixp33_ASAP7_75t_L   g18396(.A1(new_n5626), .A2(new_n18315), .B(new_n18317), .C(new_n18425), .Y(new_n18653));
  O2A1O1Ixp33_ASAP7_75t_L   g18397(.A1(new_n18319), .A2(new_n18320), .B(new_n18424), .C(new_n18653), .Y(new_n18654));
  XOR2x2_ASAP7_75t_L        g18398(.A(new_n18654), .B(new_n18652), .Y(new_n18655));
  INVx1_ASAP7_75t_L         g18399(.A(new_n18655), .Y(new_n18656));
  NOR2xp33_ASAP7_75t_L      g18400(.A(new_n7860), .B(new_n4908), .Y(new_n18657));
  AOI221xp5_ASAP7_75t_L     g18401(.A1(\b[46] ), .A2(new_n5139), .B1(\b[47] ), .B2(new_n4916), .C(new_n18657), .Y(new_n18658));
  O2A1O1Ixp33_ASAP7_75t_L   g18402(.A1(new_n4911), .A2(new_n7868), .B(new_n18658), .C(new_n4906), .Y(new_n18659));
  O2A1O1Ixp33_ASAP7_75t_L   g18403(.A1(new_n4911), .A2(new_n7868), .B(new_n18658), .C(\a[38] ), .Y(new_n18660));
  INVx1_ASAP7_75t_L         g18404(.A(new_n18660), .Y(new_n18661));
  O2A1O1Ixp33_ASAP7_75t_L   g18405(.A1(new_n18659), .A2(new_n4906), .B(new_n18661), .C(new_n18656), .Y(new_n18662));
  O2A1O1Ixp33_ASAP7_75t_L   g18406(.A1(new_n18659), .A2(new_n4906), .B(new_n18661), .C(new_n18655), .Y(new_n18663));
  INVx1_ASAP7_75t_L         g18407(.A(new_n18663), .Y(new_n18664));
  O2A1O1Ixp33_ASAP7_75t_L   g18408(.A1(new_n18311), .A2(new_n18201), .B(new_n18426), .C(new_n18433), .Y(new_n18665));
  OAI211xp5_ASAP7_75t_L     g18409(.A1(new_n18656), .A2(new_n18662), .B(new_n18665), .C(new_n18664), .Y(new_n18666));
  INVx1_ASAP7_75t_L         g18410(.A(new_n18662), .Y(new_n18667));
  INVx1_ASAP7_75t_L         g18411(.A(new_n18665), .Y(new_n18668));
  A2O1A1Ixp33_ASAP7_75t_L   g18412(.A1(new_n18667), .A2(new_n18655), .B(new_n18663), .C(new_n18668), .Y(new_n18669));
  NAND2xp33_ASAP7_75t_L     g18413(.A(new_n18666), .B(new_n18669), .Y(new_n18670));
  NOR2xp33_ASAP7_75t_L      g18414(.A(new_n8779), .B(new_n4147), .Y(new_n18671));
  AOI221xp5_ASAP7_75t_L     g18415(.A1(\b[49] ), .A2(new_n4402), .B1(\b[50] ), .B2(new_n4155), .C(new_n18671), .Y(new_n18672));
  O2A1O1Ixp33_ASAP7_75t_L   g18416(.A1(new_n4150), .A2(new_n8789), .B(new_n18672), .C(new_n4145), .Y(new_n18673));
  INVx1_ASAP7_75t_L         g18417(.A(new_n18673), .Y(new_n18674));
  O2A1O1Ixp33_ASAP7_75t_L   g18418(.A1(new_n4150), .A2(new_n8789), .B(new_n18672), .C(\a[35] ), .Y(new_n18675));
  AOI21xp33_ASAP7_75t_L     g18419(.A1(new_n18674), .A2(\a[35] ), .B(new_n18675), .Y(new_n18676));
  NAND2xp33_ASAP7_75t_L     g18420(.A(new_n18676), .B(new_n18670), .Y(new_n18677));
  INVx1_ASAP7_75t_L         g18421(.A(new_n18670), .Y(new_n18678));
  O2A1O1Ixp33_ASAP7_75t_L   g18422(.A1(new_n18445), .A2(new_n4145), .B(new_n18447), .C(new_n18442), .Y(new_n18679));
  A2O1A1Ixp33_ASAP7_75t_L   g18423(.A1(new_n18440), .A2(new_n18439), .B(new_n18679), .C(new_n18677), .Y(new_n18680));
  A2O1A1O1Ixp25_ASAP7_75t_L g18424(.A1(new_n18674), .A2(\a[35] ), .B(new_n18675), .C(new_n18678), .D(new_n18680), .Y(new_n18681));
  O2A1O1Ixp33_ASAP7_75t_L   g18425(.A1(new_n18442), .A2(new_n18448), .B(new_n18441), .C(new_n18681), .Y(new_n18682));
  A2O1A1O1Ixp25_ASAP7_75t_L g18426(.A1(new_n18674), .A2(\a[35] ), .B(new_n18675), .C(new_n18678), .D(new_n18681), .Y(new_n18683));
  A2O1A1Ixp33_ASAP7_75t_L   g18427(.A1(new_n18683), .A2(new_n18677), .B(new_n18682), .C(new_n18530), .Y(new_n18684));
  AO221x2_ASAP7_75t_L       g18428(.A1(new_n18528), .A2(new_n18529), .B1(new_n18683), .B2(new_n18677), .C(new_n18682), .Y(new_n18685));
  NAND3xp33_ASAP7_75t_L     g18429(.A(new_n18523), .B(new_n18684), .C(new_n18685), .Y(new_n18686));
  AND3x1_ASAP7_75t_L        g18430(.A(new_n18686), .B(new_n18685), .C(new_n18684), .Y(new_n18687));
  A2O1A1Ixp33_ASAP7_75t_L   g18431(.A1(new_n18523), .A2(new_n18686), .B(new_n18687), .C(new_n18517), .Y(new_n18688));
  INVx1_ASAP7_75t_L         g18432(.A(new_n18688), .Y(new_n18689));
  AOI21xp33_ASAP7_75t_L     g18433(.A1(new_n18686), .A2(new_n18523), .B(new_n18687), .Y(new_n18690));
  OAI21xp33_ASAP7_75t_L     g18434(.A1(new_n18516), .A2(new_n18514), .B(new_n18690), .Y(new_n18691));
  INVx1_ASAP7_75t_L         g18435(.A(new_n18691), .Y(new_n18692));
  OAI21xp33_ASAP7_75t_L     g18436(.A1(new_n18689), .A2(new_n18692), .B(new_n18508), .Y(new_n18693));
  INVx1_ASAP7_75t_L         g18437(.A(new_n18503), .Y(new_n18694));
  A2O1A1O1Ixp25_ASAP7_75t_L g18438(.A1(new_n18296), .A2(new_n18499), .B(new_n18478), .C(new_n18299), .D(new_n18694), .Y(new_n18695));
  O2A1O1Ixp33_ASAP7_75t_L   g18439(.A1(new_n18695), .A2(new_n18506), .B(new_n18688), .C(new_n18692), .Y(new_n18696));
  NAND2xp33_ASAP7_75t_L     g18440(.A(new_n18688), .B(new_n18696), .Y(new_n18697));
  INVx1_ASAP7_75t_L         g18441(.A(new_n18281), .Y(new_n18698));
  A2O1A1Ixp33_ASAP7_75t_L   g18442(.A1(new_n12986), .A2(new_n1513), .B(new_n18280), .C(new_n1501), .Y(new_n18699));
  O2A1O1Ixp33_ASAP7_75t_L   g18443(.A1(new_n18698), .A2(new_n1501), .B(new_n18699), .C(new_n18485), .Y(new_n18700));
  O2A1O1Ixp33_ASAP7_75t_L   g18444(.A1(new_n18290), .A2(new_n18284), .B(new_n18482), .C(new_n18700), .Y(new_n18701));
  AND3x1_ASAP7_75t_L        g18445(.A(new_n18693), .B(new_n18701), .C(new_n18697), .Y(new_n18702));
  A2O1A1Ixp33_ASAP7_75t_L   g18446(.A1(new_n18505), .A2(new_n18694), .B(new_n18695), .C(new_n18691), .Y(new_n18703));
  A2O1A1O1Ixp25_ASAP7_75t_L g18447(.A1(new_n18686), .A2(new_n18523), .B(new_n18687), .C(new_n18517), .D(new_n18703), .Y(new_n18704));
  O2A1O1Ixp33_ASAP7_75t_L   g18448(.A1(new_n18507), .A2(new_n18704), .B(new_n18697), .C(new_n18701), .Y(new_n18705));
  NOR2xp33_ASAP7_75t_L      g18449(.A(new_n18705), .B(new_n18702), .Y(new_n18706));
  A2O1A1Ixp33_ASAP7_75t_L   g18450(.A1(new_n18496), .A2(new_n18493), .B(new_n18490), .C(new_n18706), .Y(new_n18707));
  INVx1_ASAP7_75t_L         g18451(.A(new_n18707), .Y(new_n18708));
  NOR3xp33_ASAP7_75t_L      g18452(.A(new_n18495), .B(new_n18706), .C(new_n18490), .Y(new_n18709));
  NOR2xp33_ASAP7_75t_L      g18453(.A(new_n18708), .B(new_n18709), .Y(\f[84] ));
  OAI21xp33_ASAP7_75t_L     g18454(.A1(new_n18514), .A2(new_n18690), .B(new_n18515), .Y(new_n18711));
  NOR2xp33_ASAP7_75t_L      g18455(.A(new_n12956), .B(new_n1962), .Y(new_n18712));
  AOI21xp33_ASAP7_75t_L     g18456(.A1(new_n2093), .A2(\b[62] ), .B(new_n18712), .Y(new_n18713));
  A2O1A1O1Ixp25_ASAP7_75t_L g18457(.A1(\b[62] ), .A2(new_n1949), .B(new_n1945), .C(new_n1954), .D(new_n18712), .Y(new_n18714));
  A2O1A1Ixp33_ASAP7_75t_L   g18458(.A1(new_n12993), .A2(new_n18713), .B(new_n18714), .C(\a[23] ), .Y(new_n18715));
  O2A1O1Ixp33_ASAP7_75t_L   g18459(.A1(new_n1956), .A2(new_n12993), .B(new_n18713), .C(\a[23] ), .Y(new_n18716));
  INVx1_ASAP7_75t_L         g18460(.A(new_n18716), .Y(new_n18717));
  AND2x2_ASAP7_75t_L        g18461(.A(new_n18715), .B(new_n18717), .Y(new_n18718));
  XOR2x2_ASAP7_75t_L        g18462(.A(new_n18718), .B(new_n18711), .Y(new_n18719));
  INVx1_ASAP7_75t_L         g18463(.A(new_n18519), .Y(new_n18720));
  NOR2xp33_ASAP7_75t_L      g18464(.A(new_n12258), .B(new_n2415), .Y(new_n18721));
  AOI221xp5_ASAP7_75t_L     g18465(.A1(\b[59] ), .A2(new_n2577), .B1(\b[60] ), .B2(new_n2421), .C(new_n18721), .Y(new_n18722));
  O2A1O1Ixp33_ASAP7_75t_L   g18466(.A1(new_n2425), .A2(new_n14764), .B(new_n18722), .C(new_n2413), .Y(new_n18723));
  NOR2xp33_ASAP7_75t_L      g18467(.A(new_n2413), .B(new_n18723), .Y(new_n18724));
  O2A1O1Ixp33_ASAP7_75t_L   g18468(.A1(new_n2425), .A2(new_n14764), .B(new_n18722), .C(\a[26] ), .Y(new_n18725));
  NOR2xp33_ASAP7_75t_L      g18469(.A(new_n18725), .B(new_n18724), .Y(new_n18726));
  OA211x2_ASAP7_75t_L       g18470(.A1(new_n18720), .A2(new_n18522), .B(new_n18686), .C(new_n18726), .Y(new_n18727));
  O2A1O1Ixp33_ASAP7_75t_L   g18471(.A1(new_n18720), .A2(new_n18522), .B(new_n18686), .C(new_n18726), .Y(new_n18728));
  A2O1A1Ixp33_ASAP7_75t_L   g18472(.A1(new_n18460), .A2(new_n18457), .B(new_n18526), .C(new_n18684), .Y(new_n18729));
  NAND2xp33_ASAP7_75t_L     g18473(.A(\b[57] ), .B(new_n2936), .Y(new_n18730));
  OAI221xp5_ASAP7_75t_L     g18474(.A1(new_n2930), .A2(new_n11303), .B1(new_n10332), .B2(new_n3133), .C(new_n18730), .Y(new_n18731));
  AOI21xp33_ASAP7_75t_L     g18475(.A1(new_n11314), .A2(new_n2932), .B(new_n18731), .Y(new_n18732));
  NAND2xp33_ASAP7_75t_L     g18476(.A(\a[29] ), .B(new_n18732), .Y(new_n18733));
  A2O1A1Ixp33_ASAP7_75t_L   g18477(.A1(new_n11314), .A2(new_n2932), .B(new_n18731), .C(new_n2928), .Y(new_n18734));
  NAND2xp33_ASAP7_75t_L     g18478(.A(new_n18734), .B(new_n18733), .Y(new_n18735));
  XOR2x2_ASAP7_75t_L        g18479(.A(new_n18735), .B(new_n18729), .Y(new_n18736));
  NOR2xp33_ASAP7_75t_L      g18480(.A(new_n10309), .B(new_n3510), .Y(new_n18737));
  AOI221xp5_ASAP7_75t_L     g18481(.A1(\b[53] ), .A2(new_n3708), .B1(\b[54] ), .B2(new_n3499), .C(new_n18737), .Y(new_n18738));
  O2A1O1Ixp33_ASAP7_75t_L   g18482(.A1(new_n3513), .A2(new_n15849), .B(new_n18738), .C(new_n3493), .Y(new_n18739));
  NOR2xp33_ASAP7_75t_L      g18483(.A(new_n3493), .B(new_n18739), .Y(new_n18740));
  O2A1O1Ixp33_ASAP7_75t_L   g18484(.A1(new_n3513), .A2(new_n15849), .B(new_n18738), .C(\a[32] ), .Y(new_n18741));
  NOR2xp33_ASAP7_75t_L      g18485(.A(new_n18741), .B(new_n18740), .Y(new_n18742));
  INVx1_ASAP7_75t_L         g18486(.A(new_n18742), .Y(new_n18743));
  O2A1O1Ixp33_ASAP7_75t_L   g18487(.A1(new_n18670), .A2(new_n18676), .B(new_n18680), .C(new_n18743), .Y(new_n18744));
  A2O1A1Ixp33_ASAP7_75t_L   g18488(.A1(\a[35] ), .A2(new_n18674), .B(new_n18675), .C(new_n18678), .Y(new_n18745));
  AND3x1_ASAP7_75t_L        g18489(.A(new_n18680), .B(new_n18743), .C(new_n18745), .Y(new_n18746));
  NAND2xp33_ASAP7_75t_L     g18490(.A(\a[47] ), .B(new_n18420), .Y(new_n18747));
  A2O1A1Ixp33_ASAP7_75t_L   g18491(.A1(new_n18747), .A2(new_n18335), .B(new_n18418), .C(new_n18415), .Y(new_n18748));
  INVx1_ASAP7_75t_L         g18492(.A(new_n18532), .Y(new_n18749));
  INVx1_ASAP7_75t_L         g18493(.A(new_n18610), .Y(new_n18750));
  NOR2xp33_ASAP7_75t_L      g18494(.A(new_n2703), .B(new_n11354), .Y(new_n18751));
  AOI221xp5_ASAP7_75t_L     g18495(.A1(\b[28] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[27] ), .C(new_n18751), .Y(new_n18752));
  O2A1O1Ixp33_ASAP7_75t_L   g18496(.A1(new_n11053), .A2(new_n3087), .B(new_n18752), .C(new_n11048), .Y(new_n18753));
  INVx1_ASAP7_75t_L         g18497(.A(new_n18753), .Y(new_n18754));
  O2A1O1Ixp33_ASAP7_75t_L   g18498(.A1(new_n11053), .A2(new_n3087), .B(new_n18752), .C(\a[59] ), .Y(new_n18755));
  NOR2xp33_ASAP7_75t_L      g18499(.A(new_n1895), .B(new_n13030), .Y(new_n18756));
  A2O1A1O1Ixp25_ASAP7_75t_L g18500(.A1(new_n13028), .A2(\b[20] ), .B(new_n18358), .C(new_n18537), .D(new_n18535), .Y(new_n18757));
  A2O1A1Ixp33_ASAP7_75t_L   g18501(.A1(new_n13028), .A2(\b[22] ), .B(new_n18756), .C(new_n18757), .Y(new_n18758));
  O2A1O1Ixp33_ASAP7_75t_L   g18502(.A1(new_n12669), .A2(new_n12671), .B(\b[22] ), .C(new_n18756), .Y(new_n18759));
  INVx1_ASAP7_75t_L         g18503(.A(new_n18759), .Y(new_n18760));
  O2A1O1Ixp33_ASAP7_75t_L   g18504(.A1(new_n18359), .A2(new_n18538), .B(new_n18534), .C(new_n18760), .Y(new_n18761));
  INVx1_ASAP7_75t_L         g18505(.A(new_n18761), .Y(new_n18762));
  NAND2xp33_ASAP7_75t_L     g18506(.A(new_n18758), .B(new_n18762), .Y(new_n18763));
  NOR2xp33_ASAP7_75t_L      g18507(.A(new_n2205), .B(new_n12318), .Y(new_n18764));
  AOI221xp5_ASAP7_75t_L     g18508(.A1(new_n11995), .A2(\b[25] ), .B1(new_n13314), .B2(\b[23] ), .C(new_n18764), .Y(new_n18765));
  INVx1_ASAP7_75t_L         g18509(.A(new_n18765), .Y(new_n18766));
  A2O1A1Ixp33_ASAP7_75t_L   g18510(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n18765), .Y(new_n18767));
  A2O1A1O1Ixp25_ASAP7_75t_L g18511(.A1(new_n2384), .A2(new_n2382), .B(new_n18766), .C(new_n18767), .D(new_n11987), .Y(new_n18768));
  O2A1O1Ixp33_ASAP7_75t_L   g18512(.A1(new_n11998), .A2(new_n2385), .B(new_n18765), .C(\a[62] ), .Y(new_n18769));
  NOR2xp33_ASAP7_75t_L      g18513(.A(new_n18768), .B(new_n18769), .Y(new_n18770));
  NOR2xp33_ASAP7_75t_L      g18514(.A(new_n18763), .B(new_n18770), .Y(new_n18771));
  AOI211xp5_ASAP7_75t_L     g18515(.A1(new_n18758), .A2(new_n18762), .B(new_n18768), .C(new_n18769), .Y(new_n18772));
  NOR2xp33_ASAP7_75t_L      g18516(.A(new_n18772), .B(new_n18771), .Y(new_n18773));
  INVx1_ASAP7_75t_L         g18517(.A(new_n18773), .Y(new_n18774));
  O2A1O1Ixp33_ASAP7_75t_L   g18518(.A1(new_n18552), .A2(new_n18558), .B(new_n18550), .C(new_n18774), .Y(new_n18775));
  INVx1_ASAP7_75t_L         g18519(.A(new_n18775), .Y(new_n18776));
  A2O1A1O1Ixp25_ASAP7_75t_L g18520(.A1(new_n18359), .A2(new_n18111), .B(new_n18370), .C(new_n18553), .D(new_n18549), .Y(new_n18777));
  NAND2xp33_ASAP7_75t_L     g18521(.A(new_n18774), .B(new_n18777), .Y(new_n18778));
  AND2x2_ASAP7_75t_L        g18522(.A(new_n18776), .B(new_n18778), .Y(new_n18779));
  A2O1A1Ixp33_ASAP7_75t_L   g18523(.A1(new_n18754), .A2(\a[59] ), .B(new_n18755), .C(new_n18779), .Y(new_n18780));
  NOR2xp33_ASAP7_75t_L      g18524(.A(new_n11048), .B(new_n18753), .Y(new_n18781));
  OR3x1_ASAP7_75t_L         g18525(.A(new_n18779), .B(new_n18781), .C(new_n18755), .Y(new_n18782));
  AND2x2_ASAP7_75t_L        g18526(.A(new_n18780), .B(new_n18782), .Y(new_n18783));
  INVx1_ASAP7_75t_L         g18527(.A(new_n18783), .Y(new_n18784));
  O2A1O1Ixp33_ASAP7_75t_L   g18528(.A1(new_n18569), .A2(new_n18571), .B(new_n18566), .C(new_n18784), .Y(new_n18785));
  INVx1_ASAP7_75t_L         g18529(.A(new_n18785), .Y(new_n18786));
  A2O1A1O1Ixp25_ASAP7_75t_L g18530(.A1(new_n18564), .A2(\a[59] ), .B(new_n18565), .C(new_n18560), .D(new_n18574), .Y(new_n18787));
  NAND2xp33_ASAP7_75t_L     g18531(.A(new_n18787), .B(new_n18784), .Y(new_n18788));
  NAND2xp33_ASAP7_75t_L     g18532(.A(new_n18788), .B(new_n18786), .Y(new_n18789));
  NOR2xp33_ASAP7_75t_L      g18533(.A(new_n3456), .B(new_n10388), .Y(new_n18790));
  AOI221xp5_ASAP7_75t_L     g18534(.A1(new_n10086), .A2(\b[31] ), .B1(new_n11361), .B2(\b[29] ), .C(new_n18790), .Y(new_n18791));
  O2A1O1Ixp33_ASAP7_75t_L   g18535(.A1(new_n10088), .A2(new_n3681), .B(new_n18791), .C(new_n10083), .Y(new_n18792));
  O2A1O1Ixp33_ASAP7_75t_L   g18536(.A1(new_n10088), .A2(new_n3681), .B(new_n18791), .C(\a[56] ), .Y(new_n18793));
  INVx1_ASAP7_75t_L         g18537(.A(new_n18793), .Y(new_n18794));
  O2A1O1Ixp33_ASAP7_75t_L   g18538(.A1(new_n18792), .A2(new_n10083), .B(new_n18794), .C(new_n18789), .Y(new_n18795));
  INVx1_ASAP7_75t_L         g18539(.A(new_n18789), .Y(new_n18796));
  O2A1O1Ixp33_ASAP7_75t_L   g18540(.A1(new_n18792), .A2(new_n10083), .B(new_n18794), .C(new_n18796), .Y(new_n18797));
  INVx1_ASAP7_75t_L         g18541(.A(new_n18797), .Y(new_n18798));
  O2A1O1Ixp33_ASAP7_75t_L   g18542(.A1(new_n18577), .A2(new_n18585), .B(new_n18590), .C(new_n18583), .Y(new_n18799));
  OAI211xp5_ASAP7_75t_L     g18543(.A1(new_n18789), .A2(new_n18795), .B(new_n18798), .C(new_n18799), .Y(new_n18800));
  INVx1_ASAP7_75t_L         g18544(.A(new_n18795), .Y(new_n18801));
  INVx1_ASAP7_75t_L         g18545(.A(new_n18799), .Y(new_n18802));
  A2O1A1Ixp33_ASAP7_75t_L   g18546(.A1(new_n18801), .A2(new_n18796), .B(new_n18797), .C(new_n18802), .Y(new_n18803));
  NAND2xp33_ASAP7_75t_L     g18547(.A(new_n18803), .B(new_n18800), .Y(new_n18804));
  NOR2xp33_ASAP7_75t_L      g18548(.A(new_n4101), .B(new_n10400), .Y(new_n18805));
  AOI221xp5_ASAP7_75t_L     g18549(.A1(new_n9102), .A2(\b[34] ), .B1(new_n10398), .B2(\b[32] ), .C(new_n18805), .Y(new_n18806));
  O2A1O1Ixp33_ASAP7_75t_L   g18550(.A1(new_n9104), .A2(new_n4352), .B(new_n18806), .C(new_n9099), .Y(new_n18807));
  O2A1O1Ixp33_ASAP7_75t_L   g18551(.A1(new_n9104), .A2(new_n4352), .B(new_n18806), .C(\a[53] ), .Y(new_n18808));
  INVx1_ASAP7_75t_L         g18552(.A(new_n18808), .Y(new_n18809));
  O2A1O1Ixp33_ASAP7_75t_L   g18553(.A1(new_n18807), .A2(new_n9099), .B(new_n18809), .C(new_n18804), .Y(new_n18810));
  INVx1_ASAP7_75t_L         g18554(.A(new_n18807), .Y(new_n18811));
  A2O1A1Ixp33_ASAP7_75t_L   g18555(.A1(\a[53] ), .A2(new_n18811), .B(new_n18808), .C(new_n18804), .Y(new_n18812));
  OA21x2_ASAP7_75t_L        g18556(.A1(new_n18804), .A2(new_n18810), .B(new_n18812), .Y(new_n18813));
  O2A1O1Ixp33_ASAP7_75t_L   g18557(.A1(new_n18400), .A2(new_n18404), .B(new_n18391), .C(new_n18600), .Y(new_n18814));
  INVx1_ASAP7_75t_L         g18558(.A(new_n18603), .Y(new_n18815));
  AOI21xp33_ASAP7_75t_L     g18559(.A1(new_n18815), .A2(new_n18594), .B(new_n18814), .Y(new_n18816));
  NAND2xp33_ASAP7_75t_L     g18560(.A(new_n18816), .B(new_n18813), .Y(new_n18817));
  O2A1O1Ixp33_ASAP7_75t_L   g18561(.A1(new_n18804), .A2(new_n18810), .B(new_n18812), .C(new_n18816), .Y(new_n18818));
  INVx1_ASAP7_75t_L         g18562(.A(new_n18818), .Y(new_n18819));
  NOR2xp33_ASAP7_75t_L      g18563(.A(new_n4613), .B(new_n10065), .Y(new_n18820));
  AOI221xp5_ASAP7_75t_L     g18564(.A1(new_n8175), .A2(\b[37] ), .B1(new_n8484), .B2(\b[35] ), .C(new_n18820), .Y(new_n18821));
  O2A1O1Ixp33_ASAP7_75t_L   g18565(.A1(new_n8176), .A2(new_n5083), .B(new_n18821), .C(new_n8172), .Y(new_n18822));
  O2A1O1Ixp33_ASAP7_75t_L   g18566(.A1(new_n8176), .A2(new_n5083), .B(new_n18821), .C(\a[50] ), .Y(new_n18823));
  INVx1_ASAP7_75t_L         g18567(.A(new_n18823), .Y(new_n18824));
  OAI21xp33_ASAP7_75t_L     g18568(.A1(new_n8172), .A2(new_n18822), .B(new_n18824), .Y(new_n18825));
  AOI21xp33_ASAP7_75t_L     g18569(.A1(new_n18817), .A2(new_n18819), .B(new_n18825), .Y(new_n18826));
  NAND2xp33_ASAP7_75t_L     g18570(.A(new_n18819), .B(new_n18817), .Y(new_n18827));
  O2A1O1Ixp33_ASAP7_75t_L   g18571(.A1(new_n18822), .A2(new_n8172), .B(new_n18824), .C(new_n18827), .Y(new_n18828));
  NOR2xp33_ASAP7_75t_L      g18572(.A(new_n18826), .B(new_n18828), .Y(new_n18829));
  A2O1A1Ixp33_ASAP7_75t_L   g18573(.A1(new_n18749), .A2(new_n18612), .B(new_n18750), .C(new_n18829), .Y(new_n18830));
  INVx1_ASAP7_75t_L         g18574(.A(new_n18830), .Y(new_n18831));
  NAND2xp33_ASAP7_75t_L     g18575(.A(\b[39] ), .B(new_n7333), .Y(new_n18832));
  OAI221xp5_ASAP7_75t_L     g18576(.A1(new_n7318), .A2(new_n5855), .B1(new_n5311), .B2(new_n7614), .C(new_n18832), .Y(new_n18833));
  A2O1A1Ixp33_ASAP7_75t_L   g18577(.A1(new_n6651), .A2(new_n7322), .B(new_n18833), .C(\a[47] ), .Y(new_n18834));
  AOI211xp5_ASAP7_75t_L     g18578(.A1(new_n6651), .A2(new_n7322), .B(new_n18833), .C(new_n7316), .Y(new_n18835));
  A2O1A1O1Ixp25_ASAP7_75t_L g18579(.A1(new_n7322), .A2(new_n6651), .B(new_n18833), .C(new_n18834), .D(new_n18835), .Y(new_n18836));
  INVx1_ASAP7_75t_L         g18580(.A(new_n18829), .Y(new_n18837));
  A2O1A1Ixp33_ASAP7_75t_L   g18581(.A1(new_n18612), .A2(new_n18749), .B(new_n18750), .C(new_n18837), .Y(new_n18838));
  O2A1O1Ixp33_ASAP7_75t_L   g18582(.A1(new_n18837), .A2(new_n18831), .B(new_n18838), .C(new_n18836), .Y(new_n18839));
  NAND2xp33_ASAP7_75t_L     g18583(.A(new_n18829), .B(new_n18830), .Y(new_n18840));
  AND2x2_ASAP7_75t_L        g18584(.A(new_n18836), .B(new_n18840), .Y(new_n18841));
  A2O1A1O1Ixp25_ASAP7_75t_L g18585(.A1(new_n18616), .A2(new_n18610), .B(new_n18831), .C(new_n18841), .D(new_n18839), .Y(new_n18842));
  A2O1A1Ixp33_ASAP7_75t_L   g18586(.A1(new_n18629), .A2(new_n18748), .B(new_n18623), .C(new_n18842), .Y(new_n18843));
  O2A1O1Ixp33_ASAP7_75t_L   g18587(.A1(new_n18419), .A2(new_n18626), .B(new_n18629), .C(new_n18623), .Y(new_n18844));
  A2O1A1Ixp33_ASAP7_75t_L   g18588(.A1(new_n18841), .A2(new_n18838), .B(new_n18839), .C(new_n18844), .Y(new_n18845));
  NAND2xp33_ASAP7_75t_L     g18589(.A(new_n18845), .B(new_n18843), .Y(new_n18846));
  NOR2xp33_ASAP7_75t_L      g18590(.A(new_n6378), .B(new_n7304), .Y(new_n18847));
  AOI221xp5_ASAP7_75t_L     g18591(.A1(\b[41] ), .A2(new_n6742), .B1(\b[43] ), .B2(new_n6442), .C(new_n18847), .Y(new_n18848));
  O2A1O1Ixp33_ASAP7_75t_L   g18592(.A1(new_n6443), .A2(new_n6679), .B(new_n18848), .C(new_n6439), .Y(new_n18849));
  O2A1O1Ixp33_ASAP7_75t_L   g18593(.A1(new_n6443), .A2(new_n6679), .B(new_n18848), .C(\a[44] ), .Y(new_n18850));
  INVx1_ASAP7_75t_L         g18594(.A(new_n18850), .Y(new_n18851));
  O2A1O1Ixp33_ASAP7_75t_L   g18595(.A1(new_n18849), .A2(new_n6439), .B(new_n18851), .C(new_n18846), .Y(new_n18852));
  INVx1_ASAP7_75t_L         g18596(.A(new_n18849), .Y(new_n18853));
  A2O1A1Ixp33_ASAP7_75t_L   g18597(.A1(\a[44] ), .A2(new_n18853), .B(new_n18850), .C(new_n18846), .Y(new_n18854));
  O2A1O1Ixp33_ASAP7_75t_L   g18598(.A1(new_n6439), .A2(new_n18634), .B(new_n18636), .C(new_n18637), .Y(new_n18855));
  O2A1O1Ixp33_ASAP7_75t_L   g18599(.A1(new_n17928), .A2(new_n17925), .B(new_n18177), .C(new_n18176), .Y(new_n18856));
  INVx1_ASAP7_75t_L         g18600(.A(new_n18856), .Y(new_n18857));
  A2O1A1Ixp33_ASAP7_75t_L   g18601(.A1(new_n18325), .A2(\a[44] ), .B(new_n18326), .C(new_n18423), .Y(new_n18858));
  A2O1A1Ixp33_ASAP7_75t_L   g18602(.A1(new_n18641), .A2(new_n18857), .B(new_n18642), .C(new_n18858), .Y(new_n18859));
  A2O1A1O1Ixp25_ASAP7_75t_L g18603(.A1(new_n18628), .A2(new_n18630), .B(new_n18855), .C(new_n18859), .D(new_n18637), .Y(new_n18860));
  OAI211xp5_ASAP7_75t_L     g18604(.A1(new_n18846), .A2(new_n18852), .B(new_n18860), .C(new_n18854), .Y(new_n18861));
  OAI21xp33_ASAP7_75t_L     g18605(.A1(new_n18846), .A2(new_n18852), .B(new_n18854), .Y(new_n18862));
  A2O1A1Ixp33_ASAP7_75t_L   g18606(.A1(new_n18640), .A2(new_n18859), .B(new_n18637), .C(new_n18862), .Y(new_n18863));
  NAND2xp33_ASAP7_75t_L     g18607(.A(new_n18863), .B(new_n18861), .Y(new_n18864));
  NOR2xp33_ASAP7_75t_L      g18608(.A(new_n7249), .B(new_n5640), .Y(new_n18865));
  AOI221xp5_ASAP7_75t_L     g18609(.A1(\b[44] ), .A2(new_n5920), .B1(\b[46] ), .B2(new_n5629), .C(new_n18865), .Y(new_n18866));
  O2A1O1Ixp33_ASAP7_75t_L   g18610(.A1(new_n5630), .A2(new_n7279), .B(new_n18866), .C(new_n5626), .Y(new_n18867));
  O2A1O1Ixp33_ASAP7_75t_L   g18611(.A1(new_n5630), .A2(new_n7279), .B(new_n18866), .C(\a[41] ), .Y(new_n18868));
  INVx1_ASAP7_75t_L         g18612(.A(new_n18868), .Y(new_n18869));
  O2A1O1Ixp33_ASAP7_75t_L   g18613(.A1(new_n18867), .A2(new_n5626), .B(new_n18869), .C(new_n18864), .Y(new_n18870));
  INVx1_ASAP7_75t_L         g18614(.A(new_n18867), .Y(new_n18871));
  A2O1A1Ixp33_ASAP7_75t_L   g18615(.A1(\a[41] ), .A2(new_n18871), .B(new_n18868), .C(new_n18864), .Y(new_n18872));
  OAI21xp33_ASAP7_75t_L     g18616(.A1(new_n18864), .A2(new_n18870), .B(new_n18872), .Y(new_n18873));
  O2A1O1Ixp33_ASAP7_75t_L   g18617(.A1(new_n18648), .A2(new_n5626), .B(new_n18650), .C(new_n18645), .Y(new_n18874));
  INVx1_ASAP7_75t_L         g18618(.A(new_n18648), .Y(new_n18875));
  A2O1A1Ixp33_ASAP7_75t_L   g18619(.A1(\a[41] ), .A2(new_n18875), .B(new_n18649), .C(new_n18645), .Y(new_n18876));
  O2A1O1Ixp33_ASAP7_75t_L   g18620(.A1(new_n18645), .A2(new_n18874), .B(new_n18876), .C(new_n18654), .Y(new_n18877));
  NOR2xp33_ASAP7_75t_L      g18621(.A(new_n18874), .B(new_n18877), .Y(new_n18878));
  XOR2x2_ASAP7_75t_L        g18622(.A(new_n18878), .B(new_n18873), .Y(new_n18879));
  NOR2xp33_ASAP7_75t_L      g18623(.A(new_n8427), .B(new_n4908), .Y(new_n18880));
  AOI221xp5_ASAP7_75t_L     g18624(.A1(\b[47] ), .A2(new_n5139), .B1(\b[48] ), .B2(new_n4916), .C(new_n18880), .Y(new_n18881));
  O2A1O1Ixp33_ASAP7_75t_L   g18625(.A1(new_n4911), .A2(new_n14802), .B(new_n18881), .C(new_n4906), .Y(new_n18882));
  O2A1O1Ixp33_ASAP7_75t_L   g18626(.A1(new_n4911), .A2(new_n14802), .B(new_n18881), .C(\a[38] ), .Y(new_n18883));
  INVx1_ASAP7_75t_L         g18627(.A(new_n18883), .Y(new_n18884));
  OAI21xp33_ASAP7_75t_L     g18628(.A1(new_n4906), .A2(new_n18882), .B(new_n18884), .Y(new_n18885));
  OR2x4_ASAP7_75t_L         g18629(.A(new_n18885), .B(new_n18879), .Y(new_n18886));
  INVx1_ASAP7_75t_L         g18630(.A(new_n18882), .Y(new_n18887));
  A2O1A1Ixp33_ASAP7_75t_L   g18631(.A1(\a[38] ), .A2(new_n18887), .B(new_n18883), .C(new_n18879), .Y(new_n18888));
  O2A1O1Ixp33_ASAP7_75t_L   g18632(.A1(new_n18655), .A2(new_n18663), .B(new_n18668), .C(new_n18662), .Y(new_n18889));
  AND3x1_ASAP7_75t_L        g18633(.A(new_n18886), .B(new_n18889), .C(new_n18888), .Y(new_n18890));
  O2A1O1Ixp33_ASAP7_75t_L   g18634(.A1(new_n18882), .A2(new_n4906), .B(new_n18884), .C(new_n18879), .Y(new_n18891));
  O2A1O1Ixp33_ASAP7_75t_L   g18635(.A1(new_n18879), .A2(new_n18891), .B(new_n18888), .C(new_n18889), .Y(new_n18892));
  NOR2xp33_ASAP7_75t_L      g18636(.A(new_n18892), .B(new_n18890), .Y(new_n18893));
  NOR2xp33_ASAP7_75t_L      g18637(.A(new_n8779), .B(new_n4142), .Y(new_n18894));
  AOI221xp5_ASAP7_75t_L     g18638(.A1(\b[50] ), .A2(new_n4402), .B1(\b[52] ), .B2(new_n4156), .C(new_n18894), .Y(new_n18895));
  INVx1_ASAP7_75t_L         g18639(.A(new_n18895), .Y(new_n18896));
  A2O1A1Ixp33_ASAP7_75t_L   g18640(.A1(new_n9367), .A2(new_n4151), .B(new_n18896), .C(\a[35] ), .Y(new_n18897));
  O2A1O1Ixp33_ASAP7_75t_L   g18641(.A1(new_n4150), .A2(new_n17363), .B(new_n18895), .C(\a[35] ), .Y(new_n18898));
  A2O1A1Ixp33_ASAP7_75t_L   g18642(.A1(\a[35] ), .A2(new_n18897), .B(new_n18898), .C(new_n18893), .Y(new_n18899));
  NAND2xp33_ASAP7_75t_L     g18643(.A(new_n18893), .B(new_n18899), .Y(new_n18900));
  A2O1A1Ixp33_ASAP7_75t_L   g18644(.A1(new_n18897), .A2(\a[35] ), .B(new_n18898), .C(new_n18899), .Y(new_n18901));
  NAND2xp33_ASAP7_75t_L     g18645(.A(new_n18900), .B(new_n18901), .Y(new_n18902));
  OAI21xp33_ASAP7_75t_L     g18646(.A1(new_n18744), .A2(new_n18746), .B(new_n18902), .Y(new_n18903));
  OR3x1_ASAP7_75t_L         g18647(.A(new_n18902), .B(new_n18744), .C(new_n18746), .Y(new_n18904));
  NAND3xp33_ASAP7_75t_L     g18648(.A(new_n18736), .B(new_n18903), .C(new_n18904), .Y(new_n18905));
  NAND2xp33_ASAP7_75t_L     g18649(.A(new_n18736), .B(new_n18905), .Y(new_n18906));
  INVx1_ASAP7_75t_L         g18650(.A(new_n18736), .Y(new_n18907));
  NAND3xp33_ASAP7_75t_L     g18651(.A(new_n18907), .B(new_n18903), .C(new_n18904), .Y(new_n18908));
  AND2x2_ASAP7_75t_L        g18652(.A(new_n18908), .B(new_n18906), .Y(new_n18909));
  OR3x1_ASAP7_75t_L         g18653(.A(new_n18909), .B(new_n18727), .C(new_n18728), .Y(new_n18910));
  OAI21xp33_ASAP7_75t_L     g18654(.A1(new_n18728), .A2(new_n18727), .B(new_n18909), .Y(new_n18911));
  AO21x2_ASAP7_75t_L        g18655(.A1(new_n18911), .A2(new_n18910), .B(new_n18719), .Y(new_n18912));
  NAND3xp33_ASAP7_75t_L     g18656(.A(new_n18910), .B(new_n18719), .C(new_n18911), .Y(new_n18913));
  O2A1O1Ixp33_ASAP7_75t_L   g18657(.A1(new_n18298), .A2(new_n18500), .B(new_n18694), .C(new_n18704), .Y(new_n18914));
  NAND3xp33_ASAP7_75t_L     g18658(.A(new_n18912), .B(new_n18914), .C(new_n18913), .Y(new_n18915));
  O2A1O1Ixp33_ASAP7_75t_L   g18659(.A1(new_n18257), .A2(new_n18246), .B(new_n18297), .C(new_n18500), .Y(new_n18916));
  INVx1_ASAP7_75t_L         g18660(.A(new_n18916), .Y(new_n18917));
  O2A1O1Ixp33_ASAP7_75t_L   g18661(.A1(new_n18727), .A2(new_n18728), .B(new_n18909), .C(new_n18719), .Y(new_n18918));
  A2O1A1Ixp33_ASAP7_75t_L   g18662(.A1(new_n18918), .A2(new_n18910), .B(new_n18719), .C(new_n18913), .Y(new_n18919));
  A2O1A1Ixp33_ASAP7_75t_L   g18663(.A1(new_n18694), .A2(new_n18917), .B(new_n18704), .C(new_n18919), .Y(new_n18920));
  NAND2xp33_ASAP7_75t_L     g18664(.A(new_n18915), .B(new_n18920), .Y(new_n18921));
  A2O1A1O1Ixp25_ASAP7_75t_L g18665(.A1(new_n18697), .A2(new_n18693), .B(new_n18701), .C(new_n18707), .D(new_n18921), .Y(new_n18922));
  A2O1A1Ixp33_ASAP7_75t_L   g18666(.A1(new_n18697), .A2(new_n18693), .B(new_n18701), .C(new_n18707), .Y(new_n18923));
  AOI21xp33_ASAP7_75t_L     g18667(.A1(new_n18920), .A2(new_n18915), .B(new_n18923), .Y(new_n18924));
  NOR2xp33_ASAP7_75t_L      g18668(.A(new_n18922), .B(new_n18924), .Y(\f[85] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18669(.A1(new_n18514), .A2(new_n18690), .B(new_n18515), .C(new_n18718), .Y(new_n18926));
  AOI21xp33_ASAP7_75t_L     g18670(.A1(new_n18918), .A2(new_n18910), .B(new_n18926), .Y(new_n18927));
  NOR2xp33_ASAP7_75t_L      g18671(.A(new_n12956), .B(new_n2089), .Y(new_n18928));
  A2O1A1Ixp33_ASAP7_75t_L   g18672(.A1(new_n12986), .A2(new_n1964), .B(new_n18928), .C(\a[23] ), .Y(new_n18929));
  A2O1A1O1Ixp25_ASAP7_75t_L g18673(.A1(new_n1964), .A2(new_n14172), .B(new_n2093), .C(\b[63] ), .D(new_n1952), .Y(new_n18930));
  A2O1A1O1Ixp25_ASAP7_75t_L g18674(.A1(new_n12986), .A2(new_n1964), .B(new_n18928), .C(new_n18929), .D(new_n18930), .Y(new_n18931));
  INVx1_ASAP7_75t_L         g18675(.A(new_n18728), .Y(new_n18932));
  A2O1A1O1Ixp25_ASAP7_75t_L g18676(.A1(new_n18908), .A2(new_n18906), .B(new_n18727), .C(new_n18932), .D(new_n18931), .Y(new_n18933));
  INVx1_ASAP7_75t_L         g18677(.A(new_n18931), .Y(new_n18934));
  A2O1A1O1Ixp25_ASAP7_75t_L g18678(.A1(new_n18908), .A2(new_n18906), .B(new_n18727), .C(new_n18932), .D(new_n18934), .Y(new_n18935));
  INVx1_ASAP7_75t_L         g18679(.A(new_n18935), .Y(new_n18936));
  NAND2xp33_ASAP7_75t_L     g18680(.A(new_n18735), .B(new_n18729), .Y(new_n18937));
  NAND2xp33_ASAP7_75t_L     g18681(.A(\b[61] ), .B(new_n2421), .Y(new_n18938));
  OAI221xp5_ASAP7_75t_L     g18682(.A1(new_n2415), .A2(new_n12603), .B1(new_n11626), .B2(new_n2572), .C(new_n18938), .Y(new_n18939));
  A2O1A1Ixp33_ASAP7_75t_L   g18683(.A1(new_n13559), .A2(new_n2417), .B(new_n18939), .C(\a[26] ), .Y(new_n18940));
  NAND2xp33_ASAP7_75t_L     g18684(.A(\a[26] ), .B(new_n18940), .Y(new_n18941));
  A2O1A1Ixp33_ASAP7_75t_L   g18685(.A1(new_n13559), .A2(new_n2417), .B(new_n18939), .C(new_n2413), .Y(new_n18942));
  NAND4xp25_ASAP7_75t_L     g18686(.A(new_n18905), .B(new_n18941), .C(new_n18942), .D(new_n18937), .Y(new_n18943));
  INVx1_ASAP7_75t_L         g18687(.A(new_n18905), .Y(new_n18944));
  NAND2xp33_ASAP7_75t_L     g18688(.A(new_n18942), .B(new_n18941), .Y(new_n18945));
  A2O1A1Ixp33_ASAP7_75t_L   g18689(.A1(new_n18735), .A2(new_n18729), .B(new_n18944), .C(new_n18945), .Y(new_n18946));
  NAND2xp33_ASAP7_75t_L     g18690(.A(new_n18943), .B(new_n18946), .Y(new_n18947));
  NOR2xp33_ASAP7_75t_L      g18691(.A(new_n11303), .B(new_n2925), .Y(new_n18948));
  AOI221xp5_ASAP7_75t_L     g18692(.A1(\b[57] ), .A2(new_n3129), .B1(\b[59] ), .B2(new_n2938), .C(new_n18948), .Y(new_n18949));
  O2A1O1Ixp33_ASAP7_75t_L   g18693(.A1(new_n2940), .A2(new_n11597), .B(new_n18949), .C(new_n2928), .Y(new_n18950));
  O2A1O1Ixp33_ASAP7_75t_L   g18694(.A1(new_n2940), .A2(new_n11597), .B(new_n18949), .C(\a[29] ), .Y(new_n18951));
  INVx1_ASAP7_75t_L         g18695(.A(new_n18951), .Y(new_n18952));
  OAI21xp33_ASAP7_75t_L     g18696(.A1(new_n2928), .A2(new_n18950), .B(new_n18952), .Y(new_n18953));
  O2A1O1Ixp33_ASAP7_75t_L   g18697(.A1(new_n18670), .A2(new_n18676), .B(new_n18680), .C(new_n18742), .Y(new_n18954));
  O2A1O1Ixp33_ASAP7_75t_L   g18698(.A1(new_n18744), .A2(new_n18746), .B(new_n18902), .C(new_n18954), .Y(new_n18955));
  O2A1O1Ixp33_ASAP7_75t_L   g18699(.A1(new_n2928), .A2(new_n18950), .B(new_n18952), .C(new_n18955), .Y(new_n18956));
  INVx1_ASAP7_75t_L         g18700(.A(new_n18956), .Y(new_n18957));
  O2A1O1Ixp33_ASAP7_75t_L   g18701(.A1(new_n18683), .A2(new_n18742), .B(new_n18903), .C(new_n18953), .Y(new_n18958));
  NOR2xp33_ASAP7_75t_L      g18702(.A(new_n10332), .B(new_n3510), .Y(new_n18959));
  AOI221xp5_ASAP7_75t_L     g18703(.A1(\b[54] ), .A2(new_n3708), .B1(\b[55] ), .B2(new_n3499), .C(new_n18959), .Y(new_n18960));
  O2A1O1Ixp33_ASAP7_75t_L   g18704(.A1(new_n3513), .A2(new_n10339), .B(new_n18960), .C(new_n3493), .Y(new_n18961));
  O2A1O1Ixp33_ASAP7_75t_L   g18705(.A1(new_n3513), .A2(new_n10339), .B(new_n18960), .C(\a[32] ), .Y(new_n18962));
  INVx1_ASAP7_75t_L         g18706(.A(new_n18962), .Y(new_n18963));
  A2O1A1O1Ixp25_ASAP7_75t_L g18707(.A1(new_n18897), .A2(\a[35] ), .B(new_n18898), .C(new_n18893), .D(new_n18892), .Y(new_n18964));
  OAI211xp5_ASAP7_75t_L     g18708(.A1(new_n3493), .A2(new_n18961), .B(new_n18964), .C(new_n18963), .Y(new_n18965));
  O2A1O1Ixp33_ASAP7_75t_L   g18709(.A1(new_n3493), .A2(new_n18961), .B(new_n18963), .C(new_n18964), .Y(new_n18966));
  INVx1_ASAP7_75t_L         g18710(.A(new_n18966), .Y(new_n18967));
  NAND2xp33_ASAP7_75t_L     g18711(.A(new_n18965), .B(new_n18967), .Y(new_n18968));
  INVx1_ASAP7_75t_L         g18712(.A(new_n18968), .Y(new_n18969));
  INVx1_ASAP7_75t_L         g18713(.A(new_n18878), .Y(new_n18970));
  NAND2xp33_ASAP7_75t_L     g18714(.A(\a[44] ), .B(new_n18853), .Y(new_n18971));
  A2O1A1Ixp33_ASAP7_75t_L   g18715(.A1(new_n18971), .A2(new_n18851), .B(new_n18846), .C(new_n18843), .Y(new_n18972));
  NOR2xp33_ASAP7_75t_L      g18716(.A(new_n6378), .B(new_n6741), .Y(new_n18973));
  AOI221xp5_ASAP7_75t_L     g18717(.A1(\b[44] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[43] ), .C(new_n18973), .Y(new_n18974));
  O2A1O1Ixp33_ASAP7_75t_L   g18718(.A1(new_n6443), .A2(new_n6951), .B(new_n18974), .C(new_n6439), .Y(new_n18975));
  INVx1_ASAP7_75t_L         g18719(.A(new_n18975), .Y(new_n18976));
  O2A1O1Ixp33_ASAP7_75t_L   g18720(.A1(new_n6443), .A2(new_n6951), .B(new_n18974), .C(\a[44] ), .Y(new_n18977));
  AOI21xp33_ASAP7_75t_L     g18721(.A1(new_n18976), .A2(\a[44] ), .B(new_n18977), .Y(new_n18978));
  O2A1O1Ixp33_ASAP7_75t_L   g18722(.A1(new_n18750), .A2(new_n18615), .B(new_n18829), .C(new_n18839), .Y(new_n18979));
  A2O1A1O1Ixp25_ASAP7_75t_L g18723(.A1(new_n18801), .A2(new_n18796), .B(new_n18797), .C(new_n18802), .D(new_n18810), .Y(new_n18980));
  NOR2xp33_ASAP7_75t_L      g18724(.A(new_n4344), .B(new_n10400), .Y(new_n18981));
  AOI221xp5_ASAP7_75t_L     g18725(.A1(new_n9102), .A2(\b[35] ), .B1(new_n10398), .B2(\b[33] ), .C(new_n18981), .Y(new_n18982));
  INVx1_ASAP7_75t_L         g18726(.A(new_n18982), .Y(new_n18983));
  A2O1A1Ixp33_ASAP7_75t_L   g18727(.A1(new_n7773), .A2(new_n9437), .B(new_n18983), .C(\a[53] ), .Y(new_n18984));
  O2A1O1Ixp33_ASAP7_75t_L   g18728(.A1(new_n9104), .A2(new_n4589), .B(new_n18982), .C(\a[53] ), .Y(new_n18985));
  AO21x2_ASAP7_75t_L        g18729(.A1(\a[53] ), .A2(new_n18984), .B(new_n18985), .Y(new_n18986));
  INVx1_ASAP7_75t_L         g18730(.A(new_n18787), .Y(new_n18987));
  INVx1_ASAP7_75t_L         g18731(.A(new_n18771), .Y(new_n18988));
  NOR2xp33_ASAP7_75t_L      g18732(.A(new_n2045), .B(new_n13030), .Y(new_n18989));
  O2A1O1Ixp33_ASAP7_75t_L   g18733(.A1(new_n12669), .A2(new_n12671), .B(\b[23] ), .C(new_n18989), .Y(new_n18990));
  A2O1A1Ixp33_ASAP7_75t_L   g18734(.A1(new_n13028), .A2(\b[22] ), .B(new_n18756), .C(new_n18990), .Y(new_n18991));
  A2O1A1Ixp33_ASAP7_75t_L   g18735(.A1(\b[23] ), .A2(new_n13028), .B(new_n18989), .C(new_n18759), .Y(new_n18992));
  NAND2xp33_ASAP7_75t_L     g18736(.A(new_n18992), .B(new_n18991), .Y(new_n18993));
  NOR2xp33_ASAP7_75t_L      g18737(.A(new_n2377), .B(new_n12318), .Y(new_n18994));
  AOI221xp5_ASAP7_75t_L     g18738(.A1(new_n11995), .A2(\b[26] ), .B1(new_n13314), .B2(\b[24] ), .C(new_n18994), .Y(new_n18995));
  INVx1_ASAP7_75t_L         g18739(.A(new_n18995), .Y(new_n18996));
  A2O1A1Ixp33_ASAP7_75t_L   g18740(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n18995), .Y(new_n18997));
  A2O1A1O1Ixp25_ASAP7_75t_L g18741(.A1(new_n2706), .A2(new_n2707), .B(new_n18996), .C(new_n18997), .D(new_n11987), .Y(new_n18998));
  O2A1O1Ixp33_ASAP7_75t_L   g18742(.A1(new_n11998), .A2(new_n2708), .B(new_n18995), .C(\a[62] ), .Y(new_n18999));
  NOR2xp33_ASAP7_75t_L      g18743(.A(new_n18998), .B(new_n18999), .Y(new_n19000));
  XOR2x2_ASAP7_75t_L        g18744(.A(new_n18993), .B(new_n19000), .Y(new_n19001));
  INVx1_ASAP7_75t_L         g18745(.A(new_n19001), .Y(new_n19002));
  O2A1O1Ixp33_ASAP7_75t_L   g18746(.A1(new_n18760), .A2(new_n18757), .B(new_n18988), .C(new_n19002), .Y(new_n19003));
  INVx1_ASAP7_75t_L         g18747(.A(new_n19003), .Y(new_n19004));
  O2A1O1Ixp33_ASAP7_75t_L   g18748(.A1(new_n18768), .A2(new_n18769), .B(new_n18758), .C(new_n18761), .Y(new_n19005));
  NAND2xp33_ASAP7_75t_L     g18749(.A(new_n19005), .B(new_n19002), .Y(new_n19006));
  AND2x2_ASAP7_75t_L        g18750(.A(new_n19006), .B(new_n19004), .Y(new_n19007));
  INVx1_ASAP7_75t_L         g18751(.A(new_n19007), .Y(new_n19008));
  NOR2xp33_ASAP7_75t_L      g18752(.A(new_n2879), .B(new_n11354), .Y(new_n19009));
  AOI221xp5_ASAP7_75t_L     g18753(.A1(\b[29] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[28] ), .C(new_n19009), .Y(new_n19010));
  O2A1O1Ixp33_ASAP7_75t_L   g18754(.A1(new_n11053), .A2(new_n3104), .B(new_n19010), .C(new_n11048), .Y(new_n19011));
  O2A1O1Ixp33_ASAP7_75t_L   g18755(.A1(new_n11053), .A2(new_n3104), .B(new_n19010), .C(\a[59] ), .Y(new_n19012));
  INVx1_ASAP7_75t_L         g18756(.A(new_n19012), .Y(new_n19013));
  O2A1O1Ixp33_ASAP7_75t_L   g18757(.A1(new_n19011), .A2(new_n11048), .B(new_n19013), .C(new_n19008), .Y(new_n19014));
  INVx1_ASAP7_75t_L         g18758(.A(new_n19014), .Y(new_n19015));
  O2A1O1Ixp33_ASAP7_75t_L   g18759(.A1(new_n19011), .A2(new_n11048), .B(new_n19013), .C(new_n19007), .Y(new_n19016));
  AOI21xp33_ASAP7_75t_L     g18760(.A1(new_n19015), .A2(new_n19007), .B(new_n19016), .Y(new_n19017));
  O2A1O1Ixp33_ASAP7_75t_L   g18761(.A1(new_n18755), .A2(new_n18781), .B(new_n18778), .C(new_n18775), .Y(new_n19018));
  NAND2xp33_ASAP7_75t_L     g18762(.A(new_n19018), .B(new_n19017), .Y(new_n19019));
  INVx1_ASAP7_75t_L         g18763(.A(new_n19018), .Y(new_n19020));
  A2O1A1Ixp33_ASAP7_75t_L   g18764(.A1(new_n19015), .A2(new_n19007), .B(new_n19016), .C(new_n19020), .Y(new_n19021));
  AND2x2_ASAP7_75t_L        g18765(.A(new_n19021), .B(new_n19019), .Y(new_n19022));
  NOR2xp33_ASAP7_75t_L      g18766(.A(new_n3674), .B(new_n10388), .Y(new_n19023));
  AOI221xp5_ASAP7_75t_L     g18767(.A1(new_n10086), .A2(\b[32] ), .B1(new_n11361), .B2(\b[30] ), .C(new_n19023), .Y(new_n19024));
  O2A1O1Ixp33_ASAP7_75t_L   g18768(.A1(new_n10088), .A2(new_n3897), .B(new_n19024), .C(new_n10083), .Y(new_n19025));
  NOR2xp33_ASAP7_75t_L      g18769(.A(new_n10083), .B(new_n19025), .Y(new_n19026));
  O2A1O1Ixp33_ASAP7_75t_L   g18770(.A1(new_n10088), .A2(new_n3897), .B(new_n19024), .C(\a[56] ), .Y(new_n19027));
  OR3x1_ASAP7_75t_L         g18771(.A(new_n19022), .B(new_n19026), .C(new_n19027), .Y(new_n19028));
  INVx1_ASAP7_75t_L         g18772(.A(new_n19024), .Y(new_n19029));
  A2O1A1Ixp33_ASAP7_75t_L   g18773(.A1(new_n3900), .A2(new_n10386), .B(new_n19029), .C(\a[56] ), .Y(new_n19030));
  A2O1A1Ixp33_ASAP7_75t_L   g18774(.A1(\a[56] ), .A2(new_n19030), .B(new_n19027), .C(new_n19022), .Y(new_n19031));
  AND2x2_ASAP7_75t_L        g18775(.A(new_n19031), .B(new_n19028), .Y(new_n19032));
  A2O1A1Ixp33_ASAP7_75t_L   g18776(.A1(new_n18783), .A2(new_n18987), .B(new_n18795), .C(new_n19032), .Y(new_n19033));
  INVx1_ASAP7_75t_L         g18777(.A(new_n19032), .Y(new_n19034));
  NAND3xp33_ASAP7_75t_L     g18778(.A(new_n19034), .B(new_n18801), .C(new_n18786), .Y(new_n19035));
  NAND3xp33_ASAP7_75t_L     g18779(.A(new_n19035), .B(new_n19033), .C(new_n18986), .Y(new_n19036));
  AO21x2_ASAP7_75t_L        g18780(.A1(new_n19033), .A2(new_n19035), .B(new_n18986), .Y(new_n19037));
  NAND2xp33_ASAP7_75t_L     g18781(.A(new_n19036), .B(new_n19037), .Y(new_n19038));
  NOR2xp33_ASAP7_75t_L      g18782(.A(new_n18980), .B(new_n19038), .Y(new_n19039));
  INVx1_ASAP7_75t_L         g18783(.A(new_n19039), .Y(new_n19040));
  NAND2xp33_ASAP7_75t_L     g18784(.A(new_n18980), .B(new_n19038), .Y(new_n19041));
  AND2x2_ASAP7_75t_L        g18785(.A(new_n19041), .B(new_n19040), .Y(new_n19042));
  NOR2xp33_ASAP7_75t_L      g18786(.A(new_n5074), .B(new_n10065), .Y(new_n19043));
  AOI221xp5_ASAP7_75t_L     g18787(.A1(new_n8175), .A2(\b[38] ), .B1(new_n8484), .B2(\b[36] ), .C(new_n19043), .Y(new_n19044));
  O2A1O1Ixp33_ASAP7_75t_L   g18788(.A1(new_n8176), .A2(new_n5318), .B(new_n19044), .C(new_n8172), .Y(new_n19045));
  INVx1_ASAP7_75t_L         g18789(.A(new_n19045), .Y(new_n19046));
  O2A1O1Ixp33_ASAP7_75t_L   g18790(.A1(new_n8176), .A2(new_n5318), .B(new_n19044), .C(\a[50] ), .Y(new_n19047));
  A2O1A1Ixp33_ASAP7_75t_L   g18791(.A1(\a[50] ), .A2(new_n19046), .B(new_n19047), .C(new_n19042), .Y(new_n19048));
  INVx1_ASAP7_75t_L         g18792(.A(new_n19047), .Y(new_n19049));
  O2A1O1Ixp33_ASAP7_75t_L   g18793(.A1(new_n19045), .A2(new_n8172), .B(new_n19049), .C(new_n19042), .Y(new_n19050));
  AO21x2_ASAP7_75t_L        g18794(.A1(new_n19042), .A2(new_n19048), .B(new_n19050), .Y(new_n19051));
  A2O1A1Ixp33_ASAP7_75t_L   g18795(.A1(new_n18825), .A2(new_n18817), .B(new_n18818), .C(new_n19051), .Y(new_n19052));
  INVx1_ASAP7_75t_L         g18796(.A(new_n18828), .Y(new_n19053));
  O2A1O1Ixp33_ASAP7_75t_L   g18797(.A1(new_n18813), .A2(new_n18816), .B(new_n19053), .C(new_n19051), .Y(new_n19054));
  NOR2xp33_ASAP7_75t_L      g18798(.A(new_n6110), .B(new_n7318), .Y(new_n19055));
  AOI221xp5_ASAP7_75t_L     g18799(.A1(new_n7333), .A2(\b[40] ), .B1(new_n7609), .B2(\b[39] ), .C(new_n19055), .Y(new_n19056));
  O2A1O1Ixp33_ASAP7_75t_L   g18800(.A1(new_n7321), .A2(new_n6117), .B(new_n19056), .C(new_n7316), .Y(new_n19057));
  NOR2xp33_ASAP7_75t_L      g18801(.A(new_n7316), .B(new_n19057), .Y(new_n19058));
  O2A1O1Ixp33_ASAP7_75t_L   g18802(.A1(new_n7321), .A2(new_n6117), .B(new_n19056), .C(\a[47] ), .Y(new_n19059));
  NOR2xp33_ASAP7_75t_L      g18803(.A(new_n19059), .B(new_n19058), .Y(new_n19060));
  A2O1A1Ixp33_ASAP7_75t_L   g18804(.A1(new_n19052), .A2(new_n19051), .B(new_n19054), .C(new_n19060), .Y(new_n19061));
  A2O1A1O1Ixp25_ASAP7_75t_L g18805(.A1(new_n19048), .A2(new_n19042), .B(new_n19050), .C(new_n19052), .D(new_n19054), .Y(new_n19062));
  INVx1_ASAP7_75t_L         g18806(.A(new_n19057), .Y(new_n19063));
  A2O1A1Ixp33_ASAP7_75t_L   g18807(.A1(\a[47] ), .A2(new_n19063), .B(new_n19059), .C(new_n19062), .Y(new_n19064));
  AND2x2_ASAP7_75t_L        g18808(.A(new_n19061), .B(new_n19064), .Y(new_n19065));
  XNOR2x2_ASAP7_75t_L       g18809(.A(new_n18979), .B(new_n19065), .Y(new_n19066));
  XNOR2x2_ASAP7_75t_L       g18810(.A(new_n18978), .B(new_n19066), .Y(new_n19067));
  XNOR2x2_ASAP7_75t_L       g18811(.A(new_n18972), .B(new_n19067), .Y(new_n19068));
  NOR2xp33_ASAP7_75t_L      g18812(.A(new_n7552), .B(new_n5641), .Y(new_n19069));
  AOI221xp5_ASAP7_75t_L     g18813(.A1(\b[45] ), .A2(new_n5920), .B1(\b[46] ), .B2(new_n5623), .C(new_n19069), .Y(new_n19070));
  O2A1O1Ixp33_ASAP7_75t_L   g18814(.A1(new_n5630), .A2(new_n7560), .B(new_n19070), .C(new_n5626), .Y(new_n19071));
  INVx1_ASAP7_75t_L         g18815(.A(new_n19071), .Y(new_n19072));
  O2A1O1Ixp33_ASAP7_75t_L   g18816(.A1(new_n5630), .A2(new_n7560), .B(new_n19070), .C(\a[41] ), .Y(new_n19073));
  A2O1A1Ixp33_ASAP7_75t_L   g18817(.A1(\a[41] ), .A2(new_n19072), .B(new_n19073), .C(new_n19068), .Y(new_n19074));
  INVx1_ASAP7_75t_L         g18818(.A(new_n19073), .Y(new_n19075));
  O2A1O1Ixp33_ASAP7_75t_L   g18819(.A1(new_n19071), .A2(new_n5626), .B(new_n19075), .C(new_n19068), .Y(new_n19076));
  AOI21xp33_ASAP7_75t_L     g18820(.A1(new_n19074), .A2(new_n19068), .B(new_n19076), .Y(new_n19077));
  O2A1O1Ixp33_ASAP7_75t_L   g18821(.A1(new_n18846), .A2(new_n18852), .B(new_n18854), .C(new_n18860), .Y(new_n19078));
  A2O1A1O1Ixp25_ASAP7_75t_L g18822(.A1(new_n18871), .A2(\a[41] ), .B(new_n18868), .C(new_n18861), .D(new_n19078), .Y(new_n19079));
  XNOR2x2_ASAP7_75t_L       g18823(.A(new_n19079), .B(new_n19077), .Y(new_n19080));
  NOR2xp33_ASAP7_75t_L      g18824(.A(new_n8427), .B(new_n4903), .Y(new_n19081));
  AOI221xp5_ASAP7_75t_L     g18825(.A1(\b[48] ), .A2(new_n5139), .B1(\b[50] ), .B2(new_n4917), .C(new_n19081), .Y(new_n19082));
  O2A1O1Ixp33_ASAP7_75t_L   g18826(.A1(new_n4911), .A2(new_n8764), .B(new_n19082), .C(new_n4906), .Y(new_n19083));
  INVx1_ASAP7_75t_L         g18827(.A(new_n19082), .Y(new_n19084));
  A2O1A1Ixp33_ASAP7_75t_L   g18828(.A1(new_n8763), .A2(new_n4912), .B(new_n19084), .C(new_n4906), .Y(new_n19085));
  OA211x2_ASAP7_75t_L       g18829(.A1(new_n4906), .A2(new_n19083), .B(new_n19080), .C(new_n19085), .Y(new_n19086));
  O2A1O1Ixp33_ASAP7_75t_L   g18830(.A1(new_n19083), .A2(new_n4906), .B(new_n19085), .C(new_n19080), .Y(new_n19087));
  NOR2xp33_ASAP7_75t_L      g18831(.A(new_n19087), .B(new_n19086), .Y(new_n19088));
  A2O1A1Ixp33_ASAP7_75t_L   g18832(.A1(new_n18970), .A2(new_n18873), .B(new_n18891), .C(new_n19088), .Y(new_n19089));
  A2O1A1Ixp33_ASAP7_75t_L   g18833(.A1(new_n18970), .A2(new_n18873), .B(new_n18891), .C(new_n19089), .Y(new_n19090));
  O2A1O1Ixp33_ASAP7_75t_L   g18834(.A1(new_n18874), .A2(new_n18877), .B(new_n18873), .C(new_n18891), .Y(new_n19091));
  NAND2xp33_ASAP7_75t_L     g18835(.A(new_n19091), .B(new_n19088), .Y(new_n19092));
  NAND2xp33_ASAP7_75t_L     g18836(.A(new_n19092), .B(new_n19090), .Y(new_n19093));
  NOR2xp33_ASAP7_75t_L      g18837(.A(new_n9355), .B(new_n4142), .Y(new_n19094));
  AOI221xp5_ASAP7_75t_L     g18838(.A1(\b[51] ), .A2(new_n4402), .B1(\b[53] ), .B2(new_n4156), .C(new_n19094), .Y(new_n19095));
  O2A1O1Ixp33_ASAP7_75t_L   g18839(.A1(new_n4150), .A2(new_n9691), .B(new_n19095), .C(new_n4145), .Y(new_n19096));
  INVx1_ASAP7_75t_L         g18840(.A(new_n19096), .Y(new_n19097));
  O2A1O1Ixp33_ASAP7_75t_L   g18841(.A1(new_n4150), .A2(new_n9691), .B(new_n19095), .C(\a[35] ), .Y(new_n19098));
  A2O1A1Ixp33_ASAP7_75t_L   g18842(.A1(new_n19097), .A2(\a[35] ), .B(new_n19098), .C(new_n19093), .Y(new_n19099));
  INVx1_ASAP7_75t_L         g18843(.A(new_n19098), .Y(new_n19100));
  O2A1O1Ixp33_ASAP7_75t_L   g18844(.A1(new_n4145), .A2(new_n19096), .B(new_n19100), .C(new_n19093), .Y(new_n19101));
  A2O1A1Ixp33_ASAP7_75t_L   g18845(.A1(new_n19099), .A2(new_n19093), .B(new_n19101), .C(new_n18969), .Y(new_n19102));
  INVx1_ASAP7_75t_L         g18846(.A(new_n19102), .Y(new_n19103));
  A2O1A1Ixp33_ASAP7_75t_L   g18847(.A1(new_n19099), .A2(new_n19093), .B(new_n19101), .C(new_n18968), .Y(new_n19104));
  OAI21xp33_ASAP7_75t_L     g18848(.A1(new_n18968), .A2(new_n19103), .B(new_n19104), .Y(new_n19105));
  INVx1_ASAP7_75t_L         g18849(.A(new_n19105), .Y(new_n19106));
  A2O1A1Ixp33_ASAP7_75t_L   g18850(.A1(new_n18957), .A2(new_n18953), .B(new_n18958), .C(new_n19106), .Y(new_n19107));
  INVx1_ASAP7_75t_L         g18851(.A(new_n18950), .Y(new_n19108));
  A2O1A1O1Ixp25_ASAP7_75t_L g18852(.A1(new_n19108), .A2(\a[29] ), .B(new_n18951), .C(new_n18957), .D(new_n18958), .Y(new_n19109));
  AOI21xp33_ASAP7_75t_L     g18853(.A1(new_n19097), .A2(\a[35] ), .B(new_n19098), .Y(new_n19110));
  XNOR2x2_ASAP7_75t_L       g18854(.A(new_n19110), .B(new_n19093), .Y(new_n19111));
  NOR2xp33_ASAP7_75t_L      g18855(.A(new_n18968), .B(new_n19111), .Y(new_n19112));
  A2O1A1Ixp33_ASAP7_75t_L   g18856(.A1(new_n19111), .A2(new_n19102), .B(new_n19112), .C(new_n19109), .Y(new_n19113));
  NAND2xp33_ASAP7_75t_L     g18857(.A(new_n19113), .B(new_n19107), .Y(new_n19114));
  XNOR2x2_ASAP7_75t_L       g18858(.A(new_n19114), .B(new_n18947), .Y(new_n19115));
  O2A1O1Ixp33_ASAP7_75t_L   g18859(.A1(new_n18931), .A2(new_n18933), .B(new_n18936), .C(new_n19115), .Y(new_n19116));
  A2O1A1O1Ixp25_ASAP7_75t_L g18860(.A1(new_n12603), .A2(new_n14444), .B(new_n1956), .C(new_n2089), .D(new_n12956), .Y(new_n19117));
  INVx1_ASAP7_75t_L         g18861(.A(new_n18933), .Y(new_n19118));
  A2O1A1O1Ixp25_ASAP7_75t_L g18862(.A1(new_n18929), .A2(new_n19117), .B(new_n18930), .C(new_n19118), .D(new_n18935), .Y(new_n19119));
  AND2x2_ASAP7_75t_L        g18863(.A(new_n19115), .B(new_n19119), .Y(new_n19120));
  NOR2xp33_ASAP7_75t_L      g18864(.A(new_n19116), .B(new_n19120), .Y(new_n19121));
  NOR2xp33_ASAP7_75t_L      g18865(.A(new_n18927), .B(new_n19121), .Y(new_n19122));
  A2O1A1O1Ixp25_ASAP7_75t_L g18866(.A1(new_n18493), .A2(new_n18496), .B(new_n18490), .C(new_n18706), .D(new_n18705), .Y(new_n19123));
  A2O1A1Ixp33_ASAP7_75t_L   g18867(.A1(new_n18910), .A2(new_n18918), .B(new_n18926), .C(new_n19121), .Y(new_n19124));
  OAI21xp33_ASAP7_75t_L     g18868(.A1(new_n19121), .A2(new_n19122), .B(new_n19124), .Y(new_n19125));
  INVx1_ASAP7_75t_L         g18869(.A(new_n19125), .Y(new_n19126));
  O2A1O1Ixp33_ASAP7_75t_L   g18870(.A1(new_n18921), .A2(new_n19123), .B(new_n18920), .C(new_n19126), .Y(new_n19127));
  INVx1_ASAP7_75t_L         g18871(.A(new_n18705), .Y(new_n19128));
  A2O1A1Ixp33_ASAP7_75t_L   g18872(.A1(new_n18707), .A2(new_n19128), .B(new_n18921), .C(new_n18920), .Y(new_n19129));
  O2A1O1Ixp33_ASAP7_75t_L   g18873(.A1(new_n19116), .A2(new_n19120), .B(new_n18927), .C(new_n19129), .Y(new_n19130));
  O2A1O1Ixp33_ASAP7_75t_L   g18874(.A1(new_n19122), .A2(new_n18927), .B(new_n19130), .C(new_n19127), .Y(\f[86] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18875(.A1(new_n18935), .A2(new_n18934), .B(new_n19115), .C(new_n18933), .Y(new_n19132));
  NOR2xp33_ASAP7_75t_L      g18876(.A(new_n12956), .B(new_n2415), .Y(new_n19133));
  AOI221xp5_ASAP7_75t_L     g18877(.A1(\b[61] ), .A2(new_n2577), .B1(\b[62] ), .B2(new_n2421), .C(new_n19133), .Y(new_n19134));
  O2A1O1Ixp33_ASAP7_75t_L   g18878(.A1(new_n2425), .A2(new_n17815), .B(new_n19134), .C(new_n2413), .Y(new_n19135));
  INVx1_ASAP7_75t_L         g18879(.A(new_n19135), .Y(new_n19136));
  O2A1O1Ixp33_ASAP7_75t_L   g18880(.A1(new_n2425), .A2(new_n17815), .B(new_n19134), .C(\a[26] ), .Y(new_n19137));
  AOI21xp33_ASAP7_75t_L     g18881(.A1(new_n19136), .A2(\a[26] ), .B(new_n19137), .Y(new_n19138));
  INVx1_ASAP7_75t_L         g18882(.A(new_n19138), .Y(new_n19139));
  NAND2xp33_ASAP7_75t_L     g18883(.A(new_n18937), .B(new_n18905), .Y(new_n19140));
  NOR2xp33_ASAP7_75t_L      g18884(.A(new_n18945), .B(new_n19140), .Y(new_n19141));
  A2O1A1O1Ixp25_ASAP7_75t_L g18885(.A1(new_n19107), .A2(new_n19113), .B(new_n19141), .C(new_n18946), .D(new_n19138), .Y(new_n19142));
  INVx1_ASAP7_75t_L         g18886(.A(new_n19142), .Y(new_n19143));
  A2O1A1O1Ixp25_ASAP7_75t_L g18887(.A1(new_n19107), .A2(new_n19113), .B(new_n19141), .C(new_n18946), .D(new_n19139), .Y(new_n19144));
  INVx1_ASAP7_75t_L         g18888(.A(new_n18955), .Y(new_n19145));
  O2A1O1Ixp33_ASAP7_75t_L   g18889(.A1(new_n18968), .A2(new_n19103), .B(new_n19104), .C(new_n19109), .Y(new_n19146));
  OAI22xp33_ASAP7_75t_L     g18890(.A1(new_n3133), .A2(new_n11303), .B1(new_n11591), .B2(new_n2925), .Y(new_n19147));
  AOI221xp5_ASAP7_75t_L     g18891(.A1(new_n2938), .A2(\b[60] ), .B1(new_n2932), .B2(new_n13839), .C(new_n19147), .Y(new_n19148));
  XNOR2x2_ASAP7_75t_L       g18892(.A(new_n2928), .B(new_n19148), .Y(new_n19149));
  A2O1A1Ixp33_ASAP7_75t_L   g18893(.A1(new_n19145), .A2(new_n18953), .B(new_n19146), .C(new_n19149), .Y(new_n19150));
  O2A1O1Ixp33_ASAP7_75t_L   g18894(.A1(new_n2928), .A2(new_n18950), .B(new_n18952), .C(new_n19145), .Y(new_n19151));
  O2A1O1Ixp33_ASAP7_75t_L   g18895(.A1(new_n18958), .A2(new_n19151), .B(new_n19105), .C(new_n18956), .Y(new_n19152));
  INVx1_ASAP7_75t_L         g18896(.A(new_n19149), .Y(new_n19153));
  NAND2xp33_ASAP7_75t_L     g18897(.A(new_n19153), .B(new_n19152), .Y(new_n19154));
  NAND2xp33_ASAP7_75t_L     g18898(.A(new_n19150), .B(new_n19154), .Y(new_n19155));
  OAI22xp33_ASAP7_75t_L     g18899(.A1(new_n3703), .A2(new_n10309), .B1(new_n10332), .B2(new_n3509), .Y(new_n19156));
  AOI221xp5_ASAP7_75t_L     g18900(.A1(new_n3503), .A2(\b[57] ), .B1(new_n3505), .B2(new_n10991), .C(new_n19156), .Y(new_n19157));
  XNOR2x2_ASAP7_75t_L       g18901(.A(new_n3493), .B(new_n19157), .Y(new_n19158));
  A2O1A1O1Ixp25_ASAP7_75t_L g18902(.A1(new_n19093), .A2(new_n19099), .B(new_n19101), .C(new_n18965), .D(new_n18966), .Y(new_n19159));
  NAND2xp33_ASAP7_75t_L     g18903(.A(new_n19158), .B(new_n19159), .Y(new_n19160));
  INVx1_ASAP7_75t_L         g18904(.A(new_n19158), .Y(new_n19161));
  A2O1A1Ixp33_ASAP7_75t_L   g18905(.A1(new_n19111), .A2(new_n18965), .B(new_n18966), .C(new_n19161), .Y(new_n19162));
  A2O1A1Ixp33_ASAP7_75t_L   g18906(.A1(new_n19092), .A2(new_n19091), .B(new_n19110), .C(new_n19089), .Y(new_n19163));
  AO21x2_ASAP7_75t_L        g18907(.A1(new_n19068), .A2(new_n19074), .B(new_n19076), .Y(new_n19164));
  O2A1O1Ixp33_ASAP7_75t_L   g18908(.A1(new_n19078), .A2(new_n18870), .B(new_n19164), .C(new_n19087), .Y(new_n19165));
  A2O1A1O1Ixp25_ASAP7_75t_L g18909(.A1(new_n18838), .A2(new_n18840), .B(new_n18836), .C(new_n18830), .D(new_n19065), .Y(new_n19166));
  INVx1_ASAP7_75t_L         g18910(.A(new_n19166), .Y(new_n19167));
  O2A1O1Ixp33_ASAP7_75t_L   g18911(.A1(new_n18761), .A2(new_n18771), .B(new_n19001), .C(new_n19014), .Y(new_n19168));
  INVx1_ASAP7_75t_L         g18912(.A(new_n18991), .Y(new_n19169));
  INVx1_ASAP7_75t_L         g18913(.A(new_n19000), .Y(new_n19170));
  NOR2xp33_ASAP7_75t_L      g18914(.A(new_n2703), .B(new_n12318), .Y(new_n19171));
  AOI221xp5_ASAP7_75t_L     g18915(.A1(new_n11995), .A2(\b[27] ), .B1(new_n13314), .B2(\b[25] ), .C(new_n19171), .Y(new_n19172));
  O2A1O1Ixp33_ASAP7_75t_L   g18916(.A1(new_n11998), .A2(new_n2889), .B(new_n19172), .C(new_n11987), .Y(new_n19173));
  NOR2xp33_ASAP7_75t_L      g18917(.A(new_n11987), .B(new_n19173), .Y(new_n19174));
  O2A1O1Ixp33_ASAP7_75t_L   g18918(.A1(new_n11998), .A2(new_n2889), .B(new_n19172), .C(\a[62] ), .Y(new_n19175));
  NOR2xp33_ASAP7_75t_L      g18919(.A(new_n2188), .B(new_n13030), .Y(new_n19176));
  A2O1A1Ixp33_ASAP7_75t_L   g18920(.A1(new_n13028), .A2(\b[24] ), .B(new_n19176), .C(new_n1952), .Y(new_n19177));
  INVx1_ASAP7_75t_L         g18921(.A(new_n19177), .Y(new_n19178));
  O2A1O1Ixp33_ASAP7_75t_L   g18922(.A1(new_n12669), .A2(new_n12671), .B(\b[24] ), .C(new_n19176), .Y(new_n19179));
  NAND2xp33_ASAP7_75t_L     g18923(.A(\a[23] ), .B(new_n19179), .Y(new_n19180));
  INVx1_ASAP7_75t_L         g18924(.A(new_n19180), .Y(new_n19181));
  NOR2xp33_ASAP7_75t_L      g18925(.A(new_n19178), .B(new_n19181), .Y(new_n19182));
  A2O1A1Ixp33_ASAP7_75t_L   g18926(.A1(new_n13028), .A2(\b[23] ), .B(new_n18989), .C(new_n19182), .Y(new_n19183));
  OAI21xp33_ASAP7_75t_L     g18927(.A1(new_n19178), .A2(new_n19181), .B(new_n18990), .Y(new_n19184));
  AND2x2_ASAP7_75t_L        g18928(.A(new_n19184), .B(new_n19183), .Y(new_n19185));
  INVx1_ASAP7_75t_L         g18929(.A(new_n19185), .Y(new_n19186));
  INVx1_ASAP7_75t_L         g18930(.A(new_n19175), .Y(new_n19187));
  O2A1O1Ixp33_ASAP7_75t_L   g18931(.A1(new_n11987), .A2(new_n19173), .B(new_n19187), .C(new_n19186), .Y(new_n19188));
  INVx1_ASAP7_75t_L         g18932(.A(new_n19188), .Y(new_n19189));
  NOR2xp33_ASAP7_75t_L      g18933(.A(new_n19186), .B(new_n19188), .Y(new_n19190));
  O2A1O1Ixp33_ASAP7_75t_L   g18934(.A1(new_n19174), .A2(new_n19175), .B(new_n19189), .C(new_n19190), .Y(new_n19191));
  A2O1A1Ixp33_ASAP7_75t_L   g18935(.A1(new_n18992), .A2(new_n19170), .B(new_n19169), .C(new_n19191), .Y(new_n19192));
  O2A1O1Ixp33_ASAP7_75t_L   g18936(.A1(new_n18998), .A2(new_n18999), .B(new_n18992), .C(new_n19169), .Y(new_n19193));
  O2A1O1Ixp33_ASAP7_75t_L   g18937(.A1(new_n11987), .A2(new_n19173), .B(new_n19187), .C(new_n19185), .Y(new_n19194));
  A2O1A1Ixp33_ASAP7_75t_L   g18938(.A1(new_n19189), .A2(new_n19185), .B(new_n19194), .C(new_n19193), .Y(new_n19195));
  AND2x2_ASAP7_75t_L        g18939(.A(new_n19195), .B(new_n19192), .Y(new_n19196));
  NOR2xp33_ASAP7_75t_L      g18940(.A(new_n3079), .B(new_n11354), .Y(new_n19197));
  AOI221xp5_ASAP7_75t_L     g18941(.A1(\b[30] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[29] ), .C(new_n19197), .Y(new_n19198));
  O2A1O1Ixp33_ASAP7_75t_L   g18942(.A1(new_n11053), .A2(new_n3464), .B(new_n19198), .C(new_n11048), .Y(new_n19199));
  O2A1O1Ixp33_ASAP7_75t_L   g18943(.A1(new_n11053), .A2(new_n3464), .B(new_n19198), .C(\a[59] ), .Y(new_n19200));
  INVx1_ASAP7_75t_L         g18944(.A(new_n19200), .Y(new_n19201));
  O2A1O1Ixp33_ASAP7_75t_L   g18945(.A1(new_n19199), .A2(new_n11048), .B(new_n19201), .C(new_n19196), .Y(new_n19202));
  INVx1_ASAP7_75t_L         g18946(.A(new_n19202), .Y(new_n19203));
  OAI211xp5_ASAP7_75t_L     g18947(.A1(new_n11048), .A2(new_n19199), .B(new_n19196), .C(new_n19201), .Y(new_n19204));
  AND2x2_ASAP7_75t_L        g18948(.A(new_n19204), .B(new_n19203), .Y(new_n19205));
  XNOR2x2_ASAP7_75t_L       g18949(.A(new_n19168), .B(new_n19205), .Y(new_n19206));
  NOR2xp33_ASAP7_75t_L      g18950(.A(new_n3891), .B(new_n10388), .Y(new_n19207));
  AOI221xp5_ASAP7_75t_L     g18951(.A1(new_n10086), .A2(\b[33] ), .B1(new_n11361), .B2(\b[31] ), .C(new_n19207), .Y(new_n19208));
  O2A1O1Ixp33_ASAP7_75t_L   g18952(.A1(new_n10088), .A2(new_n4108), .B(new_n19208), .C(new_n10083), .Y(new_n19209));
  INVx1_ASAP7_75t_L         g18953(.A(new_n19209), .Y(new_n19210));
  O2A1O1Ixp33_ASAP7_75t_L   g18954(.A1(new_n10088), .A2(new_n4108), .B(new_n19208), .C(\a[56] ), .Y(new_n19211));
  AOI21xp33_ASAP7_75t_L     g18955(.A1(new_n19210), .A2(\a[56] ), .B(new_n19211), .Y(new_n19212));
  O2A1O1Ixp33_ASAP7_75t_L   g18956(.A1(new_n19017), .A2(new_n19018), .B(new_n19031), .C(new_n19212), .Y(new_n19213));
  INVx1_ASAP7_75t_L         g18957(.A(new_n19021), .Y(new_n19214));
  O2A1O1Ixp33_ASAP7_75t_L   g18958(.A1(new_n19026), .A2(new_n19027), .B(new_n19019), .C(new_n19214), .Y(new_n19215));
  AND2x2_ASAP7_75t_L        g18959(.A(new_n19212), .B(new_n19215), .Y(new_n19216));
  NOR2xp33_ASAP7_75t_L      g18960(.A(new_n19216), .B(new_n19213), .Y(new_n19217));
  XOR2x2_ASAP7_75t_L        g18961(.A(new_n19206), .B(new_n19217), .Y(new_n19218));
  NOR2xp33_ASAP7_75t_L      g18962(.A(new_n4581), .B(new_n10400), .Y(new_n19219));
  AOI221xp5_ASAP7_75t_L     g18963(.A1(new_n9102), .A2(\b[36] ), .B1(new_n10398), .B2(\b[34] ), .C(new_n19219), .Y(new_n19220));
  O2A1O1Ixp33_ASAP7_75t_L   g18964(.A1(new_n9104), .A2(new_n4622), .B(new_n19220), .C(new_n9099), .Y(new_n19221));
  INVx1_ASAP7_75t_L         g18965(.A(new_n19221), .Y(new_n19222));
  O2A1O1Ixp33_ASAP7_75t_L   g18966(.A1(new_n9104), .A2(new_n4622), .B(new_n19220), .C(\a[53] ), .Y(new_n19223));
  A2O1A1Ixp33_ASAP7_75t_L   g18967(.A1(\a[53] ), .A2(new_n19222), .B(new_n19223), .C(new_n19218), .Y(new_n19224));
  INVx1_ASAP7_75t_L         g18968(.A(new_n19223), .Y(new_n19225));
  O2A1O1Ixp33_ASAP7_75t_L   g18969(.A1(new_n19221), .A2(new_n9099), .B(new_n19225), .C(new_n19218), .Y(new_n19226));
  AO21x2_ASAP7_75t_L        g18970(.A1(new_n19218), .A2(new_n19224), .B(new_n19226), .Y(new_n19227));
  A2O1A1Ixp33_ASAP7_75t_L   g18971(.A1(new_n18801), .A2(new_n18786), .B(new_n19034), .C(new_n19036), .Y(new_n19228));
  INVx1_ASAP7_75t_L         g18972(.A(new_n19228), .Y(new_n19229));
  XNOR2x2_ASAP7_75t_L       g18973(.A(new_n19229), .B(new_n19227), .Y(new_n19230));
  INVx1_ASAP7_75t_L         g18974(.A(new_n19230), .Y(new_n19231));
  NOR2xp33_ASAP7_75t_L      g18975(.A(new_n5311), .B(new_n10065), .Y(new_n19232));
  AOI221xp5_ASAP7_75t_L     g18976(.A1(new_n8175), .A2(\b[39] ), .B1(new_n8484), .B2(\b[37] ), .C(new_n19232), .Y(new_n19233));
  O2A1O1Ixp33_ASAP7_75t_L   g18977(.A1(new_n8176), .A2(new_n5578), .B(new_n19233), .C(new_n8172), .Y(new_n19234));
  INVx1_ASAP7_75t_L         g18978(.A(new_n19234), .Y(new_n19235));
  O2A1O1Ixp33_ASAP7_75t_L   g18979(.A1(new_n8176), .A2(new_n5578), .B(new_n19233), .C(\a[50] ), .Y(new_n19236));
  A2O1A1Ixp33_ASAP7_75t_L   g18980(.A1(\a[50] ), .A2(new_n19235), .B(new_n19236), .C(new_n19230), .Y(new_n19237));
  INVx1_ASAP7_75t_L         g18981(.A(new_n19237), .Y(new_n19238));
  INVx1_ASAP7_75t_L         g18982(.A(new_n19236), .Y(new_n19239));
  O2A1O1Ixp33_ASAP7_75t_L   g18983(.A1(new_n19234), .A2(new_n8172), .B(new_n19239), .C(new_n19230), .Y(new_n19240));
  INVx1_ASAP7_75t_L         g18984(.A(new_n19240), .Y(new_n19241));
  A2O1A1O1Ixp25_ASAP7_75t_L g18985(.A1(new_n19046), .A2(\a[50] ), .B(new_n19047), .C(new_n19041), .D(new_n19039), .Y(new_n19242));
  OAI211xp5_ASAP7_75t_L     g18986(.A1(new_n19231), .A2(new_n19238), .B(new_n19241), .C(new_n19242), .Y(new_n19243));
  INVx1_ASAP7_75t_L         g18987(.A(new_n19242), .Y(new_n19244));
  A2O1A1Ixp33_ASAP7_75t_L   g18988(.A1(new_n19237), .A2(new_n19230), .B(new_n19240), .C(new_n19244), .Y(new_n19245));
  NAND2xp33_ASAP7_75t_L     g18989(.A(new_n19245), .B(new_n19243), .Y(new_n19246));
  NOR2xp33_ASAP7_75t_L      g18990(.A(new_n6110), .B(new_n7312), .Y(new_n19247));
  AOI221xp5_ASAP7_75t_L     g18991(.A1(\b[40] ), .A2(new_n7609), .B1(\b[42] ), .B2(new_n7334), .C(new_n19247), .Y(new_n19248));
  O2A1O1Ixp33_ASAP7_75t_L   g18992(.A1(new_n7321), .A2(new_n6386), .B(new_n19248), .C(new_n7316), .Y(new_n19249));
  O2A1O1Ixp33_ASAP7_75t_L   g18993(.A1(new_n7321), .A2(new_n6386), .B(new_n19248), .C(\a[47] ), .Y(new_n19250));
  INVx1_ASAP7_75t_L         g18994(.A(new_n19250), .Y(new_n19251));
  O2A1O1Ixp33_ASAP7_75t_L   g18995(.A1(new_n19249), .A2(new_n7316), .B(new_n19251), .C(new_n19246), .Y(new_n19252));
  INVx1_ASAP7_75t_L         g18996(.A(new_n19246), .Y(new_n19253));
  O2A1O1Ixp33_ASAP7_75t_L   g18997(.A1(new_n19249), .A2(new_n7316), .B(new_n19251), .C(new_n19253), .Y(new_n19254));
  INVx1_ASAP7_75t_L         g18998(.A(new_n19254), .Y(new_n19255));
  OAI21xp33_ASAP7_75t_L     g18999(.A1(new_n19246), .A2(new_n19252), .B(new_n19255), .Y(new_n19256));
  O2A1O1Ixp33_ASAP7_75t_L   g19000(.A1(new_n19062), .A2(new_n19060), .B(new_n19052), .C(new_n19256), .Y(new_n19257));
  INVx1_ASAP7_75t_L         g19001(.A(new_n18822), .Y(new_n19258));
  A2O1A1O1Ixp25_ASAP7_75t_L g19002(.A1(new_n19258), .A2(\a[50] ), .B(new_n18823), .C(new_n18817), .D(new_n18818), .Y(new_n19259));
  A2O1A1Ixp33_ASAP7_75t_L   g19003(.A1(new_n19048), .A2(new_n19042), .B(new_n19050), .C(new_n19259), .Y(new_n19260));
  A2O1A1Ixp33_ASAP7_75t_L   g19004(.A1(new_n19259), .A2(new_n19260), .B(new_n19060), .C(new_n19052), .Y(new_n19261));
  O2A1O1Ixp33_ASAP7_75t_L   g19005(.A1(new_n19246), .A2(new_n19252), .B(new_n19255), .C(new_n19261), .Y(new_n19262));
  NOR2xp33_ASAP7_75t_L      g19006(.A(new_n19262), .B(new_n19257), .Y(new_n19263));
  NOR2xp33_ASAP7_75t_L      g19007(.A(new_n6671), .B(new_n6741), .Y(new_n19264));
  AOI221xp5_ASAP7_75t_L     g19008(.A1(\b[45] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[44] ), .C(new_n19264), .Y(new_n19265));
  O2A1O1Ixp33_ASAP7_75t_L   g19009(.A1(new_n6443), .A2(new_n7255), .B(new_n19265), .C(new_n6439), .Y(new_n19266));
  O2A1O1Ixp33_ASAP7_75t_L   g19010(.A1(new_n6443), .A2(new_n7255), .B(new_n19265), .C(\a[44] ), .Y(new_n19267));
  INVx1_ASAP7_75t_L         g19011(.A(new_n19267), .Y(new_n19268));
  O2A1O1Ixp33_ASAP7_75t_L   g19012(.A1(new_n19266), .A2(new_n6439), .B(new_n19268), .C(new_n19263), .Y(new_n19269));
  INVx1_ASAP7_75t_L         g19013(.A(new_n19269), .Y(new_n19270));
  OAI211xp5_ASAP7_75t_L     g19014(.A1(new_n6439), .A2(new_n19266), .B(new_n19263), .C(new_n19268), .Y(new_n19271));
  NAND2xp33_ASAP7_75t_L     g19015(.A(new_n19271), .B(new_n19270), .Y(new_n19272));
  OAI211xp5_ASAP7_75t_L     g19016(.A1(new_n18978), .A2(new_n19066), .B(new_n19272), .C(new_n19167), .Y(new_n19273));
  O2A1O1Ixp33_ASAP7_75t_L   g19017(.A1(new_n18978), .A2(new_n19066), .B(new_n19167), .C(new_n19272), .Y(new_n19274));
  INVx1_ASAP7_75t_L         g19018(.A(new_n19274), .Y(new_n19275));
  NAND2xp33_ASAP7_75t_L     g19019(.A(new_n19273), .B(new_n19275), .Y(new_n19276));
  NOR2xp33_ASAP7_75t_L      g19020(.A(new_n7860), .B(new_n5641), .Y(new_n19277));
  AOI221xp5_ASAP7_75t_L     g19021(.A1(\b[46] ), .A2(new_n5920), .B1(\b[47] ), .B2(new_n5623), .C(new_n19277), .Y(new_n19278));
  O2A1O1Ixp33_ASAP7_75t_L   g19022(.A1(new_n5630), .A2(new_n7868), .B(new_n19278), .C(new_n5626), .Y(new_n19279));
  O2A1O1Ixp33_ASAP7_75t_L   g19023(.A1(new_n5630), .A2(new_n7868), .B(new_n19278), .C(\a[41] ), .Y(new_n19280));
  INVx1_ASAP7_75t_L         g19024(.A(new_n19280), .Y(new_n19281));
  O2A1O1Ixp33_ASAP7_75t_L   g19025(.A1(new_n19279), .A2(new_n5626), .B(new_n19281), .C(new_n19276), .Y(new_n19282));
  INVx1_ASAP7_75t_L         g19026(.A(new_n19279), .Y(new_n19283));
  A2O1A1Ixp33_ASAP7_75t_L   g19027(.A1(\a[41] ), .A2(new_n19283), .B(new_n19280), .C(new_n19276), .Y(new_n19284));
  OAI21xp33_ASAP7_75t_L     g19028(.A1(new_n19276), .A2(new_n19282), .B(new_n19284), .Y(new_n19285));
  INVx1_ASAP7_75t_L         g19029(.A(new_n18852), .Y(new_n19286));
  A2O1A1Ixp33_ASAP7_75t_L   g19030(.A1(new_n19286), .A2(new_n18843), .B(new_n19067), .C(new_n19074), .Y(new_n19287));
  NOR2xp33_ASAP7_75t_L      g19031(.A(new_n19287), .B(new_n19285), .Y(new_n19288));
  NAND2xp33_ASAP7_75t_L     g19032(.A(new_n19287), .B(new_n19285), .Y(new_n19289));
  INVx1_ASAP7_75t_L         g19033(.A(new_n19289), .Y(new_n19290));
  NOR2xp33_ASAP7_75t_L      g19034(.A(new_n19288), .B(new_n19290), .Y(new_n19291));
  NOR2xp33_ASAP7_75t_L      g19035(.A(new_n8779), .B(new_n4908), .Y(new_n19292));
  AOI221xp5_ASAP7_75t_L     g19036(.A1(\b[49] ), .A2(new_n5139), .B1(\b[50] ), .B2(new_n4916), .C(new_n19292), .Y(new_n19293));
  O2A1O1Ixp33_ASAP7_75t_L   g19037(.A1(new_n4911), .A2(new_n8789), .B(new_n19293), .C(new_n4906), .Y(new_n19294));
  INVx1_ASAP7_75t_L         g19038(.A(new_n19294), .Y(new_n19295));
  O2A1O1Ixp33_ASAP7_75t_L   g19039(.A1(new_n4911), .A2(new_n8789), .B(new_n19293), .C(\a[38] ), .Y(new_n19296));
  A2O1A1Ixp33_ASAP7_75t_L   g19040(.A1(\a[38] ), .A2(new_n19295), .B(new_n19296), .C(new_n19291), .Y(new_n19297));
  INVx1_ASAP7_75t_L         g19041(.A(new_n19293), .Y(new_n19298));
  NOR2xp33_ASAP7_75t_L      g19042(.A(new_n4906), .B(new_n19294), .Y(new_n19299));
  A2O1A1O1Ixp25_ASAP7_75t_L g19043(.A1(new_n8790), .A2(new_n4912), .B(new_n19298), .C(new_n19295), .D(new_n19299), .Y(new_n19300));
  O2A1O1Ixp33_ASAP7_75t_L   g19044(.A1(new_n19288), .A2(new_n19290), .B(new_n19300), .C(new_n19165), .Y(new_n19301));
  INVx1_ASAP7_75t_L         g19045(.A(new_n19300), .Y(new_n19302));
  O2A1O1Ixp33_ASAP7_75t_L   g19046(.A1(new_n19299), .A2(new_n19296), .B(new_n19291), .C(new_n19301), .Y(new_n19303));
  OAI21xp33_ASAP7_75t_L     g19047(.A1(new_n19291), .A2(new_n19302), .B(new_n19303), .Y(new_n19304));
  A2O1A1Ixp33_ASAP7_75t_L   g19048(.A1(new_n19297), .A2(new_n19301), .B(new_n19165), .C(new_n19304), .Y(new_n19305));
  NOR2xp33_ASAP7_75t_L      g19049(.A(new_n9709), .B(new_n4147), .Y(new_n19306));
  AOI221xp5_ASAP7_75t_L     g19050(.A1(\b[52] ), .A2(new_n4402), .B1(\b[53] ), .B2(new_n4155), .C(new_n19306), .Y(new_n19307));
  O2A1O1Ixp33_ASAP7_75t_L   g19051(.A1(new_n4150), .A2(new_n9718), .B(new_n19307), .C(new_n4145), .Y(new_n19308));
  INVx1_ASAP7_75t_L         g19052(.A(new_n19308), .Y(new_n19309));
  O2A1O1Ixp33_ASAP7_75t_L   g19053(.A1(new_n4150), .A2(new_n9718), .B(new_n19307), .C(\a[35] ), .Y(new_n19310));
  AOI21xp33_ASAP7_75t_L     g19054(.A1(new_n19309), .A2(\a[35] ), .B(new_n19310), .Y(new_n19311));
  XNOR2x2_ASAP7_75t_L       g19055(.A(new_n19311), .B(new_n19305), .Y(new_n19312));
  NAND2xp33_ASAP7_75t_L     g19056(.A(new_n19163), .B(new_n19312), .Y(new_n19313));
  OR2x4_ASAP7_75t_L         g19057(.A(new_n19163), .B(new_n19312), .Y(new_n19314));
  NAND4xp25_ASAP7_75t_L     g19058(.A(new_n19314), .B(new_n19160), .C(new_n19162), .D(new_n19313), .Y(new_n19315));
  AO22x1_ASAP7_75t_L        g19059(.A1(new_n19160), .A2(new_n19162), .B1(new_n19313), .B2(new_n19314), .Y(new_n19316));
  NAND3xp33_ASAP7_75t_L     g19060(.A(new_n19155), .B(new_n19315), .C(new_n19316), .Y(new_n19317));
  AND3x1_ASAP7_75t_L        g19061(.A(new_n19317), .B(new_n19316), .C(new_n19315), .Y(new_n19318));
  AOI21xp33_ASAP7_75t_L     g19062(.A1(new_n19317), .A2(new_n19155), .B(new_n19318), .Y(new_n19319));
  A2O1A1Ixp33_ASAP7_75t_L   g19063(.A1(new_n19143), .A2(new_n19139), .B(new_n19144), .C(new_n19319), .Y(new_n19320));
  A2O1A1O1Ixp25_ASAP7_75t_L g19064(.A1(new_n19136), .A2(\a[26] ), .B(new_n19137), .C(new_n19143), .D(new_n19144), .Y(new_n19321));
  A2O1A1Ixp33_ASAP7_75t_L   g19065(.A1(new_n19155), .A2(new_n19317), .B(new_n19318), .C(new_n19321), .Y(new_n19322));
  NAND2xp33_ASAP7_75t_L     g19066(.A(new_n19320), .B(new_n19322), .Y(new_n19323));
  XNOR2x2_ASAP7_75t_L       g19067(.A(new_n19132), .B(new_n19323), .Y(new_n19324));
  A2O1A1Ixp33_ASAP7_75t_L   g19068(.A1(new_n18929), .A2(new_n19117), .B(new_n18930), .C(new_n19118), .Y(new_n19325));
  A2O1A1Ixp33_ASAP7_75t_L   g19069(.A1(new_n18910), .A2(new_n18932), .B(new_n18933), .C(new_n19325), .Y(new_n19326));
  A2O1A1Ixp33_ASAP7_75t_L   g19070(.A1(new_n19326), .A2(new_n19115), .B(new_n18933), .C(new_n19323), .Y(new_n19327));
  INVx1_ASAP7_75t_L         g19071(.A(new_n18920), .Y(new_n19328));
  O2A1O1Ixp33_ASAP7_75t_L   g19072(.A1(new_n19328), .A2(new_n18922), .B(new_n19125), .C(new_n19122), .Y(new_n19329));
  INVx1_ASAP7_75t_L         g19073(.A(new_n19132), .Y(new_n19330));
  A2O1A1Ixp33_ASAP7_75t_L   g19074(.A1(new_n19320), .A2(new_n19322), .B(new_n19330), .C(new_n19329), .Y(new_n19331));
  A2O1A1O1Ixp25_ASAP7_75t_L g19075(.A1(new_n19326), .A2(new_n19115), .B(new_n18933), .C(new_n19327), .D(new_n19331), .Y(new_n19332));
  O2A1O1Ixp33_ASAP7_75t_L   g19076(.A1(new_n19122), .A2(new_n19127), .B(new_n19324), .C(new_n19332), .Y(\f[87] ));
  INVx1_ASAP7_75t_L         g19077(.A(new_n19144), .Y(new_n19334));
  A2O1A1Ixp33_ASAP7_75t_L   g19078(.A1(new_n19138), .A2(new_n19334), .B(new_n19319), .C(new_n19143), .Y(new_n19335));
  INVx1_ASAP7_75t_L         g19079(.A(new_n19335), .Y(new_n19336));
  NOR2xp33_ASAP7_75t_L      g19080(.A(new_n11626), .B(new_n2925), .Y(new_n19337));
  AOI221xp5_ASAP7_75t_L     g19081(.A1(\b[59] ), .A2(new_n3129), .B1(\b[61] ), .B2(new_n2938), .C(new_n19337), .Y(new_n19338));
  O2A1O1Ixp33_ASAP7_75t_L   g19082(.A1(new_n2940), .A2(new_n14764), .B(new_n19338), .C(new_n2928), .Y(new_n19339));
  INVx1_ASAP7_75t_L         g19083(.A(new_n19339), .Y(new_n19340));
  O2A1O1Ixp33_ASAP7_75t_L   g19084(.A1(new_n2940), .A2(new_n14764), .B(new_n19338), .C(\a[29] ), .Y(new_n19341));
  AOI21xp33_ASAP7_75t_L     g19085(.A1(new_n19340), .A2(\a[29] ), .B(new_n19341), .Y(new_n19342));
  O2A1O1Ixp33_ASAP7_75t_L   g19086(.A1(new_n19158), .A2(new_n19159), .B(new_n19315), .C(new_n19342), .Y(new_n19343));
  INVx1_ASAP7_75t_L         g19087(.A(new_n19343), .Y(new_n19344));
  O2A1O1Ixp33_ASAP7_75t_L   g19088(.A1(new_n19158), .A2(new_n19159), .B(new_n19315), .C(new_n19343), .Y(new_n19345));
  A2O1A1O1Ixp25_ASAP7_75t_L g19089(.A1(new_n19340), .A2(\a[29] ), .B(new_n19341), .C(new_n19344), .D(new_n19345), .Y(new_n19346));
  A2O1A1Ixp33_ASAP7_75t_L   g19090(.A1(new_n19102), .A2(new_n18967), .B(new_n19158), .C(new_n19315), .Y(new_n19347));
  NAND2xp33_ASAP7_75t_L     g19091(.A(new_n19342), .B(new_n19347), .Y(new_n19348));
  A2O1A1O1Ixp25_ASAP7_75t_L g19092(.A1(new_n19297), .A2(new_n19301), .B(new_n19165), .C(new_n19304), .D(new_n19311), .Y(new_n19349));
  NAND2xp33_ASAP7_75t_L     g19093(.A(\b[57] ), .B(new_n3499), .Y(new_n19350));
  OAI221xp5_ASAP7_75t_L     g19094(.A1(new_n3510), .A2(new_n11303), .B1(new_n10332), .B2(new_n3703), .C(new_n19350), .Y(new_n19351));
  AOI21xp33_ASAP7_75t_L     g19095(.A1(new_n11314), .A2(new_n3505), .B(new_n19351), .Y(new_n19352));
  NAND2xp33_ASAP7_75t_L     g19096(.A(\a[32] ), .B(new_n19352), .Y(new_n19353));
  A2O1A1Ixp33_ASAP7_75t_L   g19097(.A1(new_n11314), .A2(new_n3505), .B(new_n19351), .C(new_n3493), .Y(new_n19354));
  NAND2xp33_ASAP7_75t_L     g19098(.A(new_n19354), .B(new_n19353), .Y(new_n19355));
  A2O1A1Ixp33_ASAP7_75t_L   g19099(.A1(new_n19312), .A2(new_n19163), .B(new_n19349), .C(new_n19355), .Y(new_n19356));
  A2O1A1Ixp33_ASAP7_75t_L   g19100(.A1(\a[35] ), .A2(new_n19309), .B(new_n19310), .C(new_n19305), .Y(new_n19357));
  NAND4xp25_ASAP7_75t_L     g19101(.A(new_n19313), .B(new_n19353), .C(new_n19354), .D(new_n19357), .Y(new_n19358));
  NAND2xp33_ASAP7_75t_L     g19102(.A(new_n19218), .B(new_n19224), .Y(new_n19359));
  A2O1A1Ixp33_ASAP7_75t_L   g19103(.A1(new_n19222), .A2(\a[53] ), .B(new_n19223), .C(new_n19224), .Y(new_n19360));
  A2O1A1Ixp33_ASAP7_75t_L   g19104(.A1(new_n19360), .A2(new_n19359), .B(new_n19229), .C(new_n19224), .Y(new_n19361));
  INVx1_ASAP7_75t_L         g19105(.A(new_n19213), .Y(new_n19362));
  NAND2xp33_ASAP7_75t_L     g19106(.A(new_n19206), .B(new_n19217), .Y(new_n19363));
  INVx1_ASAP7_75t_L         g19107(.A(new_n19194), .Y(new_n19364));
  A2O1A1Ixp33_ASAP7_75t_L   g19108(.A1(new_n19364), .A2(new_n19186), .B(new_n19193), .C(new_n19189), .Y(new_n19365));
  NOR2xp33_ASAP7_75t_L      g19109(.A(new_n2205), .B(new_n13030), .Y(new_n19366));
  A2O1A1O1Ixp25_ASAP7_75t_L g19110(.A1(new_n13028), .A2(\b[23] ), .B(new_n18989), .C(new_n19180), .D(new_n19178), .Y(new_n19367));
  A2O1A1Ixp33_ASAP7_75t_L   g19111(.A1(new_n13028), .A2(\b[25] ), .B(new_n19366), .C(new_n19367), .Y(new_n19368));
  O2A1O1Ixp33_ASAP7_75t_L   g19112(.A1(new_n12669), .A2(new_n12671), .B(\b[25] ), .C(new_n19366), .Y(new_n19369));
  INVx1_ASAP7_75t_L         g19113(.A(new_n19369), .Y(new_n19370));
  O2A1O1Ixp33_ASAP7_75t_L   g19114(.A1(new_n18990), .A2(new_n19181), .B(new_n19177), .C(new_n19370), .Y(new_n19371));
  INVx1_ASAP7_75t_L         g19115(.A(new_n19371), .Y(new_n19372));
  NAND2xp33_ASAP7_75t_L     g19116(.A(new_n19368), .B(new_n19372), .Y(new_n19373));
  NOR2xp33_ASAP7_75t_L      g19117(.A(new_n2879), .B(new_n12318), .Y(new_n19374));
  AOI221xp5_ASAP7_75t_L     g19118(.A1(new_n11995), .A2(\b[28] ), .B1(new_n13314), .B2(\b[26] ), .C(new_n19374), .Y(new_n19375));
  INVx1_ASAP7_75t_L         g19119(.A(new_n19375), .Y(new_n19376));
  A2O1A1Ixp33_ASAP7_75t_L   g19120(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n19375), .Y(new_n19377));
  O2A1O1Ixp33_ASAP7_75t_L   g19121(.A1(new_n19376), .A2(new_n3085), .B(new_n19377), .C(new_n11987), .Y(new_n19378));
  O2A1O1Ixp33_ASAP7_75t_L   g19122(.A1(new_n11998), .A2(new_n3087), .B(new_n19375), .C(\a[62] ), .Y(new_n19379));
  NOR2xp33_ASAP7_75t_L      g19123(.A(new_n19378), .B(new_n19379), .Y(new_n19380));
  NOR2xp33_ASAP7_75t_L      g19124(.A(new_n19373), .B(new_n19380), .Y(new_n19381));
  INVx1_ASAP7_75t_L         g19125(.A(new_n19381), .Y(new_n19382));
  NAND2xp33_ASAP7_75t_L     g19126(.A(new_n19373), .B(new_n19380), .Y(new_n19383));
  AND2x2_ASAP7_75t_L        g19127(.A(new_n19383), .B(new_n19382), .Y(new_n19384));
  NAND2xp33_ASAP7_75t_L     g19128(.A(new_n19365), .B(new_n19384), .Y(new_n19385));
  O2A1O1Ixp33_ASAP7_75t_L   g19129(.A1(new_n19186), .A2(new_n19188), .B(new_n19364), .C(new_n19193), .Y(new_n19386));
  O2A1O1Ixp33_ASAP7_75t_L   g19130(.A1(new_n19174), .A2(new_n19175), .B(new_n19185), .C(new_n19386), .Y(new_n19387));
  INVx1_ASAP7_75t_L         g19131(.A(new_n19384), .Y(new_n19388));
  NAND2xp33_ASAP7_75t_L     g19132(.A(new_n19387), .B(new_n19388), .Y(new_n19389));
  AND2x2_ASAP7_75t_L        g19133(.A(new_n19385), .B(new_n19389), .Y(new_n19390));
  NOR2xp33_ASAP7_75t_L      g19134(.A(new_n3098), .B(new_n11354), .Y(new_n19391));
  AOI221xp5_ASAP7_75t_L     g19135(.A1(\b[31] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[30] ), .C(new_n19391), .Y(new_n19392));
  O2A1O1Ixp33_ASAP7_75t_L   g19136(.A1(new_n11053), .A2(new_n3681), .B(new_n19392), .C(new_n11048), .Y(new_n19393));
  INVx1_ASAP7_75t_L         g19137(.A(new_n19393), .Y(new_n19394));
  O2A1O1Ixp33_ASAP7_75t_L   g19138(.A1(new_n11053), .A2(new_n3681), .B(new_n19392), .C(\a[59] ), .Y(new_n19395));
  A2O1A1Ixp33_ASAP7_75t_L   g19139(.A1(\a[59] ), .A2(new_n19394), .B(new_n19395), .C(new_n19390), .Y(new_n19396));
  NAND2xp33_ASAP7_75t_L     g19140(.A(new_n19390), .B(new_n19396), .Y(new_n19397));
  INVx1_ASAP7_75t_L         g19141(.A(new_n19390), .Y(new_n19398));
  A2O1A1Ixp33_ASAP7_75t_L   g19142(.A1(\a[59] ), .A2(new_n19394), .B(new_n19395), .C(new_n19398), .Y(new_n19399));
  AND2x2_ASAP7_75t_L        g19143(.A(new_n19399), .B(new_n19397), .Y(new_n19400));
  O2A1O1Ixp33_ASAP7_75t_L   g19144(.A1(new_n19014), .A2(new_n19003), .B(new_n19204), .C(new_n19202), .Y(new_n19401));
  NAND2xp33_ASAP7_75t_L     g19145(.A(new_n19401), .B(new_n19400), .Y(new_n19402));
  INVx1_ASAP7_75t_L         g19146(.A(new_n19396), .Y(new_n19403));
  O2A1O1Ixp33_ASAP7_75t_L   g19147(.A1(new_n19398), .A2(new_n19403), .B(new_n19399), .C(new_n19401), .Y(new_n19404));
  INVx1_ASAP7_75t_L         g19148(.A(new_n19404), .Y(new_n19405));
  AND2x2_ASAP7_75t_L        g19149(.A(new_n19405), .B(new_n19402), .Y(new_n19406));
  INVx1_ASAP7_75t_L         g19150(.A(new_n19406), .Y(new_n19407));
  NOR2xp33_ASAP7_75t_L      g19151(.A(new_n4101), .B(new_n10388), .Y(new_n19408));
  AOI221xp5_ASAP7_75t_L     g19152(.A1(new_n10086), .A2(\b[34] ), .B1(new_n11361), .B2(\b[32] ), .C(new_n19408), .Y(new_n19409));
  O2A1O1Ixp33_ASAP7_75t_L   g19153(.A1(new_n10088), .A2(new_n4352), .B(new_n19409), .C(new_n10083), .Y(new_n19410));
  O2A1O1Ixp33_ASAP7_75t_L   g19154(.A1(new_n10088), .A2(new_n4352), .B(new_n19409), .C(\a[56] ), .Y(new_n19411));
  INVx1_ASAP7_75t_L         g19155(.A(new_n19411), .Y(new_n19412));
  O2A1O1Ixp33_ASAP7_75t_L   g19156(.A1(new_n19410), .A2(new_n10083), .B(new_n19412), .C(new_n19407), .Y(new_n19413));
  INVx1_ASAP7_75t_L         g19157(.A(new_n19413), .Y(new_n19414));
  O2A1O1Ixp33_ASAP7_75t_L   g19158(.A1(new_n19410), .A2(new_n10083), .B(new_n19412), .C(new_n19406), .Y(new_n19415));
  AOI21xp33_ASAP7_75t_L     g19159(.A1(new_n19414), .A2(new_n19406), .B(new_n19415), .Y(new_n19416));
  NAND3xp33_ASAP7_75t_L     g19160(.A(new_n19416), .B(new_n19363), .C(new_n19362), .Y(new_n19417));
  A2O1A1Ixp33_ASAP7_75t_L   g19161(.A1(new_n19031), .A2(new_n19021), .B(new_n19212), .C(new_n19363), .Y(new_n19418));
  A2O1A1Ixp33_ASAP7_75t_L   g19162(.A1(new_n19414), .A2(new_n19406), .B(new_n19415), .C(new_n19418), .Y(new_n19419));
  AND2x2_ASAP7_75t_L        g19163(.A(new_n19419), .B(new_n19417), .Y(new_n19420));
  NOR2xp33_ASAP7_75t_L      g19164(.A(new_n4613), .B(new_n10400), .Y(new_n19421));
  AOI221xp5_ASAP7_75t_L     g19165(.A1(new_n9102), .A2(\b[37] ), .B1(new_n10398), .B2(\b[35] ), .C(new_n19421), .Y(new_n19422));
  INVx1_ASAP7_75t_L         g19166(.A(new_n19422), .Y(new_n19423));
  O2A1O1Ixp33_ASAP7_75t_L   g19167(.A1(new_n9104), .A2(new_n5083), .B(new_n19422), .C(new_n9099), .Y(new_n19424));
  INVx1_ASAP7_75t_L         g19168(.A(new_n19424), .Y(new_n19425));
  NOR2xp33_ASAP7_75t_L      g19169(.A(new_n9099), .B(new_n19424), .Y(new_n19426));
  A2O1A1O1Ixp25_ASAP7_75t_L g19170(.A1(new_n9437), .A2(new_n10229), .B(new_n19423), .C(new_n19425), .D(new_n19426), .Y(new_n19427));
  XNOR2x2_ASAP7_75t_L       g19171(.A(new_n19427), .B(new_n19420), .Y(new_n19428));
  NAND2xp33_ASAP7_75t_L     g19172(.A(new_n19361), .B(new_n19428), .Y(new_n19429));
  NAND2xp33_ASAP7_75t_L     g19173(.A(new_n19361), .B(new_n19429), .Y(new_n19430));
  A2O1A1Ixp33_ASAP7_75t_L   g19174(.A1(new_n19224), .A2(new_n19218), .B(new_n19226), .C(new_n19228), .Y(new_n19431));
  NAND2xp33_ASAP7_75t_L     g19175(.A(\b[39] ), .B(new_n8169), .Y(new_n19432));
  OAI221xp5_ASAP7_75t_L     g19176(.A1(new_n8483), .A2(new_n5311), .B1(new_n5855), .B2(new_n8843), .C(new_n19432), .Y(new_n19433));
  A2O1A1Ixp33_ASAP7_75t_L   g19177(.A1(new_n6651), .A2(new_n8490), .B(new_n19433), .C(\a[50] ), .Y(new_n19434));
  AOI211xp5_ASAP7_75t_L     g19178(.A1(new_n6651), .A2(new_n8490), .B(new_n19433), .C(new_n8172), .Y(new_n19435));
  A2O1A1O1Ixp25_ASAP7_75t_L g19179(.A1(new_n8490), .A2(new_n6651), .B(new_n19433), .C(new_n19434), .D(new_n19435), .Y(new_n19436));
  INVx1_ASAP7_75t_L         g19180(.A(new_n19429), .Y(new_n19437));
  NAND2xp33_ASAP7_75t_L     g19181(.A(new_n19428), .B(new_n19429), .Y(new_n19438));
  A2O1A1O1Ixp25_ASAP7_75t_L g19182(.A1(new_n19224), .A2(new_n19431), .B(new_n19437), .C(new_n19438), .D(new_n19436), .Y(new_n19439));
  AND2x2_ASAP7_75t_L        g19183(.A(new_n19436), .B(new_n19438), .Y(new_n19440));
  AO221x2_ASAP7_75t_L       g19184(.A1(new_n19237), .A2(new_n19245), .B1(new_n19440), .B2(new_n19430), .C(new_n19439), .Y(new_n19441));
  O2A1O1Ixp33_ASAP7_75t_L   g19185(.A1(new_n19240), .A2(new_n19230), .B(new_n19244), .C(new_n19238), .Y(new_n19442));
  A2O1A1Ixp33_ASAP7_75t_L   g19186(.A1(new_n19440), .A2(new_n19430), .B(new_n19439), .C(new_n19442), .Y(new_n19443));
  NAND2xp33_ASAP7_75t_L     g19187(.A(new_n19443), .B(new_n19441), .Y(new_n19444));
  INVx1_ASAP7_75t_L         g19188(.A(new_n19444), .Y(new_n19445));
  NOR2xp33_ASAP7_75t_L      g19189(.A(new_n6378), .B(new_n7312), .Y(new_n19446));
  AOI221xp5_ASAP7_75t_L     g19190(.A1(\b[41] ), .A2(new_n7609), .B1(\b[43] ), .B2(new_n7334), .C(new_n19446), .Y(new_n19447));
  O2A1O1Ixp33_ASAP7_75t_L   g19191(.A1(new_n7321), .A2(new_n6679), .B(new_n19447), .C(new_n7316), .Y(new_n19448));
  INVx1_ASAP7_75t_L         g19192(.A(new_n19448), .Y(new_n19449));
  O2A1O1Ixp33_ASAP7_75t_L   g19193(.A1(new_n7321), .A2(new_n6679), .B(new_n19447), .C(\a[47] ), .Y(new_n19450));
  A2O1A1Ixp33_ASAP7_75t_L   g19194(.A1(\a[47] ), .A2(new_n19449), .B(new_n19450), .C(new_n19445), .Y(new_n19451));
  NAND2xp33_ASAP7_75t_L     g19195(.A(new_n19445), .B(new_n19451), .Y(new_n19452));
  A2O1A1Ixp33_ASAP7_75t_L   g19196(.A1(\a[47] ), .A2(new_n19449), .B(new_n19450), .C(new_n19444), .Y(new_n19453));
  O2A1O1Ixp33_ASAP7_75t_L   g19197(.A1(new_n19253), .A2(new_n19254), .B(new_n19261), .C(new_n19252), .Y(new_n19454));
  NAND3xp33_ASAP7_75t_L     g19198(.A(new_n19452), .B(new_n19453), .C(new_n19454), .Y(new_n19455));
  INVx1_ASAP7_75t_L         g19199(.A(new_n19451), .Y(new_n19456));
  O2A1O1Ixp33_ASAP7_75t_L   g19200(.A1(new_n19444), .A2(new_n19456), .B(new_n19453), .C(new_n19454), .Y(new_n19457));
  INVx1_ASAP7_75t_L         g19201(.A(new_n19457), .Y(new_n19458));
  NAND2xp33_ASAP7_75t_L     g19202(.A(new_n19455), .B(new_n19458), .Y(new_n19459));
  NOR2xp33_ASAP7_75t_L      g19203(.A(new_n7249), .B(new_n7304), .Y(new_n19460));
  AOI221xp5_ASAP7_75t_L     g19204(.A1(\b[44] ), .A2(new_n6742), .B1(\b[46] ), .B2(new_n6442), .C(new_n19460), .Y(new_n19461));
  O2A1O1Ixp33_ASAP7_75t_L   g19205(.A1(new_n6443), .A2(new_n7279), .B(new_n19461), .C(new_n6439), .Y(new_n19462));
  O2A1O1Ixp33_ASAP7_75t_L   g19206(.A1(new_n6443), .A2(new_n7279), .B(new_n19461), .C(\a[44] ), .Y(new_n19463));
  INVx1_ASAP7_75t_L         g19207(.A(new_n19463), .Y(new_n19464));
  O2A1O1Ixp33_ASAP7_75t_L   g19208(.A1(new_n19462), .A2(new_n6439), .B(new_n19464), .C(new_n19459), .Y(new_n19465));
  INVx1_ASAP7_75t_L         g19209(.A(new_n19462), .Y(new_n19466));
  A2O1A1Ixp33_ASAP7_75t_L   g19210(.A1(\a[44] ), .A2(new_n19466), .B(new_n19463), .C(new_n19459), .Y(new_n19467));
  OAI21xp33_ASAP7_75t_L     g19211(.A1(new_n19459), .A2(new_n19465), .B(new_n19467), .Y(new_n19468));
  NOR3xp33_ASAP7_75t_L      g19212(.A(new_n19468), .B(new_n19274), .C(new_n19269), .Y(new_n19469));
  INVx1_ASAP7_75t_L         g19213(.A(new_n18977), .Y(new_n19470));
  O2A1O1Ixp33_ASAP7_75t_L   g19214(.A1(new_n6439), .A2(new_n18975), .B(new_n19470), .C(new_n19066), .Y(new_n19471));
  O2A1O1Ixp33_ASAP7_75t_L   g19215(.A1(new_n19166), .A2(new_n19471), .B(new_n19271), .C(new_n19269), .Y(new_n19472));
  O2A1O1Ixp33_ASAP7_75t_L   g19216(.A1(new_n19459), .A2(new_n19465), .B(new_n19467), .C(new_n19472), .Y(new_n19473));
  NOR2xp33_ASAP7_75t_L      g19217(.A(new_n19473), .B(new_n19469), .Y(new_n19474));
  NOR2xp33_ASAP7_75t_L      g19218(.A(new_n7860), .B(new_n5640), .Y(new_n19475));
  AOI221xp5_ASAP7_75t_L     g19219(.A1(\b[47] ), .A2(new_n5920), .B1(\b[49] ), .B2(new_n5629), .C(new_n19475), .Y(new_n19476));
  INVx1_ASAP7_75t_L         g19220(.A(new_n19476), .Y(new_n19477));
  A2O1A1Ixp33_ASAP7_75t_L   g19221(.A1(new_n8438), .A2(new_n5637), .B(new_n19477), .C(\a[41] ), .Y(new_n19478));
  O2A1O1Ixp33_ASAP7_75t_L   g19222(.A1(new_n5630), .A2(new_n14802), .B(new_n19476), .C(\a[41] ), .Y(new_n19479));
  A2O1A1Ixp33_ASAP7_75t_L   g19223(.A1(\a[41] ), .A2(new_n19478), .B(new_n19479), .C(new_n19474), .Y(new_n19480));
  NAND2xp33_ASAP7_75t_L     g19224(.A(new_n19474), .B(new_n19480), .Y(new_n19481));
  A2O1A1Ixp33_ASAP7_75t_L   g19225(.A1(new_n19478), .A2(\a[41] ), .B(new_n19479), .C(new_n19480), .Y(new_n19482));
  NAND2xp33_ASAP7_75t_L     g19226(.A(new_n19481), .B(new_n19482), .Y(new_n19483));
  NAND2xp33_ASAP7_75t_L     g19227(.A(\a[41] ), .B(new_n19283), .Y(new_n19484));
  A2O1A1Ixp33_ASAP7_75t_L   g19228(.A1(new_n19484), .A2(new_n19281), .B(new_n19276), .C(new_n19289), .Y(new_n19485));
  NOR2xp33_ASAP7_75t_L      g19229(.A(new_n19485), .B(new_n19483), .Y(new_n19486));
  O2A1O1Ixp33_ASAP7_75t_L   g19230(.A1(new_n5626), .A2(new_n19279), .B(new_n19281), .C(new_n19282), .Y(new_n19487));
  A2O1A1O1Ixp25_ASAP7_75t_L g19231(.A1(new_n19273), .A2(new_n19275), .B(new_n19487), .C(new_n19287), .D(new_n19282), .Y(new_n19488));
  AOI21xp33_ASAP7_75t_L     g19232(.A1(new_n19482), .A2(new_n19481), .B(new_n19488), .Y(new_n19489));
  NOR2xp33_ASAP7_75t_L      g19233(.A(new_n19489), .B(new_n19486), .Y(new_n19490));
  NOR2xp33_ASAP7_75t_L      g19234(.A(new_n8779), .B(new_n4903), .Y(new_n19491));
  AOI221xp5_ASAP7_75t_L     g19235(.A1(\b[50] ), .A2(new_n5139), .B1(\b[52] ), .B2(new_n4917), .C(new_n19491), .Y(new_n19492));
  O2A1O1Ixp33_ASAP7_75t_L   g19236(.A1(new_n4911), .A2(new_n17363), .B(new_n19492), .C(new_n4906), .Y(new_n19493));
  INVx1_ASAP7_75t_L         g19237(.A(new_n19493), .Y(new_n19494));
  O2A1O1Ixp33_ASAP7_75t_L   g19238(.A1(new_n4911), .A2(new_n17363), .B(new_n19492), .C(\a[38] ), .Y(new_n19495));
  A2O1A1Ixp33_ASAP7_75t_L   g19239(.A1(\a[38] ), .A2(new_n19494), .B(new_n19495), .C(new_n19490), .Y(new_n19496));
  INVx1_ASAP7_75t_L         g19240(.A(new_n19495), .Y(new_n19497));
  O2A1O1Ixp33_ASAP7_75t_L   g19241(.A1(new_n19493), .A2(new_n4906), .B(new_n19497), .C(new_n19490), .Y(new_n19498));
  AOI21xp33_ASAP7_75t_L     g19242(.A1(new_n19496), .A2(new_n19490), .B(new_n19498), .Y(new_n19499));
  A2O1A1Ixp33_ASAP7_75t_L   g19243(.A1(new_n19302), .A2(new_n19291), .B(new_n19301), .C(new_n19499), .Y(new_n19500));
  A2O1A1Ixp33_ASAP7_75t_L   g19244(.A1(new_n19496), .A2(new_n19490), .B(new_n19498), .C(new_n19303), .Y(new_n19501));
  NAND2xp33_ASAP7_75t_L     g19245(.A(new_n19501), .B(new_n19500), .Y(new_n19502));
  NOR2xp33_ASAP7_75t_L      g19246(.A(new_n10309), .B(new_n4147), .Y(new_n19503));
  AOI221xp5_ASAP7_75t_L     g19247(.A1(\b[53] ), .A2(new_n4402), .B1(\b[54] ), .B2(new_n4155), .C(new_n19503), .Y(new_n19504));
  O2A1O1Ixp33_ASAP7_75t_L   g19248(.A1(new_n4150), .A2(new_n15849), .B(new_n19504), .C(new_n4145), .Y(new_n19505));
  INVx1_ASAP7_75t_L         g19249(.A(new_n19505), .Y(new_n19506));
  O2A1O1Ixp33_ASAP7_75t_L   g19250(.A1(new_n4150), .A2(new_n15849), .B(new_n19504), .C(\a[35] ), .Y(new_n19507));
  A2O1A1Ixp33_ASAP7_75t_L   g19251(.A1(\a[35] ), .A2(new_n19506), .B(new_n19507), .C(new_n19502), .Y(new_n19508));
  INVx1_ASAP7_75t_L         g19252(.A(new_n19504), .Y(new_n19509));
  NOR2xp33_ASAP7_75t_L      g19253(.A(new_n4145), .B(new_n19505), .Y(new_n19510));
  A2O1A1O1Ixp25_ASAP7_75t_L g19254(.A1(new_n10320), .A2(new_n4151), .B(new_n19509), .C(new_n19506), .D(new_n19510), .Y(new_n19511));
  NAND3xp33_ASAP7_75t_L     g19255(.A(new_n19500), .B(new_n19501), .C(new_n19511), .Y(new_n19512));
  NAND4xp25_ASAP7_75t_L     g19256(.A(new_n19358), .B(new_n19508), .C(new_n19512), .D(new_n19356), .Y(new_n19513));
  AO22x1_ASAP7_75t_L        g19257(.A1(new_n19512), .A2(new_n19508), .B1(new_n19356), .B2(new_n19358), .Y(new_n19514));
  NAND2xp33_ASAP7_75t_L     g19258(.A(new_n19513), .B(new_n19514), .Y(new_n19515));
  O2A1O1Ixp33_ASAP7_75t_L   g19259(.A1(new_n19342), .A2(new_n19343), .B(new_n19348), .C(new_n19515), .Y(new_n19516));
  NAND3xp33_ASAP7_75t_L     g19260(.A(new_n19346), .B(new_n19513), .C(new_n19514), .Y(new_n19517));
  AOI22xp33_ASAP7_75t_L     g19261(.A1(new_n2421), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2577), .Y(new_n19518));
  A2O1A1Ixp33_ASAP7_75t_L   g19262(.A1(new_n12990), .A2(new_n12988), .B(new_n2425), .C(new_n19518), .Y(new_n19519));
  NOR2xp33_ASAP7_75t_L      g19263(.A(new_n2413), .B(new_n19519), .Y(new_n19520));
  O2A1O1Ixp33_ASAP7_75t_L   g19264(.A1(new_n2425), .A2(new_n12993), .B(new_n19518), .C(\a[26] ), .Y(new_n19521));
  NOR2xp33_ASAP7_75t_L      g19265(.A(new_n19521), .B(new_n19520), .Y(new_n19522));
  O2A1O1Ixp33_ASAP7_75t_L   g19266(.A1(new_n19152), .A2(new_n19149), .B(new_n19317), .C(new_n19522), .Y(new_n19523));
  INVx1_ASAP7_75t_L         g19267(.A(new_n19523), .Y(new_n19524));
  INVx1_ASAP7_75t_L         g19268(.A(new_n19522), .Y(new_n19525));
  O2A1O1Ixp33_ASAP7_75t_L   g19269(.A1(new_n19152), .A2(new_n19149), .B(new_n19317), .C(new_n19525), .Y(new_n19526));
  O2A1O1Ixp33_ASAP7_75t_L   g19270(.A1(new_n19520), .A2(new_n19521), .B(new_n19524), .C(new_n19526), .Y(new_n19527));
  O2A1O1Ixp33_ASAP7_75t_L   g19271(.A1(new_n19346), .A2(new_n19516), .B(new_n19517), .C(new_n19527), .Y(new_n19528));
  A2O1A1Ixp33_ASAP7_75t_L   g19272(.A1(new_n19340), .A2(\a[29] ), .B(new_n19341), .C(new_n19344), .Y(new_n19529));
  A2O1A1Ixp33_ASAP7_75t_L   g19273(.A1(new_n19348), .A2(new_n19529), .B(new_n19516), .C(new_n19517), .Y(new_n19530));
  AOI211xp5_ASAP7_75t_L     g19274(.A1(new_n19525), .A2(new_n19524), .B(new_n19526), .C(new_n19530), .Y(new_n19531));
  NOR2xp33_ASAP7_75t_L      g19275(.A(new_n19531), .B(new_n19528), .Y(new_n19532));
  A2O1A1Ixp33_ASAP7_75t_L   g19276(.A1(new_n19129), .A2(new_n19125), .B(new_n19122), .C(new_n19324), .Y(new_n19533));
  O2A1O1Ixp33_ASAP7_75t_L   g19277(.A1(new_n19138), .A2(new_n19142), .B(new_n19334), .C(new_n19319), .Y(new_n19534));
  A2O1A1Ixp33_ASAP7_75t_L   g19278(.A1(new_n19107), .A2(new_n19113), .B(new_n19141), .C(new_n18946), .Y(new_n19535));
  A2O1A1Ixp33_ASAP7_75t_L   g19279(.A1(new_n19139), .A2(new_n19535), .B(new_n19534), .C(new_n19532), .Y(new_n19536));
  NOR3xp33_ASAP7_75t_L      g19280(.A(new_n19528), .B(new_n19531), .C(new_n19335), .Y(new_n19537));
  O2A1O1Ixp33_ASAP7_75t_L   g19281(.A1(new_n19142), .A2(new_n19534), .B(new_n19536), .C(new_n19537), .Y(new_n19538));
  A2O1A1O1Ixp25_ASAP7_75t_L g19282(.A1(new_n19320), .A2(new_n19322), .B(new_n19132), .C(new_n19533), .D(new_n19538), .Y(new_n19539));
  A2O1A1Ixp33_ASAP7_75t_L   g19283(.A1(new_n19320), .A2(new_n19322), .B(new_n19132), .C(new_n19533), .Y(new_n19540));
  NOR2xp33_ASAP7_75t_L      g19284(.A(new_n19537), .B(new_n19540), .Y(new_n19541));
  O2A1O1Ixp33_ASAP7_75t_L   g19285(.A1(new_n19532), .A2(new_n19336), .B(new_n19541), .C(new_n19539), .Y(\f[88] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19286(.A1(new_n19526), .A2(new_n19525), .B(new_n19530), .C(new_n19523), .Y(new_n19543));
  A2O1A1O1Ixp25_ASAP7_75t_L g19287(.A1(new_n19340), .A2(\a[29] ), .B(new_n19341), .C(new_n19347), .D(new_n19516), .Y(new_n19544));
  INVx1_ASAP7_75t_L         g19288(.A(new_n19544), .Y(new_n19545));
  NOR2xp33_ASAP7_75t_L      g19289(.A(new_n12956), .B(new_n2572), .Y(new_n19546));
  A2O1A1Ixp33_ASAP7_75t_L   g19290(.A1(new_n12986), .A2(new_n2417), .B(new_n19546), .C(\a[26] ), .Y(new_n19547));
  A2O1A1Ixp33_ASAP7_75t_L   g19291(.A1(new_n12986), .A2(new_n2417), .B(new_n19546), .C(new_n2413), .Y(new_n19548));
  INVx1_ASAP7_75t_L         g19292(.A(new_n19548), .Y(new_n19549));
  A2O1A1Ixp33_ASAP7_75t_L   g19293(.A1(\a[26] ), .A2(new_n19547), .B(new_n19549), .C(new_n19545), .Y(new_n19550));
  INVx1_ASAP7_75t_L         g19294(.A(new_n19550), .Y(new_n19551));
  A2O1A1Ixp33_ASAP7_75t_L   g19295(.A1(\a[26] ), .A2(new_n19547), .B(new_n19549), .C(new_n19544), .Y(new_n19552));
  NAND2xp33_ASAP7_75t_L     g19296(.A(\b[61] ), .B(new_n2936), .Y(new_n19553));
  OAI221xp5_ASAP7_75t_L     g19297(.A1(new_n2930), .A2(new_n12603), .B1(new_n11626), .B2(new_n3133), .C(new_n19553), .Y(new_n19554));
  A2O1A1Ixp33_ASAP7_75t_L   g19298(.A1(new_n13559), .A2(new_n2932), .B(new_n19554), .C(\a[29] ), .Y(new_n19555));
  NAND2xp33_ASAP7_75t_L     g19299(.A(\a[29] ), .B(new_n19555), .Y(new_n19556));
  A2O1A1Ixp33_ASAP7_75t_L   g19300(.A1(new_n13559), .A2(new_n2932), .B(new_n19554), .C(new_n2928), .Y(new_n19557));
  AND4x1_ASAP7_75t_L        g19301(.A(new_n19513), .B(new_n19356), .C(new_n19557), .D(new_n19556), .Y(new_n19558));
  AOI22xp33_ASAP7_75t_L     g19302(.A1(new_n19556), .A2(new_n19557), .B1(new_n19356), .B2(new_n19513), .Y(new_n19559));
  NOR2xp33_ASAP7_75t_L      g19303(.A(new_n11303), .B(new_n3509), .Y(new_n19560));
  AOI221xp5_ASAP7_75t_L     g19304(.A1(\b[57] ), .A2(new_n3708), .B1(\b[59] ), .B2(new_n3503), .C(new_n19560), .Y(new_n19561));
  O2A1O1Ixp33_ASAP7_75t_L   g19305(.A1(new_n3513), .A2(new_n11597), .B(new_n19561), .C(new_n3493), .Y(new_n19562));
  INVx1_ASAP7_75t_L         g19306(.A(new_n19561), .Y(new_n19563));
  A2O1A1Ixp33_ASAP7_75t_L   g19307(.A1(new_n12577), .A2(new_n3505), .B(new_n19563), .C(new_n3493), .Y(new_n19564));
  OAI21xp33_ASAP7_75t_L     g19308(.A1(new_n3493), .A2(new_n19562), .B(new_n19564), .Y(new_n19565));
  NAND2xp33_ASAP7_75t_L     g19309(.A(new_n19301), .B(new_n19297), .Y(new_n19566));
  A2O1A1Ixp33_ASAP7_75t_L   g19310(.A1(new_n19566), .A2(new_n19297), .B(new_n19499), .C(new_n19508), .Y(new_n19567));
  NOR2xp33_ASAP7_75t_L      g19311(.A(new_n19565), .B(new_n19567), .Y(new_n19568));
  INVx1_ASAP7_75t_L         g19312(.A(new_n19567), .Y(new_n19569));
  O2A1O1Ixp33_ASAP7_75t_L   g19313(.A1(new_n3493), .A2(new_n19562), .B(new_n19564), .C(new_n19569), .Y(new_n19570));
  NOR2xp33_ASAP7_75t_L      g19314(.A(new_n19568), .B(new_n19570), .Y(new_n19571));
  A2O1A1Ixp33_ASAP7_75t_L   g19315(.A1(new_n19482), .A2(new_n19481), .B(new_n19488), .C(new_n19496), .Y(new_n19572));
  NOR2xp33_ASAP7_75t_L      g19316(.A(new_n9683), .B(new_n4908), .Y(new_n19573));
  AOI221xp5_ASAP7_75t_L     g19317(.A1(\b[51] ), .A2(new_n5139), .B1(\b[52] ), .B2(new_n4916), .C(new_n19573), .Y(new_n19574));
  O2A1O1Ixp33_ASAP7_75t_L   g19318(.A1(new_n4911), .A2(new_n9691), .B(new_n19574), .C(new_n4906), .Y(new_n19575));
  INVx1_ASAP7_75t_L         g19319(.A(new_n19575), .Y(new_n19576));
  O2A1O1Ixp33_ASAP7_75t_L   g19320(.A1(new_n4911), .A2(new_n9691), .B(new_n19574), .C(\a[38] ), .Y(new_n19577));
  O2A1O1Ixp33_ASAP7_75t_L   g19321(.A1(new_n19231), .A2(new_n19238), .B(new_n19241), .C(new_n19242), .Y(new_n19578));
  A2O1A1O1Ixp25_ASAP7_75t_L g19322(.A1(new_n19431), .A2(new_n19224), .B(new_n19437), .C(new_n19440), .D(new_n19439), .Y(new_n19579));
  O2A1O1Ixp33_ASAP7_75t_L   g19323(.A1(new_n19238), .A2(new_n19578), .B(new_n19579), .C(new_n19456), .Y(new_n19580));
  NOR2xp33_ASAP7_75t_L      g19324(.A(new_n6944), .B(new_n7318), .Y(new_n19581));
  AOI221xp5_ASAP7_75t_L     g19325(.A1(new_n7333), .A2(\b[43] ), .B1(new_n7609), .B2(\b[42] ), .C(new_n19581), .Y(new_n19582));
  O2A1O1Ixp33_ASAP7_75t_L   g19326(.A1(new_n7321), .A2(new_n6951), .B(new_n19582), .C(new_n7316), .Y(new_n19583));
  INVx1_ASAP7_75t_L         g19327(.A(new_n19583), .Y(new_n19584));
  O2A1O1Ixp33_ASAP7_75t_L   g19328(.A1(new_n7321), .A2(new_n6951), .B(new_n19582), .C(\a[47] ), .Y(new_n19585));
  AOI21xp33_ASAP7_75t_L     g19329(.A1(new_n19584), .A2(\a[47] ), .B(new_n19585), .Y(new_n19586));
  NOR2xp33_ASAP7_75t_L      g19330(.A(new_n4344), .B(new_n10388), .Y(new_n19587));
  AOI221xp5_ASAP7_75t_L     g19331(.A1(new_n10086), .A2(\b[35] ), .B1(new_n11361), .B2(\b[33] ), .C(new_n19587), .Y(new_n19588));
  INVx1_ASAP7_75t_L         g19332(.A(new_n19588), .Y(new_n19589));
  A2O1A1Ixp33_ASAP7_75t_L   g19333(.A1(new_n7773), .A2(new_n10386), .B(new_n19589), .C(\a[56] ), .Y(new_n19590));
  O2A1O1Ixp33_ASAP7_75t_L   g19334(.A1(new_n10088), .A2(new_n4589), .B(new_n19588), .C(\a[56] ), .Y(new_n19591));
  AO21x2_ASAP7_75t_L        g19335(.A1(\a[56] ), .A2(new_n19590), .B(new_n19591), .Y(new_n19592));
  NOR2xp33_ASAP7_75t_L      g19336(.A(new_n3456), .B(new_n11354), .Y(new_n19593));
  AOI221xp5_ASAP7_75t_L     g19337(.A1(\b[32] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[31] ), .C(new_n19593), .Y(new_n19594));
  INVx1_ASAP7_75t_L         g19338(.A(new_n19594), .Y(new_n19595));
  A2O1A1Ixp33_ASAP7_75t_L   g19339(.A1(new_n3900), .A2(new_n11351), .B(new_n19595), .C(\a[59] ), .Y(new_n19596));
  O2A1O1Ixp33_ASAP7_75t_L   g19340(.A1(new_n11053), .A2(new_n3897), .B(new_n19594), .C(\a[59] ), .Y(new_n19597));
  AO21x2_ASAP7_75t_L        g19341(.A1(\a[59] ), .A2(new_n19596), .B(new_n19597), .Y(new_n19598));
  NOR2xp33_ASAP7_75t_L      g19342(.A(new_n2377), .B(new_n13030), .Y(new_n19599));
  O2A1O1Ixp33_ASAP7_75t_L   g19343(.A1(new_n12669), .A2(new_n12671), .B(\b[26] ), .C(new_n19599), .Y(new_n19600));
  A2O1A1Ixp33_ASAP7_75t_L   g19344(.A1(new_n13028), .A2(\b[25] ), .B(new_n19366), .C(new_n19600), .Y(new_n19601));
  A2O1A1Ixp33_ASAP7_75t_L   g19345(.A1(\b[26] ), .A2(new_n13028), .B(new_n19599), .C(new_n19369), .Y(new_n19602));
  NAND2xp33_ASAP7_75t_L     g19346(.A(new_n19602), .B(new_n19601), .Y(new_n19603));
  NAND2xp33_ASAP7_75t_L     g19347(.A(\b[29] ), .B(new_n11995), .Y(new_n19604));
  OAI221xp5_ASAP7_75t_L     g19348(.A1(new_n12318), .A2(new_n3079), .B1(new_n2879), .B2(new_n12320), .C(new_n19604), .Y(new_n19605));
  AOI21xp33_ASAP7_75t_L     g19349(.A1(new_n3873), .A2(new_n11997), .B(new_n19605), .Y(new_n19606));
  NAND2xp33_ASAP7_75t_L     g19350(.A(\a[62] ), .B(new_n19606), .Y(new_n19607));
  A2O1A1Ixp33_ASAP7_75t_L   g19351(.A1(new_n3873), .A2(new_n11997), .B(new_n19605), .C(new_n11987), .Y(new_n19608));
  AOI21xp33_ASAP7_75t_L     g19352(.A1(new_n19607), .A2(new_n19608), .B(new_n19603), .Y(new_n19609));
  INVx1_ASAP7_75t_L         g19353(.A(new_n19609), .Y(new_n19610));
  NAND3xp33_ASAP7_75t_L     g19354(.A(new_n19607), .B(new_n19603), .C(new_n19608), .Y(new_n19611));
  AND2x2_ASAP7_75t_L        g19355(.A(new_n19611), .B(new_n19610), .Y(new_n19612));
  INVx1_ASAP7_75t_L         g19356(.A(new_n19612), .Y(new_n19613));
  O2A1O1Ixp33_ASAP7_75t_L   g19357(.A1(new_n19370), .A2(new_n19367), .B(new_n19382), .C(new_n19613), .Y(new_n19614));
  INVx1_ASAP7_75t_L         g19358(.A(new_n19614), .Y(new_n19615));
  O2A1O1Ixp33_ASAP7_75t_L   g19359(.A1(new_n19378), .A2(new_n19379), .B(new_n19368), .C(new_n19371), .Y(new_n19616));
  NAND2xp33_ASAP7_75t_L     g19360(.A(new_n19616), .B(new_n19613), .Y(new_n19617));
  NAND3xp33_ASAP7_75t_L     g19361(.A(new_n19617), .B(new_n19615), .C(new_n19598), .Y(new_n19618));
  AO21x2_ASAP7_75t_L        g19362(.A1(new_n19617), .A2(new_n19615), .B(new_n19598), .Y(new_n19619));
  AND2x2_ASAP7_75t_L        g19363(.A(new_n19618), .B(new_n19619), .Y(new_n19620));
  INVx1_ASAP7_75t_L         g19364(.A(new_n19620), .Y(new_n19621));
  O2A1O1Ixp33_ASAP7_75t_L   g19365(.A1(new_n19387), .A2(new_n19388), .B(new_n19396), .C(new_n19621), .Y(new_n19622));
  AOI211xp5_ASAP7_75t_L     g19366(.A1(new_n19365), .A2(new_n19384), .B(new_n19403), .C(new_n19620), .Y(new_n19623));
  NOR2xp33_ASAP7_75t_L      g19367(.A(new_n19623), .B(new_n19622), .Y(new_n19624));
  XOR2x2_ASAP7_75t_L        g19368(.A(new_n19592), .B(new_n19624), .Y(new_n19625));
  INVx1_ASAP7_75t_L         g19369(.A(new_n19625), .Y(new_n19626));
  O2A1O1Ixp33_ASAP7_75t_L   g19370(.A1(new_n19400), .A2(new_n19401), .B(new_n19414), .C(new_n19626), .Y(new_n19627));
  INVx1_ASAP7_75t_L         g19371(.A(new_n19627), .Y(new_n19628));
  NAND3xp33_ASAP7_75t_L     g19372(.A(new_n19626), .B(new_n19414), .C(new_n19405), .Y(new_n19629));
  AND2x2_ASAP7_75t_L        g19373(.A(new_n19629), .B(new_n19628), .Y(new_n19630));
  INVx1_ASAP7_75t_L         g19374(.A(new_n19630), .Y(new_n19631));
  NOR2xp33_ASAP7_75t_L      g19375(.A(new_n5074), .B(new_n10400), .Y(new_n19632));
  AOI221xp5_ASAP7_75t_L     g19376(.A1(new_n9102), .A2(\b[38] ), .B1(new_n10398), .B2(\b[36] ), .C(new_n19632), .Y(new_n19633));
  O2A1O1Ixp33_ASAP7_75t_L   g19377(.A1(new_n9104), .A2(new_n5318), .B(new_n19633), .C(new_n9099), .Y(new_n19634));
  O2A1O1Ixp33_ASAP7_75t_L   g19378(.A1(new_n9104), .A2(new_n5318), .B(new_n19633), .C(\a[53] ), .Y(new_n19635));
  INVx1_ASAP7_75t_L         g19379(.A(new_n19635), .Y(new_n19636));
  O2A1O1Ixp33_ASAP7_75t_L   g19380(.A1(new_n19634), .A2(new_n9099), .B(new_n19636), .C(new_n19631), .Y(new_n19637));
  INVx1_ASAP7_75t_L         g19381(.A(new_n19637), .Y(new_n19638));
  O2A1O1Ixp33_ASAP7_75t_L   g19382(.A1(new_n19634), .A2(new_n9099), .B(new_n19636), .C(new_n19630), .Y(new_n19639));
  O2A1O1Ixp33_ASAP7_75t_L   g19383(.A1(new_n9104), .A2(new_n5083), .B(new_n19422), .C(\a[53] ), .Y(new_n19640));
  A2O1A1Ixp33_ASAP7_75t_L   g19384(.A1(\a[53] ), .A2(new_n19425), .B(new_n19640), .C(new_n19420), .Y(new_n19641));
  A2O1A1Ixp33_ASAP7_75t_L   g19385(.A1(new_n19363), .A2(new_n19362), .B(new_n19416), .C(new_n19641), .Y(new_n19642));
  A2O1A1Ixp33_ASAP7_75t_L   g19386(.A1(new_n19638), .A2(new_n19630), .B(new_n19639), .C(new_n19642), .Y(new_n19643));
  AO21x2_ASAP7_75t_L        g19387(.A1(new_n19630), .A2(new_n19638), .B(new_n19639), .Y(new_n19644));
  A2O1A1O1Ixp25_ASAP7_75t_L g19388(.A1(new_n19363), .A2(new_n19362), .B(new_n19416), .C(new_n19641), .D(new_n19644), .Y(new_n19645));
  A2O1A1O1Ixp25_ASAP7_75t_L g19389(.A1(new_n19638), .A2(new_n19630), .B(new_n19639), .C(new_n19643), .D(new_n19645), .Y(new_n19646));
  NOR2xp33_ASAP7_75t_L      g19390(.A(new_n5855), .B(new_n10065), .Y(new_n19647));
  AOI221xp5_ASAP7_75t_L     g19391(.A1(new_n8175), .A2(\b[41] ), .B1(new_n8484), .B2(\b[39] ), .C(new_n19647), .Y(new_n19648));
  O2A1O1Ixp33_ASAP7_75t_L   g19392(.A1(new_n8176), .A2(new_n6117), .B(new_n19648), .C(new_n8172), .Y(new_n19649));
  NOR2xp33_ASAP7_75t_L      g19393(.A(new_n8172), .B(new_n19649), .Y(new_n19650));
  O2A1O1Ixp33_ASAP7_75t_L   g19394(.A1(new_n8176), .A2(new_n6117), .B(new_n19648), .C(\a[50] ), .Y(new_n19651));
  NOR2xp33_ASAP7_75t_L      g19395(.A(new_n19651), .B(new_n19650), .Y(new_n19652));
  XNOR2x2_ASAP7_75t_L       g19396(.A(new_n19652), .B(new_n19646), .Y(new_n19653));
  A2O1A1O1Ixp25_ASAP7_75t_L g19397(.A1(new_n19430), .A2(new_n19438), .B(new_n19436), .C(new_n19429), .D(new_n19653), .Y(new_n19654));
  INVx1_ASAP7_75t_L         g19398(.A(new_n19654), .Y(new_n19655));
  A2O1A1Ixp33_ASAP7_75t_L   g19399(.A1(new_n19430), .A2(new_n19438), .B(new_n19436), .C(new_n19429), .Y(new_n19656));
  INVx1_ASAP7_75t_L         g19400(.A(new_n19656), .Y(new_n19657));
  NAND2xp33_ASAP7_75t_L     g19401(.A(new_n19657), .B(new_n19653), .Y(new_n19658));
  NAND2xp33_ASAP7_75t_L     g19402(.A(new_n19658), .B(new_n19655), .Y(new_n19659));
  XNOR2x2_ASAP7_75t_L       g19403(.A(new_n19586), .B(new_n19659), .Y(new_n19660));
  XOR2x2_ASAP7_75t_L        g19404(.A(new_n19580), .B(new_n19660), .Y(new_n19661));
  NOR2xp33_ASAP7_75t_L      g19405(.A(new_n7249), .B(new_n6741), .Y(new_n19662));
  AOI221xp5_ASAP7_75t_L     g19406(.A1(\b[47] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[46] ), .C(new_n19662), .Y(new_n19663));
  O2A1O1Ixp33_ASAP7_75t_L   g19407(.A1(new_n6443), .A2(new_n7560), .B(new_n19663), .C(new_n6439), .Y(new_n19664));
  INVx1_ASAP7_75t_L         g19408(.A(new_n19664), .Y(new_n19665));
  O2A1O1Ixp33_ASAP7_75t_L   g19409(.A1(new_n6443), .A2(new_n7560), .B(new_n19663), .C(\a[44] ), .Y(new_n19666));
  A2O1A1Ixp33_ASAP7_75t_L   g19410(.A1(\a[44] ), .A2(new_n19665), .B(new_n19666), .C(new_n19661), .Y(new_n19667));
  INVx1_ASAP7_75t_L         g19411(.A(new_n19666), .Y(new_n19668));
  O2A1O1Ixp33_ASAP7_75t_L   g19412(.A1(new_n19664), .A2(new_n6439), .B(new_n19668), .C(new_n19661), .Y(new_n19669));
  AOI21xp33_ASAP7_75t_L     g19413(.A1(new_n19667), .A2(new_n19661), .B(new_n19669), .Y(new_n19670));
  A2O1A1O1Ixp25_ASAP7_75t_L g19414(.A1(new_n19466), .A2(\a[44] ), .B(new_n19463), .C(new_n19455), .D(new_n19457), .Y(new_n19671));
  NAND2xp33_ASAP7_75t_L     g19415(.A(new_n19671), .B(new_n19670), .Y(new_n19672));
  INVx1_ASAP7_75t_L         g19416(.A(new_n19671), .Y(new_n19673));
  A2O1A1Ixp33_ASAP7_75t_L   g19417(.A1(new_n19667), .A2(new_n19661), .B(new_n19669), .C(new_n19673), .Y(new_n19674));
  AND2x2_ASAP7_75t_L        g19418(.A(new_n19674), .B(new_n19672), .Y(new_n19675));
  NOR2xp33_ASAP7_75t_L      g19419(.A(new_n8755), .B(new_n5641), .Y(new_n19676));
  AOI221xp5_ASAP7_75t_L     g19420(.A1(\b[48] ), .A2(new_n5920), .B1(\b[49] ), .B2(new_n5623), .C(new_n19676), .Y(new_n19677));
  O2A1O1Ixp33_ASAP7_75t_L   g19421(.A1(new_n5630), .A2(new_n8764), .B(new_n19677), .C(new_n5626), .Y(new_n19678));
  INVx1_ASAP7_75t_L         g19422(.A(new_n19678), .Y(new_n19679));
  O2A1O1Ixp33_ASAP7_75t_L   g19423(.A1(new_n5630), .A2(new_n8764), .B(new_n19677), .C(\a[41] ), .Y(new_n19680));
  AOI211xp5_ASAP7_75t_L     g19424(.A1(new_n19679), .A2(\a[41] ), .B(new_n19680), .C(new_n19675), .Y(new_n19681));
  A2O1A1Ixp33_ASAP7_75t_L   g19425(.A1(\a[41] ), .A2(new_n19679), .B(new_n19680), .C(new_n19675), .Y(new_n19682));
  INVx1_ASAP7_75t_L         g19426(.A(new_n19682), .Y(new_n19683));
  NOR2xp33_ASAP7_75t_L      g19427(.A(new_n19681), .B(new_n19683), .Y(new_n19684));
  A2O1A1O1Ixp25_ASAP7_75t_L g19428(.A1(new_n19478), .A2(\a[41] ), .B(new_n19479), .C(new_n19474), .D(new_n19473), .Y(new_n19685));
  INVx1_ASAP7_75t_L         g19429(.A(new_n19685), .Y(new_n19686));
  NAND2xp33_ASAP7_75t_L     g19430(.A(new_n19686), .B(new_n19684), .Y(new_n19687));
  INVx1_ASAP7_75t_L         g19431(.A(new_n19468), .Y(new_n19688));
  O2A1O1Ixp33_ASAP7_75t_L   g19432(.A1(new_n19688), .A2(new_n19472), .B(new_n19480), .C(new_n19684), .Y(new_n19689));
  AO21x2_ASAP7_75t_L        g19433(.A1(new_n19684), .A2(new_n19687), .B(new_n19689), .Y(new_n19690));
  AOI21xp33_ASAP7_75t_L     g19434(.A1(new_n19576), .A2(\a[38] ), .B(new_n19577), .Y(new_n19691));
  OAI31xp33_ASAP7_75t_L     g19435(.A1(new_n19681), .A2(new_n19686), .A3(new_n19683), .B(new_n19691), .Y(new_n19692));
  O2A1O1Ixp33_ASAP7_75t_L   g19436(.A1(new_n19681), .A2(new_n19683), .B(new_n19686), .C(new_n19692), .Y(new_n19693));
  A2O1A1O1Ixp25_ASAP7_75t_L g19437(.A1(new_n19576), .A2(\a[38] ), .B(new_n19577), .C(new_n19690), .D(new_n19693), .Y(new_n19694));
  NAND2xp33_ASAP7_75t_L     g19438(.A(new_n19572), .B(new_n19694), .Y(new_n19695));
  INVx1_ASAP7_75t_L         g19439(.A(new_n19695), .Y(new_n19696));
  A2O1A1Ixp33_ASAP7_75t_L   g19440(.A1(new_n19576), .A2(\a[38] ), .B(new_n19577), .C(new_n19690), .Y(new_n19697));
  O2A1O1Ixp33_ASAP7_75t_L   g19441(.A1(new_n19692), .A2(new_n19689), .B(new_n19697), .C(new_n19572), .Y(new_n19698));
  NOR2xp33_ASAP7_75t_L      g19442(.A(new_n19698), .B(new_n19696), .Y(new_n19699));
  NOR2xp33_ASAP7_75t_L      g19443(.A(new_n10332), .B(new_n4147), .Y(new_n19700));
  AOI221xp5_ASAP7_75t_L     g19444(.A1(\b[54] ), .A2(new_n4402), .B1(\b[55] ), .B2(new_n4155), .C(new_n19700), .Y(new_n19701));
  O2A1O1Ixp33_ASAP7_75t_L   g19445(.A1(new_n4150), .A2(new_n10339), .B(new_n19701), .C(new_n4145), .Y(new_n19702));
  O2A1O1Ixp33_ASAP7_75t_L   g19446(.A1(new_n4150), .A2(new_n10339), .B(new_n19701), .C(\a[35] ), .Y(new_n19703));
  INVx1_ASAP7_75t_L         g19447(.A(new_n19703), .Y(new_n19704));
  INVx1_ASAP7_75t_L         g19448(.A(new_n19699), .Y(new_n19705));
  O2A1O1Ixp33_ASAP7_75t_L   g19449(.A1(new_n4145), .A2(new_n19702), .B(new_n19704), .C(new_n19705), .Y(new_n19706));
  INVx1_ASAP7_75t_L         g19450(.A(new_n19706), .Y(new_n19707));
  O2A1O1Ixp33_ASAP7_75t_L   g19451(.A1(new_n4145), .A2(new_n19702), .B(new_n19704), .C(new_n19699), .Y(new_n19708));
  A2O1A1Ixp33_ASAP7_75t_L   g19452(.A1(new_n19699), .A2(new_n19707), .B(new_n19708), .C(new_n19571), .Y(new_n19709));
  NAND2xp33_ASAP7_75t_L     g19453(.A(new_n19571), .B(new_n19709), .Y(new_n19710));
  INVx1_ASAP7_75t_L         g19454(.A(new_n19708), .Y(new_n19711));
  O2A1O1Ixp33_ASAP7_75t_L   g19455(.A1(new_n19705), .A2(new_n19706), .B(new_n19711), .C(new_n19571), .Y(new_n19712));
  INVx1_ASAP7_75t_L         g19456(.A(new_n19712), .Y(new_n19713));
  OAI211xp5_ASAP7_75t_L     g19457(.A1(new_n19559), .A2(new_n19558), .B(new_n19710), .C(new_n19713), .Y(new_n19714));
  NOR2xp33_ASAP7_75t_L      g19458(.A(new_n19559), .B(new_n19558), .Y(new_n19715));
  A2O1A1Ixp33_ASAP7_75t_L   g19459(.A1(new_n19709), .A2(new_n19571), .B(new_n19712), .C(new_n19715), .Y(new_n19716));
  NAND2xp33_ASAP7_75t_L     g19460(.A(new_n19716), .B(new_n19714), .Y(new_n19717));
  O2A1O1Ixp33_ASAP7_75t_L   g19461(.A1(new_n19544), .A2(new_n19551), .B(new_n19552), .C(new_n19717), .Y(new_n19718));
  A2O1A1O1Ixp25_ASAP7_75t_L g19462(.A1(new_n2417), .A2(new_n14172), .B(new_n2577), .C(\b[63] ), .D(new_n2413), .Y(new_n19719));
  A2O1A1O1Ixp25_ASAP7_75t_L g19463(.A1(new_n12986), .A2(new_n2417), .B(new_n19546), .C(new_n19547), .D(new_n19719), .Y(new_n19720));
  INVx1_ASAP7_75t_L         g19464(.A(new_n19720), .Y(new_n19721));
  A2O1A1O1Ixp25_ASAP7_75t_L g19465(.A1(new_n19342), .A2(new_n19348), .B(new_n19515), .C(new_n19344), .D(new_n19721), .Y(new_n19722));
  O2A1O1Ixp33_ASAP7_75t_L   g19466(.A1(new_n19719), .A2(new_n19549), .B(new_n19550), .C(new_n19722), .Y(new_n19723));
  AND2x2_ASAP7_75t_L        g19467(.A(new_n19717), .B(new_n19723), .Y(new_n19724));
  NOR3xp33_ASAP7_75t_L      g19468(.A(new_n19724), .B(new_n19718), .C(new_n19543), .Y(new_n19725));
  INVx1_ASAP7_75t_L         g19469(.A(new_n19725), .Y(new_n19726));
  OAI21xp33_ASAP7_75t_L     g19470(.A1(new_n19718), .A2(new_n19724), .B(new_n19543), .Y(new_n19727));
  AND2x2_ASAP7_75t_L        g19471(.A(new_n19727), .B(new_n19726), .Y(new_n19728));
  INVx1_ASAP7_75t_L         g19472(.A(new_n19728), .Y(new_n19729));
  A2O1A1O1Ixp25_ASAP7_75t_L g19473(.A1(new_n19533), .A2(new_n19327), .B(new_n19538), .C(new_n19536), .D(new_n19729), .Y(new_n19730));
  A2O1A1Ixp33_ASAP7_75t_L   g19474(.A1(new_n19533), .A2(new_n19327), .B(new_n19538), .C(new_n19536), .Y(new_n19731));
  NOR2xp33_ASAP7_75t_L      g19475(.A(new_n19728), .B(new_n19731), .Y(new_n19732));
  NOR2xp33_ASAP7_75t_L      g19476(.A(new_n19732), .B(new_n19730), .Y(\f[89] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19477(.A1(new_n19719), .A2(new_n19549), .B(new_n19545), .C(new_n19718), .Y(new_n19734));
  A2O1A1O1Ixp25_ASAP7_75t_L g19478(.A1(new_n19571), .A2(new_n19709), .B(new_n19712), .C(new_n19715), .D(new_n19559), .Y(new_n19735));
  NAND2xp33_ASAP7_75t_L     g19479(.A(new_n19356), .B(new_n19513), .Y(new_n19736));
  INVx1_ASAP7_75t_L         g19480(.A(new_n19736), .Y(new_n19737));
  NOR2xp33_ASAP7_75t_L      g19481(.A(new_n12956), .B(new_n2930), .Y(new_n19738));
  AOI221xp5_ASAP7_75t_L     g19482(.A1(\b[61] ), .A2(new_n3129), .B1(\b[62] ), .B2(new_n2936), .C(new_n19738), .Y(new_n19739));
  O2A1O1Ixp33_ASAP7_75t_L   g19483(.A1(new_n2940), .A2(new_n17815), .B(new_n19739), .C(new_n2928), .Y(new_n19740));
  INVx1_ASAP7_75t_L         g19484(.A(new_n19740), .Y(new_n19741));
  O2A1O1Ixp33_ASAP7_75t_L   g19485(.A1(new_n2940), .A2(new_n17815), .B(new_n19739), .C(\a[29] ), .Y(new_n19742));
  AOI21xp33_ASAP7_75t_L     g19486(.A1(new_n19741), .A2(\a[29] ), .B(new_n19742), .Y(new_n19743));
  A2O1A1O1Ixp25_ASAP7_75t_L g19487(.A1(new_n19557), .A2(new_n19556), .B(new_n19737), .C(new_n19716), .D(new_n19743), .Y(new_n19744));
  A2O1A1Ixp33_ASAP7_75t_L   g19488(.A1(\a[29] ), .A2(new_n19741), .B(new_n19742), .C(new_n19735), .Y(new_n19745));
  A2O1A1O1Ixp25_ASAP7_75t_L g19489(.A1(new_n19584), .A2(\a[47] ), .B(new_n19585), .C(new_n19658), .D(new_n19654), .Y(new_n19746));
  NOR2xp33_ASAP7_75t_L      g19490(.A(new_n6110), .B(new_n10065), .Y(new_n19747));
  AOI221xp5_ASAP7_75t_L     g19491(.A1(new_n8175), .A2(\b[42] ), .B1(new_n8484), .B2(\b[40] ), .C(new_n19747), .Y(new_n19748));
  O2A1O1Ixp33_ASAP7_75t_L   g19492(.A1(new_n8176), .A2(new_n6386), .B(new_n19748), .C(new_n8172), .Y(new_n19749));
  INVx1_ASAP7_75t_L         g19493(.A(new_n19749), .Y(new_n19750));
  O2A1O1Ixp33_ASAP7_75t_L   g19494(.A1(new_n8176), .A2(new_n6386), .B(new_n19748), .C(\a[50] ), .Y(new_n19751));
  NOR2xp33_ASAP7_75t_L      g19495(.A(new_n3674), .B(new_n11354), .Y(new_n19752));
  AOI221xp5_ASAP7_75t_L     g19496(.A1(\b[33] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[32] ), .C(new_n19752), .Y(new_n19753));
  O2A1O1Ixp33_ASAP7_75t_L   g19497(.A1(new_n11053), .A2(new_n4108), .B(new_n19753), .C(new_n11048), .Y(new_n19754));
  INVx1_ASAP7_75t_L         g19498(.A(new_n19754), .Y(new_n19755));
  O2A1O1Ixp33_ASAP7_75t_L   g19499(.A1(new_n11053), .A2(new_n4108), .B(new_n19753), .C(\a[59] ), .Y(new_n19756));
  AOI21xp33_ASAP7_75t_L     g19500(.A1(new_n19755), .A2(\a[59] ), .B(new_n19756), .Y(new_n19757));
  A2O1A1O1Ixp25_ASAP7_75t_L g19501(.A1(new_n19596), .A2(\a[59] ), .B(new_n19597), .C(new_n19617), .D(new_n19614), .Y(new_n19758));
  NAND2xp33_ASAP7_75t_L     g19502(.A(new_n19757), .B(new_n19758), .Y(new_n19759));
  INVx1_ASAP7_75t_L         g19503(.A(new_n19758), .Y(new_n19760));
  A2O1A1Ixp33_ASAP7_75t_L   g19504(.A1(new_n19755), .A2(\a[59] ), .B(new_n19756), .C(new_n19760), .Y(new_n19761));
  AND2x2_ASAP7_75t_L        g19505(.A(new_n19759), .B(new_n19761), .Y(new_n19762));
  OAI22xp33_ASAP7_75t_L     g19506(.A1(new_n12320), .A2(new_n3079), .B1(new_n3098), .B2(new_n12318), .Y(new_n19763));
  AOI221xp5_ASAP7_75t_L     g19507(.A1(new_n11995), .A2(\b[30] ), .B1(new_n11997), .B2(new_n4813), .C(new_n19763), .Y(new_n19764));
  XNOR2x2_ASAP7_75t_L       g19508(.A(new_n11987), .B(new_n19764), .Y(new_n19765));
  NOR2xp33_ASAP7_75t_L      g19509(.A(new_n2703), .B(new_n13030), .Y(new_n19766));
  A2O1A1Ixp33_ASAP7_75t_L   g19510(.A1(new_n13028), .A2(\b[27] ), .B(new_n19766), .C(new_n2413), .Y(new_n19767));
  INVx1_ASAP7_75t_L         g19511(.A(new_n19767), .Y(new_n19768));
  O2A1O1Ixp33_ASAP7_75t_L   g19512(.A1(new_n12669), .A2(new_n12671), .B(\b[27] ), .C(new_n19766), .Y(new_n19769));
  NAND2xp33_ASAP7_75t_L     g19513(.A(\a[26] ), .B(new_n19769), .Y(new_n19770));
  INVx1_ASAP7_75t_L         g19514(.A(new_n19770), .Y(new_n19771));
  NOR2xp33_ASAP7_75t_L      g19515(.A(new_n19768), .B(new_n19771), .Y(new_n19772));
  A2O1A1Ixp33_ASAP7_75t_L   g19516(.A1(new_n13028), .A2(\b[26] ), .B(new_n19599), .C(new_n19772), .Y(new_n19773));
  OAI21xp33_ASAP7_75t_L     g19517(.A1(new_n19768), .A2(new_n19771), .B(new_n19600), .Y(new_n19774));
  AND2x2_ASAP7_75t_L        g19518(.A(new_n19774), .B(new_n19773), .Y(new_n19775));
  INVx1_ASAP7_75t_L         g19519(.A(new_n19775), .Y(new_n19776));
  A2O1A1O1Ixp25_ASAP7_75t_L g19520(.A1(new_n19608), .A2(new_n19607), .B(new_n19603), .C(new_n19601), .D(new_n19776), .Y(new_n19777));
  INVx1_ASAP7_75t_L         g19521(.A(new_n19777), .Y(new_n19778));
  A2O1A1O1Ixp25_ASAP7_75t_L g19522(.A1(new_n13028), .A2(\b[25] ), .B(new_n19366), .C(new_n19600), .D(new_n19609), .Y(new_n19779));
  NAND2xp33_ASAP7_75t_L     g19523(.A(new_n19776), .B(new_n19779), .Y(new_n19780));
  AND2x2_ASAP7_75t_L        g19524(.A(new_n19778), .B(new_n19780), .Y(new_n19781));
  INVx1_ASAP7_75t_L         g19525(.A(new_n19781), .Y(new_n19782));
  NOR2xp33_ASAP7_75t_L      g19526(.A(new_n19765), .B(new_n19782), .Y(new_n19783));
  NAND2xp33_ASAP7_75t_L     g19527(.A(new_n19765), .B(new_n19781), .Y(new_n19784));
  OA21x2_ASAP7_75t_L        g19528(.A1(new_n19765), .A2(new_n19783), .B(new_n19784), .Y(new_n19785));
  INVx1_ASAP7_75t_L         g19529(.A(new_n19785), .Y(new_n19786));
  NOR2xp33_ASAP7_75t_L      g19530(.A(new_n19786), .B(new_n19762), .Y(new_n19787));
  INVx1_ASAP7_75t_L         g19531(.A(new_n19762), .Y(new_n19788));
  O2A1O1Ixp33_ASAP7_75t_L   g19532(.A1(new_n19765), .A2(new_n19783), .B(new_n19784), .C(new_n19788), .Y(new_n19789));
  NOR2xp33_ASAP7_75t_L      g19533(.A(new_n19787), .B(new_n19789), .Y(new_n19790));
  NOR2xp33_ASAP7_75t_L      g19534(.A(new_n4581), .B(new_n10388), .Y(new_n19791));
  AOI221xp5_ASAP7_75t_L     g19535(.A1(new_n10086), .A2(\b[36] ), .B1(new_n11361), .B2(\b[34] ), .C(new_n19791), .Y(new_n19792));
  O2A1O1Ixp33_ASAP7_75t_L   g19536(.A1(new_n10088), .A2(new_n4622), .B(new_n19792), .C(new_n10083), .Y(new_n19793));
  INVx1_ASAP7_75t_L         g19537(.A(new_n19793), .Y(new_n19794));
  O2A1O1Ixp33_ASAP7_75t_L   g19538(.A1(new_n10088), .A2(new_n4622), .B(new_n19792), .C(\a[56] ), .Y(new_n19795));
  A2O1A1Ixp33_ASAP7_75t_L   g19539(.A1(\a[56] ), .A2(new_n19794), .B(new_n19795), .C(new_n19790), .Y(new_n19796));
  INVx1_ASAP7_75t_L         g19540(.A(new_n19795), .Y(new_n19797));
  O2A1O1Ixp33_ASAP7_75t_L   g19541(.A1(new_n19793), .A2(new_n10083), .B(new_n19797), .C(new_n19790), .Y(new_n19798));
  AO21x2_ASAP7_75t_L        g19542(.A1(new_n19790), .A2(new_n19796), .B(new_n19798), .Y(new_n19799));
  A2O1A1O1Ixp25_ASAP7_75t_L g19543(.A1(new_n19590), .A2(\a[56] ), .B(new_n19591), .C(new_n19624), .D(new_n19622), .Y(new_n19800));
  XNOR2x2_ASAP7_75t_L       g19544(.A(new_n19800), .B(new_n19799), .Y(new_n19801));
  NOR2xp33_ASAP7_75t_L      g19545(.A(new_n5311), .B(new_n10400), .Y(new_n19802));
  AOI221xp5_ASAP7_75t_L     g19546(.A1(new_n9102), .A2(\b[39] ), .B1(new_n10398), .B2(\b[37] ), .C(new_n19802), .Y(new_n19803));
  O2A1O1Ixp33_ASAP7_75t_L   g19547(.A1(new_n9104), .A2(new_n5578), .B(new_n19803), .C(new_n9099), .Y(new_n19804));
  INVx1_ASAP7_75t_L         g19548(.A(new_n19804), .Y(new_n19805));
  O2A1O1Ixp33_ASAP7_75t_L   g19549(.A1(new_n9104), .A2(new_n5578), .B(new_n19803), .C(\a[53] ), .Y(new_n19806));
  A2O1A1Ixp33_ASAP7_75t_L   g19550(.A1(\a[53] ), .A2(new_n19805), .B(new_n19806), .C(new_n19801), .Y(new_n19807));
  INVx1_ASAP7_75t_L         g19551(.A(new_n19806), .Y(new_n19808));
  O2A1O1Ixp33_ASAP7_75t_L   g19552(.A1(new_n19804), .A2(new_n9099), .B(new_n19808), .C(new_n19801), .Y(new_n19809));
  AO21x2_ASAP7_75t_L        g19553(.A1(new_n19801), .A2(new_n19807), .B(new_n19809), .Y(new_n19810));
  OR3x1_ASAP7_75t_L         g19554(.A(new_n19810), .B(new_n19627), .C(new_n19637), .Y(new_n19811));
  A2O1A1Ixp33_ASAP7_75t_L   g19555(.A1(new_n19399), .A2(new_n19397), .B(new_n19401), .C(new_n19414), .Y(new_n19812));
  A2O1A1Ixp33_ASAP7_75t_L   g19556(.A1(new_n19625), .A2(new_n19812), .B(new_n19637), .C(new_n19810), .Y(new_n19813));
  AND2x2_ASAP7_75t_L        g19557(.A(new_n19813), .B(new_n19811), .Y(new_n19814));
  A2O1A1Ixp33_ASAP7_75t_L   g19558(.A1(\a[50] ), .A2(new_n19750), .B(new_n19751), .C(new_n19814), .Y(new_n19815));
  AOI21xp33_ASAP7_75t_L     g19559(.A1(new_n19750), .A2(\a[50] ), .B(new_n19751), .Y(new_n19816));
  AND3x1_ASAP7_75t_L        g19560(.A(new_n19811), .B(new_n19816), .C(new_n19813), .Y(new_n19817));
  A2O1A1O1Ixp25_ASAP7_75t_L g19561(.A1(new_n19750), .A2(\a[50] ), .B(new_n19751), .C(new_n19815), .D(new_n19817), .Y(new_n19818));
  INVx1_ASAP7_75t_L         g19562(.A(new_n19818), .Y(new_n19819));
  O2A1O1Ixp33_ASAP7_75t_L   g19563(.A1(new_n19646), .A2(new_n19652), .B(new_n19643), .C(new_n19819), .Y(new_n19820));
  INVx1_ASAP7_75t_L         g19564(.A(new_n19642), .Y(new_n19821));
  A2O1A1Ixp33_ASAP7_75t_L   g19565(.A1(new_n19638), .A2(new_n19630), .B(new_n19639), .C(new_n19821), .Y(new_n19822));
  A2O1A1Ixp33_ASAP7_75t_L   g19566(.A1(new_n19822), .A2(new_n19821), .B(new_n19652), .C(new_n19643), .Y(new_n19823));
  NOR2xp33_ASAP7_75t_L      g19567(.A(new_n19823), .B(new_n19818), .Y(new_n19824));
  NOR2xp33_ASAP7_75t_L      g19568(.A(new_n19824), .B(new_n19820), .Y(new_n19825));
  INVx1_ASAP7_75t_L         g19569(.A(new_n19825), .Y(new_n19826));
  NOR2xp33_ASAP7_75t_L      g19570(.A(new_n7249), .B(new_n7318), .Y(new_n19827));
  AOI221xp5_ASAP7_75t_L     g19571(.A1(new_n7333), .A2(\b[44] ), .B1(new_n7609), .B2(\b[43] ), .C(new_n19827), .Y(new_n19828));
  O2A1O1Ixp33_ASAP7_75t_L   g19572(.A1(new_n7321), .A2(new_n7255), .B(new_n19828), .C(new_n7316), .Y(new_n19829));
  INVx1_ASAP7_75t_L         g19573(.A(new_n19829), .Y(new_n19830));
  O2A1O1Ixp33_ASAP7_75t_L   g19574(.A1(new_n7321), .A2(new_n7255), .B(new_n19828), .C(\a[47] ), .Y(new_n19831));
  A2O1A1Ixp33_ASAP7_75t_L   g19575(.A1(\a[47] ), .A2(new_n19830), .B(new_n19831), .C(new_n19826), .Y(new_n19832));
  AOI21xp33_ASAP7_75t_L     g19576(.A1(new_n19830), .A2(\a[47] ), .B(new_n19831), .Y(new_n19833));
  NAND2xp33_ASAP7_75t_L     g19577(.A(new_n19833), .B(new_n19825), .Y(new_n19834));
  NAND2xp33_ASAP7_75t_L     g19578(.A(new_n19834), .B(new_n19832), .Y(new_n19835));
  NAND2xp33_ASAP7_75t_L     g19579(.A(new_n19746), .B(new_n19835), .Y(new_n19836));
  O2A1O1Ixp33_ASAP7_75t_L   g19580(.A1(new_n19586), .A2(new_n19659), .B(new_n19655), .C(new_n19835), .Y(new_n19837));
  INVx1_ASAP7_75t_L         g19581(.A(new_n19837), .Y(new_n19838));
  NAND2xp33_ASAP7_75t_L     g19582(.A(new_n19836), .B(new_n19838), .Y(new_n19839));
  INVx1_ASAP7_75t_L         g19583(.A(new_n19839), .Y(new_n19840));
  NOR2xp33_ASAP7_75t_L      g19584(.A(new_n7270), .B(new_n6741), .Y(new_n19841));
  AOI221xp5_ASAP7_75t_L     g19585(.A1(\b[48] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[47] ), .C(new_n19841), .Y(new_n19842));
  O2A1O1Ixp33_ASAP7_75t_L   g19586(.A1(new_n6443), .A2(new_n7868), .B(new_n19842), .C(new_n6439), .Y(new_n19843));
  O2A1O1Ixp33_ASAP7_75t_L   g19587(.A1(new_n6443), .A2(new_n7868), .B(new_n19842), .C(\a[44] ), .Y(new_n19844));
  INVx1_ASAP7_75t_L         g19588(.A(new_n19844), .Y(new_n19845));
  O2A1O1Ixp33_ASAP7_75t_L   g19589(.A1(new_n19843), .A2(new_n6439), .B(new_n19845), .C(new_n19839), .Y(new_n19846));
  INVx1_ASAP7_75t_L         g19590(.A(new_n19846), .Y(new_n19847));
  O2A1O1Ixp33_ASAP7_75t_L   g19591(.A1(new_n19843), .A2(new_n6439), .B(new_n19845), .C(new_n19840), .Y(new_n19848));
  AOI21xp33_ASAP7_75t_L     g19592(.A1(new_n19847), .A2(new_n19840), .B(new_n19848), .Y(new_n19849));
  A2O1A1Ixp33_ASAP7_75t_L   g19593(.A1(new_n19451), .A2(new_n19441), .B(new_n19660), .C(new_n19667), .Y(new_n19850));
  XNOR2x2_ASAP7_75t_L       g19594(.A(new_n19850), .B(new_n19849), .Y(new_n19851));
  NOR2xp33_ASAP7_75t_L      g19595(.A(new_n8779), .B(new_n5641), .Y(new_n19852));
  AOI221xp5_ASAP7_75t_L     g19596(.A1(\b[49] ), .A2(new_n5920), .B1(\b[50] ), .B2(new_n5623), .C(new_n19852), .Y(new_n19853));
  INVx1_ASAP7_75t_L         g19597(.A(new_n19853), .Y(new_n19854));
  O2A1O1Ixp33_ASAP7_75t_L   g19598(.A1(new_n5630), .A2(new_n8789), .B(new_n19853), .C(new_n5626), .Y(new_n19855));
  INVx1_ASAP7_75t_L         g19599(.A(new_n19855), .Y(new_n19856));
  NOR2xp33_ASAP7_75t_L      g19600(.A(new_n5626), .B(new_n19855), .Y(new_n19857));
  A2O1A1O1Ixp25_ASAP7_75t_L g19601(.A1(new_n8790), .A2(new_n5637), .B(new_n19854), .C(new_n19856), .D(new_n19857), .Y(new_n19858));
  INVx1_ASAP7_75t_L         g19602(.A(new_n19858), .Y(new_n19859));
  A2O1A1O1Ixp25_ASAP7_75t_L g19603(.A1(new_n19667), .A2(new_n19661), .B(new_n19669), .C(new_n19673), .D(new_n19683), .Y(new_n19860));
  O2A1O1Ixp33_ASAP7_75t_L   g19604(.A1(new_n5630), .A2(new_n8789), .B(new_n19853), .C(\a[41] ), .Y(new_n19861));
  A2O1A1Ixp33_ASAP7_75t_L   g19605(.A1(\a[41] ), .A2(new_n19856), .B(new_n19861), .C(new_n19851), .Y(new_n19862));
  NOR2xp33_ASAP7_75t_L      g19606(.A(new_n19859), .B(new_n19851), .Y(new_n19863));
  INVx1_ASAP7_75t_L         g19607(.A(new_n19863), .Y(new_n19864));
  AOI21xp33_ASAP7_75t_L     g19608(.A1(new_n19864), .A2(new_n19862), .B(new_n19860), .Y(new_n19865));
  A2O1A1Ixp33_ASAP7_75t_L   g19609(.A1(new_n19674), .A2(new_n19682), .B(new_n19863), .C(new_n19862), .Y(new_n19866));
  INVx1_ASAP7_75t_L         g19610(.A(new_n19866), .Y(new_n19867));
  O2A1O1Ixp33_ASAP7_75t_L   g19611(.A1(new_n19859), .A2(new_n19851), .B(new_n19867), .C(new_n19865), .Y(new_n19868));
  INVx1_ASAP7_75t_L         g19612(.A(new_n19868), .Y(new_n19869));
  NOR2xp33_ASAP7_75t_L      g19613(.A(new_n9709), .B(new_n4908), .Y(new_n19870));
  AOI221xp5_ASAP7_75t_L     g19614(.A1(\b[52] ), .A2(new_n5139), .B1(\b[53] ), .B2(new_n4916), .C(new_n19870), .Y(new_n19871));
  O2A1O1Ixp33_ASAP7_75t_L   g19615(.A1(new_n4911), .A2(new_n9718), .B(new_n19871), .C(new_n4906), .Y(new_n19872));
  O2A1O1Ixp33_ASAP7_75t_L   g19616(.A1(new_n4911), .A2(new_n9718), .B(new_n19871), .C(\a[38] ), .Y(new_n19873));
  INVx1_ASAP7_75t_L         g19617(.A(new_n19873), .Y(new_n19874));
  OAI21xp33_ASAP7_75t_L     g19618(.A1(new_n4906), .A2(new_n19872), .B(new_n19874), .Y(new_n19875));
  NOR2xp33_ASAP7_75t_L      g19619(.A(new_n19875), .B(new_n19869), .Y(new_n19876));
  O2A1O1Ixp33_ASAP7_75t_L   g19620(.A1(new_n19872), .A2(new_n4906), .B(new_n19874), .C(new_n19868), .Y(new_n19877));
  AOI211xp5_ASAP7_75t_L     g19621(.A1(new_n19697), .A2(new_n19687), .B(new_n19877), .C(new_n19876), .Y(new_n19878));
  INVx1_ASAP7_75t_L         g19622(.A(new_n19878), .Y(new_n19879));
  OAI211xp5_ASAP7_75t_L     g19623(.A1(new_n19877), .A2(new_n19876), .B(new_n19697), .C(new_n19687), .Y(new_n19880));
  NAND2xp33_ASAP7_75t_L     g19624(.A(new_n19880), .B(new_n19879), .Y(new_n19881));
  NOR2xp33_ASAP7_75t_L      g19625(.A(new_n10978), .B(new_n4147), .Y(new_n19882));
  AOI221xp5_ASAP7_75t_L     g19626(.A1(\b[55] ), .A2(new_n4402), .B1(\b[56] ), .B2(new_n4155), .C(new_n19882), .Y(new_n19883));
  O2A1O1Ixp33_ASAP7_75t_L   g19627(.A1(new_n4150), .A2(new_n17096), .B(new_n19883), .C(new_n4145), .Y(new_n19884));
  O2A1O1Ixp33_ASAP7_75t_L   g19628(.A1(new_n4150), .A2(new_n17096), .B(new_n19883), .C(\a[35] ), .Y(new_n19885));
  INVx1_ASAP7_75t_L         g19629(.A(new_n19885), .Y(new_n19886));
  O2A1O1Ixp33_ASAP7_75t_L   g19630(.A1(new_n19884), .A2(new_n4145), .B(new_n19886), .C(new_n19881), .Y(new_n19887));
  INVx1_ASAP7_75t_L         g19631(.A(new_n19884), .Y(new_n19888));
  A2O1A1Ixp33_ASAP7_75t_L   g19632(.A1(\a[35] ), .A2(new_n19888), .B(new_n19885), .C(new_n19881), .Y(new_n19889));
  OAI21xp33_ASAP7_75t_L     g19633(.A1(new_n19881), .A2(new_n19887), .B(new_n19889), .Y(new_n19890));
  INVx1_ASAP7_75t_L         g19634(.A(new_n19702), .Y(new_n19891));
  A2O1A1O1Ixp25_ASAP7_75t_L g19635(.A1(new_n19891), .A2(\a[35] ), .B(new_n19703), .C(new_n19699), .D(new_n19696), .Y(new_n19892));
  XOR2x2_ASAP7_75t_L        g19636(.A(new_n19892), .B(new_n19890), .Y(new_n19893));
  OAI22xp33_ASAP7_75t_L     g19637(.A1(new_n3703), .A2(new_n11303), .B1(new_n11591), .B2(new_n3509), .Y(new_n19894));
  AOI221xp5_ASAP7_75t_L     g19638(.A1(new_n3503), .A2(\b[60] ), .B1(new_n3505), .B2(new_n13839), .C(new_n19894), .Y(new_n19895));
  XNOR2x2_ASAP7_75t_L       g19639(.A(new_n3493), .B(new_n19895), .Y(new_n19896));
  A2O1A1O1Ixp25_ASAP7_75t_L g19640(.A1(new_n19707), .A2(new_n19699), .B(new_n19708), .C(new_n19571), .D(new_n19570), .Y(new_n19897));
  XNOR2x2_ASAP7_75t_L       g19641(.A(new_n19896), .B(new_n19897), .Y(new_n19898));
  XNOR2x2_ASAP7_75t_L       g19642(.A(new_n19893), .B(new_n19898), .Y(new_n19899));
  O2A1O1Ixp33_ASAP7_75t_L   g19643(.A1(new_n19735), .A2(new_n19744), .B(new_n19745), .C(new_n19899), .Y(new_n19900));
  INVx1_ASAP7_75t_L         g19644(.A(new_n19900), .Y(new_n19901));
  INVx1_ASAP7_75t_L         g19645(.A(new_n19744), .Y(new_n19902));
  INVx1_ASAP7_75t_L         g19646(.A(new_n19743), .Y(new_n19903));
  A2O1A1O1Ixp25_ASAP7_75t_L g19647(.A1(new_n19557), .A2(new_n19556), .B(new_n19737), .C(new_n19716), .D(new_n19903), .Y(new_n19904));
  A2O1A1O1Ixp25_ASAP7_75t_L g19648(.A1(new_n19741), .A2(\a[29] ), .B(new_n19742), .C(new_n19902), .D(new_n19904), .Y(new_n19905));
  NAND2xp33_ASAP7_75t_L     g19649(.A(new_n19899), .B(new_n19905), .Y(new_n19906));
  NAND2xp33_ASAP7_75t_L     g19650(.A(new_n19906), .B(new_n19901), .Y(new_n19907));
  XOR2x2_ASAP7_75t_L        g19651(.A(new_n19734), .B(new_n19907), .Y(new_n19908));
  A2O1A1Ixp33_ASAP7_75t_L   g19652(.A1(new_n19731), .A2(new_n19728), .B(new_n19725), .C(new_n19908), .Y(new_n19909));
  INVx1_ASAP7_75t_L         g19653(.A(new_n19908), .Y(new_n19910));
  A2O1A1O1Ixp25_ASAP7_75t_L g19654(.A1(new_n19532), .A2(new_n19335), .B(new_n19539), .C(new_n19728), .D(new_n19725), .Y(new_n19911));
  NAND2xp33_ASAP7_75t_L     g19655(.A(new_n19910), .B(new_n19911), .Y(new_n19912));
  AND2x2_ASAP7_75t_L        g19656(.A(new_n19909), .B(new_n19912), .Y(\f[90] ));
  MAJIxp5_ASAP7_75t_L       g19657(.A(new_n19893), .B(new_n19896), .C(new_n19897), .Y(new_n19914));
  AOI22xp33_ASAP7_75t_L     g19658(.A1(new_n2936), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3129), .Y(new_n19915));
  INVx1_ASAP7_75t_L         g19659(.A(new_n19915), .Y(new_n19916));
  A2O1A1Ixp33_ASAP7_75t_L   g19660(.A1(new_n2927), .A2(new_n2929), .B(new_n2739), .C(new_n19915), .Y(new_n19917));
  O2A1O1Ixp33_ASAP7_75t_L   g19661(.A1(new_n19916), .A2(new_n17329), .B(new_n19917), .C(new_n2928), .Y(new_n19918));
  O2A1O1Ixp33_ASAP7_75t_L   g19662(.A1(new_n2940), .A2(new_n12993), .B(new_n19915), .C(\a[29] ), .Y(new_n19919));
  OAI21xp33_ASAP7_75t_L     g19663(.A1(new_n19918), .A2(new_n19919), .B(new_n19914), .Y(new_n19920));
  INVx1_ASAP7_75t_L         g19664(.A(new_n19920), .Y(new_n19921));
  NOR3xp33_ASAP7_75t_L      g19665(.A(new_n19914), .B(new_n19918), .C(new_n19919), .Y(new_n19922));
  NOR2xp33_ASAP7_75t_L      g19666(.A(new_n19922), .B(new_n19921), .Y(new_n19923));
  NOR2xp33_ASAP7_75t_L      g19667(.A(new_n12258), .B(new_n3510), .Y(new_n19924));
  AOI221xp5_ASAP7_75t_L     g19668(.A1(\b[59] ), .A2(new_n3708), .B1(\b[60] ), .B2(new_n3499), .C(new_n19924), .Y(new_n19925));
  O2A1O1Ixp33_ASAP7_75t_L   g19669(.A1(new_n3513), .A2(new_n14764), .B(new_n19925), .C(new_n3493), .Y(new_n19926));
  INVx1_ASAP7_75t_L         g19670(.A(new_n19926), .Y(new_n19927));
  O2A1O1Ixp33_ASAP7_75t_L   g19671(.A1(new_n3513), .A2(new_n14764), .B(new_n19925), .C(\a[32] ), .Y(new_n19928));
  AOI21xp33_ASAP7_75t_L     g19672(.A1(new_n19927), .A2(\a[32] ), .B(new_n19928), .Y(new_n19929));
  O2A1O1Ixp33_ASAP7_75t_L   g19673(.A1(new_n19706), .A2(new_n19696), .B(new_n19890), .C(new_n19887), .Y(new_n19930));
  AND2x2_ASAP7_75t_L        g19674(.A(new_n19929), .B(new_n19930), .Y(new_n19931));
  INVx1_ASAP7_75t_L         g19675(.A(new_n19928), .Y(new_n19932));
  O2A1O1Ixp33_ASAP7_75t_L   g19676(.A1(new_n3493), .A2(new_n19926), .B(new_n19932), .C(new_n19930), .Y(new_n19933));
  NOR2xp33_ASAP7_75t_L      g19677(.A(new_n19933), .B(new_n19931), .Y(new_n19934));
  O2A1O1Ixp33_ASAP7_75t_L   g19678(.A1(new_n19670), .A2(new_n19671), .B(new_n19682), .C(new_n19863), .Y(new_n19935));
  INVx1_ASAP7_75t_L         g19679(.A(new_n19807), .Y(new_n19936));
  O2A1O1Ixp33_ASAP7_75t_L   g19680(.A1(new_n19627), .A2(new_n19637), .B(new_n19810), .C(new_n19936), .Y(new_n19937));
  NAND2xp33_ASAP7_75t_L     g19681(.A(new_n19790), .B(new_n19796), .Y(new_n19938));
  A2O1A1Ixp33_ASAP7_75t_L   g19682(.A1(new_n19794), .A2(\a[56] ), .B(new_n19795), .C(new_n19796), .Y(new_n19939));
  A2O1A1Ixp33_ASAP7_75t_L   g19683(.A1(new_n19939), .A2(new_n19938), .B(new_n19800), .C(new_n19796), .Y(new_n19940));
  A2O1A1O1Ixp25_ASAP7_75t_L g19684(.A1(new_n19755), .A2(\a[59] ), .B(new_n19756), .C(new_n19760), .D(new_n19789), .Y(new_n19941));
  INVx1_ASAP7_75t_L         g19685(.A(new_n19941), .Y(new_n19942));
  NOR2xp33_ASAP7_75t_L      g19686(.A(new_n2879), .B(new_n13030), .Y(new_n19943));
  A2O1A1O1Ixp25_ASAP7_75t_L g19687(.A1(new_n13028), .A2(\b[26] ), .B(new_n19599), .C(new_n19770), .D(new_n19768), .Y(new_n19944));
  A2O1A1Ixp33_ASAP7_75t_L   g19688(.A1(new_n13028), .A2(\b[28] ), .B(new_n19943), .C(new_n19944), .Y(new_n19945));
  O2A1O1Ixp33_ASAP7_75t_L   g19689(.A1(new_n12669), .A2(new_n12671), .B(\b[28] ), .C(new_n19943), .Y(new_n19946));
  INVx1_ASAP7_75t_L         g19690(.A(new_n19946), .Y(new_n19947));
  O2A1O1Ixp33_ASAP7_75t_L   g19691(.A1(new_n19600), .A2(new_n19771), .B(new_n19767), .C(new_n19947), .Y(new_n19948));
  INVx1_ASAP7_75t_L         g19692(.A(new_n19948), .Y(new_n19949));
  NAND2xp33_ASAP7_75t_L     g19693(.A(new_n19945), .B(new_n19949), .Y(new_n19950));
  NOR2xp33_ASAP7_75t_L      g19694(.A(new_n3456), .B(new_n12318), .Y(new_n19951));
  AOI221xp5_ASAP7_75t_L     g19695(.A1(new_n11995), .A2(\b[31] ), .B1(new_n13314), .B2(\b[29] ), .C(new_n19951), .Y(new_n19952));
  O2A1O1Ixp33_ASAP7_75t_L   g19696(.A1(new_n11998), .A2(new_n3681), .B(new_n19952), .C(new_n11987), .Y(new_n19953));
  INVx1_ASAP7_75t_L         g19697(.A(new_n19953), .Y(new_n19954));
  O2A1O1Ixp33_ASAP7_75t_L   g19698(.A1(new_n11998), .A2(new_n3681), .B(new_n19952), .C(\a[62] ), .Y(new_n19955));
  AOI21xp33_ASAP7_75t_L     g19699(.A1(new_n19954), .A2(\a[62] ), .B(new_n19955), .Y(new_n19956));
  NAND2xp33_ASAP7_75t_L     g19700(.A(new_n19950), .B(new_n19956), .Y(new_n19957));
  INVx1_ASAP7_75t_L         g19701(.A(new_n19950), .Y(new_n19958));
  A2O1A1Ixp33_ASAP7_75t_L   g19702(.A1(new_n19954), .A2(\a[62] ), .B(new_n19955), .C(new_n19958), .Y(new_n19959));
  AND2x2_ASAP7_75t_L        g19703(.A(new_n19959), .B(new_n19957), .Y(new_n19960));
  INVx1_ASAP7_75t_L         g19704(.A(new_n19960), .Y(new_n19961));
  O2A1O1Ixp33_ASAP7_75t_L   g19705(.A1(new_n19782), .A2(new_n19765), .B(new_n19778), .C(new_n19961), .Y(new_n19962));
  INVx1_ASAP7_75t_L         g19706(.A(new_n19962), .Y(new_n19963));
  A2O1A1O1Ixp25_ASAP7_75t_L g19707(.A1(new_n19600), .A2(new_n19370), .B(new_n19609), .C(new_n19775), .D(new_n19783), .Y(new_n19964));
  NAND2xp33_ASAP7_75t_L     g19708(.A(new_n19961), .B(new_n19964), .Y(new_n19965));
  AND2x2_ASAP7_75t_L        g19709(.A(new_n19963), .B(new_n19965), .Y(new_n19966));
  INVx1_ASAP7_75t_L         g19710(.A(new_n19966), .Y(new_n19967));
  NOR2xp33_ASAP7_75t_L      g19711(.A(new_n3891), .B(new_n11354), .Y(new_n19968));
  AOI221xp5_ASAP7_75t_L     g19712(.A1(\b[34] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[33] ), .C(new_n19968), .Y(new_n19969));
  O2A1O1Ixp33_ASAP7_75t_L   g19713(.A1(new_n11053), .A2(new_n4352), .B(new_n19969), .C(new_n11048), .Y(new_n19970));
  O2A1O1Ixp33_ASAP7_75t_L   g19714(.A1(new_n11053), .A2(new_n4352), .B(new_n19969), .C(\a[59] ), .Y(new_n19971));
  INVx1_ASAP7_75t_L         g19715(.A(new_n19971), .Y(new_n19972));
  O2A1O1Ixp33_ASAP7_75t_L   g19716(.A1(new_n19970), .A2(new_n11048), .B(new_n19972), .C(new_n19967), .Y(new_n19973));
  O2A1O1Ixp33_ASAP7_75t_L   g19717(.A1(new_n19970), .A2(new_n11048), .B(new_n19972), .C(new_n19966), .Y(new_n19974));
  INVx1_ASAP7_75t_L         g19718(.A(new_n19974), .Y(new_n19975));
  O2A1O1Ixp33_ASAP7_75t_L   g19719(.A1(new_n19967), .A2(new_n19973), .B(new_n19975), .C(new_n19941), .Y(new_n19976));
  INVx1_ASAP7_75t_L         g19720(.A(new_n19976), .Y(new_n19977));
  O2A1O1Ixp33_ASAP7_75t_L   g19721(.A1(new_n19967), .A2(new_n19973), .B(new_n19975), .C(new_n19942), .Y(new_n19978));
  NOR2xp33_ASAP7_75t_L      g19722(.A(new_n4613), .B(new_n10388), .Y(new_n19979));
  AOI221xp5_ASAP7_75t_L     g19723(.A1(new_n10086), .A2(\b[37] ), .B1(new_n11361), .B2(\b[35] ), .C(new_n19979), .Y(new_n19980));
  O2A1O1Ixp33_ASAP7_75t_L   g19724(.A1(new_n10088), .A2(new_n5083), .B(new_n19980), .C(new_n10083), .Y(new_n19981));
  INVx1_ASAP7_75t_L         g19725(.A(new_n19981), .Y(new_n19982));
  O2A1O1Ixp33_ASAP7_75t_L   g19726(.A1(new_n10088), .A2(new_n5083), .B(new_n19980), .C(\a[56] ), .Y(new_n19983));
  AOI21xp33_ASAP7_75t_L     g19727(.A1(new_n19982), .A2(\a[56] ), .B(new_n19983), .Y(new_n19984));
  A2O1A1Ixp33_ASAP7_75t_L   g19728(.A1(new_n19977), .A2(new_n19942), .B(new_n19978), .C(new_n19984), .Y(new_n19985));
  O2A1O1Ixp33_ASAP7_75t_L   g19729(.A1(new_n19616), .A2(new_n19613), .B(new_n19618), .C(new_n19757), .Y(new_n19986));
  O2A1O1Ixp33_ASAP7_75t_L   g19730(.A1(new_n19986), .A2(new_n19789), .B(new_n19977), .C(new_n19978), .Y(new_n19987));
  A2O1A1Ixp33_ASAP7_75t_L   g19731(.A1(\a[56] ), .A2(new_n19982), .B(new_n19983), .C(new_n19987), .Y(new_n19988));
  AND2x2_ASAP7_75t_L        g19732(.A(new_n19985), .B(new_n19988), .Y(new_n19989));
  NAND2xp33_ASAP7_75t_L     g19733(.A(\b[39] ), .B(new_n9096), .Y(new_n19990));
  OAI221xp5_ASAP7_75t_L     g19734(.A1(new_n9440), .A2(new_n5311), .B1(new_n5855), .B2(new_n9439), .C(new_n19990), .Y(new_n19991));
  A2O1A1Ixp33_ASAP7_75t_L   g19735(.A1(new_n6651), .A2(new_n9437), .B(new_n19991), .C(\a[53] ), .Y(new_n19992));
  AOI211xp5_ASAP7_75t_L     g19736(.A1(new_n6651), .A2(new_n9437), .B(new_n19991), .C(new_n9099), .Y(new_n19993));
  A2O1A1O1Ixp25_ASAP7_75t_L g19737(.A1(new_n9437), .A2(new_n6651), .B(new_n19991), .C(new_n19992), .D(new_n19993), .Y(new_n19994));
  A2O1A1O1Ixp25_ASAP7_75t_L g19738(.A1(new_n19939), .A2(new_n19938), .B(new_n19800), .C(new_n19796), .D(new_n19989), .Y(new_n19995));
  NAND2xp33_ASAP7_75t_L     g19739(.A(new_n19940), .B(new_n19989), .Y(new_n19996));
  O2A1O1Ixp33_ASAP7_75t_L   g19740(.A1(new_n19989), .A2(new_n19995), .B(new_n19996), .C(new_n19994), .Y(new_n19997));
  INVx1_ASAP7_75t_L         g19741(.A(new_n19997), .Y(new_n19998));
  A2O1A1Ixp33_ASAP7_75t_L   g19742(.A1(new_n19988), .A2(new_n19985), .B(new_n19940), .C(new_n19994), .Y(new_n19999));
  A2O1A1Ixp33_ASAP7_75t_L   g19743(.A1(new_n19940), .A2(new_n19989), .B(new_n19999), .C(new_n19998), .Y(new_n20000));
  NOR2xp33_ASAP7_75t_L      g19744(.A(new_n19937), .B(new_n20000), .Y(new_n20001));
  INVx1_ASAP7_75t_L         g19745(.A(new_n20001), .Y(new_n20002));
  NAND2xp33_ASAP7_75t_L     g19746(.A(new_n19937), .B(new_n20000), .Y(new_n20003));
  NAND2xp33_ASAP7_75t_L     g19747(.A(new_n20003), .B(new_n20002), .Y(new_n20004));
  INVx1_ASAP7_75t_L         g19748(.A(new_n20004), .Y(new_n20005));
  NOR2xp33_ASAP7_75t_L      g19749(.A(new_n6378), .B(new_n10065), .Y(new_n20006));
  AOI221xp5_ASAP7_75t_L     g19750(.A1(new_n8175), .A2(\b[43] ), .B1(new_n8484), .B2(\b[41] ), .C(new_n20006), .Y(new_n20007));
  INVx1_ASAP7_75t_L         g19751(.A(new_n20007), .Y(new_n20008));
  A2O1A1Ixp33_ASAP7_75t_L   g19752(.A1(new_n6682), .A2(new_n8490), .B(new_n20008), .C(\a[50] ), .Y(new_n20009));
  O2A1O1Ixp33_ASAP7_75t_L   g19753(.A1(new_n8176), .A2(new_n6679), .B(new_n20007), .C(\a[50] ), .Y(new_n20010));
  A2O1A1Ixp33_ASAP7_75t_L   g19754(.A1(\a[50] ), .A2(new_n20009), .B(new_n20010), .C(new_n20005), .Y(new_n20011));
  NAND2xp33_ASAP7_75t_L     g19755(.A(new_n20005), .B(new_n20011), .Y(new_n20012));
  A2O1A1Ixp33_ASAP7_75t_L   g19756(.A1(\a[50] ), .A2(new_n20009), .B(new_n20010), .C(new_n20004), .Y(new_n20013));
  O2A1O1Ixp33_ASAP7_75t_L   g19757(.A1(new_n19646), .A2(new_n19652), .B(new_n19643), .C(new_n19818), .Y(new_n20014));
  A2O1A1O1Ixp25_ASAP7_75t_L g19758(.A1(new_n19750), .A2(\a[50] ), .B(new_n19751), .C(new_n19814), .D(new_n20014), .Y(new_n20015));
  NAND3xp33_ASAP7_75t_L     g19759(.A(new_n20012), .B(new_n20013), .C(new_n20015), .Y(new_n20016));
  AO21x2_ASAP7_75t_L        g19760(.A1(new_n20013), .A2(new_n20012), .B(new_n20015), .Y(new_n20017));
  NAND2xp33_ASAP7_75t_L     g19761(.A(new_n20016), .B(new_n20017), .Y(new_n20018));
  INVx1_ASAP7_75t_L         g19762(.A(new_n20018), .Y(new_n20019));
  NOR2xp33_ASAP7_75t_L      g19763(.A(new_n7249), .B(new_n7312), .Y(new_n20020));
  AOI221xp5_ASAP7_75t_L     g19764(.A1(\b[44] ), .A2(new_n7609), .B1(\b[46] ), .B2(new_n7334), .C(new_n20020), .Y(new_n20021));
  O2A1O1Ixp33_ASAP7_75t_L   g19765(.A1(new_n7321), .A2(new_n7279), .B(new_n20021), .C(new_n7316), .Y(new_n20022));
  O2A1O1Ixp33_ASAP7_75t_L   g19766(.A1(new_n7321), .A2(new_n7279), .B(new_n20021), .C(\a[47] ), .Y(new_n20023));
  INVx1_ASAP7_75t_L         g19767(.A(new_n20023), .Y(new_n20024));
  O2A1O1Ixp33_ASAP7_75t_L   g19768(.A1(new_n20022), .A2(new_n7316), .B(new_n20024), .C(new_n20018), .Y(new_n20025));
  INVx1_ASAP7_75t_L         g19769(.A(new_n20025), .Y(new_n20026));
  NAND2xp33_ASAP7_75t_L     g19770(.A(new_n20019), .B(new_n20026), .Y(new_n20027));
  O2A1O1Ixp33_ASAP7_75t_L   g19771(.A1(new_n20022), .A2(new_n7316), .B(new_n20024), .C(new_n20019), .Y(new_n20028));
  INVx1_ASAP7_75t_L         g19772(.A(new_n20028), .Y(new_n20029));
  A2O1A1O1Ixp25_ASAP7_75t_L g19773(.A1(new_n19830), .A2(\a[47] ), .B(new_n19831), .C(new_n19826), .D(new_n19837), .Y(new_n20030));
  NAND3xp33_ASAP7_75t_L     g19774(.A(new_n20027), .B(new_n20029), .C(new_n20030), .Y(new_n20031));
  O2A1O1Ixp33_ASAP7_75t_L   g19775(.A1(new_n20018), .A2(new_n20025), .B(new_n20029), .C(new_n20030), .Y(new_n20032));
  INVx1_ASAP7_75t_L         g19776(.A(new_n20032), .Y(new_n20033));
  AND2x2_ASAP7_75t_L        g19777(.A(new_n20031), .B(new_n20033), .Y(new_n20034));
  NOR2xp33_ASAP7_75t_L      g19778(.A(new_n7860), .B(new_n7304), .Y(new_n20035));
  AOI221xp5_ASAP7_75t_L     g19779(.A1(\b[47] ), .A2(new_n6742), .B1(\b[49] ), .B2(new_n6442), .C(new_n20035), .Y(new_n20036));
  O2A1O1Ixp33_ASAP7_75t_L   g19780(.A1(new_n6443), .A2(new_n14802), .B(new_n20036), .C(new_n6439), .Y(new_n20037));
  INVx1_ASAP7_75t_L         g19781(.A(new_n20037), .Y(new_n20038));
  O2A1O1Ixp33_ASAP7_75t_L   g19782(.A1(new_n6443), .A2(new_n14802), .B(new_n20036), .C(\a[44] ), .Y(new_n20039));
  A2O1A1Ixp33_ASAP7_75t_L   g19783(.A1(\a[44] ), .A2(new_n20038), .B(new_n20039), .C(new_n20034), .Y(new_n20040));
  INVx1_ASAP7_75t_L         g19784(.A(new_n20039), .Y(new_n20041));
  O2A1O1Ixp33_ASAP7_75t_L   g19785(.A1(new_n20037), .A2(new_n6439), .B(new_n20041), .C(new_n20034), .Y(new_n20042));
  AOI21xp33_ASAP7_75t_L     g19786(.A1(new_n20040), .A2(new_n20034), .B(new_n20042), .Y(new_n20043));
  O2A1O1Ixp33_ASAP7_75t_L   g19787(.A1(new_n19840), .A2(new_n19848), .B(new_n19850), .C(new_n19846), .Y(new_n20044));
  NAND2xp33_ASAP7_75t_L     g19788(.A(new_n20044), .B(new_n20043), .Y(new_n20045));
  INVx1_ASAP7_75t_L         g19789(.A(new_n20044), .Y(new_n20046));
  A2O1A1Ixp33_ASAP7_75t_L   g19790(.A1(new_n20040), .A2(new_n20034), .B(new_n20042), .C(new_n20046), .Y(new_n20047));
  AND2x2_ASAP7_75t_L        g19791(.A(new_n20047), .B(new_n20045), .Y(new_n20048));
  NOR2xp33_ASAP7_75t_L      g19792(.A(new_n8779), .B(new_n5640), .Y(new_n20049));
  AOI221xp5_ASAP7_75t_L     g19793(.A1(\b[50] ), .A2(new_n5920), .B1(\b[52] ), .B2(new_n5629), .C(new_n20049), .Y(new_n20050));
  O2A1O1Ixp33_ASAP7_75t_L   g19794(.A1(new_n5630), .A2(new_n17363), .B(new_n20050), .C(new_n5626), .Y(new_n20051));
  INVx1_ASAP7_75t_L         g19795(.A(new_n20051), .Y(new_n20052));
  O2A1O1Ixp33_ASAP7_75t_L   g19796(.A1(new_n5630), .A2(new_n17363), .B(new_n20050), .C(\a[41] ), .Y(new_n20053));
  A2O1A1Ixp33_ASAP7_75t_L   g19797(.A1(\a[41] ), .A2(new_n20052), .B(new_n20053), .C(new_n20048), .Y(new_n20054));
  INVx1_ASAP7_75t_L         g19798(.A(new_n20053), .Y(new_n20055));
  O2A1O1Ixp33_ASAP7_75t_L   g19799(.A1(new_n20051), .A2(new_n5626), .B(new_n20055), .C(new_n20048), .Y(new_n20056));
  AOI21xp33_ASAP7_75t_L     g19800(.A1(new_n20054), .A2(new_n20048), .B(new_n20056), .Y(new_n20057));
  A2O1A1Ixp33_ASAP7_75t_L   g19801(.A1(new_n19859), .A2(new_n19851), .B(new_n19935), .C(new_n20057), .Y(new_n20058));
  A2O1A1Ixp33_ASAP7_75t_L   g19802(.A1(new_n20054), .A2(new_n20048), .B(new_n20056), .C(new_n19867), .Y(new_n20059));
  NAND2xp33_ASAP7_75t_L     g19803(.A(new_n20059), .B(new_n20058), .Y(new_n20060));
  NOR2xp33_ASAP7_75t_L      g19804(.A(new_n10309), .B(new_n4908), .Y(new_n20061));
  AOI221xp5_ASAP7_75t_L     g19805(.A1(\b[53] ), .A2(new_n5139), .B1(\b[54] ), .B2(new_n4916), .C(new_n20061), .Y(new_n20062));
  O2A1O1Ixp33_ASAP7_75t_L   g19806(.A1(new_n4911), .A2(new_n15849), .B(new_n20062), .C(new_n4906), .Y(new_n20063));
  NOR2xp33_ASAP7_75t_L      g19807(.A(new_n4906), .B(new_n20063), .Y(new_n20064));
  O2A1O1Ixp33_ASAP7_75t_L   g19808(.A1(new_n4911), .A2(new_n15849), .B(new_n20062), .C(\a[38] ), .Y(new_n20065));
  NOR2xp33_ASAP7_75t_L      g19809(.A(new_n20065), .B(new_n20064), .Y(new_n20066));
  XNOR2x2_ASAP7_75t_L       g19810(.A(new_n20066), .B(new_n20060), .Y(new_n20067));
  A2O1A1Ixp33_ASAP7_75t_L   g19811(.A1(new_n19875), .A2(new_n19869), .B(new_n19878), .C(new_n20067), .Y(new_n20068));
  INVx1_ASAP7_75t_L         g19812(.A(new_n20068), .Y(new_n20069));
  NOR3xp33_ASAP7_75t_L      g19813(.A(new_n20067), .B(new_n19878), .C(new_n19877), .Y(new_n20070));
  NOR2xp33_ASAP7_75t_L      g19814(.A(new_n20070), .B(new_n20069), .Y(new_n20071));
  INVx1_ASAP7_75t_L         g19815(.A(new_n20071), .Y(new_n20072));
  INVx1_ASAP7_75t_L         g19816(.A(new_n11314), .Y(new_n20073));
  NOR2xp33_ASAP7_75t_L      g19817(.A(new_n11303), .B(new_n4147), .Y(new_n20074));
  AOI221xp5_ASAP7_75t_L     g19818(.A1(\b[56] ), .A2(new_n4402), .B1(\b[57] ), .B2(new_n4155), .C(new_n20074), .Y(new_n20075));
  O2A1O1Ixp33_ASAP7_75t_L   g19819(.A1(new_n4150), .A2(new_n20073), .B(new_n20075), .C(new_n4145), .Y(new_n20076));
  O2A1O1Ixp33_ASAP7_75t_L   g19820(.A1(new_n4150), .A2(new_n20073), .B(new_n20075), .C(\a[35] ), .Y(new_n20077));
  INVx1_ASAP7_75t_L         g19821(.A(new_n20077), .Y(new_n20078));
  O2A1O1Ixp33_ASAP7_75t_L   g19822(.A1(new_n20076), .A2(new_n4145), .B(new_n20078), .C(new_n20072), .Y(new_n20079));
  INVx1_ASAP7_75t_L         g19823(.A(new_n20079), .Y(new_n20080));
  O2A1O1Ixp33_ASAP7_75t_L   g19824(.A1(new_n20076), .A2(new_n4145), .B(new_n20078), .C(new_n20071), .Y(new_n20081));
  A2O1A1Ixp33_ASAP7_75t_L   g19825(.A1(new_n20071), .A2(new_n20080), .B(new_n20081), .C(new_n19934), .Y(new_n20082));
  INVx1_ASAP7_75t_L         g19826(.A(new_n20081), .Y(new_n20083));
  OAI221xp5_ASAP7_75t_L     g19827(.A1(new_n20079), .A2(new_n20072), .B1(new_n19933), .B2(new_n19931), .C(new_n20083), .Y(new_n20084));
  NAND3xp33_ASAP7_75t_L     g19828(.A(new_n19923), .B(new_n20082), .C(new_n20084), .Y(new_n20085));
  NAND2xp33_ASAP7_75t_L     g19829(.A(new_n19923), .B(new_n20085), .Y(new_n20086));
  NAND3xp33_ASAP7_75t_L     g19830(.A(new_n20085), .B(new_n20084), .C(new_n20082), .Y(new_n20087));
  INVx1_ASAP7_75t_L         g19831(.A(new_n19735), .Y(new_n20088));
  A2O1A1O1Ixp25_ASAP7_75t_L g19832(.A1(new_n19741), .A2(\a[29] ), .B(new_n19742), .C(new_n20088), .D(new_n19900), .Y(new_n20089));
  NAND3xp33_ASAP7_75t_L     g19833(.A(new_n20087), .B(new_n20089), .C(new_n20086), .Y(new_n20090));
  NAND2xp33_ASAP7_75t_L     g19834(.A(new_n20086), .B(new_n20087), .Y(new_n20091));
  A2O1A1Ixp33_ASAP7_75t_L   g19835(.A1(new_n19903), .A2(new_n20088), .B(new_n19900), .C(new_n20091), .Y(new_n20092));
  NAND2xp33_ASAP7_75t_L     g19836(.A(new_n20090), .B(new_n20092), .Y(new_n20093));
  O2A1O1Ixp33_ASAP7_75t_L   g19837(.A1(new_n19734), .A2(new_n19907), .B(new_n19909), .C(new_n20093), .Y(new_n20094));
  O2A1O1Ixp33_ASAP7_75t_L   g19838(.A1(new_n19723), .A2(new_n19717), .B(new_n19550), .C(new_n19907), .Y(new_n20095));
  A2O1A1O1Ixp25_ASAP7_75t_L g19839(.A1(new_n19727), .A2(new_n19731), .B(new_n19725), .C(new_n19908), .D(new_n20095), .Y(new_n20096));
  AND2x2_ASAP7_75t_L        g19840(.A(new_n20093), .B(new_n20096), .Y(new_n20097));
  NOR2xp33_ASAP7_75t_L      g19841(.A(new_n20094), .B(new_n20097), .Y(\f[91] ));
  NAND2xp33_ASAP7_75t_L     g19842(.A(new_n19920), .B(new_n20085), .Y(new_n20099));
  NOR2xp33_ASAP7_75t_L      g19843(.A(new_n12956), .B(new_n3133), .Y(new_n20100));
  A2O1A1Ixp33_ASAP7_75t_L   g19844(.A1(new_n12986), .A2(new_n2932), .B(new_n20100), .C(\a[29] ), .Y(new_n20101));
  A2O1A1O1Ixp25_ASAP7_75t_L g19845(.A1(new_n2932), .A2(new_n14172), .B(new_n3129), .C(\b[63] ), .D(new_n2928), .Y(new_n20102));
  A2O1A1O1Ixp25_ASAP7_75t_L g19846(.A1(new_n12986), .A2(new_n2932), .B(new_n20100), .C(new_n20101), .D(new_n20102), .Y(new_n20103));
  NAND2xp33_ASAP7_75t_L     g19847(.A(\a[32] ), .B(new_n19927), .Y(new_n20104));
  A2O1A1Ixp33_ASAP7_75t_L   g19848(.A1(new_n19932), .A2(new_n20104), .B(new_n19930), .C(new_n20082), .Y(new_n20105));
  A2O1A1Ixp33_ASAP7_75t_L   g19849(.A1(new_n12986), .A2(new_n2932), .B(new_n20100), .C(new_n2928), .Y(new_n20106));
  INVx1_ASAP7_75t_L         g19850(.A(new_n20106), .Y(new_n20107));
  A2O1A1Ixp33_ASAP7_75t_L   g19851(.A1(\a[29] ), .A2(new_n20101), .B(new_n20107), .C(new_n20105), .Y(new_n20108));
  INVx1_ASAP7_75t_L         g19852(.A(new_n20108), .Y(new_n20109));
  INVx1_ASAP7_75t_L         g19853(.A(new_n20076), .Y(new_n20110));
  NAND2xp33_ASAP7_75t_L     g19854(.A(\a[35] ), .B(new_n20110), .Y(new_n20111));
  NAND2xp33_ASAP7_75t_L     g19855(.A(new_n20071), .B(new_n20080), .Y(new_n20112));
  A2O1A1Ixp33_ASAP7_75t_L   g19856(.A1(new_n20078), .A2(new_n20111), .B(new_n20079), .C(new_n20112), .Y(new_n20113));
  A2O1A1Ixp33_ASAP7_75t_L   g19857(.A1(new_n20113), .A2(new_n19934), .B(new_n19933), .C(new_n20103), .Y(new_n20114));
  NOR2xp33_ASAP7_75t_L      g19858(.A(new_n12603), .B(new_n3510), .Y(new_n20115));
  AOI221xp5_ASAP7_75t_L     g19859(.A1(\b[60] ), .A2(new_n3708), .B1(\b[61] ), .B2(new_n3499), .C(new_n20115), .Y(new_n20116));
  O2A1O1Ixp33_ASAP7_75t_L   g19860(.A1(new_n3513), .A2(new_n12610), .B(new_n20116), .C(new_n3493), .Y(new_n20117));
  INVx1_ASAP7_75t_L         g19861(.A(new_n20117), .Y(new_n20118));
  O2A1O1Ixp33_ASAP7_75t_L   g19862(.A1(new_n3513), .A2(new_n12610), .B(new_n20116), .C(\a[32] ), .Y(new_n20119));
  A2O1A1Ixp33_ASAP7_75t_L   g19863(.A1(new_n20111), .A2(new_n20078), .B(new_n20070), .C(new_n20068), .Y(new_n20120));
  AOI211xp5_ASAP7_75t_L     g19864(.A1(\a[32] ), .A2(new_n20118), .B(new_n20119), .C(new_n20120), .Y(new_n20121));
  A2O1A1Ixp33_ASAP7_75t_L   g19865(.A1(new_n20118), .A2(\a[32] ), .B(new_n20119), .C(new_n20120), .Y(new_n20122));
  INVx1_ASAP7_75t_L         g19866(.A(new_n20122), .Y(new_n20123));
  O2A1O1Ixp33_ASAP7_75t_L   g19867(.A1(new_n19860), .A2(new_n19863), .B(new_n19862), .C(new_n20057), .Y(new_n20124));
  INVx1_ASAP7_75t_L         g19868(.A(new_n20124), .Y(new_n20125));
  A2O1A1Ixp33_ASAP7_75t_L   g19869(.A1(new_n20058), .A2(new_n20059), .B(new_n20066), .C(new_n20125), .Y(new_n20126));
  NOR2xp33_ASAP7_75t_L      g19870(.A(new_n10309), .B(new_n4903), .Y(new_n20127));
  AOI221xp5_ASAP7_75t_L     g19871(.A1(\b[54] ), .A2(new_n5139), .B1(\b[56] ), .B2(new_n4917), .C(new_n20127), .Y(new_n20128));
  INVx1_ASAP7_75t_L         g19872(.A(new_n20128), .Y(new_n20129));
  O2A1O1Ixp33_ASAP7_75t_L   g19873(.A1(new_n4911), .A2(new_n10339), .B(new_n20128), .C(new_n4906), .Y(new_n20130));
  INVx1_ASAP7_75t_L         g19874(.A(new_n20130), .Y(new_n20131));
  NOR2xp33_ASAP7_75t_L      g19875(.A(new_n4906), .B(new_n20130), .Y(new_n20132));
  A2O1A1O1Ixp25_ASAP7_75t_L g19876(.A1(new_n11579), .A2(new_n4912), .B(new_n20129), .C(new_n20131), .D(new_n20132), .Y(new_n20133));
  A2O1A1O1Ixp25_ASAP7_75t_L g19877(.A1(new_n20038), .A2(\a[44] ), .B(new_n20039), .C(new_n20031), .D(new_n20032), .Y(new_n20134));
  INVx1_ASAP7_75t_L         g19878(.A(new_n20134), .Y(new_n20135));
  NOR2xp33_ASAP7_75t_L      g19879(.A(new_n6671), .B(new_n10065), .Y(new_n20136));
  AOI221xp5_ASAP7_75t_L     g19880(.A1(new_n8175), .A2(\b[44] ), .B1(new_n8484), .B2(\b[42] ), .C(new_n20136), .Y(new_n20137));
  O2A1O1Ixp33_ASAP7_75t_L   g19881(.A1(new_n8176), .A2(new_n6951), .B(new_n20137), .C(new_n8172), .Y(new_n20138));
  INVx1_ASAP7_75t_L         g19882(.A(new_n20138), .Y(new_n20139));
  O2A1O1Ixp33_ASAP7_75t_L   g19883(.A1(new_n8176), .A2(new_n6951), .B(new_n20137), .C(\a[50] ), .Y(new_n20140));
  INVx1_ASAP7_75t_L         g19884(.A(new_n19940), .Y(new_n20141));
  INVx1_ASAP7_75t_L         g19885(.A(new_n19973), .Y(new_n20142));
  NOR2xp33_ASAP7_75t_L      g19886(.A(new_n4101), .B(new_n11354), .Y(new_n20143));
  AOI221xp5_ASAP7_75t_L     g19887(.A1(\b[35] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[34] ), .C(new_n20143), .Y(new_n20144));
  O2A1O1Ixp33_ASAP7_75t_L   g19888(.A1(new_n11053), .A2(new_n4589), .B(new_n20144), .C(new_n11048), .Y(new_n20145));
  NOR2xp33_ASAP7_75t_L      g19889(.A(new_n11048), .B(new_n20145), .Y(new_n20146));
  O2A1O1Ixp33_ASAP7_75t_L   g19890(.A1(new_n11053), .A2(new_n4589), .B(new_n20144), .C(\a[59] ), .Y(new_n20147));
  NOR2xp33_ASAP7_75t_L      g19891(.A(new_n20147), .B(new_n20146), .Y(new_n20148));
  NOR2xp33_ASAP7_75t_L      g19892(.A(new_n3079), .B(new_n13030), .Y(new_n20149));
  INVx1_ASAP7_75t_L         g19893(.A(new_n20149), .Y(new_n20150));
  O2A1O1Ixp33_ASAP7_75t_L   g19894(.A1(new_n12672), .A2(new_n3098), .B(new_n20150), .C(new_n19947), .Y(new_n20151));
  INVx1_ASAP7_75t_L         g19895(.A(new_n20151), .Y(new_n20152));
  INVx1_ASAP7_75t_L         g19896(.A(new_n19956), .Y(new_n20153));
  O2A1O1Ixp33_ASAP7_75t_L   g19897(.A1(new_n12669), .A2(new_n12671), .B(\b[29] ), .C(new_n20149), .Y(new_n20154));
  A2O1A1Ixp33_ASAP7_75t_L   g19898(.A1(new_n13028), .A2(\b[28] ), .B(new_n19943), .C(new_n20154), .Y(new_n20155));
  A2O1A1Ixp33_ASAP7_75t_L   g19899(.A1(new_n20153), .A2(new_n19945), .B(new_n19948), .C(new_n20155), .Y(new_n20156));
  A2O1A1O1Ixp25_ASAP7_75t_L g19900(.A1(new_n13028), .A2(\b[29] ), .B(new_n20149), .C(new_n19946), .D(new_n20156), .Y(new_n20157));
  O2A1O1Ixp33_ASAP7_75t_L   g19901(.A1(new_n19947), .A2(new_n19944), .B(new_n19959), .C(new_n20157), .Y(new_n20158));
  INVx1_ASAP7_75t_L         g19902(.A(new_n20155), .Y(new_n20159));
  A2O1A1O1Ixp25_ASAP7_75t_L g19903(.A1(new_n19945), .A2(new_n20153), .B(new_n19948), .C(new_n20152), .D(new_n20159), .Y(new_n20160));
  OAI22xp33_ASAP7_75t_L     g19904(.A1(new_n12320), .A2(new_n3456), .B1(new_n3674), .B2(new_n12318), .Y(new_n20161));
  AOI221xp5_ASAP7_75t_L     g19905(.A1(new_n11995), .A2(\b[32] ), .B1(new_n11997), .B2(new_n3900), .C(new_n20161), .Y(new_n20162));
  XNOR2x2_ASAP7_75t_L       g19906(.A(new_n11987), .B(new_n20162), .Y(new_n20163));
  A2O1A1Ixp33_ASAP7_75t_L   g19907(.A1(new_n20160), .A2(new_n20152), .B(new_n20158), .C(new_n20163), .Y(new_n20164));
  O2A1O1Ixp33_ASAP7_75t_L   g19908(.A1(new_n20154), .A2(new_n19947), .B(new_n20160), .C(new_n20158), .Y(new_n20165));
  INVx1_ASAP7_75t_L         g19909(.A(new_n20163), .Y(new_n20166));
  NAND2xp33_ASAP7_75t_L     g19910(.A(new_n20166), .B(new_n20165), .Y(new_n20167));
  AND2x2_ASAP7_75t_L        g19911(.A(new_n20164), .B(new_n20167), .Y(new_n20168));
  XOR2x2_ASAP7_75t_L        g19912(.A(new_n20148), .B(new_n20168), .Y(new_n20169));
  INVx1_ASAP7_75t_L         g19913(.A(new_n20169), .Y(new_n20170));
  O2A1O1Ixp33_ASAP7_75t_L   g19914(.A1(new_n19961), .A2(new_n19964), .B(new_n20142), .C(new_n20170), .Y(new_n20171));
  INVx1_ASAP7_75t_L         g19915(.A(new_n20171), .Y(new_n20172));
  INVx1_ASAP7_75t_L         g19916(.A(new_n19970), .Y(new_n20173));
  A2O1A1O1Ixp25_ASAP7_75t_L g19917(.A1(new_n20173), .A2(\a[59] ), .B(new_n19971), .C(new_n19965), .D(new_n19962), .Y(new_n20174));
  NAND2xp33_ASAP7_75t_L     g19918(.A(new_n20174), .B(new_n20170), .Y(new_n20175));
  AND2x2_ASAP7_75t_L        g19919(.A(new_n20175), .B(new_n20172), .Y(new_n20176));
  INVx1_ASAP7_75t_L         g19920(.A(new_n20176), .Y(new_n20177));
  NOR2xp33_ASAP7_75t_L      g19921(.A(new_n5074), .B(new_n10388), .Y(new_n20178));
  AOI221xp5_ASAP7_75t_L     g19922(.A1(new_n10086), .A2(\b[38] ), .B1(new_n11361), .B2(\b[36] ), .C(new_n20178), .Y(new_n20179));
  O2A1O1Ixp33_ASAP7_75t_L   g19923(.A1(new_n10088), .A2(new_n5318), .B(new_n20179), .C(new_n10083), .Y(new_n20180));
  O2A1O1Ixp33_ASAP7_75t_L   g19924(.A1(new_n10088), .A2(new_n5318), .B(new_n20179), .C(\a[56] ), .Y(new_n20181));
  INVx1_ASAP7_75t_L         g19925(.A(new_n20181), .Y(new_n20182));
  O2A1O1Ixp33_ASAP7_75t_L   g19926(.A1(new_n20180), .A2(new_n10083), .B(new_n20182), .C(new_n20177), .Y(new_n20183));
  INVx1_ASAP7_75t_L         g19927(.A(new_n20183), .Y(new_n20184));
  O2A1O1Ixp33_ASAP7_75t_L   g19928(.A1(new_n20180), .A2(new_n10083), .B(new_n20182), .C(new_n20176), .Y(new_n20185));
  AOI21xp33_ASAP7_75t_L     g19929(.A1(new_n20184), .A2(new_n20176), .B(new_n20185), .Y(new_n20186));
  INVx1_ASAP7_75t_L         g19930(.A(new_n20186), .Y(new_n20187));
  O2A1O1Ixp33_ASAP7_75t_L   g19931(.A1(new_n19987), .A2(new_n19984), .B(new_n19977), .C(new_n20186), .Y(new_n20188));
  INVx1_ASAP7_75t_L         g19932(.A(new_n20188), .Y(new_n20189));
  O2A1O1Ixp33_ASAP7_75t_L   g19933(.A1(new_n19987), .A2(new_n19984), .B(new_n19977), .C(new_n20187), .Y(new_n20190));
  NOR2xp33_ASAP7_75t_L      g19934(.A(new_n5855), .B(new_n10400), .Y(new_n20191));
  AOI221xp5_ASAP7_75t_L     g19935(.A1(new_n9102), .A2(\b[41] ), .B1(new_n10398), .B2(\b[39] ), .C(new_n20191), .Y(new_n20192));
  O2A1O1Ixp33_ASAP7_75t_L   g19936(.A1(new_n9104), .A2(new_n6117), .B(new_n20192), .C(new_n9099), .Y(new_n20193));
  INVx1_ASAP7_75t_L         g19937(.A(new_n20193), .Y(new_n20194));
  O2A1O1Ixp33_ASAP7_75t_L   g19938(.A1(new_n9104), .A2(new_n6117), .B(new_n20192), .C(\a[53] ), .Y(new_n20195));
  AOI21xp33_ASAP7_75t_L     g19939(.A1(new_n20194), .A2(\a[53] ), .B(new_n20195), .Y(new_n20196));
  A2O1A1Ixp33_ASAP7_75t_L   g19940(.A1(new_n20189), .A2(new_n20187), .B(new_n20190), .C(new_n20196), .Y(new_n20197));
  A2O1A1O1Ixp25_ASAP7_75t_L g19941(.A1(new_n20184), .A2(new_n20176), .B(new_n20185), .C(new_n20189), .D(new_n20190), .Y(new_n20198));
  A2O1A1Ixp33_ASAP7_75t_L   g19942(.A1(\a[53] ), .A2(new_n20194), .B(new_n20195), .C(new_n20198), .Y(new_n20199));
  NAND2xp33_ASAP7_75t_L     g19943(.A(new_n20197), .B(new_n20199), .Y(new_n20200));
  INVx1_ASAP7_75t_L         g19944(.A(new_n20200), .Y(new_n20201));
  O2A1O1Ixp33_ASAP7_75t_L   g19945(.A1(new_n20141), .A2(new_n19989), .B(new_n19998), .C(new_n20201), .Y(new_n20202));
  INVx1_ASAP7_75t_L         g19946(.A(new_n20202), .Y(new_n20203));
  OR3x1_ASAP7_75t_L         g19947(.A(new_n20200), .B(new_n19995), .C(new_n19997), .Y(new_n20204));
  NAND2xp33_ASAP7_75t_L     g19948(.A(new_n20204), .B(new_n20203), .Y(new_n20205));
  INVx1_ASAP7_75t_L         g19949(.A(new_n20205), .Y(new_n20206));
  A2O1A1Ixp33_ASAP7_75t_L   g19950(.A1(new_n20139), .A2(\a[50] ), .B(new_n20140), .C(new_n20206), .Y(new_n20207));
  AOI21xp33_ASAP7_75t_L     g19951(.A1(new_n20139), .A2(\a[50] ), .B(new_n20140), .Y(new_n20208));
  NAND2xp33_ASAP7_75t_L     g19952(.A(new_n20208), .B(new_n20205), .Y(new_n20209));
  NAND2xp33_ASAP7_75t_L     g19953(.A(new_n20209), .B(new_n20207), .Y(new_n20210));
  O2A1O1Ixp33_ASAP7_75t_L   g19954(.A1(new_n19937), .A2(new_n20000), .B(new_n20011), .C(new_n20210), .Y(new_n20211));
  INVx1_ASAP7_75t_L         g19955(.A(new_n20211), .Y(new_n20212));
  A2O1A1O1Ixp25_ASAP7_75t_L g19956(.A1(new_n20009), .A2(\a[50] ), .B(new_n20010), .C(new_n20003), .D(new_n20001), .Y(new_n20213));
  NAND2xp33_ASAP7_75t_L     g19957(.A(new_n20213), .B(new_n20210), .Y(new_n20214));
  AND2x2_ASAP7_75t_L        g19958(.A(new_n20214), .B(new_n20212), .Y(new_n20215));
  NOR2xp33_ASAP7_75t_L      g19959(.A(new_n7552), .B(new_n7318), .Y(new_n20216));
  AOI221xp5_ASAP7_75t_L     g19960(.A1(new_n7333), .A2(\b[46] ), .B1(new_n7609), .B2(\b[45] ), .C(new_n20216), .Y(new_n20217));
  O2A1O1Ixp33_ASAP7_75t_L   g19961(.A1(new_n7321), .A2(new_n7560), .B(new_n20217), .C(new_n7316), .Y(new_n20218));
  INVx1_ASAP7_75t_L         g19962(.A(new_n20218), .Y(new_n20219));
  O2A1O1Ixp33_ASAP7_75t_L   g19963(.A1(new_n7321), .A2(new_n7560), .B(new_n20217), .C(\a[47] ), .Y(new_n20220));
  A2O1A1Ixp33_ASAP7_75t_L   g19964(.A1(\a[47] ), .A2(new_n20219), .B(new_n20220), .C(new_n20215), .Y(new_n20221));
  INVx1_ASAP7_75t_L         g19965(.A(new_n20220), .Y(new_n20222));
  O2A1O1Ixp33_ASAP7_75t_L   g19966(.A1(new_n20218), .A2(new_n7316), .B(new_n20222), .C(new_n20215), .Y(new_n20223));
  AOI21xp33_ASAP7_75t_L     g19967(.A1(new_n20221), .A2(new_n20215), .B(new_n20223), .Y(new_n20224));
  A2O1A1Ixp33_ASAP7_75t_L   g19968(.A1(new_n20013), .A2(new_n20012), .B(new_n20015), .C(new_n20026), .Y(new_n20225));
  INVx1_ASAP7_75t_L         g19969(.A(new_n20225), .Y(new_n20226));
  NAND2xp33_ASAP7_75t_L     g19970(.A(new_n20226), .B(new_n20224), .Y(new_n20227));
  A2O1A1Ixp33_ASAP7_75t_L   g19971(.A1(new_n20221), .A2(new_n20215), .B(new_n20223), .C(new_n20225), .Y(new_n20228));
  NAND2xp33_ASAP7_75t_L     g19972(.A(new_n20228), .B(new_n20227), .Y(new_n20229));
  NOR2xp33_ASAP7_75t_L      g19973(.A(new_n7860), .B(new_n6741), .Y(new_n20230));
  AOI221xp5_ASAP7_75t_L     g19974(.A1(\b[50] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[49] ), .C(new_n20230), .Y(new_n20231));
  O2A1O1Ixp33_ASAP7_75t_L   g19975(.A1(new_n6443), .A2(new_n8764), .B(new_n20231), .C(new_n6439), .Y(new_n20232));
  O2A1O1Ixp33_ASAP7_75t_L   g19976(.A1(new_n6443), .A2(new_n8764), .B(new_n20231), .C(\a[44] ), .Y(new_n20233));
  INVx1_ASAP7_75t_L         g19977(.A(new_n20233), .Y(new_n20234));
  OAI21xp33_ASAP7_75t_L     g19978(.A1(new_n6439), .A2(new_n20232), .B(new_n20234), .Y(new_n20235));
  XNOR2x2_ASAP7_75t_L       g19979(.A(new_n20235), .B(new_n20229), .Y(new_n20236));
  NAND2xp33_ASAP7_75t_L     g19980(.A(new_n20135), .B(new_n20236), .Y(new_n20237));
  NOR2xp33_ASAP7_75t_L      g19981(.A(new_n9683), .B(new_n5641), .Y(new_n20238));
  AOI221xp5_ASAP7_75t_L     g19982(.A1(\b[51] ), .A2(new_n5920), .B1(\b[52] ), .B2(new_n5623), .C(new_n20238), .Y(new_n20239));
  O2A1O1Ixp33_ASAP7_75t_L   g19983(.A1(new_n5630), .A2(new_n9691), .B(new_n20239), .C(new_n5626), .Y(new_n20240));
  INVx1_ASAP7_75t_L         g19984(.A(new_n20240), .Y(new_n20241));
  O2A1O1Ixp33_ASAP7_75t_L   g19985(.A1(new_n5630), .A2(new_n9691), .B(new_n20239), .C(\a[41] ), .Y(new_n20242));
  AND2x2_ASAP7_75t_L        g19986(.A(new_n20135), .B(new_n20236), .Y(new_n20243));
  NAND2xp33_ASAP7_75t_L     g19987(.A(new_n20134), .B(new_n20236), .Y(new_n20244));
  A2O1A1Ixp33_ASAP7_75t_L   g19988(.A1(new_n20040), .A2(new_n20033), .B(new_n20243), .C(new_n20244), .Y(new_n20245));
  A2O1A1Ixp33_ASAP7_75t_L   g19989(.A1(new_n20241), .A2(\a[41] ), .B(new_n20242), .C(new_n20245), .Y(new_n20246));
  AOI21xp33_ASAP7_75t_L     g19990(.A1(new_n20241), .A2(\a[41] ), .B(new_n20242), .Y(new_n20247));
  NAND2xp33_ASAP7_75t_L     g19991(.A(new_n20247), .B(new_n20244), .Y(new_n20248));
  A2O1A1Ixp33_ASAP7_75t_L   g19992(.A1(new_n20135), .A2(new_n20237), .B(new_n20248), .C(new_n20246), .Y(new_n20249));
  O2A1O1Ixp33_ASAP7_75t_L   g19993(.A1(new_n20043), .A2(new_n20044), .B(new_n20054), .C(new_n20249), .Y(new_n20250));
  O2A1O1Ixp33_ASAP7_75t_L   g19994(.A1(new_n19580), .A2(new_n19660), .B(new_n19667), .C(new_n19849), .Y(new_n20251));
  INVx1_ASAP7_75t_L         g19995(.A(new_n20251), .Y(new_n20252));
  A2O1A1Ixp33_ASAP7_75t_L   g19996(.A1(new_n20252), .A2(new_n19847), .B(new_n20043), .C(new_n20054), .Y(new_n20253));
  A2O1A1O1Ixp25_ASAP7_75t_L g19997(.A1(new_n20029), .A2(new_n20027), .B(new_n20030), .C(new_n20040), .D(new_n20236), .Y(new_n20254));
  O2A1O1Ixp33_ASAP7_75t_L   g19998(.A1(new_n20248), .A2(new_n20254), .B(new_n20246), .C(new_n20253), .Y(new_n20255));
  NOR2xp33_ASAP7_75t_L      g19999(.A(new_n20255), .B(new_n20250), .Y(new_n20256));
  XNOR2x2_ASAP7_75t_L       g20000(.A(new_n20133), .B(new_n20256), .Y(new_n20257));
  XNOR2x2_ASAP7_75t_L       g20001(.A(new_n20126), .B(new_n20257), .Y(new_n20258));
  NOR2xp33_ASAP7_75t_L      g20002(.A(new_n11303), .B(new_n4142), .Y(new_n20259));
  AOI221xp5_ASAP7_75t_L     g20003(.A1(\b[57] ), .A2(new_n4402), .B1(\b[59] ), .B2(new_n4156), .C(new_n20259), .Y(new_n20260));
  O2A1O1Ixp33_ASAP7_75t_L   g20004(.A1(new_n4150), .A2(new_n11597), .B(new_n20260), .C(new_n4145), .Y(new_n20261));
  O2A1O1Ixp33_ASAP7_75t_L   g20005(.A1(new_n4150), .A2(new_n11597), .B(new_n20260), .C(\a[35] ), .Y(new_n20262));
  INVx1_ASAP7_75t_L         g20006(.A(new_n20262), .Y(new_n20263));
  O2A1O1Ixp33_ASAP7_75t_L   g20007(.A1(new_n20261), .A2(new_n4145), .B(new_n20263), .C(new_n20258), .Y(new_n20264));
  INVx1_ASAP7_75t_L         g20008(.A(new_n20261), .Y(new_n20265));
  A2O1A1Ixp33_ASAP7_75t_L   g20009(.A1(\a[35] ), .A2(new_n20265), .B(new_n20262), .C(new_n20258), .Y(new_n20266));
  OAI221xp5_ASAP7_75t_L     g20010(.A1(new_n20121), .A2(new_n20123), .B1(new_n20258), .B2(new_n20264), .C(new_n20266), .Y(new_n20267));
  INVx1_ASAP7_75t_L         g20011(.A(new_n20121), .Y(new_n20268));
  OAI21xp33_ASAP7_75t_L     g20012(.A1(new_n20258), .A2(new_n20264), .B(new_n20266), .Y(new_n20269));
  NAND3xp33_ASAP7_75t_L     g20013(.A(new_n20269), .B(new_n20122), .C(new_n20268), .Y(new_n20270));
  NAND2xp33_ASAP7_75t_L     g20014(.A(new_n20267), .B(new_n20270), .Y(new_n20271));
  O2A1O1Ixp33_ASAP7_75t_L   g20015(.A1(new_n20103), .A2(new_n20109), .B(new_n20114), .C(new_n20271), .Y(new_n20272));
  A2O1A1Ixp33_ASAP7_75t_L   g20016(.A1(new_n20101), .A2(\a[29] ), .B(new_n20107), .C(new_n20108), .Y(new_n20273));
  NAND3xp33_ASAP7_75t_L     g20017(.A(new_n20273), .B(new_n20114), .C(new_n20271), .Y(new_n20274));
  INVx1_ASAP7_75t_L         g20018(.A(new_n20274), .Y(new_n20275));
  NOR2xp33_ASAP7_75t_L      g20019(.A(new_n20272), .B(new_n20275), .Y(new_n20276));
  NAND2xp33_ASAP7_75t_L     g20020(.A(new_n20099), .B(new_n20276), .Y(new_n20277));
  INVx1_ASAP7_75t_L         g20021(.A(new_n20277), .Y(new_n20278));
  INVx1_ASAP7_75t_L         g20022(.A(new_n19907), .Y(new_n20279));
  A2O1A1Ixp33_ASAP7_75t_L   g20023(.A1(new_n19721), .A2(new_n19545), .B(new_n19718), .C(new_n20279), .Y(new_n20280));
  A2O1A1Ixp33_ASAP7_75t_L   g20024(.A1(new_n19909), .A2(new_n20280), .B(new_n20093), .C(new_n20092), .Y(new_n20281));
  INVx1_ASAP7_75t_L         g20025(.A(new_n20281), .Y(new_n20282));
  NAND2xp33_ASAP7_75t_L     g20026(.A(new_n20276), .B(new_n20277), .Y(new_n20283));
  A2O1A1O1Ixp25_ASAP7_75t_L g20027(.A1(new_n19920), .A2(new_n20085), .B(new_n20278), .C(new_n20283), .D(new_n20282), .Y(new_n20284));
  AOI21xp33_ASAP7_75t_L     g20028(.A1(new_n20277), .A2(new_n20276), .B(new_n20281), .Y(new_n20285));
  A2O1A1O1Ixp25_ASAP7_75t_L g20029(.A1(new_n20085), .A2(new_n19920), .B(new_n20278), .C(new_n20285), .D(new_n20284), .Y(\f[92] ));
  NAND2xp33_ASAP7_75t_L     g20030(.A(new_n20099), .B(new_n20277), .Y(new_n20287));
  NAND2xp33_ASAP7_75t_L     g20031(.A(new_n20283), .B(new_n20287), .Y(new_n20288));
  O2A1O1Ixp33_ASAP7_75t_L   g20032(.A1(new_n20102), .A2(new_n20107), .B(new_n20105), .C(new_n20272), .Y(new_n20289));
  A2O1A1Ixp33_ASAP7_75t_L   g20033(.A1(new_n20244), .A2(new_n20134), .B(new_n20247), .C(new_n20237), .Y(new_n20290));
  O2A1O1Ixp33_ASAP7_75t_L   g20034(.A1(new_n20232), .A2(new_n6439), .B(new_n20234), .C(new_n20229), .Y(new_n20291));
  INVx1_ASAP7_75t_L         g20035(.A(new_n20291), .Y(new_n20292));
  A2O1A1Ixp33_ASAP7_75t_L   g20036(.A1(new_n20026), .A2(new_n20017), .B(new_n20224), .C(new_n20292), .Y(new_n20293));
  A2O1A1O1Ixp25_ASAP7_75t_L g20037(.A1(new_n20139), .A2(\a[50] ), .B(new_n20140), .C(new_n20204), .D(new_n20202), .Y(new_n20294));
  INVx1_ASAP7_75t_L         g20038(.A(new_n19978), .Y(new_n20295));
  O2A1O1Ixp33_ASAP7_75t_L   g20039(.A1(new_n19941), .A2(new_n19976), .B(new_n20295), .C(new_n19984), .Y(new_n20296));
  A2O1A1O1Ixp25_ASAP7_75t_L g20040(.A1(new_n20142), .A2(new_n19966), .B(new_n19974), .C(new_n19942), .D(new_n20296), .Y(new_n20297));
  INVx1_ASAP7_75t_L         g20041(.A(new_n20297), .Y(new_n20298));
  A2O1A1Ixp33_ASAP7_75t_L   g20042(.A1(new_n20184), .A2(new_n20176), .B(new_n20185), .C(new_n20297), .Y(new_n20299));
  O2A1O1Ixp33_ASAP7_75t_L   g20043(.A1(new_n20297), .A2(new_n20188), .B(new_n20299), .C(new_n20196), .Y(new_n20300));
  A2O1A1Ixp33_ASAP7_75t_L   g20044(.A1(new_n20160), .A2(new_n20152), .B(new_n20158), .C(new_n20166), .Y(new_n20301));
  NOR2xp33_ASAP7_75t_L      g20045(.A(new_n3098), .B(new_n13030), .Y(new_n20302));
  A2O1A1Ixp33_ASAP7_75t_L   g20046(.A1(new_n13028), .A2(\b[30] ), .B(new_n20302), .C(new_n2928), .Y(new_n20303));
  O2A1O1Ixp33_ASAP7_75t_L   g20047(.A1(new_n12669), .A2(new_n12671), .B(\b[30] ), .C(new_n20302), .Y(new_n20304));
  NAND2xp33_ASAP7_75t_L     g20048(.A(\a[29] ), .B(new_n20304), .Y(new_n20305));
  NAND2xp33_ASAP7_75t_L     g20049(.A(new_n20303), .B(new_n20305), .Y(new_n20306));
  INVx1_ASAP7_75t_L         g20050(.A(new_n20306), .Y(new_n20307));
  O2A1O1Ixp33_ASAP7_75t_L   g20051(.A1(new_n3098), .A2(new_n12672), .B(new_n20150), .C(new_n20306), .Y(new_n20308));
  INVx1_ASAP7_75t_L         g20052(.A(new_n20308), .Y(new_n20309));
  O2A1O1Ixp33_ASAP7_75t_L   g20053(.A1(new_n3098), .A2(new_n12672), .B(new_n20150), .C(new_n20307), .Y(new_n20310));
  A2O1A1Ixp33_ASAP7_75t_L   g20054(.A1(new_n19773), .A2(new_n19767), .B(new_n19947), .C(new_n19959), .Y(new_n20311));
  AO21x2_ASAP7_75t_L        g20055(.A1(new_n20307), .A2(new_n20309), .B(new_n20310), .Y(new_n20312));
  A2O1A1Ixp33_ASAP7_75t_L   g20056(.A1(new_n20311), .A2(new_n20152), .B(new_n20159), .C(new_n20312), .Y(new_n20313));
  A2O1A1O1Ixp25_ASAP7_75t_L g20057(.A1(new_n19949), .A2(new_n19959), .B(new_n20151), .C(new_n20155), .D(new_n20312), .Y(new_n20314));
  A2O1A1O1Ixp25_ASAP7_75t_L g20058(.A1(new_n20309), .A2(new_n20307), .B(new_n20310), .C(new_n20313), .D(new_n20314), .Y(new_n20315));
  NAND2xp33_ASAP7_75t_L     g20059(.A(\b[33] ), .B(new_n11995), .Y(new_n20316));
  OAI221xp5_ASAP7_75t_L     g20060(.A1(new_n12318), .A2(new_n3891), .B1(new_n3674), .B2(new_n12320), .C(new_n20316), .Y(new_n20317));
  A2O1A1Ixp33_ASAP7_75t_L   g20061(.A1(new_n4831), .A2(new_n11997), .B(new_n20317), .C(\a[62] ), .Y(new_n20318));
  NAND2xp33_ASAP7_75t_L     g20062(.A(\a[62] ), .B(new_n20318), .Y(new_n20319));
  A2O1A1Ixp33_ASAP7_75t_L   g20063(.A1(new_n4831), .A2(new_n11997), .B(new_n20317), .C(new_n11987), .Y(new_n20320));
  NAND2xp33_ASAP7_75t_L     g20064(.A(new_n20320), .B(new_n20319), .Y(new_n20321));
  XOR2x2_ASAP7_75t_L        g20065(.A(new_n20321), .B(new_n20315), .Y(new_n20322));
  NOR2xp33_ASAP7_75t_L      g20066(.A(new_n4344), .B(new_n11354), .Y(new_n20323));
  AOI221xp5_ASAP7_75t_L     g20067(.A1(\b[36] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[35] ), .C(new_n20323), .Y(new_n20324));
  O2A1O1Ixp33_ASAP7_75t_L   g20068(.A1(new_n11053), .A2(new_n4622), .B(new_n20324), .C(new_n11048), .Y(new_n20325));
  O2A1O1Ixp33_ASAP7_75t_L   g20069(.A1(new_n11053), .A2(new_n4622), .B(new_n20324), .C(\a[59] ), .Y(new_n20326));
  INVx1_ASAP7_75t_L         g20070(.A(new_n20326), .Y(new_n20327));
  O2A1O1Ixp33_ASAP7_75t_L   g20071(.A1(new_n20325), .A2(new_n11048), .B(new_n20327), .C(new_n20322), .Y(new_n20328));
  INVx1_ASAP7_75t_L         g20072(.A(new_n20328), .Y(new_n20329));
  OAI211xp5_ASAP7_75t_L     g20073(.A1(new_n11048), .A2(new_n20325), .B(new_n20322), .C(new_n20327), .Y(new_n20330));
  AND2x2_ASAP7_75t_L        g20074(.A(new_n20330), .B(new_n20329), .Y(new_n20331));
  INVx1_ASAP7_75t_L         g20075(.A(new_n20331), .Y(new_n20332));
  O2A1O1Ixp33_ASAP7_75t_L   g20076(.A1(new_n20148), .A2(new_n20168), .B(new_n20301), .C(new_n20332), .Y(new_n20333));
  A2O1A1Ixp33_ASAP7_75t_L   g20077(.A1(new_n20167), .A2(new_n20164), .B(new_n20148), .C(new_n20301), .Y(new_n20334));
  NOR2xp33_ASAP7_75t_L      g20078(.A(new_n20334), .B(new_n20331), .Y(new_n20335));
  NOR2xp33_ASAP7_75t_L      g20079(.A(new_n20335), .B(new_n20333), .Y(new_n20336));
  NOR2xp33_ASAP7_75t_L      g20080(.A(new_n5311), .B(new_n10388), .Y(new_n20337));
  AOI221xp5_ASAP7_75t_L     g20081(.A1(new_n10086), .A2(\b[39] ), .B1(new_n11361), .B2(\b[37] ), .C(new_n20337), .Y(new_n20338));
  O2A1O1Ixp33_ASAP7_75t_L   g20082(.A1(new_n10088), .A2(new_n5578), .B(new_n20338), .C(new_n10083), .Y(new_n20339));
  INVx1_ASAP7_75t_L         g20083(.A(new_n20339), .Y(new_n20340));
  O2A1O1Ixp33_ASAP7_75t_L   g20084(.A1(new_n10088), .A2(new_n5578), .B(new_n20338), .C(\a[56] ), .Y(new_n20341));
  A2O1A1Ixp33_ASAP7_75t_L   g20085(.A1(\a[56] ), .A2(new_n20340), .B(new_n20341), .C(new_n20336), .Y(new_n20342));
  INVx1_ASAP7_75t_L         g20086(.A(new_n20341), .Y(new_n20343));
  O2A1O1Ixp33_ASAP7_75t_L   g20087(.A1(new_n20339), .A2(new_n10083), .B(new_n20343), .C(new_n20336), .Y(new_n20344));
  AOI21xp33_ASAP7_75t_L     g20088(.A1(new_n20342), .A2(new_n20336), .B(new_n20344), .Y(new_n20345));
  O2A1O1Ixp33_ASAP7_75t_L   g20089(.A1(new_n19962), .A2(new_n19973), .B(new_n20169), .C(new_n20183), .Y(new_n20346));
  NAND2xp33_ASAP7_75t_L     g20090(.A(new_n20345), .B(new_n20346), .Y(new_n20347));
  INVx1_ASAP7_75t_L         g20091(.A(new_n20174), .Y(new_n20348));
  INVx1_ASAP7_75t_L         g20092(.A(new_n20345), .Y(new_n20349));
  A2O1A1Ixp33_ASAP7_75t_L   g20093(.A1(new_n20169), .A2(new_n20348), .B(new_n20183), .C(new_n20349), .Y(new_n20350));
  AND2x2_ASAP7_75t_L        g20094(.A(new_n20350), .B(new_n20347), .Y(new_n20351));
  NOR2xp33_ASAP7_75t_L      g20095(.A(new_n6110), .B(new_n10400), .Y(new_n20352));
  AOI221xp5_ASAP7_75t_L     g20096(.A1(new_n9102), .A2(\b[42] ), .B1(new_n10398), .B2(\b[40] ), .C(new_n20352), .Y(new_n20353));
  O2A1O1Ixp33_ASAP7_75t_L   g20097(.A1(new_n9104), .A2(new_n6386), .B(new_n20353), .C(new_n9099), .Y(new_n20354));
  INVx1_ASAP7_75t_L         g20098(.A(new_n20354), .Y(new_n20355));
  O2A1O1Ixp33_ASAP7_75t_L   g20099(.A1(new_n9104), .A2(new_n6386), .B(new_n20353), .C(\a[53] ), .Y(new_n20356));
  A2O1A1Ixp33_ASAP7_75t_L   g20100(.A1(\a[53] ), .A2(new_n20355), .B(new_n20356), .C(new_n20351), .Y(new_n20357));
  INVx1_ASAP7_75t_L         g20101(.A(new_n20356), .Y(new_n20358));
  O2A1O1Ixp33_ASAP7_75t_L   g20102(.A1(new_n20354), .A2(new_n9099), .B(new_n20358), .C(new_n20351), .Y(new_n20359));
  AOI21xp33_ASAP7_75t_L     g20103(.A1(new_n20357), .A2(new_n20351), .B(new_n20359), .Y(new_n20360));
  A2O1A1Ixp33_ASAP7_75t_L   g20104(.A1(new_n20298), .A2(new_n20187), .B(new_n20300), .C(new_n20360), .Y(new_n20361));
  O2A1O1Ixp33_ASAP7_75t_L   g20105(.A1(new_n19976), .A2(new_n20296), .B(new_n20187), .C(new_n20300), .Y(new_n20362));
  A2O1A1Ixp33_ASAP7_75t_L   g20106(.A1(new_n20351), .A2(new_n20357), .B(new_n20359), .C(new_n20362), .Y(new_n20363));
  AND2x2_ASAP7_75t_L        g20107(.A(new_n20363), .B(new_n20361), .Y(new_n20364));
  INVx1_ASAP7_75t_L         g20108(.A(new_n20364), .Y(new_n20365));
  NOR2xp33_ASAP7_75t_L      g20109(.A(new_n6944), .B(new_n10065), .Y(new_n20366));
  AOI221xp5_ASAP7_75t_L     g20110(.A1(new_n8175), .A2(\b[45] ), .B1(new_n8484), .B2(\b[43] ), .C(new_n20366), .Y(new_n20367));
  O2A1O1Ixp33_ASAP7_75t_L   g20111(.A1(new_n8176), .A2(new_n7255), .B(new_n20367), .C(new_n8172), .Y(new_n20368));
  INVx1_ASAP7_75t_L         g20112(.A(new_n20368), .Y(new_n20369));
  O2A1O1Ixp33_ASAP7_75t_L   g20113(.A1(new_n8176), .A2(new_n7255), .B(new_n20367), .C(\a[50] ), .Y(new_n20370));
  A2O1A1Ixp33_ASAP7_75t_L   g20114(.A1(\a[50] ), .A2(new_n20369), .B(new_n20370), .C(new_n20365), .Y(new_n20371));
  AOI21xp33_ASAP7_75t_L     g20115(.A1(new_n20369), .A2(\a[50] ), .B(new_n20370), .Y(new_n20372));
  NAND2xp33_ASAP7_75t_L     g20116(.A(new_n20372), .B(new_n20364), .Y(new_n20373));
  AND2x2_ASAP7_75t_L        g20117(.A(new_n20373), .B(new_n20371), .Y(new_n20374));
  INVx1_ASAP7_75t_L         g20118(.A(new_n20374), .Y(new_n20375));
  NAND2xp33_ASAP7_75t_L     g20119(.A(new_n20294), .B(new_n20375), .Y(new_n20376));
  O2A1O1Ixp33_ASAP7_75t_L   g20120(.A1(new_n20208), .A2(new_n20205), .B(new_n20203), .C(new_n20375), .Y(new_n20377));
  INVx1_ASAP7_75t_L         g20121(.A(new_n20377), .Y(new_n20378));
  AND2x2_ASAP7_75t_L        g20122(.A(new_n20376), .B(new_n20378), .Y(new_n20379));
  INVx1_ASAP7_75t_L         g20123(.A(new_n20379), .Y(new_n20380));
  NOR2xp33_ASAP7_75t_L      g20124(.A(new_n7860), .B(new_n7318), .Y(new_n20381));
  AOI221xp5_ASAP7_75t_L     g20125(.A1(new_n7333), .A2(\b[47] ), .B1(new_n7609), .B2(\b[46] ), .C(new_n20381), .Y(new_n20382));
  O2A1O1Ixp33_ASAP7_75t_L   g20126(.A1(new_n7321), .A2(new_n7868), .B(new_n20382), .C(new_n7316), .Y(new_n20383));
  O2A1O1Ixp33_ASAP7_75t_L   g20127(.A1(new_n7321), .A2(new_n7868), .B(new_n20382), .C(\a[47] ), .Y(new_n20384));
  INVx1_ASAP7_75t_L         g20128(.A(new_n20384), .Y(new_n20385));
  O2A1O1Ixp33_ASAP7_75t_L   g20129(.A1(new_n20383), .A2(new_n7316), .B(new_n20385), .C(new_n20380), .Y(new_n20386));
  INVx1_ASAP7_75t_L         g20130(.A(new_n20386), .Y(new_n20387));
  O2A1O1Ixp33_ASAP7_75t_L   g20131(.A1(new_n20383), .A2(new_n7316), .B(new_n20385), .C(new_n20379), .Y(new_n20388));
  AOI21xp33_ASAP7_75t_L     g20132(.A1(new_n20387), .A2(new_n20379), .B(new_n20388), .Y(new_n20389));
  A2O1A1O1Ixp25_ASAP7_75t_L g20133(.A1(new_n20219), .A2(\a[47] ), .B(new_n20220), .C(new_n20214), .D(new_n20211), .Y(new_n20390));
  AND2x2_ASAP7_75t_L        g20134(.A(new_n20390), .B(new_n20389), .Y(new_n20391));
  O2A1O1Ixp33_ASAP7_75t_L   g20135(.A1(new_n20213), .A2(new_n20210), .B(new_n20221), .C(new_n20389), .Y(new_n20392));
  NOR2xp33_ASAP7_75t_L      g20136(.A(new_n20392), .B(new_n20391), .Y(new_n20393));
  NOR2xp33_ASAP7_75t_L      g20137(.A(new_n8427), .B(new_n6741), .Y(new_n20394));
  AOI221xp5_ASAP7_75t_L     g20138(.A1(\b[51] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[50] ), .C(new_n20394), .Y(new_n20395));
  O2A1O1Ixp33_ASAP7_75t_L   g20139(.A1(new_n6443), .A2(new_n8789), .B(new_n20395), .C(new_n6439), .Y(new_n20396));
  INVx1_ASAP7_75t_L         g20140(.A(new_n20396), .Y(new_n20397));
  O2A1O1Ixp33_ASAP7_75t_L   g20141(.A1(new_n6443), .A2(new_n8789), .B(new_n20395), .C(\a[44] ), .Y(new_n20398));
  A2O1A1Ixp33_ASAP7_75t_L   g20142(.A1(\a[44] ), .A2(new_n20397), .B(new_n20398), .C(new_n20393), .Y(new_n20399));
  AOI21xp33_ASAP7_75t_L     g20143(.A1(new_n20397), .A2(\a[44] ), .B(new_n20398), .Y(new_n20400));
  INVx1_ASAP7_75t_L         g20144(.A(new_n20400), .Y(new_n20401));
  NOR2xp33_ASAP7_75t_L      g20145(.A(new_n20401), .B(new_n20393), .Y(new_n20402));
  O2A1O1Ixp33_ASAP7_75t_L   g20146(.A1(new_n20224), .A2(new_n20226), .B(new_n20292), .C(new_n20402), .Y(new_n20403));
  NAND2xp33_ASAP7_75t_L     g20147(.A(new_n20399), .B(new_n20403), .Y(new_n20404));
  A2O1A1Ixp33_ASAP7_75t_L   g20148(.A1(new_n20292), .A2(new_n20228), .B(new_n20402), .C(new_n20399), .Y(new_n20405));
  O2A1O1Ixp33_ASAP7_75t_L   g20149(.A1(new_n20391), .A2(new_n20392), .B(new_n20400), .C(new_n20405), .Y(new_n20406));
  NOR2xp33_ASAP7_75t_L      g20150(.A(new_n9709), .B(new_n5641), .Y(new_n20407));
  AOI221xp5_ASAP7_75t_L     g20151(.A1(\b[52] ), .A2(new_n5920), .B1(\b[53] ), .B2(new_n5623), .C(new_n20407), .Y(new_n20408));
  O2A1O1Ixp33_ASAP7_75t_L   g20152(.A1(new_n5630), .A2(new_n9718), .B(new_n20408), .C(new_n5626), .Y(new_n20409));
  O2A1O1Ixp33_ASAP7_75t_L   g20153(.A1(new_n5630), .A2(new_n9718), .B(new_n20408), .C(\a[41] ), .Y(new_n20410));
  INVx1_ASAP7_75t_L         g20154(.A(new_n20410), .Y(new_n20411));
  OAI21xp33_ASAP7_75t_L     g20155(.A1(new_n5626), .A2(new_n20409), .B(new_n20411), .Y(new_n20412));
  AOI211xp5_ASAP7_75t_L     g20156(.A1(new_n20404), .A2(new_n20293), .B(new_n20412), .C(new_n20406), .Y(new_n20413));
  INVx1_ASAP7_75t_L         g20157(.A(new_n20228), .Y(new_n20414));
  O2A1O1Ixp33_ASAP7_75t_L   g20158(.A1(new_n20414), .A2(new_n20291), .B(new_n20404), .C(new_n20406), .Y(new_n20415));
  O2A1O1Ixp33_ASAP7_75t_L   g20159(.A1(new_n20409), .A2(new_n5626), .B(new_n20411), .C(new_n20415), .Y(new_n20416));
  NOR2xp33_ASAP7_75t_L      g20160(.A(new_n20413), .B(new_n20416), .Y(new_n20417));
  XNOR2x2_ASAP7_75t_L       g20161(.A(new_n20290), .B(new_n20417), .Y(new_n20418));
  NOR2xp33_ASAP7_75t_L      g20162(.A(new_n10332), .B(new_n4903), .Y(new_n20419));
  AOI221xp5_ASAP7_75t_L     g20163(.A1(\b[55] ), .A2(new_n5139), .B1(\b[57] ), .B2(new_n4917), .C(new_n20419), .Y(new_n20420));
  O2A1O1Ixp33_ASAP7_75t_L   g20164(.A1(new_n4911), .A2(new_n17096), .B(new_n20420), .C(new_n4906), .Y(new_n20421));
  O2A1O1Ixp33_ASAP7_75t_L   g20165(.A1(new_n4911), .A2(new_n17096), .B(new_n20420), .C(\a[38] ), .Y(new_n20422));
  INVx1_ASAP7_75t_L         g20166(.A(new_n20422), .Y(new_n20423));
  O2A1O1Ixp33_ASAP7_75t_L   g20167(.A1(new_n20421), .A2(new_n4906), .B(new_n20423), .C(new_n20418), .Y(new_n20424));
  INVx1_ASAP7_75t_L         g20168(.A(new_n20418), .Y(new_n20425));
  O2A1O1Ixp33_ASAP7_75t_L   g20169(.A1(new_n20421), .A2(new_n4906), .B(new_n20423), .C(new_n20425), .Y(new_n20426));
  INVx1_ASAP7_75t_L         g20170(.A(new_n20426), .Y(new_n20427));
  O2A1O1Ixp33_ASAP7_75t_L   g20171(.A1(new_n4911), .A2(new_n10339), .B(new_n20128), .C(\a[38] ), .Y(new_n20428));
  O2A1O1Ixp33_ASAP7_75t_L   g20172(.A1(new_n20428), .A2(new_n20132), .B(new_n20256), .C(new_n20250), .Y(new_n20429));
  OAI211xp5_ASAP7_75t_L     g20173(.A1(new_n20418), .A2(new_n20424), .B(new_n20427), .C(new_n20429), .Y(new_n20430));
  INVx1_ASAP7_75t_L         g20174(.A(new_n20424), .Y(new_n20431));
  INVx1_ASAP7_75t_L         g20175(.A(new_n20429), .Y(new_n20432));
  A2O1A1Ixp33_ASAP7_75t_L   g20176(.A1(new_n20431), .A2(new_n20425), .B(new_n20426), .C(new_n20432), .Y(new_n20433));
  NOR2xp33_ASAP7_75t_L      g20177(.A(new_n11591), .B(new_n4142), .Y(new_n20434));
  AOI221xp5_ASAP7_75t_L     g20178(.A1(\b[58] ), .A2(new_n4402), .B1(\b[60] ), .B2(new_n4156), .C(new_n20434), .Y(new_n20435));
  INVx1_ASAP7_75t_L         g20179(.A(new_n20435), .Y(new_n20436));
  A2O1A1Ixp33_ASAP7_75t_L   g20180(.A1(new_n13839), .A2(new_n4151), .B(new_n20436), .C(\a[35] ), .Y(new_n20437));
  O2A1O1Ixp33_ASAP7_75t_L   g20181(.A1(new_n4150), .A2(new_n11634), .B(new_n20435), .C(\a[35] ), .Y(new_n20438));
  AO21x2_ASAP7_75t_L        g20182(.A1(\a[35] ), .A2(new_n20437), .B(new_n20438), .Y(new_n20439));
  NAND3xp33_ASAP7_75t_L     g20183(.A(new_n20430), .B(new_n20433), .C(new_n20439), .Y(new_n20440));
  NAND3xp33_ASAP7_75t_L     g20184(.A(new_n20440), .B(new_n20433), .C(new_n20430), .Y(new_n20441));
  NAND2xp33_ASAP7_75t_L     g20185(.A(new_n20433), .B(new_n20430), .Y(new_n20442));
  A2O1A1Ixp33_ASAP7_75t_L   g20186(.A1(\a[35] ), .A2(new_n20437), .B(new_n20438), .C(new_n20442), .Y(new_n20443));
  NAND2xp33_ASAP7_75t_L     g20187(.A(new_n20443), .B(new_n20441), .Y(new_n20444));
  INVx1_ASAP7_75t_L         g20188(.A(new_n20066), .Y(new_n20445));
  A2O1A1O1Ixp25_ASAP7_75t_L g20189(.A1(new_n20445), .A2(new_n20060), .B(new_n20124), .C(new_n20257), .D(new_n20264), .Y(new_n20446));
  INVx1_ASAP7_75t_L         g20190(.A(new_n20446), .Y(new_n20447));
  NOR2xp33_ASAP7_75t_L      g20191(.A(new_n20447), .B(new_n20444), .Y(new_n20448));
  O2A1O1Ixp33_ASAP7_75t_L   g20192(.A1(new_n4150), .A2(new_n11634), .B(new_n20435), .C(new_n4145), .Y(new_n20449));
  INVx1_ASAP7_75t_L         g20193(.A(new_n20438), .Y(new_n20450));
  O2A1O1Ixp33_ASAP7_75t_L   g20194(.A1(new_n20449), .A2(new_n4145), .B(new_n20450), .C(new_n20442), .Y(new_n20451));
  O2A1O1Ixp33_ASAP7_75t_L   g20195(.A1(new_n20442), .A2(new_n20451), .B(new_n20443), .C(new_n20446), .Y(new_n20452));
  NOR2xp33_ASAP7_75t_L      g20196(.A(new_n20452), .B(new_n20448), .Y(new_n20453));
  INVx1_ASAP7_75t_L         g20197(.A(new_n20453), .Y(new_n20454));
  NAND2xp33_ASAP7_75t_L     g20198(.A(new_n20122), .B(new_n20270), .Y(new_n20455));
  NAND2xp33_ASAP7_75t_L     g20199(.A(new_n20122), .B(new_n20268), .Y(new_n20456));
  O2A1O1Ixp33_ASAP7_75t_L   g20200(.A1(new_n20258), .A2(new_n20264), .B(new_n20266), .C(new_n20456), .Y(new_n20457));
  A2O1A1O1Ixp25_ASAP7_75t_L g20201(.A1(new_n20118), .A2(\a[32] ), .B(new_n20119), .C(new_n20120), .D(new_n20457), .Y(new_n20458));
  NOR2xp33_ASAP7_75t_L      g20202(.A(new_n12956), .B(new_n3510), .Y(new_n20459));
  AOI221xp5_ASAP7_75t_L     g20203(.A1(\b[61] ), .A2(new_n3708), .B1(\b[62] ), .B2(new_n3499), .C(new_n20459), .Y(new_n20460));
  O2A1O1Ixp33_ASAP7_75t_L   g20204(.A1(new_n3513), .A2(new_n17815), .B(new_n20460), .C(new_n3493), .Y(new_n20461));
  O2A1O1Ixp33_ASAP7_75t_L   g20205(.A1(new_n3513), .A2(new_n17815), .B(new_n20460), .C(\a[32] ), .Y(new_n20462));
  INVx1_ASAP7_75t_L         g20206(.A(new_n20462), .Y(new_n20463));
  O2A1O1Ixp33_ASAP7_75t_L   g20207(.A1(new_n20461), .A2(new_n3493), .B(new_n20463), .C(new_n20458), .Y(new_n20464));
  INVx1_ASAP7_75t_L         g20208(.A(new_n20464), .Y(new_n20465));
  O2A1O1Ixp33_ASAP7_75t_L   g20209(.A1(new_n20461), .A2(new_n3493), .B(new_n20463), .C(new_n20455), .Y(new_n20466));
  AOI21xp33_ASAP7_75t_L     g20210(.A1(new_n20465), .A2(new_n20455), .B(new_n20466), .Y(new_n20467));
  NAND2xp33_ASAP7_75t_L     g20211(.A(new_n20454), .B(new_n20467), .Y(new_n20468));
  A2O1A1Ixp33_ASAP7_75t_L   g20212(.A1(new_n20465), .A2(new_n20455), .B(new_n20466), .C(new_n20453), .Y(new_n20469));
  AND2x2_ASAP7_75t_L        g20213(.A(new_n20469), .B(new_n20468), .Y(new_n20470));
  XNOR2x2_ASAP7_75t_L       g20214(.A(new_n20289), .B(new_n20470), .Y(new_n20471));
  A2O1A1Ixp33_ASAP7_75t_L   g20215(.A1(new_n20281), .A2(new_n20288), .B(new_n20278), .C(new_n20471), .Y(new_n20472));
  INVx1_ASAP7_75t_L         g20216(.A(new_n20472), .Y(new_n20473));
  A2O1A1Ixp33_ASAP7_75t_L   g20217(.A1(new_n20287), .A2(new_n20283), .B(new_n20282), .C(new_n20277), .Y(new_n20474));
  NOR2xp33_ASAP7_75t_L      g20218(.A(new_n20471), .B(new_n20474), .Y(new_n20475));
  NOR2xp33_ASAP7_75t_L      g20219(.A(new_n20473), .B(new_n20475), .Y(\f[93] ));
  O2A1O1Ixp33_ASAP7_75t_L   g20220(.A1(new_n20455), .A2(new_n20466), .B(new_n20453), .C(new_n20464), .Y(new_n20477));
  INVx1_ASAP7_75t_L         g20221(.A(new_n20467), .Y(new_n20478));
  AOI22xp33_ASAP7_75t_L     g20222(.A1(new_n3499), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3708), .Y(new_n20479));
  INVx1_ASAP7_75t_L         g20223(.A(new_n20479), .Y(new_n20480));
  A2O1A1Ixp33_ASAP7_75t_L   g20224(.A1(new_n3500), .A2(new_n3501), .B(new_n3302), .C(new_n20479), .Y(new_n20481));
  O2A1O1Ixp33_ASAP7_75t_L   g20225(.A1(new_n20480), .A2(new_n17329), .B(new_n20481), .C(new_n3493), .Y(new_n20482));
  O2A1O1Ixp33_ASAP7_75t_L   g20226(.A1(new_n3513), .A2(new_n12993), .B(new_n20479), .C(\a[32] ), .Y(new_n20483));
  NOR2xp33_ASAP7_75t_L      g20227(.A(new_n20483), .B(new_n20482), .Y(new_n20484));
  A2O1A1O1Ixp25_ASAP7_75t_L g20228(.A1(new_n20442), .A2(new_n20443), .B(new_n20446), .C(new_n20440), .D(new_n20484), .Y(new_n20485));
  A2O1A1Ixp33_ASAP7_75t_L   g20229(.A1(new_n20443), .A2(new_n20442), .B(new_n20446), .C(new_n20440), .Y(new_n20486));
  NOR3xp33_ASAP7_75t_L      g20230(.A(new_n20486), .B(new_n20482), .C(new_n20483), .Y(new_n20487));
  NOR2xp33_ASAP7_75t_L      g20231(.A(new_n20485), .B(new_n20487), .Y(new_n20488));
  INVx1_ASAP7_75t_L         g20232(.A(new_n20392), .Y(new_n20489));
  INVx1_ASAP7_75t_L         g20233(.A(new_n20357), .Y(new_n20490));
  NOR2xp33_ASAP7_75t_L      g20234(.A(new_n5570), .B(new_n10388), .Y(new_n20491));
  AOI221xp5_ASAP7_75t_L     g20235(.A1(new_n10086), .A2(\b[40] ), .B1(new_n11361), .B2(\b[38] ), .C(new_n20491), .Y(new_n20492));
  O2A1O1Ixp33_ASAP7_75t_L   g20236(.A1(new_n10088), .A2(new_n5862), .B(new_n20492), .C(new_n10083), .Y(new_n20493));
  INVx1_ASAP7_75t_L         g20237(.A(new_n20493), .Y(new_n20494));
  O2A1O1Ixp33_ASAP7_75t_L   g20238(.A1(new_n10088), .A2(new_n5862), .B(new_n20492), .C(\a[56] ), .Y(new_n20495));
  A2O1A1Ixp33_ASAP7_75t_L   g20239(.A1(new_n20313), .A2(new_n20312), .B(new_n20314), .C(new_n20321), .Y(new_n20496));
  NOR2xp33_ASAP7_75t_L      g20240(.A(new_n3456), .B(new_n13030), .Y(new_n20497));
  INVx1_ASAP7_75t_L         g20241(.A(new_n20303), .Y(new_n20498));
  A2O1A1O1Ixp25_ASAP7_75t_L g20242(.A1(new_n13028), .A2(\b[29] ), .B(new_n20149), .C(new_n20305), .D(new_n20498), .Y(new_n20499));
  A2O1A1Ixp33_ASAP7_75t_L   g20243(.A1(new_n13028), .A2(\b[31] ), .B(new_n20497), .C(new_n20499), .Y(new_n20500));
  INVx1_ASAP7_75t_L         g20244(.A(new_n20154), .Y(new_n20501));
  O2A1O1Ixp33_ASAP7_75t_L   g20245(.A1(new_n12669), .A2(new_n12671), .B(\b[31] ), .C(new_n20497), .Y(new_n20502));
  A2O1A1Ixp33_ASAP7_75t_L   g20246(.A1(new_n20305), .A2(new_n20501), .B(new_n20498), .C(new_n20502), .Y(new_n20503));
  NAND2xp33_ASAP7_75t_L     g20247(.A(new_n20503), .B(new_n20500), .Y(new_n20504));
  NOR2xp33_ASAP7_75t_L      g20248(.A(new_n4101), .B(new_n12318), .Y(new_n20505));
  AOI221xp5_ASAP7_75t_L     g20249(.A1(new_n11995), .A2(\b[34] ), .B1(new_n13314), .B2(\b[32] ), .C(new_n20505), .Y(new_n20506));
  O2A1O1Ixp33_ASAP7_75t_L   g20250(.A1(new_n11998), .A2(new_n4352), .B(new_n20506), .C(new_n11987), .Y(new_n20507));
  O2A1O1Ixp33_ASAP7_75t_L   g20251(.A1(new_n11998), .A2(new_n4352), .B(new_n20506), .C(\a[62] ), .Y(new_n20508));
  INVx1_ASAP7_75t_L         g20252(.A(new_n20508), .Y(new_n20509));
  OAI211xp5_ASAP7_75t_L     g20253(.A1(new_n11987), .A2(new_n20507), .B(new_n20509), .C(new_n20504), .Y(new_n20510));
  INVx1_ASAP7_75t_L         g20254(.A(new_n20504), .Y(new_n20511));
  INVx1_ASAP7_75t_L         g20255(.A(new_n20507), .Y(new_n20512));
  A2O1A1Ixp33_ASAP7_75t_L   g20256(.A1(new_n20512), .A2(\a[62] ), .B(new_n20508), .C(new_n20511), .Y(new_n20513));
  NAND2xp33_ASAP7_75t_L     g20257(.A(new_n20510), .B(new_n20513), .Y(new_n20514));
  INVx1_ASAP7_75t_L         g20258(.A(new_n20514), .Y(new_n20515));
  NOR2xp33_ASAP7_75t_L      g20259(.A(new_n4581), .B(new_n11354), .Y(new_n20516));
  AOI221xp5_ASAP7_75t_L     g20260(.A1(\b[37] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[36] ), .C(new_n20516), .Y(new_n20517));
  O2A1O1Ixp33_ASAP7_75t_L   g20261(.A1(new_n11053), .A2(new_n5083), .B(new_n20517), .C(new_n11048), .Y(new_n20518));
  NOR2xp33_ASAP7_75t_L      g20262(.A(new_n11048), .B(new_n20518), .Y(new_n20519));
  O2A1O1Ixp33_ASAP7_75t_L   g20263(.A1(new_n11053), .A2(new_n5083), .B(new_n20517), .C(\a[59] ), .Y(new_n20520));
  NOR2xp33_ASAP7_75t_L      g20264(.A(new_n20520), .B(new_n20519), .Y(new_n20521));
  A2O1A1O1Ixp25_ASAP7_75t_L g20265(.A1(new_n20320), .A2(new_n20319), .B(new_n20315), .C(new_n20313), .D(new_n20514), .Y(new_n20522));
  A2O1A1O1Ixp25_ASAP7_75t_L g20266(.A1(new_n20320), .A2(new_n20319), .B(new_n20315), .C(new_n20313), .D(new_n20515), .Y(new_n20523));
  INVx1_ASAP7_75t_L         g20267(.A(new_n20523), .Y(new_n20524));
  O2A1O1Ixp33_ASAP7_75t_L   g20268(.A1(new_n20514), .A2(new_n20522), .B(new_n20524), .C(new_n20521), .Y(new_n20525));
  A2O1A1Ixp33_ASAP7_75t_L   g20269(.A1(new_n20319), .A2(new_n20320), .B(new_n20315), .C(new_n20313), .Y(new_n20526));
  NOR2xp33_ASAP7_75t_L      g20270(.A(new_n20514), .B(new_n20526), .Y(new_n20527));
  NOR3xp33_ASAP7_75t_L      g20271(.A(new_n20527), .B(new_n20520), .C(new_n20519), .Y(new_n20528));
  A2O1A1O1Ixp25_ASAP7_75t_L g20272(.A1(new_n20496), .A2(new_n20313), .B(new_n20515), .C(new_n20528), .D(new_n20525), .Y(new_n20529));
  A2O1A1Ixp33_ASAP7_75t_L   g20273(.A1(new_n20330), .A2(new_n20334), .B(new_n20328), .C(new_n20529), .Y(new_n20530));
  A2O1A1Ixp33_ASAP7_75t_L   g20274(.A1(new_n20331), .A2(new_n20334), .B(new_n20328), .C(new_n20530), .Y(new_n20531));
  NAND2xp33_ASAP7_75t_L     g20275(.A(new_n20529), .B(new_n20530), .Y(new_n20532));
  NAND2xp33_ASAP7_75t_L     g20276(.A(new_n20532), .B(new_n20531), .Y(new_n20533));
  AOI21xp33_ASAP7_75t_L     g20277(.A1(new_n20494), .A2(\a[56] ), .B(new_n20495), .Y(new_n20534));
  NAND2xp33_ASAP7_75t_L     g20278(.A(new_n20534), .B(new_n20532), .Y(new_n20535));
  O2A1O1Ixp33_ASAP7_75t_L   g20279(.A1(new_n20328), .A2(new_n20333), .B(new_n20530), .C(new_n20535), .Y(new_n20536));
  A2O1A1O1Ixp25_ASAP7_75t_L g20280(.A1(new_n20494), .A2(\a[56] ), .B(new_n20495), .C(new_n20533), .D(new_n20536), .Y(new_n20537));
  INVx1_ASAP7_75t_L         g20281(.A(new_n20537), .Y(new_n20538));
  A2O1A1O1Ixp25_ASAP7_75t_L g20282(.A1(new_n20172), .A2(new_n20184), .B(new_n20345), .C(new_n20342), .D(new_n20538), .Y(new_n20539));
  INVx1_ASAP7_75t_L         g20283(.A(new_n20539), .Y(new_n20540));
  INVx1_ASAP7_75t_L         g20284(.A(new_n20336), .Y(new_n20541));
  O2A1O1Ixp33_ASAP7_75t_L   g20285(.A1(new_n20339), .A2(new_n10083), .B(new_n20343), .C(new_n20541), .Y(new_n20542));
  O2A1O1Ixp33_ASAP7_75t_L   g20286(.A1(new_n20171), .A2(new_n20183), .B(new_n20349), .C(new_n20542), .Y(new_n20543));
  NAND2xp33_ASAP7_75t_L     g20287(.A(new_n20538), .B(new_n20543), .Y(new_n20544));
  AND2x2_ASAP7_75t_L        g20288(.A(new_n20544), .B(new_n20540), .Y(new_n20545));
  INVx1_ASAP7_75t_L         g20289(.A(new_n20545), .Y(new_n20546));
  NOR2xp33_ASAP7_75t_L      g20290(.A(new_n6378), .B(new_n10400), .Y(new_n20547));
  AOI221xp5_ASAP7_75t_L     g20291(.A1(new_n9102), .A2(\b[43] ), .B1(new_n10398), .B2(\b[41] ), .C(new_n20547), .Y(new_n20548));
  O2A1O1Ixp33_ASAP7_75t_L   g20292(.A1(new_n9104), .A2(new_n6679), .B(new_n20548), .C(new_n9099), .Y(new_n20549));
  O2A1O1Ixp33_ASAP7_75t_L   g20293(.A1(new_n9104), .A2(new_n6679), .B(new_n20548), .C(\a[53] ), .Y(new_n20550));
  INVx1_ASAP7_75t_L         g20294(.A(new_n20550), .Y(new_n20551));
  O2A1O1Ixp33_ASAP7_75t_L   g20295(.A1(new_n20549), .A2(new_n9099), .B(new_n20551), .C(new_n20546), .Y(new_n20552));
  INVx1_ASAP7_75t_L         g20296(.A(new_n20552), .Y(new_n20553));
  O2A1O1Ixp33_ASAP7_75t_L   g20297(.A1(new_n20549), .A2(new_n9099), .B(new_n20551), .C(new_n20545), .Y(new_n20554));
  AO21x2_ASAP7_75t_L        g20298(.A1(new_n20545), .A2(new_n20553), .B(new_n20554), .Y(new_n20555));
  INVx1_ASAP7_75t_L         g20299(.A(new_n20351), .Y(new_n20556));
  INVx1_ASAP7_75t_L         g20300(.A(new_n20359), .Y(new_n20557));
  O2A1O1Ixp33_ASAP7_75t_L   g20301(.A1(new_n20556), .A2(new_n20490), .B(new_n20557), .C(new_n20362), .Y(new_n20558));
  OR3x1_ASAP7_75t_L         g20302(.A(new_n20555), .B(new_n20490), .C(new_n20558), .Y(new_n20559));
  A2O1A1Ixp33_ASAP7_75t_L   g20303(.A1(new_n20557), .A2(new_n20556), .B(new_n20362), .C(new_n20357), .Y(new_n20560));
  A2O1A1Ixp33_ASAP7_75t_L   g20304(.A1(new_n20553), .A2(new_n20545), .B(new_n20554), .C(new_n20560), .Y(new_n20561));
  NAND2xp33_ASAP7_75t_L     g20305(.A(new_n20561), .B(new_n20559), .Y(new_n20562));
  INVx1_ASAP7_75t_L         g20306(.A(new_n20562), .Y(new_n20563));
  NOR2xp33_ASAP7_75t_L      g20307(.A(new_n7249), .B(new_n10065), .Y(new_n20564));
  AOI221xp5_ASAP7_75t_L     g20308(.A1(new_n8175), .A2(\b[46] ), .B1(new_n8484), .B2(\b[44] ), .C(new_n20564), .Y(new_n20565));
  O2A1O1Ixp33_ASAP7_75t_L   g20309(.A1(new_n8176), .A2(new_n7279), .B(new_n20565), .C(new_n8172), .Y(new_n20566));
  O2A1O1Ixp33_ASAP7_75t_L   g20310(.A1(new_n8176), .A2(new_n7279), .B(new_n20565), .C(\a[50] ), .Y(new_n20567));
  INVx1_ASAP7_75t_L         g20311(.A(new_n20567), .Y(new_n20568));
  O2A1O1Ixp33_ASAP7_75t_L   g20312(.A1(new_n20566), .A2(new_n8172), .B(new_n20568), .C(new_n20562), .Y(new_n20569));
  INVx1_ASAP7_75t_L         g20313(.A(new_n20569), .Y(new_n20570));
  NAND2xp33_ASAP7_75t_L     g20314(.A(new_n20563), .B(new_n20570), .Y(new_n20571));
  O2A1O1Ixp33_ASAP7_75t_L   g20315(.A1(new_n20566), .A2(new_n8172), .B(new_n20568), .C(new_n20563), .Y(new_n20572));
  INVx1_ASAP7_75t_L         g20316(.A(new_n20572), .Y(new_n20573));
  A2O1A1O1Ixp25_ASAP7_75t_L g20317(.A1(new_n20369), .A2(\a[50] ), .B(new_n20370), .C(new_n20365), .D(new_n20377), .Y(new_n20574));
  NAND3xp33_ASAP7_75t_L     g20318(.A(new_n20574), .B(new_n20573), .C(new_n20571), .Y(new_n20575));
  O2A1O1Ixp33_ASAP7_75t_L   g20319(.A1(new_n20562), .A2(new_n20569), .B(new_n20573), .C(new_n20574), .Y(new_n20576));
  INVx1_ASAP7_75t_L         g20320(.A(new_n20576), .Y(new_n20577));
  AND2x2_ASAP7_75t_L        g20321(.A(new_n20575), .B(new_n20577), .Y(new_n20578));
  NOR2xp33_ASAP7_75t_L      g20322(.A(new_n7860), .B(new_n7312), .Y(new_n20579));
  AOI221xp5_ASAP7_75t_L     g20323(.A1(\b[47] ), .A2(new_n7609), .B1(\b[49] ), .B2(new_n7334), .C(new_n20579), .Y(new_n20580));
  INVx1_ASAP7_75t_L         g20324(.A(new_n20580), .Y(new_n20581));
  A2O1A1Ixp33_ASAP7_75t_L   g20325(.A1(new_n8438), .A2(new_n7322), .B(new_n20581), .C(\a[47] ), .Y(new_n20582));
  O2A1O1Ixp33_ASAP7_75t_L   g20326(.A1(new_n7321), .A2(new_n14802), .B(new_n20580), .C(\a[47] ), .Y(new_n20583));
  A2O1A1Ixp33_ASAP7_75t_L   g20327(.A1(\a[47] ), .A2(new_n20582), .B(new_n20583), .C(new_n20578), .Y(new_n20584));
  NAND2xp33_ASAP7_75t_L     g20328(.A(new_n20578), .B(new_n20584), .Y(new_n20585));
  A2O1A1Ixp33_ASAP7_75t_L   g20329(.A1(new_n20582), .A2(\a[47] ), .B(new_n20583), .C(new_n20584), .Y(new_n20586));
  AND4x1_ASAP7_75t_L        g20330(.A(new_n20489), .B(new_n20387), .C(new_n20586), .D(new_n20585), .Y(new_n20587));
  AND2x2_ASAP7_75t_L        g20331(.A(new_n20585), .B(new_n20586), .Y(new_n20588));
  O2A1O1Ixp33_ASAP7_75t_L   g20332(.A1(new_n20389), .A2(new_n20390), .B(new_n20387), .C(new_n20588), .Y(new_n20589));
  NOR2xp33_ASAP7_75t_L      g20333(.A(new_n20587), .B(new_n20589), .Y(new_n20590));
  NOR2xp33_ASAP7_75t_L      g20334(.A(new_n8779), .B(new_n7304), .Y(new_n20591));
  AOI221xp5_ASAP7_75t_L     g20335(.A1(\b[50] ), .A2(new_n6742), .B1(\b[52] ), .B2(new_n6442), .C(new_n20591), .Y(new_n20592));
  O2A1O1Ixp33_ASAP7_75t_L   g20336(.A1(new_n6443), .A2(new_n17363), .B(new_n20592), .C(new_n6439), .Y(new_n20593));
  INVx1_ASAP7_75t_L         g20337(.A(new_n20593), .Y(new_n20594));
  O2A1O1Ixp33_ASAP7_75t_L   g20338(.A1(new_n6443), .A2(new_n17363), .B(new_n20592), .C(\a[44] ), .Y(new_n20595));
  A2O1A1Ixp33_ASAP7_75t_L   g20339(.A1(\a[44] ), .A2(new_n20594), .B(new_n20595), .C(new_n20590), .Y(new_n20596));
  INVx1_ASAP7_75t_L         g20340(.A(new_n20595), .Y(new_n20597));
  O2A1O1Ixp33_ASAP7_75t_L   g20341(.A1(new_n20593), .A2(new_n6439), .B(new_n20597), .C(new_n20590), .Y(new_n20598));
  AOI21xp33_ASAP7_75t_L     g20342(.A1(new_n20596), .A2(new_n20590), .B(new_n20598), .Y(new_n20599));
  A2O1A1Ixp33_ASAP7_75t_L   g20343(.A1(new_n20401), .A2(new_n20393), .B(new_n20403), .C(new_n20599), .Y(new_n20600));
  INVx1_ASAP7_75t_L         g20344(.A(new_n20405), .Y(new_n20601));
  A2O1A1Ixp33_ASAP7_75t_L   g20345(.A1(new_n20596), .A2(new_n20590), .B(new_n20598), .C(new_n20601), .Y(new_n20602));
  NAND2xp33_ASAP7_75t_L     g20346(.A(new_n20602), .B(new_n20600), .Y(new_n20603));
  NOR2xp33_ASAP7_75t_L      g20347(.A(new_n10309), .B(new_n5641), .Y(new_n20604));
  AOI221xp5_ASAP7_75t_L     g20348(.A1(\b[53] ), .A2(new_n5920), .B1(\b[54] ), .B2(new_n5623), .C(new_n20604), .Y(new_n20605));
  O2A1O1Ixp33_ASAP7_75t_L   g20349(.A1(new_n5630), .A2(new_n15849), .B(new_n20605), .C(new_n5626), .Y(new_n20606));
  NOR2xp33_ASAP7_75t_L      g20350(.A(new_n5626), .B(new_n20606), .Y(new_n20607));
  O2A1O1Ixp33_ASAP7_75t_L   g20351(.A1(new_n5630), .A2(new_n15849), .B(new_n20605), .C(\a[41] ), .Y(new_n20608));
  NOR2xp33_ASAP7_75t_L      g20352(.A(new_n20608), .B(new_n20607), .Y(new_n20609));
  XNOR2x2_ASAP7_75t_L       g20353(.A(new_n20609), .B(new_n20603), .Y(new_n20610));
  A2O1A1Ixp33_ASAP7_75t_L   g20354(.A1(new_n20417), .A2(new_n20290), .B(new_n20416), .C(new_n20610), .Y(new_n20611));
  O2A1O1Ixp33_ASAP7_75t_L   g20355(.A1(new_n20134), .A2(new_n20243), .B(new_n20244), .C(new_n20247), .Y(new_n20612));
  O2A1O1Ixp33_ASAP7_75t_L   g20356(.A1(new_n20612), .A2(new_n20243), .B(new_n20417), .C(new_n20416), .Y(new_n20613));
  INVx1_ASAP7_75t_L         g20357(.A(new_n20610), .Y(new_n20614));
  NAND2xp33_ASAP7_75t_L     g20358(.A(new_n20613), .B(new_n20614), .Y(new_n20615));
  NAND2xp33_ASAP7_75t_L     g20359(.A(new_n20611), .B(new_n20615), .Y(new_n20616));
  INVx1_ASAP7_75t_L         g20360(.A(new_n20616), .Y(new_n20617));
  NOR2xp33_ASAP7_75t_L      g20361(.A(new_n11303), .B(new_n4908), .Y(new_n20618));
  AOI221xp5_ASAP7_75t_L     g20362(.A1(\b[56] ), .A2(new_n5139), .B1(\b[57] ), .B2(new_n4916), .C(new_n20618), .Y(new_n20619));
  O2A1O1Ixp33_ASAP7_75t_L   g20363(.A1(new_n4911), .A2(new_n20073), .B(new_n20619), .C(new_n4906), .Y(new_n20620));
  O2A1O1Ixp33_ASAP7_75t_L   g20364(.A1(new_n4911), .A2(new_n20073), .B(new_n20619), .C(\a[38] ), .Y(new_n20621));
  INVx1_ASAP7_75t_L         g20365(.A(new_n20621), .Y(new_n20622));
  O2A1O1Ixp33_ASAP7_75t_L   g20366(.A1(new_n20620), .A2(new_n4906), .B(new_n20622), .C(new_n20616), .Y(new_n20623));
  INVx1_ASAP7_75t_L         g20367(.A(new_n20623), .Y(new_n20624));
  O2A1O1Ixp33_ASAP7_75t_L   g20368(.A1(new_n20620), .A2(new_n4906), .B(new_n20622), .C(new_n20617), .Y(new_n20625));
  AOI21xp33_ASAP7_75t_L     g20369(.A1(new_n20624), .A2(new_n20617), .B(new_n20625), .Y(new_n20626));
  O2A1O1Ixp33_ASAP7_75t_L   g20370(.A1(new_n20425), .A2(new_n20426), .B(new_n20432), .C(new_n20424), .Y(new_n20627));
  NAND2xp33_ASAP7_75t_L     g20371(.A(new_n20627), .B(new_n20626), .Y(new_n20628));
  A2O1A1O1Ixp25_ASAP7_75t_L g20372(.A1(new_n20427), .A2(new_n20418), .B(new_n20429), .C(new_n20431), .D(new_n20626), .Y(new_n20629));
  INVx1_ASAP7_75t_L         g20373(.A(new_n20629), .Y(new_n20630));
  AND2x2_ASAP7_75t_L        g20374(.A(new_n20628), .B(new_n20630), .Y(new_n20631));
  NOR2xp33_ASAP7_75t_L      g20375(.A(new_n12258), .B(new_n4147), .Y(new_n20632));
  AOI221xp5_ASAP7_75t_L     g20376(.A1(\b[59] ), .A2(new_n4402), .B1(\b[60] ), .B2(new_n4155), .C(new_n20632), .Y(new_n20633));
  O2A1O1Ixp33_ASAP7_75t_L   g20377(.A1(new_n4150), .A2(new_n14764), .B(new_n20633), .C(new_n4145), .Y(new_n20634));
  INVx1_ASAP7_75t_L         g20378(.A(new_n20634), .Y(new_n20635));
  O2A1O1Ixp33_ASAP7_75t_L   g20379(.A1(new_n4150), .A2(new_n14764), .B(new_n20633), .C(\a[35] ), .Y(new_n20636));
  A2O1A1Ixp33_ASAP7_75t_L   g20380(.A1(\a[35] ), .A2(new_n20635), .B(new_n20636), .C(new_n20631), .Y(new_n20637));
  NOR2xp33_ASAP7_75t_L      g20381(.A(new_n4145), .B(new_n20634), .Y(new_n20638));
  OR3x1_ASAP7_75t_L         g20382(.A(new_n20631), .B(new_n20638), .C(new_n20636), .Y(new_n20639));
  NAND3xp33_ASAP7_75t_L     g20383(.A(new_n20639), .B(new_n20637), .C(new_n20488), .Y(new_n20640));
  NAND2xp33_ASAP7_75t_L     g20384(.A(new_n20488), .B(new_n20640), .Y(new_n20641));
  NAND3xp33_ASAP7_75t_L     g20385(.A(new_n20640), .B(new_n20639), .C(new_n20637), .Y(new_n20642));
  NAND2xp33_ASAP7_75t_L     g20386(.A(new_n20641), .B(new_n20642), .Y(new_n20643));
  A2O1A1Ixp33_ASAP7_75t_L   g20387(.A1(new_n20478), .A2(new_n20453), .B(new_n20464), .C(new_n20643), .Y(new_n20644));
  INVx1_ASAP7_75t_L         g20388(.A(new_n20644), .Y(new_n20645));
  INVx1_ASAP7_75t_L         g20389(.A(new_n20642), .Y(new_n20646));
  A2O1A1Ixp33_ASAP7_75t_L   g20390(.A1(new_n20640), .A2(new_n20488), .B(new_n20646), .C(new_n20477), .Y(new_n20647));
  O2A1O1Ixp33_ASAP7_75t_L   g20391(.A1(new_n20109), .A2(new_n20272), .B(new_n20470), .C(new_n20473), .Y(new_n20648));
  O2A1O1Ixp33_ASAP7_75t_L   g20392(.A1(new_n20477), .A2(new_n20645), .B(new_n20647), .C(new_n20648), .Y(new_n20649));
  OAI21xp33_ASAP7_75t_L     g20393(.A1(new_n20109), .A2(new_n20272), .B(new_n20470), .Y(new_n20650));
  O2A1O1Ixp33_ASAP7_75t_L   g20394(.A1(new_n20454), .A2(new_n20467), .B(new_n20465), .C(new_n20643), .Y(new_n20651));
  A2O1A1O1Ixp25_ASAP7_75t_L g20395(.A1(new_n20640), .A2(new_n20488), .B(new_n20646), .C(new_n20644), .D(new_n20651), .Y(new_n20652));
  AND3x1_ASAP7_75t_L        g20396(.A(new_n20472), .B(new_n20652), .C(new_n20650), .Y(new_n20653));
  NOR2xp33_ASAP7_75t_L      g20397(.A(new_n20653), .B(new_n20649), .Y(\f[94] ));
  O2A1O1Ixp33_ASAP7_75t_L   g20398(.A1(new_n20638), .A2(new_n20636), .B(new_n20628), .C(new_n20629), .Y(new_n20655));
  INVx1_ASAP7_75t_L         g20399(.A(new_n20655), .Y(new_n20656));
  NOR2xp33_ASAP7_75t_L      g20400(.A(new_n12956), .B(new_n3703), .Y(new_n20657));
  A2O1A1Ixp33_ASAP7_75t_L   g20401(.A1(new_n12986), .A2(new_n3505), .B(new_n20657), .C(\a[32] ), .Y(new_n20658));
  INVx1_ASAP7_75t_L         g20402(.A(new_n20658), .Y(new_n20659));
  A2O1A1Ixp33_ASAP7_75t_L   g20403(.A1(new_n12986), .A2(new_n3505), .B(new_n20657), .C(new_n3493), .Y(new_n20660));
  O2A1O1Ixp33_ASAP7_75t_L   g20404(.A1(new_n20659), .A2(new_n3493), .B(new_n20660), .C(new_n20655), .Y(new_n20661));
  INVx1_ASAP7_75t_L         g20405(.A(new_n20661), .Y(new_n20662));
  O2A1O1Ixp33_ASAP7_75t_L   g20406(.A1(new_n20659), .A2(new_n3493), .B(new_n20660), .C(new_n20656), .Y(new_n20663));
  INVx1_ASAP7_75t_L         g20407(.A(new_n20613), .Y(new_n20664));
  A2O1A1O1Ixp25_ASAP7_75t_L g20408(.A1(new_n20221), .A2(new_n20215), .B(new_n20223), .C(new_n20225), .D(new_n20291), .Y(new_n20665));
  O2A1O1Ixp33_ASAP7_75t_L   g20409(.A1(new_n20665), .A2(new_n20402), .B(new_n20399), .C(new_n20599), .Y(new_n20666));
  INVx1_ASAP7_75t_L         g20410(.A(new_n20666), .Y(new_n20667));
  NOR2xp33_ASAP7_75t_L      g20411(.A(new_n10309), .B(new_n5640), .Y(new_n20668));
  AOI221xp5_ASAP7_75t_L     g20412(.A1(\b[54] ), .A2(new_n5920), .B1(\b[56] ), .B2(new_n5629), .C(new_n20668), .Y(new_n20669));
  INVx1_ASAP7_75t_L         g20413(.A(new_n20669), .Y(new_n20670));
  A2O1A1Ixp33_ASAP7_75t_L   g20414(.A1(new_n11579), .A2(new_n5637), .B(new_n20670), .C(\a[41] ), .Y(new_n20671));
  O2A1O1Ixp33_ASAP7_75t_L   g20415(.A1(new_n5630), .A2(new_n10339), .B(new_n20669), .C(new_n5626), .Y(new_n20672));
  NOR2xp33_ASAP7_75t_L      g20416(.A(new_n5626), .B(new_n20672), .Y(new_n20673));
  A2O1A1O1Ixp25_ASAP7_75t_L g20417(.A1(new_n11579), .A2(new_n5637), .B(new_n20670), .C(new_n20671), .D(new_n20673), .Y(new_n20674));
  A2O1A1O1Ixp25_ASAP7_75t_L g20418(.A1(new_n20582), .A2(\a[47] ), .B(new_n20583), .C(new_n20575), .D(new_n20576), .Y(new_n20675));
  INVx1_ASAP7_75t_L         g20419(.A(new_n20675), .Y(new_n20676));
  NOR2xp33_ASAP7_75t_L      g20420(.A(new_n6671), .B(new_n10400), .Y(new_n20677));
  AOI221xp5_ASAP7_75t_L     g20421(.A1(new_n9102), .A2(\b[44] ), .B1(new_n10398), .B2(\b[42] ), .C(new_n20677), .Y(new_n20678));
  O2A1O1Ixp33_ASAP7_75t_L   g20422(.A1(new_n9104), .A2(new_n6951), .B(new_n20678), .C(new_n9099), .Y(new_n20679));
  INVx1_ASAP7_75t_L         g20423(.A(new_n20679), .Y(new_n20680));
  O2A1O1Ixp33_ASAP7_75t_L   g20424(.A1(new_n9104), .A2(new_n6951), .B(new_n20678), .C(\a[53] ), .Y(new_n20681));
  NOR2xp33_ASAP7_75t_L      g20425(.A(new_n20328), .B(new_n20333), .Y(new_n20682));
  NOR2xp33_ASAP7_75t_L      g20426(.A(new_n5855), .B(new_n10388), .Y(new_n20683));
  AOI221xp5_ASAP7_75t_L     g20427(.A1(new_n10086), .A2(\b[41] ), .B1(new_n11361), .B2(\b[39] ), .C(new_n20683), .Y(new_n20684));
  O2A1O1Ixp33_ASAP7_75t_L   g20428(.A1(new_n10088), .A2(new_n6117), .B(new_n20684), .C(new_n10083), .Y(new_n20685));
  INVx1_ASAP7_75t_L         g20429(.A(new_n20685), .Y(new_n20686));
  O2A1O1Ixp33_ASAP7_75t_L   g20430(.A1(new_n10088), .A2(new_n6117), .B(new_n20684), .C(\a[56] ), .Y(new_n20687));
  OAI22xp33_ASAP7_75t_L     g20431(.A1(new_n12320), .A2(new_n4101), .B1(new_n4344), .B2(new_n12318), .Y(new_n20688));
  AOI221xp5_ASAP7_75t_L     g20432(.A1(new_n11995), .A2(\b[35] ), .B1(new_n11997), .B2(new_n7773), .C(new_n20688), .Y(new_n20689));
  XNOR2x2_ASAP7_75t_L       g20433(.A(new_n11987), .B(new_n20689), .Y(new_n20690));
  INVx1_ASAP7_75t_L         g20434(.A(new_n20690), .Y(new_n20691));
  INVx1_ASAP7_75t_L         g20435(.A(new_n20502), .Y(new_n20692));
  NOR2xp33_ASAP7_75t_L      g20436(.A(new_n3674), .B(new_n13030), .Y(new_n20693));
  INVx1_ASAP7_75t_L         g20437(.A(new_n20693), .Y(new_n20694));
  O2A1O1Ixp33_ASAP7_75t_L   g20438(.A1(new_n12672), .A2(new_n3891), .B(new_n20694), .C(new_n20692), .Y(new_n20695));
  A2O1A1Ixp33_ASAP7_75t_L   g20439(.A1(new_n20309), .A2(new_n20303), .B(new_n20692), .C(new_n20513), .Y(new_n20696));
  O2A1O1Ixp33_ASAP7_75t_L   g20440(.A1(new_n12669), .A2(new_n12671), .B(\b[32] ), .C(new_n20693), .Y(new_n20697));
  A2O1A1Ixp33_ASAP7_75t_L   g20441(.A1(new_n13028), .A2(\b[31] ), .B(new_n20497), .C(new_n20697), .Y(new_n20698));
  O2A1O1Ixp33_ASAP7_75t_L   g20442(.A1(new_n20692), .A2(new_n20499), .B(new_n20513), .C(new_n20695), .Y(new_n20699));
  NAND2xp33_ASAP7_75t_L     g20443(.A(new_n20698), .B(new_n20699), .Y(new_n20700));
  NAND2xp33_ASAP7_75t_L     g20444(.A(new_n20696), .B(new_n20700), .Y(new_n20701));
  A2O1A1Ixp33_ASAP7_75t_L   g20445(.A1(new_n20513), .A2(new_n20503), .B(new_n20695), .C(new_n20698), .Y(new_n20702));
  O2A1O1Ixp33_ASAP7_75t_L   g20446(.A1(new_n20695), .A2(new_n20702), .B(new_n20701), .C(new_n20690), .Y(new_n20703));
  INVx1_ASAP7_75t_L         g20447(.A(new_n20703), .Y(new_n20704));
  O2A1O1Ixp33_ASAP7_75t_L   g20448(.A1(new_n20695), .A2(new_n20702), .B(new_n20701), .C(new_n20691), .Y(new_n20705));
  NOR2xp33_ASAP7_75t_L      g20449(.A(new_n4613), .B(new_n11354), .Y(new_n20706));
  AOI221xp5_ASAP7_75t_L     g20450(.A1(\b[38] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[37] ), .C(new_n20706), .Y(new_n20707));
  O2A1O1Ixp33_ASAP7_75t_L   g20451(.A1(new_n11053), .A2(new_n5318), .B(new_n20707), .C(new_n11048), .Y(new_n20708));
  NOR2xp33_ASAP7_75t_L      g20452(.A(new_n11048), .B(new_n20708), .Y(new_n20709));
  O2A1O1Ixp33_ASAP7_75t_L   g20453(.A1(new_n11053), .A2(new_n5318), .B(new_n20707), .C(\a[59] ), .Y(new_n20710));
  NOR2xp33_ASAP7_75t_L      g20454(.A(new_n20710), .B(new_n20709), .Y(new_n20711));
  A2O1A1Ixp33_ASAP7_75t_L   g20455(.A1(new_n20704), .A2(new_n20691), .B(new_n20705), .C(new_n20711), .Y(new_n20712));
  A2O1A1O1Ixp25_ASAP7_75t_L g20456(.A1(new_n13028), .A2(\b[32] ), .B(new_n20693), .C(new_n20502), .D(new_n20702), .Y(new_n20713));
  INVx1_ASAP7_75t_L         g20457(.A(new_n20697), .Y(new_n20714));
  A2O1A1Ixp33_ASAP7_75t_L   g20458(.A1(new_n20502), .A2(new_n20714), .B(new_n20702), .C(new_n20701), .Y(new_n20715));
  NOR2xp33_ASAP7_75t_L      g20459(.A(new_n20690), .B(new_n20715), .Y(new_n20716));
  A2O1A1O1Ixp25_ASAP7_75t_L g20460(.A1(new_n20700), .A2(new_n20696), .B(new_n20713), .C(new_n20704), .D(new_n20716), .Y(new_n20717));
  OAI21xp33_ASAP7_75t_L     g20461(.A1(new_n20709), .A2(new_n20710), .B(new_n20717), .Y(new_n20718));
  AND2x2_ASAP7_75t_L        g20462(.A(new_n20712), .B(new_n20718), .Y(new_n20719));
  INVx1_ASAP7_75t_L         g20463(.A(new_n20719), .Y(new_n20720));
  A2O1A1Ixp33_ASAP7_75t_L   g20464(.A1(new_n20515), .A2(new_n20526), .B(new_n20525), .C(new_n20720), .Y(new_n20721));
  INVx1_ASAP7_75t_L         g20465(.A(new_n20527), .Y(new_n20722));
  A2O1A1Ixp33_ASAP7_75t_L   g20466(.A1(new_n20496), .A2(new_n20313), .B(new_n20522), .C(new_n20722), .Y(new_n20723));
  O2A1O1Ixp33_ASAP7_75t_L   g20467(.A1(new_n20520), .A2(new_n20519), .B(new_n20723), .C(new_n20522), .Y(new_n20724));
  NAND2xp33_ASAP7_75t_L     g20468(.A(new_n20724), .B(new_n20719), .Y(new_n20725));
  AND2x2_ASAP7_75t_L        g20469(.A(new_n20725), .B(new_n20721), .Y(new_n20726));
  A2O1A1Ixp33_ASAP7_75t_L   g20470(.A1(new_n20686), .A2(\a[56] ), .B(new_n20687), .C(new_n20726), .Y(new_n20727));
  INVx1_ASAP7_75t_L         g20471(.A(new_n20727), .Y(new_n20728));
  NOR2xp33_ASAP7_75t_L      g20472(.A(new_n10083), .B(new_n20685), .Y(new_n20729));
  NOR3xp33_ASAP7_75t_L      g20473(.A(new_n20726), .B(new_n20687), .C(new_n20729), .Y(new_n20730));
  NOR2xp33_ASAP7_75t_L      g20474(.A(new_n20730), .B(new_n20728), .Y(new_n20731));
  INVx1_ASAP7_75t_L         g20475(.A(new_n20731), .Y(new_n20732));
  A2O1A1O1Ixp25_ASAP7_75t_L g20476(.A1(new_n20532), .A2(new_n20682), .B(new_n20534), .C(new_n20530), .D(new_n20732), .Y(new_n20733));
  INVx1_ASAP7_75t_L         g20477(.A(new_n20733), .Y(new_n20734));
  A2O1A1Ixp33_ASAP7_75t_L   g20478(.A1(new_n20531), .A2(new_n20532), .B(new_n20534), .C(new_n20530), .Y(new_n20735));
  INVx1_ASAP7_75t_L         g20479(.A(new_n20735), .Y(new_n20736));
  NAND2xp33_ASAP7_75t_L     g20480(.A(new_n20736), .B(new_n20732), .Y(new_n20737));
  AND2x2_ASAP7_75t_L        g20481(.A(new_n20737), .B(new_n20734), .Y(new_n20738));
  A2O1A1Ixp33_ASAP7_75t_L   g20482(.A1(new_n20680), .A2(\a[53] ), .B(new_n20681), .C(new_n20738), .Y(new_n20739));
  NOR2xp33_ASAP7_75t_L      g20483(.A(new_n9099), .B(new_n20679), .Y(new_n20740));
  OR3x1_ASAP7_75t_L         g20484(.A(new_n20738), .B(new_n20740), .C(new_n20681), .Y(new_n20741));
  AND2x2_ASAP7_75t_L        g20485(.A(new_n20739), .B(new_n20741), .Y(new_n20742));
  INVx1_ASAP7_75t_L         g20486(.A(new_n20742), .Y(new_n20743));
  O2A1O1Ixp33_ASAP7_75t_L   g20487(.A1(new_n20543), .A2(new_n20538), .B(new_n20553), .C(new_n20743), .Y(new_n20744));
  INVx1_ASAP7_75t_L         g20488(.A(new_n20744), .Y(new_n20745));
  NAND3xp33_ASAP7_75t_L     g20489(.A(new_n20743), .B(new_n20553), .C(new_n20540), .Y(new_n20746));
  AND2x2_ASAP7_75t_L        g20490(.A(new_n20746), .B(new_n20745), .Y(new_n20747));
  INVx1_ASAP7_75t_L         g20491(.A(new_n20747), .Y(new_n20748));
  NOR2xp33_ASAP7_75t_L      g20492(.A(new_n7270), .B(new_n10065), .Y(new_n20749));
  AOI221xp5_ASAP7_75t_L     g20493(.A1(new_n8175), .A2(\b[47] ), .B1(new_n8484), .B2(\b[45] ), .C(new_n20749), .Y(new_n20750));
  O2A1O1Ixp33_ASAP7_75t_L   g20494(.A1(new_n8176), .A2(new_n7560), .B(new_n20750), .C(new_n8172), .Y(new_n20751));
  O2A1O1Ixp33_ASAP7_75t_L   g20495(.A1(new_n8176), .A2(new_n7560), .B(new_n20750), .C(\a[50] ), .Y(new_n20752));
  INVx1_ASAP7_75t_L         g20496(.A(new_n20752), .Y(new_n20753));
  O2A1O1Ixp33_ASAP7_75t_L   g20497(.A1(new_n20751), .A2(new_n8172), .B(new_n20753), .C(new_n20748), .Y(new_n20754));
  INVx1_ASAP7_75t_L         g20498(.A(new_n20754), .Y(new_n20755));
  O2A1O1Ixp33_ASAP7_75t_L   g20499(.A1(new_n20751), .A2(new_n8172), .B(new_n20753), .C(new_n20747), .Y(new_n20756));
  AOI21xp33_ASAP7_75t_L     g20500(.A1(new_n20755), .A2(new_n20747), .B(new_n20756), .Y(new_n20757));
  O2A1O1Ixp33_ASAP7_75t_L   g20501(.A1(new_n20490), .A2(new_n20558), .B(new_n20555), .C(new_n20569), .Y(new_n20758));
  NAND2xp33_ASAP7_75t_L     g20502(.A(new_n20758), .B(new_n20757), .Y(new_n20759));
  INVx1_ASAP7_75t_L         g20503(.A(new_n20758), .Y(new_n20760));
  A2O1A1Ixp33_ASAP7_75t_L   g20504(.A1(new_n20755), .A2(new_n20747), .B(new_n20756), .C(new_n20760), .Y(new_n20761));
  AND2x2_ASAP7_75t_L        g20505(.A(new_n20761), .B(new_n20759), .Y(new_n20762));
  NOR2xp33_ASAP7_75t_L      g20506(.A(new_n8755), .B(new_n7318), .Y(new_n20763));
  AOI221xp5_ASAP7_75t_L     g20507(.A1(new_n7333), .A2(\b[49] ), .B1(new_n7609), .B2(\b[48] ), .C(new_n20763), .Y(new_n20764));
  O2A1O1Ixp33_ASAP7_75t_L   g20508(.A1(new_n7321), .A2(new_n8764), .B(new_n20764), .C(new_n7316), .Y(new_n20765));
  INVx1_ASAP7_75t_L         g20509(.A(new_n20765), .Y(new_n20766));
  O2A1O1Ixp33_ASAP7_75t_L   g20510(.A1(new_n7321), .A2(new_n8764), .B(new_n20764), .C(\a[47] ), .Y(new_n20767));
  AOI211xp5_ASAP7_75t_L     g20511(.A1(new_n20766), .A2(\a[47] ), .B(new_n20767), .C(new_n20762), .Y(new_n20768));
  A2O1A1Ixp33_ASAP7_75t_L   g20512(.A1(\a[47] ), .A2(new_n20766), .B(new_n20767), .C(new_n20762), .Y(new_n20769));
  INVx1_ASAP7_75t_L         g20513(.A(new_n20769), .Y(new_n20770));
  NOR2xp33_ASAP7_75t_L      g20514(.A(new_n20768), .B(new_n20770), .Y(new_n20771));
  NAND2xp33_ASAP7_75t_L     g20515(.A(new_n20676), .B(new_n20771), .Y(new_n20772));
  NOR2xp33_ASAP7_75t_L      g20516(.A(new_n8779), .B(new_n6741), .Y(new_n20773));
  AOI221xp5_ASAP7_75t_L     g20517(.A1(\b[53] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[52] ), .C(new_n20773), .Y(new_n20774));
  O2A1O1Ixp33_ASAP7_75t_L   g20518(.A1(new_n6443), .A2(new_n9691), .B(new_n20774), .C(new_n6439), .Y(new_n20775));
  INVx1_ASAP7_75t_L         g20519(.A(new_n20775), .Y(new_n20776));
  O2A1O1Ixp33_ASAP7_75t_L   g20520(.A1(new_n6443), .A2(new_n9691), .B(new_n20774), .C(\a[44] ), .Y(new_n20777));
  A2O1A1O1Ixp25_ASAP7_75t_L g20521(.A1(new_n20573), .A2(new_n20571), .B(new_n20574), .C(new_n20584), .D(new_n20771), .Y(new_n20778));
  INVx1_ASAP7_75t_L         g20522(.A(new_n20778), .Y(new_n20779));
  NAND2xp33_ASAP7_75t_L     g20523(.A(new_n20675), .B(new_n20771), .Y(new_n20780));
  NAND2xp33_ASAP7_75t_L     g20524(.A(new_n20780), .B(new_n20779), .Y(new_n20781));
  A2O1A1Ixp33_ASAP7_75t_L   g20525(.A1(new_n20776), .A2(\a[44] ), .B(new_n20777), .C(new_n20781), .Y(new_n20782));
  AOI21xp33_ASAP7_75t_L     g20526(.A1(new_n20776), .A2(\a[44] ), .B(new_n20777), .Y(new_n20783));
  NAND2xp33_ASAP7_75t_L     g20527(.A(new_n20783), .B(new_n20780), .Y(new_n20784));
  A2O1A1Ixp33_ASAP7_75t_L   g20528(.A1(new_n20676), .A2(new_n20772), .B(new_n20784), .C(new_n20782), .Y(new_n20785));
  A2O1A1O1Ixp25_ASAP7_75t_L g20529(.A1(new_n20489), .A2(new_n20387), .B(new_n20588), .C(new_n20596), .D(new_n20785), .Y(new_n20786));
  A2O1A1Ixp33_ASAP7_75t_L   g20530(.A1(new_n20489), .A2(new_n20387), .B(new_n20588), .C(new_n20596), .Y(new_n20787));
  O2A1O1Ixp33_ASAP7_75t_L   g20531(.A1(new_n20784), .A2(new_n20778), .B(new_n20782), .C(new_n20787), .Y(new_n20788));
  NOR2xp33_ASAP7_75t_L      g20532(.A(new_n20788), .B(new_n20786), .Y(new_n20789));
  XNOR2x2_ASAP7_75t_L       g20533(.A(new_n20674), .B(new_n20789), .Y(new_n20790));
  INVx1_ASAP7_75t_L         g20534(.A(new_n20790), .Y(new_n20791));
  A2O1A1O1Ixp25_ASAP7_75t_L g20535(.A1(new_n20602), .A2(new_n20600), .B(new_n20609), .C(new_n20667), .D(new_n20791), .Y(new_n20792));
  INVx1_ASAP7_75t_L         g20536(.A(new_n20792), .Y(new_n20793));
  O2A1O1Ixp33_ASAP7_75t_L   g20537(.A1(new_n20607), .A2(new_n20608), .B(new_n20603), .C(new_n20666), .Y(new_n20794));
  NAND2xp33_ASAP7_75t_L     g20538(.A(new_n20794), .B(new_n20791), .Y(new_n20795));
  NAND2xp33_ASAP7_75t_L     g20539(.A(new_n20795), .B(new_n20793), .Y(new_n20796));
  NOR2xp33_ASAP7_75t_L      g20540(.A(new_n11591), .B(new_n4908), .Y(new_n20797));
  AOI221xp5_ASAP7_75t_L     g20541(.A1(\b[57] ), .A2(new_n5139), .B1(\b[58] ), .B2(new_n4916), .C(new_n20797), .Y(new_n20798));
  O2A1O1Ixp33_ASAP7_75t_L   g20542(.A1(new_n4911), .A2(new_n11597), .B(new_n20798), .C(new_n4906), .Y(new_n20799));
  O2A1O1Ixp33_ASAP7_75t_L   g20543(.A1(new_n4911), .A2(new_n11597), .B(new_n20798), .C(\a[38] ), .Y(new_n20800));
  INVx1_ASAP7_75t_L         g20544(.A(new_n20800), .Y(new_n20801));
  O2A1O1Ixp33_ASAP7_75t_L   g20545(.A1(new_n20799), .A2(new_n4906), .B(new_n20801), .C(new_n20796), .Y(new_n20802));
  INVx1_ASAP7_75t_L         g20546(.A(new_n20799), .Y(new_n20803));
  A2O1A1Ixp33_ASAP7_75t_L   g20547(.A1(\a[38] ), .A2(new_n20803), .B(new_n20800), .C(new_n20796), .Y(new_n20804));
  OAI21xp33_ASAP7_75t_L     g20548(.A1(new_n20796), .A2(new_n20802), .B(new_n20804), .Y(new_n20805));
  AOI211xp5_ASAP7_75t_L     g20549(.A1(new_n20664), .A2(new_n20610), .B(new_n20623), .C(new_n20805), .Y(new_n20806));
  A2O1A1O1Ixp25_ASAP7_75t_L g20550(.A1(new_n20290), .A2(new_n20417), .B(new_n20416), .C(new_n20610), .D(new_n20623), .Y(new_n20807));
  O2A1O1Ixp33_ASAP7_75t_L   g20551(.A1(new_n20796), .A2(new_n20802), .B(new_n20804), .C(new_n20807), .Y(new_n20808));
  NOR2xp33_ASAP7_75t_L      g20552(.A(new_n20808), .B(new_n20806), .Y(new_n20809));
  NOR2xp33_ASAP7_75t_L      g20553(.A(new_n12258), .B(new_n4142), .Y(new_n20810));
  AOI221xp5_ASAP7_75t_L     g20554(.A1(\b[60] ), .A2(new_n4402), .B1(\b[62] ), .B2(new_n4156), .C(new_n20810), .Y(new_n20811));
  O2A1O1Ixp33_ASAP7_75t_L   g20555(.A1(new_n4150), .A2(new_n12610), .B(new_n20811), .C(new_n4145), .Y(new_n20812));
  INVx1_ASAP7_75t_L         g20556(.A(new_n20812), .Y(new_n20813));
  O2A1O1Ixp33_ASAP7_75t_L   g20557(.A1(new_n4150), .A2(new_n12610), .B(new_n20811), .C(\a[35] ), .Y(new_n20814));
  A2O1A1Ixp33_ASAP7_75t_L   g20558(.A1(\a[35] ), .A2(new_n20813), .B(new_n20814), .C(new_n20809), .Y(new_n20815));
  INVx1_ASAP7_75t_L         g20559(.A(new_n20814), .Y(new_n20816));
  O2A1O1Ixp33_ASAP7_75t_L   g20560(.A1(new_n20812), .A2(new_n4145), .B(new_n20816), .C(new_n20809), .Y(new_n20817));
  AOI21xp33_ASAP7_75t_L     g20561(.A1(new_n20815), .A2(new_n20809), .B(new_n20817), .Y(new_n20818));
  A2O1A1Ixp33_ASAP7_75t_L   g20562(.A1(new_n20662), .A2(new_n20656), .B(new_n20663), .C(new_n20818), .Y(new_n20819));
  INVx1_ASAP7_75t_L         g20563(.A(new_n20663), .Y(new_n20820));
  A2O1A1Ixp33_ASAP7_75t_L   g20564(.A1(new_n20637), .A2(new_n20630), .B(new_n20661), .C(new_n20820), .Y(new_n20821));
  INVx1_ASAP7_75t_L         g20565(.A(new_n20821), .Y(new_n20822));
  A2O1A1Ixp33_ASAP7_75t_L   g20566(.A1(new_n20809), .A2(new_n20815), .B(new_n20817), .C(new_n20822), .Y(new_n20823));
  A2O1A1Ixp33_ASAP7_75t_L   g20567(.A1(new_n20257), .A2(new_n20126), .B(new_n20264), .C(new_n20444), .Y(new_n20824));
  A2O1A1Ixp33_ASAP7_75t_L   g20568(.A1(new_n20824), .A2(new_n20440), .B(new_n20484), .C(new_n20640), .Y(new_n20825));
  XNOR2x2_ASAP7_75t_L       g20569(.A(new_n20821), .B(new_n20818), .Y(new_n20826));
  NAND2xp33_ASAP7_75t_L     g20570(.A(new_n20825), .B(new_n20826), .Y(new_n20827));
  INVx1_ASAP7_75t_L         g20571(.A(new_n20827), .Y(new_n20828));
  A2O1A1O1Ixp25_ASAP7_75t_L g20572(.A1(new_n20257), .A2(new_n20126), .B(new_n20264), .C(new_n20444), .D(new_n20451), .Y(new_n20829));
  O2A1O1Ixp33_ASAP7_75t_L   g20573(.A1(new_n20829), .A2(new_n20484), .B(new_n20640), .C(new_n20826), .Y(new_n20830));
  INVx1_ASAP7_75t_L         g20574(.A(new_n20830), .Y(new_n20831));
  A2O1A1Ixp33_ASAP7_75t_L   g20575(.A1(new_n20823), .A2(new_n20819), .B(new_n20828), .C(new_n20831), .Y(new_n20832));
  A2O1A1Ixp33_ASAP7_75t_L   g20576(.A1(new_n20472), .A2(new_n20650), .B(new_n20652), .C(new_n20644), .Y(new_n20833));
  AOI211xp5_ASAP7_75t_L     g20577(.A1(new_n20826), .A2(new_n20827), .B(new_n20830), .C(new_n20833), .Y(new_n20834));
  O2A1O1Ixp33_ASAP7_75t_L   g20578(.A1(new_n20645), .A2(new_n20649), .B(new_n20832), .C(new_n20834), .Y(\f[95] ));
  O2A1O1Ixp33_ASAP7_75t_L   g20579(.A1(new_n20830), .A2(new_n20826), .B(new_n20833), .C(new_n20828), .Y(new_n20836));
  A2O1A1O1Ixp25_ASAP7_75t_L g20580(.A1(new_n3505), .A2(new_n14172), .B(new_n3708), .C(\b[63] ), .D(new_n3493), .Y(new_n20837));
  A2O1A1O1Ixp25_ASAP7_75t_L g20581(.A1(new_n12986), .A2(new_n3505), .B(new_n20657), .C(new_n20658), .D(new_n20837), .Y(new_n20838));
  A2O1A1Ixp33_ASAP7_75t_L   g20582(.A1(new_n20809), .A2(new_n20815), .B(new_n20817), .C(new_n20821), .Y(new_n20839));
  A2O1A1O1Ixp25_ASAP7_75t_L g20583(.A1(new_n20755), .A2(new_n20747), .B(new_n20756), .C(new_n20760), .D(new_n20770), .Y(new_n20840));
  NOR2xp33_ASAP7_75t_L      g20584(.A(new_n3891), .B(new_n13030), .Y(new_n20841));
  A2O1A1Ixp33_ASAP7_75t_L   g20585(.A1(new_n13028), .A2(\b[33] ), .B(new_n20841), .C(new_n3493), .Y(new_n20842));
  O2A1O1Ixp33_ASAP7_75t_L   g20586(.A1(new_n12669), .A2(new_n12671), .B(\b[33] ), .C(new_n20841), .Y(new_n20843));
  NAND2xp33_ASAP7_75t_L     g20587(.A(\a[32] ), .B(new_n20843), .Y(new_n20844));
  NAND2xp33_ASAP7_75t_L     g20588(.A(new_n20842), .B(new_n20844), .Y(new_n20845));
  O2A1O1Ixp33_ASAP7_75t_L   g20589(.A1(new_n3891), .A2(new_n12672), .B(new_n20694), .C(new_n20845), .Y(new_n20846));
  A2O1A1Ixp33_ASAP7_75t_L   g20590(.A1(new_n13028), .A2(\b[32] ), .B(new_n20693), .C(new_n20845), .Y(new_n20847));
  OAI21xp33_ASAP7_75t_L     g20591(.A1(new_n20845), .A2(new_n20846), .B(new_n20847), .Y(new_n20848));
  A2O1A1Ixp33_ASAP7_75t_L   g20592(.A1(new_n20697), .A2(new_n20692), .B(new_n20699), .C(new_n20848), .Y(new_n20849));
  O2A1O1Ixp33_ASAP7_75t_L   g20593(.A1(new_n20845), .A2(new_n20846), .B(new_n20847), .C(new_n20702), .Y(new_n20850));
  A2O1A1O1Ixp25_ASAP7_75t_L g20594(.A1(new_n20697), .A2(new_n20692), .B(new_n20699), .C(new_n20849), .D(new_n20850), .Y(new_n20851));
  NAND2xp33_ASAP7_75t_L     g20595(.A(\b[36] ), .B(new_n11995), .Y(new_n20852));
  OAI221xp5_ASAP7_75t_L     g20596(.A1(new_n12318), .A2(new_n4581), .B1(new_n4344), .B2(new_n12320), .C(new_n20852), .Y(new_n20853));
  A2O1A1Ixp33_ASAP7_75t_L   g20597(.A1(new_n4621), .A2(new_n11997), .B(new_n20853), .C(\a[62] ), .Y(new_n20854));
  NAND2xp33_ASAP7_75t_L     g20598(.A(\a[62] ), .B(new_n20854), .Y(new_n20855));
  A2O1A1Ixp33_ASAP7_75t_L   g20599(.A1(new_n4621), .A2(new_n11997), .B(new_n20853), .C(new_n11987), .Y(new_n20856));
  NAND2xp33_ASAP7_75t_L     g20600(.A(new_n20856), .B(new_n20855), .Y(new_n20857));
  XOR2x2_ASAP7_75t_L        g20601(.A(new_n20857), .B(new_n20851), .Y(new_n20858));
  INVx1_ASAP7_75t_L         g20602(.A(new_n20858), .Y(new_n20859));
  NOR2xp33_ASAP7_75t_L      g20603(.A(new_n5074), .B(new_n11354), .Y(new_n20860));
  AOI221xp5_ASAP7_75t_L     g20604(.A1(\b[39] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[38] ), .C(new_n20860), .Y(new_n20861));
  O2A1O1Ixp33_ASAP7_75t_L   g20605(.A1(new_n11053), .A2(new_n5578), .B(new_n20861), .C(new_n11048), .Y(new_n20862));
  INVx1_ASAP7_75t_L         g20606(.A(new_n20862), .Y(new_n20863));
  O2A1O1Ixp33_ASAP7_75t_L   g20607(.A1(new_n11053), .A2(new_n5578), .B(new_n20861), .C(\a[59] ), .Y(new_n20864));
  A2O1A1Ixp33_ASAP7_75t_L   g20608(.A1(\a[59] ), .A2(new_n20863), .B(new_n20864), .C(new_n20859), .Y(new_n20865));
  AOI21xp33_ASAP7_75t_L     g20609(.A1(new_n20863), .A2(\a[59] ), .B(new_n20864), .Y(new_n20866));
  NAND2xp33_ASAP7_75t_L     g20610(.A(new_n20866), .B(new_n20858), .Y(new_n20867));
  NAND2xp33_ASAP7_75t_L     g20611(.A(new_n20867), .B(new_n20865), .Y(new_n20868));
  O2A1O1Ixp33_ASAP7_75t_L   g20612(.A1(new_n20717), .A2(new_n20711), .B(new_n20704), .C(new_n20868), .Y(new_n20869));
  INVx1_ASAP7_75t_L         g20613(.A(new_n20869), .Y(new_n20870));
  OAI211xp5_ASAP7_75t_L     g20614(.A1(new_n20717), .A2(new_n20711), .B(new_n20868), .C(new_n20704), .Y(new_n20871));
  AND2x2_ASAP7_75t_L        g20615(.A(new_n20871), .B(new_n20870), .Y(new_n20872));
  INVx1_ASAP7_75t_L         g20616(.A(new_n20872), .Y(new_n20873));
  NOR2xp33_ASAP7_75t_L      g20617(.A(new_n6110), .B(new_n10388), .Y(new_n20874));
  AOI221xp5_ASAP7_75t_L     g20618(.A1(new_n10086), .A2(\b[42] ), .B1(new_n11361), .B2(\b[40] ), .C(new_n20874), .Y(new_n20875));
  O2A1O1Ixp33_ASAP7_75t_L   g20619(.A1(new_n10088), .A2(new_n6386), .B(new_n20875), .C(new_n10083), .Y(new_n20876));
  O2A1O1Ixp33_ASAP7_75t_L   g20620(.A1(new_n10088), .A2(new_n6386), .B(new_n20875), .C(\a[56] ), .Y(new_n20877));
  INVx1_ASAP7_75t_L         g20621(.A(new_n20877), .Y(new_n20878));
  O2A1O1Ixp33_ASAP7_75t_L   g20622(.A1(new_n20876), .A2(new_n10083), .B(new_n20878), .C(new_n20873), .Y(new_n20879));
  INVx1_ASAP7_75t_L         g20623(.A(new_n20879), .Y(new_n20880));
  O2A1O1Ixp33_ASAP7_75t_L   g20624(.A1(new_n20876), .A2(new_n10083), .B(new_n20878), .C(new_n20872), .Y(new_n20881));
  AOI21xp33_ASAP7_75t_L     g20625(.A1(new_n20880), .A2(new_n20872), .B(new_n20881), .Y(new_n20882));
  A2O1A1Ixp33_ASAP7_75t_L   g20626(.A1(new_n20712), .A2(new_n20718), .B(new_n20724), .C(new_n20727), .Y(new_n20883));
  INVx1_ASAP7_75t_L         g20627(.A(new_n20883), .Y(new_n20884));
  NAND2xp33_ASAP7_75t_L     g20628(.A(new_n20884), .B(new_n20882), .Y(new_n20885));
  O2A1O1Ixp33_ASAP7_75t_L   g20629(.A1(new_n20724), .A2(new_n20719), .B(new_n20727), .C(new_n20882), .Y(new_n20886));
  INVx1_ASAP7_75t_L         g20630(.A(new_n20886), .Y(new_n20887));
  AND2x2_ASAP7_75t_L        g20631(.A(new_n20885), .B(new_n20887), .Y(new_n20888));
  INVx1_ASAP7_75t_L         g20632(.A(new_n20888), .Y(new_n20889));
  NOR2xp33_ASAP7_75t_L      g20633(.A(new_n6944), .B(new_n10400), .Y(new_n20890));
  AOI221xp5_ASAP7_75t_L     g20634(.A1(new_n9102), .A2(\b[45] ), .B1(new_n10398), .B2(\b[43] ), .C(new_n20890), .Y(new_n20891));
  O2A1O1Ixp33_ASAP7_75t_L   g20635(.A1(new_n9104), .A2(new_n7255), .B(new_n20891), .C(new_n9099), .Y(new_n20892));
  O2A1O1Ixp33_ASAP7_75t_L   g20636(.A1(new_n9104), .A2(new_n7255), .B(new_n20891), .C(\a[53] ), .Y(new_n20893));
  INVx1_ASAP7_75t_L         g20637(.A(new_n20893), .Y(new_n20894));
  O2A1O1Ixp33_ASAP7_75t_L   g20638(.A1(new_n20892), .A2(new_n9099), .B(new_n20894), .C(new_n20889), .Y(new_n20895));
  INVx1_ASAP7_75t_L         g20639(.A(new_n20895), .Y(new_n20896));
  O2A1O1Ixp33_ASAP7_75t_L   g20640(.A1(new_n20892), .A2(new_n9099), .B(new_n20894), .C(new_n20888), .Y(new_n20897));
  AOI21xp33_ASAP7_75t_L     g20641(.A1(new_n20896), .A2(new_n20888), .B(new_n20897), .Y(new_n20898));
  O2A1O1Ixp33_ASAP7_75t_L   g20642(.A1(new_n20681), .A2(new_n20740), .B(new_n20737), .C(new_n20733), .Y(new_n20899));
  NAND2xp33_ASAP7_75t_L     g20643(.A(new_n20899), .B(new_n20898), .Y(new_n20900));
  O2A1O1Ixp33_ASAP7_75t_L   g20644(.A1(new_n20736), .A2(new_n20732), .B(new_n20739), .C(new_n20898), .Y(new_n20901));
  INVx1_ASAP7_75t_L         g20645(.A(new_n20901), .Y(new_n20902));
  AND2x2_ASAP7_75t_L        g20646(.A(new_n20900), .B(new_n20902), .Y(new_n20903));
  INVx1_ASAP7_75t_L         g20647(.A(new_n20903), .Y(new_n20904));
  NOR2xp33_ASAP7_75t_L      g20648(.A(new_n7552), .B(new_n10065), .Y(new_n20905));
  AOI221xp5_ASAP7_75t_L     g20649(.A1(new_n8175), .A2(\b[48] ), .B1(new_n8484), .B2(\b[46] ), .C(new_n20905), .Y(new_n20906));
  O2A1O1Ixp33_ASAP7_75t_L   g20650(.A1(new_n8176), .A2(new_n7868), .B(new_n20906), .C(new_n8172), .Y(new_n20907));
  O2A1O1Ixp33_ASAP7_75t_L   g20651(.A1(new_n8176), .A2(new_n7868), .B(new_n20906), .C(\a[50] ), .Y(new_n20908));
  INVx1_ASAP7_75t_L         g20652(.A(new_n20908), .Y(new_n20909));
  O2A1O1Ixp33_ASAP7_75t_L   g20653(.A1(new_n20907), .A2(new_n8172), .B(new_n20909), .C(new_n20904), .Y(new_n20910));
  INVx1_ASAP7_75t_L         g20654(.A(new_n20910), .Y(new_n20911));
  O2A1O1Ixp33_ASAP7_75t_L   g20655(.A1(new_n20907), .A2(new_n8172), .B(new_n20909), .C(new_n20903), .Y(new_n20912));
  AOI21xp33_ASAP7_75t_L     g20656(.A1(new_n20911), .A2(new_n20903), .B(new_n20912), .Y(new_n20913));
  O2A1O1Ixp33_ASAP7_75t_L   g20657(.A1(new_n20539), .A2(new_n20552), .B(new_n20742), .C(new_n20754), .Y(new_n20914));
  AND2x2_ASAP7_75t_L        g20658(.A(new_n20914), .B(new_n20913), .Y(new_n20915));
  A2O1A1O1Ixp25_ASAP7_75t_L g20659(.A1(new_n20553), .A2(new_n20540), .B(new_n20743), .C(new_n20755), .D(new_n20913), .Y(new_n20916));
  NOR2xp33_ASAP7_75t_L      g20660(.A(new_n20916), .B(new_n20915), .Y(new_n20917));
  NOR2xp33_ASAP7_75t_L      g20661(.A(new_n8779), .B(new_n7318), .Y(new_n20918));
  AOI221xp5_ASAP7_75t_L     g20662(.A1(new_n7333), .A2(\b[50] ), .B1(new_n7609), .B2(\b[49] ), .C(new_n20918), .Y(new_n20919));
  O2A1O1Ixp33_ASAP7_75t_L   g20663(.A1(new_n7321), .A2(new_n8789), .B(new_n20919), .C(new_n7316), .Y(new_n20920));
  INVx1_ASAP7_75t_L         g20664(.A(new_n20920), .Y(new_n20921));
  O2A1O1Ixp33_ASAP7_75t_L   g20665(.A1(new_n7321), .A2(new_n8789), .B(new_n20919), .C(\a[47] ), .Y(new_n20922));
  A2O1A1Ixp33_ASAP7_75t_L   g20666(.A1(\a[47] ), .A2(new_n20921), .B(new_n20922), .C(new_n20917), .Y(new_n20923));
  INVx1_ASAP7_75t_L         g20667(.A(new_n20919), .Y(new_n20924));
  NOR2xp33_ASAP7_75t_L      g20668(.A(new_n7316), .B(new_n20920), .Y(new_n20925));
  A2O1A1O1Ixp25_ASAP7_75t_L g20669(.A1(new_n8790), .A2(new_n7322), .B(new_n20924), .C(new_n20921), .D(new_n20925), .Y(new_n20926));
  INVx1_ASAP7_75t_L         g20670(.A(new_n20926), .Y(new_n20927));
  NOR2xp33_ASAP7_75t_L      g20671(.A(new_n20927), .B(new_n20917), .Y(new_n20928));
  O2A1O1Ixp33_ASAP7_75t_L   g20672(.A1(new_n20757), .A2(new_n20758), .B(new_n20769), .C(new_n20928), .Y(new_n20929));
  NAND2xp33_ASAP7_75t_L     g20673(.A(new_n20914), .B(new_n20913), .Y(new_n20930));
  INVx1_ASAP7_75t_L         g20674(.A(new_n20916), .Y(new_n20931));
  O2A1O1Ixp33_ASAP7_75t_L   g20675(.A1(new_n20925), .A2(new_n20922), .B(new_n20917), .C(new_n20929), .Y(new_n20932));
  A2O1A1Ixp33_ASAP7_75t_L   g20676(.A1(new_n20931), .A2(new_n20930), .B(new_n20927), .C(new_n20932), .Y(new_n20933));
  A2O1A1Ixp33_ASAP7_75t_L   g20677(.A1(new_n20923), .A2(new_n20929), .B(new_n20840), .C(new_n20933), .Y(new_n20934));
  INVx1_ASAP7_75t_L         g20678(.A(new_n20934), .Y(new_n20935));
  NOR2xp33_ASAP7_75t_L      g20679(.A(new_n9355), .B(new_n6741), .Y(new_n20936));
  AOI221xp5_ASAP7_75t_L     g20680(.A1(\b[54] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[53] ), .C(new_n20936), .Y(new_n20937));
  O2A1O1Ixp33_ASAP7_75t_L   g20681(.A1(new_n6443), .A2(new_n9718), .B(new_n20937), .C(new_n6439), .Y(new_n20938));
  O2A1O1Ixp33_ASAP7_75t_L   g20682(.A1(new_n6443), .A2(new_n9718), .B(new_n20937), .C(\a[44] ), .Y(new_n20939));
  INVx1_ASAP7_75t_L         g20683(.A(new_n20939), .Y(new_n20940));
  OAI211xp5_ASAP7_75t_L     g20684(.A1(new_n6439), .A2(new_n20938), .B(new_n20935), .C(new_n20940), .Y(new_n20941));
  O2A1O1Ixp33_ASAP7_75t_L   g20685(.A1(new_n20938), .A2(new_n6439), .B(new_n20940), .C(new_n20935), .Y(new_n20942));
  INVx1_ASAP7_75t_L         g20686(.A(new_n20942), .Y(new_n20943));
  AND2x2_ASAP7_75t_L        g20687(.A(new_n20941), .B(new_n20943), .Y(new_n20944));
  INVx1_ASAP7_75t_L         g20688(.A(new_n20944), .Y(new_n20945));
  A2O1A1O1Ixp25_ASAP7_75t_L g20689(.A1(new_n20779), .A2(new_n20780), .B(new_n20783), .C(new_n20772), .D(new_n20945), .Y(new_n20946));
  INVx1_ASAP7_75t_L         g20690(.A(new_n20946), .Y(new_n20947));
  NAND3xp33_ASAP7_75t_L     g20691(.A(new_n20945), .B(new_n20782), .C(new_n20772), .Y(new_n20948));
  NAND2xp33_ASAP7_75t_L     g20692(.A(new_n20948), .B(new_n20947), .Y(new_n20949));
  NOR2xp33_ASAP7_75t_L      g20693(.A(new_n10332), .B(new_n5640), .Y(new_n20950));
  AOI221xp5_ASAP7_75t_L     g20694(.A1(\b[55] ), .A2(new_n5920), .B1(\b[57] ), .B2(new_n5629), .C(new_n20950), .Y(new_n20951));
  O2A1O1Ixp33_ASAP7_75t_L   g20695(.A1(new_n5630), .A2(new_n17096), .B(new_n20951), .C(new_n5626), .Y(new_n20952));
  O2A1O1Ixp33_ASAP7_75t_L   g20696(.A1(new_n5630), .A2(new_n17096), .B(new_n20951), .C(\a[41] ), .Y(new_n20953));
  INVx1_ASAP7_75t_L         g20697(.A(new_n20953), .Y(new_n20954));
  O2A1O1Ixp33_ASAP7_75t_L   g20698(.A1(new_n20952), .A2(new_n5626), .B(new_n20954), .C(new_n20949), .Y(new_n20955));
  INVx1_ASAP7_75t_L         g20699(.A(new_n20949), .Y(new_n20956));
  O2A1O1Ixp33_ASAP7_75t_L   g20700(.A1(new_n20952), .A2(new_n5626), .B(new_n20954), .C(new_n20956), .Y(new_n20957));
  INVx1_ASAP7_75t_L         g20701(.A(new_n20957), .Y(new_n20958));
  O2A1O1Ixp33_ASAP7_75t_L   g20702(.A1(new_n5630), .A2(new_n10339), .B(new_n20669), .C(\a[41] ), .Y(new_n20959));
  O2A1O1Ixp33_ASAP7_75t_L   g20703(.A1(new_n20959), .A2(new_n20673), .B(new_n20789), .C(new_n20786), .Y(new_n20960));
  OAI211xp5_ASAP7_75t_L     g20704(.A1(new_n20949), .A2(new_n20955), .B(new_n20958), .C(new_n20960), .Y(new_n20961));
  INVx1_ASAP7_75t_L         g20705(.A(new_n20955), .Y(new_n20962));
  INVx1_ASAP7_75t_L         g20706(.A(new_n20960), .Y(new_n20963));
  A2O1A1Ixp33_ASAP7_75t_L   g20707(.A1(new_n20962), .A2(new_n20956), .B(new_n20957), .C(new_n20963), .Y(new_n20964));
  NAND2xp33_ASAP7_75t_L     g20708(.A(new_n20964), .B(new_n20961), .Y(new_n20965));
  NOR2xp33_ASAP7_75t_L      g20709(.A(new_n11626), .B(new_n4908), .Y(new_n20966));
  AOI221xp5_ASAP7_75t_L     g20710(.A1(\b[58] ), .A2(new_n5139), .B1(\b[59] ), .B2(new_n4916), .C(new_n20966), .Y(new_n20967));
  O2A1O1Ixp33_ASAP7_75t_L   g20711(.A1(new_n4911), .A2(new_n11634), .B(new_n20967), .C(new_n4906), .Y(new_n20968));
  NOR2xp33_ASAP7_75t_L      g20712(.A(new_n4906), .B(new_n20968), .Y(new_n20969));
  O2A1O1Ixp33_ASAP7_75t_L   g20713(.A1(new_n4911), .A2(new_n11634), .B(new_n20967), .C(\a[38] ), .Y(new_n20970));
  OAI211xp5_ASAP7_75t_L     g20714(.A1(new_n20969), .A2(new_n20970), .B(new_n20961), .C(new_n20964), .Y(new_n20971));
  INVx1_ASAP7_75t_L         g20715(.A(new_n20971), .Y(new_n20972));
  INVx1_ASAP7_75t_L         g20716(.A(new_n20968), .Y(new_n20973));
  A2O1A1Ixp33_ASAP7_75t_L   g20717(.A1(\a[38] ), .A2(new_n20973), .B(new_n20970), .C(new_n20965), .Y(new_n20974));
  OAI21xp33_ASAP7_75t_L     g20718(.A1(new_n20965), .A2(new_n20972), .B(new_n20974), .Y(new_n20975));
  A2O1A1O1Ixp25_ASAP7_75t_L g20719(.A1(new_n20803), .A2(\a[38] ), .B(new_n20800), .C(new_n20795), .D(new_n20792), .Y(new_n20976));
  INVx1_ASAP7_75t_L         g20720(.A(new_n20976), .Y(new_n20977));
  NOR2xp33_ASAP7_75t_L      g20721(.A(new_n20977), .B(new_n20975), .Y(new_n20978));
  O2A1O1Ixp33_ASAP7_75t_L   g20722(.A1(new_n20965), .A2(new_n20972), .B(new_n20974), .C(new_n20976), .Y(new_n20979));
  NOR2xp33_ASAP7_75t_L      g20723(.A(new_n20979), .B(new_n20978), .Y(new_n20980));
  INVx1_ASAP7_75t_L         g20724(.A(new_n20980), .Y(new_n20981));
  NOR2xp33_ASAP7_75t_L      g20725(.A(new_n12603), .B(new_n4142), .Y(new_n20982));
  AOI221xp5_ASAP7_75t_L     g20726(.A1(\b[61] ), .A2(new_n4402), .B1(\b[63] ), .B2(new_n4156), .C(new_n20982), .Y(new_n20983));
  O2A1O1Ixp33_ASAP7_75t_L   g20727(.A1(new_n4150), .A2(new_n17815), .B(new_n20983), .C(new_n4145), .Y(new_n20984));
  INVx1_ASAP7_75t_L         g20728(.A(new_n20984), .Y(new_n20985));
  O2A1O1Ixp33_ASAP7_75t_L   g20729(.A1(new_n4150), .A2(new_n17815), .B(new_n20983), .C(\a[35] ), .Y(new_n20986));
  INVx1_ASAP7_75t_L         g20730(.A(new_n20808), .Y(new_n20987));
  NAND2xp33_ASAP7_75t_L     g20731(.A(\a[35] ), .B(new_n20813), .Y(new_n20988));
  AOI21xp33_ASAP7_75t_L     g20732(.A1(new_n20985), .A2(\a[35] ), .B(new_n20986), .Y(new_n20989));
  A2O1A1O1Ixp25_ASAP7_75t_L g20733(.A1(new_n20988), .A2(new_n20816), .B(new_n20806), .C(new_n20987), .D(new_n20989), .Y(new_n20990));
  INVx1_ASAP7_75t_L         g20734(.A(new_n20990), .Y(new_n20991));
  A2O1A1O1Ixp25_ASAP7_75t_L g20735(.A1(new_n20988), .A2(new_n20816), .B(new_n20806), .C(new_n20987), .D(new_n20990), .Y(new_n20992));
  A2O1A1O1Ixp25_ASAP7_75t_L g20736(.A1(new_n20985), .A2(\a[35] ), .B(new_n20986), .C(new_n20991), .D(new_n20992), .Y(new_n20993));
  NAND2xp33_ASAP7_75t_L     g20737(.A(new_n20981), .B(new_n20993), .Y(new_n20994));
  A2O1A1Ixp33_ASAP7_75t_L   g20738(.A1(new_n20988), .A2(new_n20816), .B(new_n20806), .C(new_n20987), .Y(new_n20995));
  INVx1_ASAP7_75t_L         g20739(.A(new_n20995), .Y(new_n20996));
  A2O1A1Ixp33_ASAP7_75t_L   g20740(.A1(\a[35] ), .A2(new_n20985), .B(new_n20986), .C(new_n20996), .Y(new_n20997));
  INVx1_ASAP7_75t_L         g20741(.A(new_n20997), .Y(new_n20998));
  A2O1A1Ixp33_ASAP7_75t_L   g20742(.A1(new_n20995), .A2(new_n20991), .B(new_n20998), .C(new_n20980), .Y(new_n20999));
  NAND2xp33_ASAP7_75t_L     g20743(.A(new_n20999), .B(new_n20994), .Y(new_n21000));
  O2A1O1Ixp33_ASAP7_75t_L   g20744(.A1(new_n20655), .A2(new_n20838), .B(new_n20839), .C(new_n21000), .Y(new_n21001));
  A2O1A1Ixp33_ASAP7_75t_L   g20745(.A1(new_n20655), .A2(new_n20820), .B(new_n20818), .C(new_n20662), .Y(new_n21002));
  AOI21xp33_ASAP7_75t_L     g20746(.A1(new_n20994), .A2(new_n20999), .B(new_n21002), .Y(new_n21003));
  NOR2xp33_ASAP7_75t_L      g20747(.A(new_n21003), .B(new_n21001), .Y(new_n21004));
  XNOR2x2_ASAP7_75t_L       g20748(.A(new_n21004), .B(new_n20836), .Y(\f[96] ));
  INVx1_ASAP7_75t_L         g20749(.A(new_n21001), .Y(new_n21006));
  AOI22xp33_ASAP7_75t_L     g20750(.A1(new_n4155), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4402), .Y(new_n21007));
  INVx1_ASAP7_75t_L         g20751(.A(new_n21007), .Y(new_n21008));
  A2O1A1Ixp33_ASAP7_75t_L   g20752(.A1(new_n4144), .A2(new_n4146), .B(new_n3926), .C(new_n21007), .Y(new_n21009));
  O2A1O1Ixp33_ASAP7_75t_L   g20753(.A1(new_n21008), .A2(new_n17329), .B(new_n21009), .C(new_n4145), .Y(new_n21010));
  O2A1O1Ixp33_ASAP7_75t_L   g20754(.A1(new_n4150), .A2(new_n12993), .B(new_n21007), .C(\a[35] ), .Y(new_n21011));
  NOR2xp33_ASAP7_75t_L      g20755(.A(new_n21011), .B(new_n21010), .Y(new_n21012));
  A2O1A1O1Ixp25_ASAP7_75t_L g20756(.A1(new_n20965), .A2(new_n20974), .B(new_n20976), .C(new_n20971), .D(new_n21012), .Y(new_n21013));
  A2O1A1Ixp33_ASAP7_75t_L   g20757(.A1(new_n20974), .A2(new_n20965), .B(new_n20976), .C(new_n20971), .Y(new_n21014));
  INVx1_ASAP7_75t_L         g20758(.A(new_n21012), .Y(new_n21015));
  NOR2xp33_ASAP7_75t_L      g20759(.A(new_n21015), .B(new_n21014), .Y(new_n21016));
  NOR2xp33_ASAP7_75t_L      g20760(.A(new_n21013), .B(new_n21016), .Y(new_n21017));
  A2O1A1O1Ixp25_ASAP7_75t_L g20761(.A1(new_n20503), .A2(new_n20513), .B(new_n20695), .C(new_n20698), .D(new_n20848), .Y(new_n21018));
  A2O1A1Ixp33_ASAP7_75t_L   g20762(.A1(new_n20849), .A2(new_n20848), .B(new_n21018), .C(new_n20857), .Y(new_n21019));
  NOR2xp33_ASAP7_75t_L      g20763(.A(new_n4101), .B(new_n13030), .Y(new_n21020));
  INVx1_ASAP7_75t_L         g20764(.A(new_n20842), .Y(new_n21021));
  A2O1A1O1Ixp25_ASAP7_75t_L g20765(.A1(new_n13028), .A2(\b[32] ), .B(new_n20693), .C(new_n20844), .D(new_n21021), .Y(new_n21022));
  A2O1A1Ixp33_ASAP7_75t_L   g20766(.A1(new_n13028), .A2(\b[34] ), .B(new_n21020), .C(new_n21022), .Y(new_n21023));
  O2A1O1Ixp33_ASAP7_75t_L   g20767(.A1(new_n12669), .A2(new_n12671), .B(\b[34] ), .C(new_n21020), .Y(new_n21024));
  INVx1_ASAP7_75t_L         g20768(.A(new_n21024), .Y(new_n21025));
  O2A1O1Ixp33_ASAP7_75t_L   g20769(.A1(new_n20697), .A2(new_n20845), .B(new_n20842), .C(new_n21025), .Y(new_n21026));
  INVx1_ASAP7_75t_L         g20770(.A(new_n21026), .Y(new_n21027));
  NAND2xp33_ASAP7_75t_L     g20771(.A(new_n21023), .B(new_n21027), .Y(new_n21028));
  NOR2xp33_ASAP7_75t_L      g20772(.A(new_n4613), .B(new_n12318), .Y(new_n21029));
  AOI221xp5_ASAP7_75t_L     g20773(.A1(new_n11995), .A2(\b[37] ), .B1(new_n13314), .B2(\b[35] ), .C(new_n21029), .Y(new_n21030));
  O2A1O1Ixp33_ASAP7_75t_L   g20774(.A1(new_n11998), .A2(new_n5083), .B(new_n21030), .C(new_n11987), .Y(new_n21031));
  INVx1_ASAP7_75t_L         g20775(.A(new_n21031), .Y(new_n21032));
  O2A1O1Ixp33_ASAP7_75t_L   g20776(.A1(new_n11998), .A2(new_n5083), .B(new_n21030), .C(\a[62] ), .Y(new_n21033));
  AOI21xp33_ASAP7_75t_L     g20777(.A1(new_n21032), .A2(\a[62] ), .B(new_n21033), .Y(new_n21034));
  NAND2xp33_ASAP7_75t_L     g20778(.A(new_n21028), .B(new_n21034), .Y(new_n21035));
  INVx1_ASAP7_75t_L         g20779(.A(new_n21033), .Y(new_n21036));
  O2A1O1Ixp33_ASAP7_75t_L   g20780(.A1(new_n21031), .A2(new_n11987), .B(new_n21036), .C(new_n21028), .Y(new_n21037));
  INVx1_ASAP7_75t_L         g20781(.A(new_n21037), .Y(new_n21038));
  NAND2xp33_ASAP7_75t_L     g20782(.A(new_n21038), .B(new_n21035), .Y(new_n21039));
  A2O1A1O1Ixp25_ASAP7_75t_L g20783(.A1(new_n20856), .A2(new_n20855), .B(new_n20851), .C(new_n20849), .D(new_n21039), .Y(new_n21040));
  NOR2xp33_ASAP7_75t_L      g20784(.A(new_n5311), .B(new_n11354), .Y(new_n21041));
  AOI221xp5_ASAP7_75t_L     g20785(.A1(\b[40] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[39] ), .C(new_n21041), .Y(new_n21042));
  O2A1O1Ixp33_ASAP7_75t_L   g20786(.A1(new_n11053), .A2(new_n5862), .B(new_n21042), .C(new_n11048), .Y(new_n21043));
  INVx1_ASAP7_75t_L         g20787(.A(new_n21043), .Y(new_n21044));
  O2A1O1Ixp33_ASAP7_75t_L   g20788(.A1(new_n11053), .A2(new_n5862), .B(new_n21042), .C(\a[59] ), .Y(new_n21045));
  AOI21xp33_ASAP7_75t_L     g20789(.A1(new_n21044), .A2(\a[59] ), .B(new_n21045), .Y(new_n21046));
  A2O1A1O1Ixp25_ASAP7_75t_L g20790(.A1(new_n13028), .A2(\b[31] ), .B(new_n20497), .C(new_n20697), .D(new_n20699), .Y(new_n21047));
  O2A1O1Ixp33_ASAP7_75t_L   g20791(.A1(new_n20845), .A2(new_n20846), .B(new_n20847), .C(new_n21047), .Y(new_n21048));
  INVx1_ASAP7_75t_L         g20792(.A(new_n20851), .Y(new_n21049));
  A2O1A1Ixp33_ASAP7_75t_L   g20793(.A1(new_n21049), .A2(new_n20857), .B(new_n21048), .C(new_n21039), .Y(new_n21050));
  O2A1O1Ixp33_ASAP7_75t_L   g20794(.A1(new_n21039), .A2(new_n21040), .B(new_n21050), .C(new_n21046), .Y(new_n21051));
  INVx1_ASAP7_75t_L         g20795(.A(new_n21040), .Y(new_n21052));
  NAND3xp33_ASAP7_75t_L     g20796(.A(new_n21052), .B(new_n21038), .C(new_n21035), .Y(new_n21053));
  AND2x2_ASAP7_75t_L        g20797(.A(new_n21046), .B(new_n21053), .Y(new_n21054));
  A2O1A1O1Ixp25_ASAP7_75t_L g20798(.A1(new_n21019), .A2(new_n20849), .B(new_n21040), .C(new_n21054), .D(new_n21051), .Y(new_n21055));
  INVx1_ASAP7_75t_L         g20799(.A(new_n21055), .Y(new_n21056));
  O2A1O1Ixp33_ASAP7_75t_L   g20800(.A1(new_n20858), .A2(new_n20866), .B(new_n20870), .C(new_n21056), .Y(new_n21057));
  INVx1_ASAP7_75t_L         g20801(.A(new_n21057), .Y(new_n21058));
  A2O1A1O1Ixp25_ASAP7_75t_L g20802(.A1(new_n20863), .A2(\a[59] ), .B(new_n20864), .C(new_n20859), .D(new_n20869), .Y(new_n21059));
  A2O1A1Ixp33_ASAP7_75t_L   g20803(.A1(new_n21054), .A2(new_n21050), .B(new_n21051), .C(new_n21059), .Y(new_n21060));
  AND2x2_ASAP7_75t_L        g20804(.A(new_n21060), .B(new_n21058), .Y(new_n21061));
  INVx1_ASAP7_75t_L         g20805(.A(new_n21061), .Y(new_n21062));
  NOR2xp33_ASAP7_75t_L      g20806(.A(new_n6378), .B(new_n10388), .Y(new_n21063));
  AOI221xp5_ASAP7_75t_L     g20807(.A1(new_n10086), .A2(\b[43] ), .B1(new_n11361), .B2(\b[41] ), .C(new_n21063), .Y(new_n21064));
  O2A1O1Ixp33_ASAP7_75t_L   g20808(.A1(new_n10088), .A2(new_n6679), .B(new_n21064), .C(new_n10083), .Y(new_n21065));
  O2A1O1Ixp33_ASAP7_75t_L   g20809(.A1(new_n10088), .A2(new_n6679), .B(new_n21064), .C(\a[56] ), .Y(new_n21066));
  INVx1_ASAP7_75t_L         g20810(.A(new_n21066), .Y(new_n21067));
  O2A1O1Ixp33_ASAP7_75t_L   g20811(.A1(new_n21065), .A2(new_n10083), .B(new_n21067), .C(new_n21062), .Y(new_n21068));
  INVx1_ASAP7_75t_L         g20812(.A(new_n21068), .Y(new_n21069));
  O2A1O1Ixp33_ASAP7_75t_L   g20813(.A1(new_n21065), .A2(new_n10083), .B(new_n21067), .C(new_n21061), .Y(new_n21070));
  AOI21xp33_ASAP7_75t_L     g20814(.A1(new_n21069), .A2(new_n21061), .B(new_n21070), .Y(new_n21071));
  O2A1O1Ixp33_ASAP7_75t_L   g20815(.A1(new_n20881), .A2(new_n20872), .B(new_n20883), .C(new_n20879), .Y(new_n21072));
  NAND2xp33_ASAP7_75t_L     g20816(.A(new_n21072), .B(new_n21071), .Y(new_n21073));
  O2A1O1Ixp33_ASAP7_75t_L   g20817(.A1(new_n20882), .A2(new_n20884), .B(new_n20880), .C(new_n21071), .Y(new_n21074));
  INVx1_ASAP7_75t_L         g20818(.A(new_n21074), .Y(new_n21075));
  AND2x2_ASAP7_75t_L        g20819(.A(new_n21073), .B(new_n21075), .Y(new_n21076));
  INVx1_ASAP7_75t_L         g20820(.A(new_n21076), .Y(new_n21077));
  NOR2xp33_ASAP7_75t_L      g20821(.A(new_n7249), .B(new_n10400), .Y(new_n21078));
  AOI221xp5_ASAP7_75t_L     g20822(.A1(new_n9102), .A2(\b[46] ), .B1(new_n10398), .B2(\b[44] ), .C(new_n21078), .Y(new_n21079));
  O2A1O1Ixp33_ASAP7_75t_L   g20823(.A1(new_n9104), .A2(new_n7279), .B(new_n21079), .C(new_n9099), .Y(new_n21080));
  O2A1O1Ixp33_ASAP7_75t_L   g20824(.A1(new_n9104), .A2(new_n7279), .B(new_n21079), .C(\a[53] ), .Y(new_n21081));
  INVx1_ASAP7_75t_L         g20825(.A(new_n21081), .Y(new_n21082));
  O2A1O1Ixp33_ASAP7_75t_L   g20826(.A1(new_n21080), .A2(new_n9099), .B(new_n21082), .C(new_n21077), .Y(new_n21083));
  INVx1_ASAP7_75t_L         g20827(.A(new_n21083), .Y(new_n21084));
  O2A1O1Ixp33_ASAP7_75t_L   g20828(.A1(new_n21080), .A2(new_n9099), .B(new_n21082), .C(new_n21076), .Y(new_n21085));
  AOI21xp33_ASAP7_75t_L     g20829(.A1(new_n21084), .A2(new_n21076), .B(new_n21085), .Y(new_n21086));
  A2O1A1Ixp33_ASAP7_75t_L   g20830(.A1(new_n20734), .A2(new_n20739), .B(new_n20898), .C(new_n20896), .Y(new_n21087));
  INVx1_ASAP7_75t_L         g20831(.A(new_n21087), .Y(new_n21088));
  NAND2xp33_ASAP7_75t_L     g20832(.A(new_n21088), .B(new_n21086), .Y(new_n21089));
  O2A1O1Ixp33_ASAP7_75t_L   g20833(.A1(new_n20898), .A2(new_n20899), .B(new_n20896), .C(new_n21086), .Y(new_n21090));
  INVx1_ASAP7_75t_L         g20834(.A(new_n21090), .Y(new_n21091));
  AND2x2_ASAP7_75t_L        g20835(.A(new_n21089), .B(new_n21091), .Y(new_n21092));
  NOR2xp33_ASAP7_75t_L      g20836(.A(new_n7860), .B(new_n10065), .Y(new_n21093));
  AOI221xp5_ASAP7_75t_L     g20837(.A1(new_n8175), .A2(\b[49] ), .B1(new_n8484), .B2(\b[47] ), .C(new_n21093), .Y(new_n21094));
  O2A1O1Ixp33_ASAP7_75t_L   g20838(.A1(new_n8176), .A2(new_n14802), .B(new_n21094), .C(new_n8172), .Y(new_n21095));
  INVx1_ASAP7_75t_L         g20839(.A(new_n21095), .Y(new_n21096));
  O2A1O1Ixp33_ASAP7_75t_L   g20840(.A1(new_n8176), .A2(new_n14802), .B(new_n21094), .C(\a[50] ), .Y(new_n21097));
  A2O1A1Ixp33_ASAP7_75t_L   g20841(.A1(\a[50] ), .A2(new_n21096), .B(new_n21097), .C(new_n21092), .Y(new_n21098));
  INVx1_ASAP7_75t_L         g20842(.A(new_n21097), .Y(new_n21099));
  O2A1O1Ixp33_ASAP7_75t_L   g20843(.A1(new_n21095), .A2(new_n8172), .B(new_n21099), .C(new_n21092), .Y(new_n21100));
  A2O1A1Ixp33_ASAP7_75t_L   g20844(.A1(new_n20745), .A2(new_n20755), .B(new_n20913), .C(new_n20911), .Y(new_n21101));
  AOI211xp5_ASAP7_75t_L     g20845(.A1(new_n21092), .A2(new_n21098), .B(new_n21100), .C(new_n21101), .Y(new_n21102));
  AOI21xp33_ASAP7_75t_L     g20846(.A1(new_n21098), .A2(new_n21092), .B(new_n21100), .Y(new_n21103));
  O2A1O1Ixp33_ASAP7_75t_L   g20847(.A1(new_n20913), .A2(new_n20914), .B(new_n20911), .C(new_n21103), .Y(new_n21104));
  NOR2xp33_ASAP7_75t_L      g20848(.A(new_n21104), .B(new_n21102), .Y(new_n21105));
  NOR2xp33_ASAP7_75t_L      g20849(.A(new_n8779), .B(new_n7312), .Y(new_n21106));
  AOI221xp5_ASAP7_75t_L     g20850(.A1(\b[50] ), .A2(new_n7609), .B1(\b[52] ), .B2(new_n7334), .C(new_n21106), .Y(new_n21107));
  O2A1O1Ixp33_ASAP7_75t_L   g20851(.A1(new_n7321), .A2(new_n17363), .B(new_n21107), .C(new_n7316), .Y(new_n21108));
  INVx1_ASAP7_75t_L         g20852(.A(new_n21108), .Y(new_n21109));
  O2A1O1Ixp33_ASAP7_75t_L   g20853(.A1(new_n7321), .A2(new_n17363), .B(new_n21107), .C(\a[47] ), .Y(new_n21110));
  A2O1A1Ixp33_ASAP7_75t_L   g20854(.A1(\a[47] ), .A2(new_n21109), .B(new_n21110), .C(new_n21105), .Y(new_n21111));
  INVx1_ASAP7_75t_L         g20855(.A(new_n21110), .Y(new_n21112));
  O2A1O1Ixp33_ASAP7_75t_L   g20856(.A1(new_n21108), .A2(new_n7316), .B(new_n21112), .C(new_n21105), .Y(new_n21113));
  AOI21xp33_ASAP7_75t_L     g20857(.A1(new_n21111), .A2(new_n21105), .B(new_n21113), .Y(new_n21114));
  A2O1A1Ixp33_ASAP7_75t_L   g20858(.A1(new_n20927), .A2(new_n20917), .B(new_n20929), .C(new_n21114), .Y(new_n21115));
  A2O1A1Ixp33_ASAP7_75t_L   g20859(.A1(new_n21105), .A2(new_n21111), .B(new_n21113), .C(new_n20932), .Y(new_n21116));
  NAND2xp33_ASAP7_75t_L     g20860(.A(new_n21115), .B(new_n21116), .Y(new_n21117));
  NOR2xp33_ASAP7_75t_L      g20861(.A(new_n9683), .B(new_n6741), .Y(new_n21118));
  AOI221xp5_ASAP7_75t_L     g20862(.A1(\b[55] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[54] ), .C(new_n21118), .Y(new_n21119));
  O2A1O1Ixp33_ASAP7_75t_L   g20863(.A1(new_n6443), .A2(new_n15849), .B(new_n21119), .C(new_n6439), .Y(new_n21120));
  NOR2xp33_ASAP7_75t_L      g20864(.A(new_n6439), .B(new_n21120), .Y(new_n21121));
  O2A1O1Ixp33_ASAP7_75t_L   g20865(.A1(new_n6443), .A2(new_n15849), .B(new_n21119), .C(\a[44] ), .Y(new_n21122));
  NOR2xp33_ASAP7_75t_L      g20866(.A(new_n21122), .B(new_n21121), .Y(new_n21123));
  XNOR2x2_ASAP7_75t_L       g20867(.A(new_n21123), .B(new_n21117), .Y(new_n21124));
  INVx1_ASAP7_75t_L         g20868(.A(new_n21124), .Y(new_n21125));
  A2O1A1O1Ixp25_ASAP7_75t_L g20869(.A1(new_n20782), .A2(new_n20772), .B(new_n20945), .C(new_n20943), .D(new_n21125), .Y(new_n21126));
  INVx1_ASAP7_75t_L         g20870(.A(new_n21126), .Y(new_n21127));
  A2O1A1Ixp33_ASAP7_75t_L   g20871(.A1(new_n20772), .A2(new_n20782), .B(new_n20945), .C(new_n20943), .Y(new_n21128));
  INVx1_ASAP7_75t_L         g20872(.A(new_n21128), .Y(new_n21129));
  NAND2xp33_ASAP7_75t_L     g20873(.A(new_n21125), .B(new_n21129), .Y(new_n21130));
  AND2x2_ASAP7_75t_L        g20874(.A(new_n21127), .B(new_n21130), .Y(new_n21131));
  INVx1_ASAP7_75t_L         g20875(.A(new_n21131), .Y(new_n21132));
  NOR2xp33_ASAP7_75t_L      g20876(.A(new_n11303), .B(new_n5641), .Y(new_n21133));
  AOI221xp5_ASAP7_75t_L     g20877(.A1(\b[56] ), .A2(new_n5920), .B1(\b[57] ), .B2(new_n5623), .C(new_n21133), .Y(new_n21134));
  O2A1O1Ixp33_ASAP7_75t_L   g20878(.A1(new_n5630), .A2(new_n20073), .B(new_n21134), .C(new_n5626), .Y(new_n21135));
  O2A1O1Ixp33_ASAP7_75t_L   g20879(.A1(new_n5630), .A2(new_n20073), .B(new_n21134), .C(\a[41] ), .Y(new_n21136));
  INVx1_ASAP7_75t_L         g20880(.A(new_n21136), .Y(new_n21137));
  O2A1O1Ixp33_ASAP7_75t_L   g20881(.A1(new_n21135), .A2(new_n5626), .B(new_n21137), .C(new_n21132), .Y(new_n21138));
  INVx1_ASAP7_75t_L         g20882(.A(new_n21138), .Y(new_n21139));
  O2A1O1Ixp33_ASAP7_75t_L   g20883(.A1(new_n21135), .A2(new_n5626), .B(new_n21137), .C(new_n21131), .Y(new_n21140));
  AOI21xp33_ASAP7_75t_L     g20884(.A1(new_n21139), .A2(new_n21131), .B(new_n21140), .Y(new_n21141));
  O2A1O1Ixp33_ASAP7_75t_L   g20885(.A1(new_n20956), .A2(new_n20957), .B(new_n20963), .C(new_n20955), .Y(new_n21142));
  NAND2xp33_ASAP7_75t_L     g20886(.A(new_n21142), .B(new_n21141), .Y(new_n21143));
  INVx1_ASAP7_75t_L         g20887(.A(new_n21142), .Y(new_n21144));
  A2O1A1Ixp33_ASAP7_75t_L   g20888(.A1(new_n21139), .A2(new_n21131), .B(new_n21140), .C(new_n21144), .Y(new_n21145));
  AND2x2_ASAP7_75t_L        g20889(.A(new_n21145), .B(new_n21143), .Y(new_n21146));
  NOR2xp33_ASAP7_75t_L      g20890(.A(new_n12258), .B(new_n4908), .Y(new_n21147));
  AOI221xp5_ASAP7_75t_L     g20891(.A1(\b[59] ), .A2(new_n5139), .B1(\b[60] ), .B2(new_n4916), .C(new_n21147), .Y(new_n21148));
  O2A1O1Ixp33_ASAP7_75t_L   g20892(.A1(new_n4911), .A2(new_n14764), .B(new_n21148), .C(new_n4906), .Y(new_n21149));
  INVx1_ASAP7_75t_L         g20893(.A(new_n21149), .Y(new_n21150));
  O2A1O1Ixp33_ASAP7_75t_L   g20894(.A1(new_n4911), .A2(new_n14764), .B(new_n21148), .C(\a[38] ), .Y(new_n21151));
  A2O1A1Ixp33_ASAP7_75t_L   g20895(.A1(\a[38] ), .A2(new_n21150), .B(new_n21151), .C(new_n21146), .Y(new_n21152));
  NOR2xp33_ASAP7_75t_L      g20896(.A(new_n4906), .B(new_n21149), .Y(new_n21153));
  OR3x1_ASAP7_75t_L         g20897(.A(new_n21146), .B(new_n21153), .C(new_n21151), .Y(new_n21154));
  NAND3xp33_ASAP7_75t_L     g20898(.A(new_n21017), .B(new_n21152), .C(new_n21154), .Y(new_n21155));
  NAND3xp33_ASAP7_75t_L     g20899(.A(new_n21155), .B(new_n21154), .C(new_n21152), .Y(new_n21156));
  INVx1_ASAP7_75t_L         g20900(.A(new_n21156), .Y(new_n21157));
  A2O1A1Ixp33_ASAP7_75t_L   g20901(.A1(new_n20997), .A2(new_n20996), .B(new_n20981), .C(new_n20991), .Y(new_n21158));
  A2O1A1Ixp33_ASAP7_75t_L   g20902(.A1(new_n21155), .A2(new_n21017), .B(new_n21157), .C(new_n21158), .Y(new_n21159));
  AO21x2_ASAP7_75t_L        g20903(.A1(new_n21017), .A2(new_n21155), .B(new_n21157), .Y(new_n21160));
  O2A1O1Ixp33_ASAP7_75t_L   g20904(.A1(new_n20981), .A2(new_n20993), .B(new_n20991), .C(new_n21160), .Y(new_n21161));
  A2O1A1O1Ixp25_ASAP7_75t_L g20905(.A1(new_n21155), .A2(new_n21017), .B(new_n21157), .C(new_n21159), .D(new_n21161), .Y(new_n21162));
  O2A1O1Ixp33_ASAP7_75t_L   g20906(.A1(new_n21003), .A2(new_n20836), .B(new_n21006), .C(new_n21162), .Y(new_n21163));
  A2O1A1Ixp33_ASAP7_75t_L   g20907(.A1(new_n20833), .A2(new_n20832), .B(new_n20828), .C(new_n21004), .Y(new_n21164));
  AND3x1_ASAP7_75t_L        g20908(.A(new_n21164), .B(new_n21162), .C(new_n21006), .Y(new_n21165));
  NOR2xp33_ASAP7_75t_L      g20909(.A(new_n21163), .B(new_n21165), .Y(\f[97] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20910(.A1(new_n21164), .A2(new_n21006), .B(new_n21162), .C(new_n21159), .Y(new_n21167));
  O2A1O1Ixp33_ASAP7_75t_L   g20911(.A1(new_n20802), .A2(new_n20792), .B(new_n20975), .C(new_n20972), .Y(new_n21168));
  INVx1_ASAP7_75t_L         g20912(.A(new_n21145), .Y(new_n21169));
  O2A1O1Ixp33_ASAP7_75t_L   g20913(.A1(new_n21153), .A2(new_n21151), .B(new_n21143), .C(new_n21169), .Y(new_n21170));
  INVx1_ASAP7_75t_L         g20914(.A(new_n21170), .Y(new_n21171));
  NOR2xp33_ASAP7_75t_L      g20915(.A(new_n12956), .B(new_n4397), .Y(new_n21172));
  A2O1A1Ixp33_ASAP7_75t_L   g20916(.A1(new_n12986), .A2(new_n4151), .B(new_n21172), .C(\a[35] ), .Y(new_n21173));
  INVx1_ASAP7_75t_L         g20917(.A(new_n21173), .Y(new_n21174));
  A2O1A1Ixp33_ASAP7_75t_L   g20918(.A1(new_n12986), .A2(new_n4151), .B(new_n21172), .C(new_n4145), .Y(new_n21175));
  O2A1O1Ixp33_ASAP7_75t_L   g20919(.A1(new_n21174), .A2(new_n4145), .B(new_n21175), .C(new_n21170), .Y(new_n21176));
  INVx1_ASAP7_75t_L         g20920(.A(new_n21176), .Y(new_n21177));
  O2A1O1Ixp33_ASAP7_75t_L   g20921(.A1(new_n21174), .A2(new_n4145), .B(new_n21175), .C(new_n21171), .Y(new_n21178));
  INVx1_ASAP7_75t_L         g20922(.A(new_n21123), .Y(new_n21179));
  O2A1O1Ixp33_ASAP7_75t_L   g20923(.A1(new_n20928), .A2(new_n20840), .B(new_n20923), .C(new_n21114), .Y(new_n21180));
  NOR2xp33_ASAP7_75t_L      g20924(.A(new_n10309), .B(new_n7304), .Y(new_n21181));
  AOI221xp5_ASAP7_75t_L     g20925(.A1(\b[54] ), .A2(new_n6742), .B1(\b[56] ), .B2(new_n6442), .C(new_n21181), .Y(new_n21182));
  INVx1_ASAP7_75t_L         g20926(.A(new_n21182), .Y(new_n21183));
  A2O1A1Ixp33_ASAP7_75t_L   g20927(.A1(new_n11579), .A2(new_n6450), .B(new_n21183), .C(\a[44] ), .Y(new_n21184));
  O2A1O1Ixp33_ASAP7_75t_L   g20928(.A1(new_n6443), .A2(new_n10339), .B(new_n21182), .C(\a[44] ), .Y(new_n21185));
  AO21x2_ASAP7_75t_L        g20929(.A1(\a[44] ), .A2(new_n21184), .B(new_n21185), .Y(new_n21186));
  A2O1A1O1Ixp25_ASAP7_75t_L g20930(.A1(new_n21096), .A2(\a[50] ), .B(new_n21097), .C(new_n21089), .D(new_n21090), .Y(new_n21187));
  INVx1_ASAP7_75t_L         g20931(.A(new_n21187), .Y(new_n21188));
  NOR2xp33_ASAP7_75t_L      g20932(.A(new_n6671), .B(new_n10388), .Y(new_n21189));
  AOI221xp5_ASAP7_75t_L     g20933(.A1(new_n10086), .A2(\b[44] ), .B1(new_n11361), .B2(\b[42] ), .C(new_n21189), .Y(new_n21190));
  O2A1O1Ixp33_ASAP7_75t_L   g20934(.A1(new_n10088), .A2(new_n6951), .B(new_n21190), .C(new_n10083), .Y(new_n21191));
  INVx1_ASAP7_75t_L         g20935(.A(new_n21191), .Y(new_n21192));
  O2A1O1Ixp33_ASAP7_75t_L   g20936(.A1(new_n10088), .A2(new_n6951), .B(new_n21190), .C(\a[56] ), .Y(new_n21193));
  NOR2xp33_ASAP7_75t_L      g20937(.A(new_n4344), .B(new_n13030), .Y(new_n21194));
  O2A1O1Ixp33_ASAP7_75t_L   g20938(.A1(new_n12669), .A2(new_n12671), .B(\b[35] ), .C(new_n21194), .Y(new_n21195));
  INVx1_ASAP7_75t_L         g20939(.A(new_n21194), .Y(new_n21196));
  O2A1O1Ixp33_ASAP7_75t_L   g20940(.A1(new_n12672), .A2(new_n4581), .B(new_n21196), .C(new_n21025), .Y(new_n21197));
  O2A1O1Ixp33_ASAP7_75t_L   g20941(.A1(new_n21028), .A2(new_n21034), .B(new_n21027), .C(new_n21197), .Y(new_n21198));
  INVx1_ASAP7_75t_L         g20942(.A(new_n21198), .Y(new_n21199));
  A2O1A1O1Ixp25_ASAP7_75t_L g20943(.A1(new_n13028), .A2(\b[34] ), .B(new_n21020), .C(new_n21195), .D(new_n21199), .Y(new_n21200));
  O2A1O1Ixp33_ASAP7_75t_L   g20944(.A1(new_n21025), .A2(new_n21022), .B(new_n21038), .C(new_n21200), .Y(new_n21201));
  A2O1A1Ixp33_ASAP7_75t_L   g20945(.A1(new_n13028), .A2(\b[34] ), .B(new_n21020), .C(new_n21195), .Y(new_n21202));
  INVx1_ASAP7_75t_L         g20946(.A(new_n21202), .Y(new_n21203));
  INVx1_ASAP7_75t_L         g20947(.A(new_n21197), .Y(new_n21204));
  O2A1O1Ixp33_ASAP7_75t_L   g20948(.A1(new_n21026), .A2(new_n21037), .B(new_n21204), .C(new_n21203), .Y(new_n21205));
  INVx1_ASAP7_75t_L         g20949(.A(new_n21205), .Y(new_n21206));
  A2O1A1O1Ixp25_ASAP7_75t_L g20950(.A1(new_n13028), .A2(\b[35] ), .B(new_n21194), .C(new_n21024), .D(new_n21206), .Y(new_n21207));
  A2O1A1O1Ixp25_ASAP7_75t_L g20951(.A1(\a[62] ), .A2(new_n21032), .B(new_n21033), .C(new_n21023), .D(new_n21026), .Y(new_n21208));
  INVx1_ASAP7_75t_L         g20952(.A(new_n21207), .Y(new_n21209));
  OAI22xp33_ASAP7_75t_L     g20953(.A1(new_n12320), .A2(new_n4613), .B1(new_n5074), .B2(new_n12318), .Y(new_n21210));
  AOI221xp5_ASAP7_75t_L     g20954(.A1(new_n11995), .A2(\b[38] ), .B1(new_n11997), .B2(new_n6083), .C(new_n21210), .Y(new_n21211));
  XNOR2x2_ASAP7_75t_L       g20955(.A(new_n11987), .B(new_n21211), .Y(new_n21212));
  O2A1O1Ixp33_ASAP7_75t_L   g20956(.A1(new_n21208), .A2(new_n21200), .B(new_n21209), .C(new_n21212), .Y(new_n21213));
  INVx1_ASAP7_75t_L         g20957(.A(new_n21213), .Y(new_n21214));
  A2O1A1Ixp33_ASAP7_75t_L   g20958(.A1(new_n21202), .A2(new_n21198), .B(new_n21208), .C(new_n21209), .Y(new_n21215));
  NOR2xp33_ASAP7_75t_L      g20959(.A(new_n21212), .B(new_n21215), .Y(new_n21216));
  O2A1O1Ixp33_ASAP7_75t_L   g20960(.A1(new_n21201), .A2(new_n21207), .B(new_n21214), .C(new_n21216), .Y(new_n21217));
  NOR2xp33_ASAP7_75t_L      g20961(.A(new_n5570), .B(new_n11354), .Y(new_n21218));
  AOI221xp5_ASAP7_75t_L     g20962(.A1(\b[41] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[40] ), .C(new_n21218), .Y(new_n21219));
  O2A1O1Ixp33_ASAP7_75t_L   g20963(.A1(new_n11053), .A2(new_n6117), .B(new_n21219), .C(new_n11048), .Y(new_n21220));
  NOR2xp33_ASAP7_75t_L      g20964(.A(new_n11048), .B(new_n21220), .Y(new_n21221));
  O2A1O1Ixp33_ASAP7_75t_L   g20965(.A1(new_n11053), .A2(new_n6117), .B(new_n21219), .C(\a[59] ), .Y(new_n21222));
  NOR2xp33_ASAP7_75t_L      g20966(.A(new_n21222), .B(new_n21221), .Y(new_n21223));
  XNOR2x2_ASAP7_75t_L       g20967(.A(new_n21223), .B(new_n21217), .Y(new_n21224));
  A2O1A1O1Ixp25_ASAP7_75t_L g20968(.A1(new_n21050), .A2(new_n21039), .B(new_n21046), .C(new_n21052), .D(new_n21224), .Y(new_n21225));
  INVx1_ASAP7_75t_L         g20969(.A(new_n21225), .Y(new_n21226));
  A2O1A1Ixp33_ASAP7_75t_L   g20970(.A1(new_n21019), .A2(new_n20849), .B(new_n21040), .C(new_n21053), .Y(new_n21227));
  A2O1A1O1Ixp25_ASAP7_75t_L g20971(.A1(new_n21044), .A2(\a[59] ), .B(new_n21045), .C(new_n21227), .D(new_n21040), .Y(new_n21228));
  NAND2xp33_ASAP7_75t_L     g20972(.A(new_n21228), .B(new_n21224), .Y(new_n21229));
  AND2x2_ASAP7_75t_L        g20973(.A(new_n21229), .B(new_n21226), .Y(new_n21230));
  A2O1A1Ixp33_ASAP7_75t_L   g20974(.A1(new_n21192), .A2(\a[56] ), .B(new_n21193), .C(new_n21230), .Y(new_n21231));
  AOI21xp33_ASAP7_75t_L     g20975(.A1(new_n21192), .A2(\a[56] ), .B(new_n21193), .Y(new_n21232));
  INVx1_ASAP7_75t_L         g20976(.A(new_n21230), .Y(new_n21233));
  NAND2xp33_ASAP7_75t_L     g20977(.A(new_n21232), .B(new_n21233), .Y(new_n21234));
  AND2x2_ASAP7_75t_L        g20978(.A(new_n21231), .B(new_n21234), .Y(new_n21235));
  INVx1_ASAP7_75t_L         g20979(.A(new_n21235), .Y(new_n21236));
  O2A1O1Ixp33_ASAP7_75t_L   g20980(.A1(new_n21059), .A2(new_n21056), .B(new_n21069), .C(new_n21236), .Y(new_n21237));
  INVx1_ASAP7_75t_L         g20981(.A(new_n21237), .Y(new_n21238));
  A2O1A1Ixp33_ASAP7_75t_L   g20982(.A1(new_n20870), .A2(new_n20865), .B(new_n21056), .C(new_n21069), .Y(new_n21239));
  INVx1_ASAP7_75t_L         g20983(.A(new_n21239), .Y(new_n21240));
  NAND2xp33_ASAP7_75t_L     g20984(.A(new_n21240), .B(new_n21236), .Y(new_n21241));
  AND2x2_ASAP7_75t_L        g20985(.A(new_n21241), .B(new_n21238), .Y(new_n21242));
  INVx1_ASAP7_75t_L         g20986(.A(new_n21242), .Y(new_n21243));
  NOR2xp33_ASAP7_75t_L      g20987(.A(new_n7270), .B(new_n10400), .Y(new_n21244));
  AOI221xp5_ASAP7_75t_L     g20988(.A1(new_n9102), .A2(\b[47] ), .B1(new_n10398), .B2(\b[45] ), .C(new_n21244), .Y(new_n21245));
  O2A1O1Ixp33_ASAP7_75t_L   g20989(.A1(new_n9104), .A2(new_n7560), .B(new_n21245), .C(new_n9099), .Y(new_n21246));
  O2A1O1Ixp33_ASAP7_75t_L   g20990(.A1(new_n9104), .A2(new_n7560), .B(new_n21245), .C(\a[53] ), .Y(new_n21247));
  INVx1_ASAP7_75t_L         g20991(.A(new_n21247), .Y(new_n21248));
  O2A1O1Ixp33_ASAP7_75t_L   g20992(.A1(new_n21246), .A2(new_n9099), .B(new_n21248), .C(new_n21243), .Y(new_n21249));
  INVx1_ASAP7_75t_L         g20993(.A(new_n21249), .Y(new_n21250));
  O2A1O1Ixp33_ASAP7_75t_L   g20994(.A1(new_n21246), .A2(new_n9099), .B(new_n21248), .C(new_n21242), .Y(new_n21251));
  AOI21xp33_ASAP7_75t_L     g20995(.A1(new_n21250), .A2(new_n21242), .B(new_n21251), .Y(new_n21252));
  A2O1A1Ixp33_ASAP7_75t_L   g20996(.A1(new_n20887), .A2(new_n20880), .B(new_n21071), .C(new_n21084), .Y(new_n21253));
  INVx1_ASAP7_75t_L         g20997(.A(new_n21253), .Y(new_n21254));
  NAND2xp33_ASAP7_75t_L     g20998(.A(new_n21254), .B(new_n21252), .Y(new_n21255));
  O2A1O1Ixp33_ASAP7_75t_L   g20999(.A1(new_n21071), .A2(new_n21072), .B(new_n21084), .C(new_n21252), .Y(new_n21256));
  INVx1_ASAP7_75t_L         g21000(.A(new_n21256), .Y(new_n21257));
  AND2x2_ASAP7_75t_L        g21001(.A(new_n21255), .B(new_n21257), .Y(new_n21258));
  NOR2xp33_ASAP7_75t_L      g21002(.A(new_n8427), .B(new_n10065), .Y(new_n21259));
  AOI221xp5_ASAP7_75t_L     g21003(.A1(new_n8175), .A2(\b[50] ), .B1(new_n8484), .B2(\b[48] ), .C(new_n21259), .Y(new_n21260));
  O2A1O1Ixp33_ASAP7_75t_L   g21004(.A1(new_n8176), .A2(new_n8764), .B(new_n21260), .C(new_n8172), .Y(new_n21261));
  INVx1_ASAP7_75t_L         g21005(.A(new_n21261), .Y(new_n21262));
  O2A1O1Ixp33_ASAP7_75t_L   g21006(.A1(new_n8176), .A2(new_n8764), .B(new_n21260), .C(\a[50] ), .Y(new_n21263));
  AOI211xp5_ASAP7_75t_L     g21007(.A1(new_n21262), .A2(\a[50] ), .B(new_n21263), .C(new_n21258), .Y(new_n21264));
  A2O1A1Ixp33_ASAP7_75t_L   g21008(.A1(\a[50] ), .A2(new_n21262), .B(new_n21263), .C(new_n21258), .Y(new_n21265));
  INVx1_ASAP7_75t_L         g21009(.A(new_n21265), .Y(new_n21266));
  NOR2xp33_ASAP7_75t_L      g21010(.A(new_n21264), .B(new_n21266), .Y(new_n21267));
  NAND2xp33_ASAP7_75t_L     g21011(.A(new_n21188), .B(new_n21267), .Y(new_n21268));
  NOR2xp33_ASAP7_75t_L      g21012(.A(new_n9683), .B(new_n7318), .Y(new_n21269));
  AOI221xp5_ASAP7_75t_L     g21013(.A1(new_n7333), .A2(\b[52] ), .B1(new_n7609), .B2(\b[51] ), .C(new_n21269), .Y(new_n21270));
  O2A1O1Ixp33_ASAP7_75t_L   g21014(.A1(new_n7321), .A2(new_n9691), .B(new_n21270), .C(new_n7316), .Y(new_n21271));
  INVx1_ASAP7_75t_L         g21015(.A(new_n21271), .Y(new_n21272));
  O2A1O1Ixp33_ASAP7_75t_L   g21016(.A1(new_n7321), .A2(new_n9691), .B(new_n21270), .C(\a[47] ), .Y(new_n21273));
  O2A1O1Ixp33_ASAP7_75t_L   g21017(.A1(new_n21086), .A2(new_n21088), .B(new_n21098), .C(new_n21267), .Y(new_n21274));
  INVx1_ASAP7_75t_L         g21018(.A(new_n21274), .Y(new_n21275));
  NAND2xp33_ASAP7_75t_L     g21019(.A(new_n21187), .B(new_n21267), .Y(new_n21276));
  NAND2xp33_ASAP7_75t_L     g21020(.A(new_n21276), .B(new_n21275), .Y(new_n21277));
  A2O1A1Ixp33_ASAP7_75t_L   g21021(.A1(new_n21272), .A2(\a[47] ), .B(new_n21273), .C(new_n21277), .Y(new_n21278));
  AOI21xp33_ASAP7_75t_L     g21022(.A1(new_n21272), .A2(\a[47] ), .B(new_n21273), .Y(new_n21279));
  NAND2xp33_ASAP7_75t_L     g21023(.A(new_n21279), .B(new_n21276), .Y(new_n21280));
  A2O1A1Ixp33_ASAP7_75t_L   g21024(.A1(new_n21188), .A2(new_n21268), .B(new_n21280), .C(new_n21278), .Y(new_n21281));
  A2O1A1O1Ixp25_ASAP7_75t_L g21025(.A1(new_n20931), .A2(new_n20911), .B(new_n21103), .C(new_n21111), .D(new_n21281), .Y(new_n21282));
  A2O1A1Ixp33_ASAP7_75t_L   g21026(.A1(new_n20931), .A2(new_n20911), .B(new_n21103), .C(new_n21111), .Y(new_n21283));
  O2A1O1Ixp33_ASAP7_75t_L   g21027(.A1(new_n21280), .A2(new_n21274), .B(new_n21278), .C(new_n21283), .Y(new_n21284));
  NOR2xp33_ASAP7_75t_L      g21028(.A(new_n21284), .B(new_n21282), .Y(new_n21285));
  XOR2x2_ASAP7_75t_L        g21029(.A(new_n21186), .B(new_n21285), .Y(new_n21286));
  A2O1A1Ixp33_ASAP7_75t_L   g21030(.A1(new_n21179), .A2(new_n21117), .B(new_n21180), .C(new_n21286), .Y(new_n21287));
  O2A1O1Ixp33_ASAP7_75t_L   g21031(.A1(new_n21121), .A2(new_n21122), .B(new_n21117), .C(new_n21180), .Y(new_n21288));
  INVx1_ASAP7_75t_L         g21032(.A(new_n21286), .Y(new_n21289));
  NAND2xp33_ASAP7_75t_L     g21033(.A(new_n21288), .B(new_n21289), .Y(new_n21290));
  AND2x2_ASAP7_75t_L        g21034(.A(new_n21287), .B(new_n21290), .Y(new_n21291));
  INVx1_ASAP7_75t_L         g21035(.A(new_n21291), .Y(new_n21292));
  NOR2xp33_ASAP7_75t_L      g21036(.A(new_n11591), .B(new_n5641), .Y(new_n21293));
  AOI221xp5_ASAP7_75t_L     g21037(.A1(\b[57] ), .A2(new_n5920), .B1(\b[58] ), .B2(new_n5623), .C(new_n21293), .Y(new_n21294));
  O2A1O1Ixp33_ASAP7_75t_L   g21038(.A1(new_n5630), .A2(new_n11597), .B(new_n21294), .C(new_n5626), .Y(new_n21295));
  O2A1O1Ixp33_ASAP7_75t_L   g21039(.A1(new_n5630), .A2(new_n11597), .B(new_n21294), .C(\a[41] ), .Y(new_n21296));
  INVx1_ASAP7_75t_L         g21040(.A(new_n21296), .Y(new_n21297));
  O2A1O1Ixp33_ASAP7_75t_L   g21041(.A1(new_n21295), .A2(new_n5626), .B(new_n21297), .C(new_n21292), .Y(new_n21298));
  INVx1_ASAP7_75t_L         g21042(.A(new_n21298), .Y(new_n21299));
  O2A1O1Ixp33_ASAP7_75t_L   g21043(.A1(new_n21295), .A2(new_n5626), .B(new_n21297), .C(new_n21291), .Y(new_n21300));
  AOI21xp33_ASAP7_75t_L     g21044(.A1(new_n21299), .A2(new_n21291), .B(new_n21300), .Y(new_n21301));
  O2A1O1Ixp33_ASAP7_75t_L   g21045(.A1(new_n20942), .A2(new_n20946), .B(new_n21124), .C(new_n21138), .Y(new_n21302));
  NAND2xp33_ASAP7_75t_L     g21046(.A(new_n21301), .B(new_n21302), .Y(new_n21303));
  O2A1O1Ixp33_ASAP7_75t_L   g21047(.A1(new_n21129), .A2(new_n21125), .B(new_n21139), .C(new_n21301), .Y(new_n21304));
  INVx1_ASAP7_75t_L         g21048(.A(new_n21304), .Y(new_n21305));
  AND2x2_ASAP7_75t_L        g21049(.A(new_n21303), .B(new_n21305), .Y(new_n21306));
  INVx1_ASAP7_75t_L         g21050(.A(new_n21306), .Y(new_n21307));
  NOR2xp33_ASAP7_75t_L      g21051(.A(new_n12603), .B(new_n4908), .Y(new_n21308));
  AOI221xp5_ASAP7_75t_L     g21052(.A1(\b[60] ), .A2(new_n5139), .B1(\b[61] ), .B2(new_n4916), .C(new_n21308), .Y(new_n21309));
  O2A1O1Ixp33_ASAP7_75t_L   g21053(.A1(new_n4911), .A2(new_n12610), .B(new_n21309), .C(new_n4906), .Y(new_n21310));
  O2A1O1Ixp33_ASAP7_75t_L   g21054(.A1(new_n4911), .A2(new_n12610), .B(new_n21309), .C(\a[38] ), .Y(new_n21311));
  INVx1_ASAP7_75t_L         g21055(.A(new_n21311), .Y(new_n21312));
  O2A1O1Ixp33_ASAP7_75t_L   g21056(.A1(new_n21310), .A2(new_n4906), .B(new_n21312), .C(new_n21307), .Y(new_n21313));
  INVx1_ASAP7_75t_L         g21057(.A(new_n21313), .Y(new_n21314));
  O2A1O1Ixp33_ASAP7_75t_L   g21058(.A1(new_n21310), .A2(new_n4906), .B(new_n21312), .C(new_n21306), .Y(new_n21315));
  AOI21xp33_ASAP7_75t_L     g21059(.A1(new_n21314), .A2(new_n21306), .B(new_n21315), .Y(new_n21316));
  A2O1A1Ixp33_ASAP7_75t_L   g21060(.A1(new_n21177), .A2(new_n21171), .B(new_n21178), .C(new_n21316), .Y(new_n21317));
  INVx1_ASAP7_75t_L         g21061(.A(new_n21178), .Y(new_n21318));
  A2O1A1Ixp33_ASAP7_75t_L   g21062(.A1(new_n21152), .A2(new_n21145), .B(new_n21176), .C(new_n21318), .Y(new_n21319));
  INVx1_ASAP7_75t_L         g21063(.A(new_n21319), .Y(new_n21320));
  A2O1A1Ixp33_ASAP7_75t_L   g21064(.A1(new_n21306), .A2(new_n21314), .B(new_n21315), .C(new_n21320), .Y(new_n21321));
  AND2x2_ASAP7_75t_L        g21065(.A(new_n21317), .B(new_n21321), .Y(new_n21322));
  O2A1O1Ixp33_ASAP7_75t_L   g21066(.A1(new_n21168), .A2(new_n21012), .B(new_n21155), .C(new_n21322), .Y(new_n21323));
  A2O1A1Ixp33_ASAP7_75t_L   g21067(.A1(new_n20975), .A2(new_n20977), .B(new_n20972), .C(new_n21015), .Y(new_n21324));
  AND3x1_ASAP7_75t_L        g21068(.A(new_n21322), .B(new_n21155), .C(new_n21324), .Y(new_n21325));
  NOR2xp33_ASAP7_75t_L      g21069(.A(new_n21323), .B(new_n21325), .Y(new_n21326));
  XOR2x2_ASAP7_75t_L        g21070(.A(new_n21326), .B(new_n21167), .Y(\f[98] ));
  NOR2xp33_ASAP7_75t_L      g21071(.A(new_n10332), .B(new_n7304), .Y(new_n21328));
  AOI221xp5_ASAP7_75t_L     g21072(.A1(\b[55] ), .A2(new_n6742), .B1(\b[57] ), .B2(new_n6442), .C(new_n21328), .Y(new_n21329));
  O2A1O1Ixp33_ASAP7_75t_L   g21073(.A1(new_n6443), .A2(new_n17096), .B(new_n21329), .C(new_n6439), .Y(new_n21330));
  INVx1_ASAP7_75t_L         g21074(.A(new_n21330), .Y(new_n21331));
  O2A1O1Ixp33_ASAP7_75t_L   g21075(.A1(new_n6443), .A2(new_n17096), .B(new_n21329), .C(\a[44] ), .Y(new_n21332));
  AOI21xp33_ASAP7_75t_L     g21076(.A1(new_n21331), .A2(\a[44] ), .B(new_n21332), .Y(new_n21333));
  NOR2xp33_ASAP7_75t_L      g21077(.A(new_n9709), .B(new_n7318), .Y(new_n21334));
  AOI221xp5_ASAP7_75t_L     g21078(.A1(new_n7333), .A2(\b[53] ), .B1(new_n7609), .B2(\b[52] ), .C(new_n21334), .Y(new_n21335));
  O2A1O1Ixp33_ASAP7_75t_L   g21079(.A1(new_n7321), .A2(new_n9718), .B(new_n21335), .C(new_n7316), .Y(new_n21336));
  INVx1_ASAP7_75t_L         g21080(.A(new_n21336), .Y(new_n21337));
  O2A1O1Ixp33_ASAP7_75t_L   g21081(.A1(new_n7321), .A2(new_n9718), .B(new_n21335), .C(\a[47] ), .Y(new_n21338));
  AO21x2_ASAP7_75t_L        g21082(.A1(\a[47] ), .A2(new_n21337), .B(new_n21338), .Y(new_n21339));
  NOR2xp33_ASAP7_75t_L      g21083(.A(new_n7552), .B(new_n10400), .Y(new_n21340));
  AOI221xp5_ASAP7_75t_L     g21084(.A1(new_n9102), .A2(\b[48] ), .B1(new_n10398), .B2(\b[46] ), .C(new_n21340), .Y(new_n21341));
  O2A1O1Ixp33_ASAP7_75t_L   g21085(.A1(new_n9104), .A2(new_n7868), .B(new_n21341), .C(new_n9099), .Y(new_n21342));
  INVx1_ASAP7_75t_L         g21086(.A(new_n21342), .Y(new_n21343));
  O2A1O1Ixp33_ASAP7_75t_L   g21087(.A1(new_n9104), .A2(new_n7868), .B(new_n21341), .C(\a[53] ), .Y(new_n21344));
  NOR2xp33_ASAP7_75t_L      g21088(.A(new_n6944), .B(new_n10388), .Y(new_n21345));
  AOI221xp5_ASAP7_75t_L     g21089(.A1(new_n10086), .A2(\b[45] ), .B1(new_n11361), .B2(\b[43] ), .C(new_n21345), .Y(new_n21346));
  INVx1_ASAP7_75t_L         g21090(.A(new_n21346), .Y(new_n21347));
  A2O1A1Ixp33_ASAP7_75t_L   g21091(.A1(new_n7256), .A2(new_n10386), .B(new_n21347), .C(\a[56] ), .Y(new_n21348));
  O2A1O1Ixp33_ASAP7_75t_L   g21092(.A1(new_n10088), .A2(new_n7255), .B(new_n21346), .C(\a[56] ), .Y(new_n21349));
  NOR2xp33_ASAP7_75t_L      g21093(.A(new_n5855), .B(new_n11354), .Y(new_n21350));
  AOI221xp5_ASAP7_75t_L     g21094(.A1(\b[42] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[41] ), .C(new_n21350), .Y(new_n21351));
  O2A1O1Ixp33_ASAP7_75t_L   g21095(.A1(new_n11053), .A2(new_n6386), .B(new_n21351), .C(new_n11048), .Y(new_n21352));
  INVx1_ASAP7_75t_L         g21096(.A(new_n21352), .Y(new_n21353));
  O2A1O1Ixp33_ASAP7_75t_L   g21097(.A1(new_n11053), .A2(new_n6386), .B(new_n21351), .C(\a[59] ), .Y(new_n21354));
  NOR2xp33_ASAP7_75t_L      g21098(.A(new_n4581), .B(new_n13030), .Y(new_n21355));
  O2A1O1Ixp33_ASAP7_75t_L   g21099(.A1(new_n4581), .A2(new_n12672), .B(new_n21196), .C(new_n4145), .Y(new_n21356));
  AOI211xp5_ASAP7_75t_L     g21100(.A1(new_n13028), .A2(\b[35] ), .B(new_n21194), .C(\a[35] ), .Y(new_n21357));
  NOR2xp33_ASAP7_75t_L      g21101(.A(new_n21357), .B(new_n21356), .Y(new_n21358));
  INVx1_ASAP7_75t_L         g21102(.A(new_n21358), .Y(new_n21359));
  A2O1A1Ixp33_ASAP7_75t_L   g21103(.A1(new_n13028), .A2(\b[36] ), .B(new_n21355), .C(new_n21359), .Y(new_n21360));
  O2A1O1Ixp33_ASAP7_75t_L   g21104(.A1(new_n12669), .A2(new_n12671), .B(\b[36] ), .C(new_n21355), .Y(new_n21361));
  NAND2xp33_ASAP7_75t_L     g21105(.A(new_n21361), .B(new_n21358), .Y(new_n21362));
  AND2x2_ASAP7_75t_L        g21106(.A(new_n21362), .B(new_n21360), .Y(new_n21363));
  INVx1_ASAP7_75t_L         g21107(.A(new_n21363), .Y(new_n21364));
  O2A1O1Ixp33_ASAP7_75t_L   g21108(.A1(new_n21197), .A2(new_n21208), .B(new_n21202), .C(new_n21364), .Y(new_n21365));
  NOR2xp33_ASAP7_75t_L      g21109(.A(new_n21363), .B(new_n21206), .Y(new_n21366));
  NOR2xp33_ASAP7_75t_L      g21110(.A(new_n21365), .B(new_n21366), .Y(new_n21367));
  NOR2xp33_ASAP7_75t_L      g21111(.A(new_n5311), .B(new_n12318), .Y(new_n21368));
  AOI221xp5_ASAP7_75t_L     g21112(.A1(new_n11995), .A2(\b[39] ), .B1(new_n13314), .B2(\b[37] ), .C(new_n21368), .Y(new_n21369));
  INVx1_ASAP7_75t_L         g21113(.A(new_n21369), .Y(new_n21370));
  O2A1O1Ixp33_ASAP7_75t_L   g21114(.A1(new_n11998), .A2(new_n5578), .B(new_n21369), .C(new_n11987), .Y(new_n21371));
  INVx1_ASAP7_75t_L         g21115(.A(new_n21371), .Y(new_n21372));
  NOR2xp33_ASAP7_75t_L      g21116(.A(new_n11987), .B(new_n21371), .Y(new_n21373));
  A2O1A1O1Ixp25_ASAP7_75t_L g21117(.A1(new_n11997), .A2(new_n11869), .B(new_n21370), .C(new_n21372), .D(new_n21373), .Y(new_n21374));
  XNOR2x2_ASAP7_75t_L       g21118(.A(new_n21374), .B(new_n21367), .Y(new_n21375));
  A2O1A1Ixp33_ASAP7_75t_L   g21119(.A1(\a[59] ), .A2(new_n21353), .B(new_n21354), .C(new_n21375), .Y(new_n21376));
  AND2x2_ASAP7_75t_L        g21120(.A(new_n21375), .B(new_n21376), .Y(new_n21377));
  A2O1A1O1Ixp25_ASAP7_75t_L g21121(.A1(new_n21353), .A2(\a[59] ), .B(new_n21354), .C(new_n21376), .D(new_n21377), .Y(new_n21378));
  INVx1_ASAP7_75t_L         g21122(.A(new_n21378), .Y(new_n21379));
  O2A1O1Ixp33_ASAP7_75t_L   g21123(.A1(new_n21217), .A2(new_n21223), .B(new_n21214), .C(new_n21378), .Y(new_n21380));
  INVx1_ASAP7_75t_L         g21124(.A(new_n21380), .Y(new_n21381));
  O2A1O1Ixp33_ASAP7_75t_L   g21125(.A1(new_n21217), .A2(new_n21223), .B(new_n21214), .C(new_n21379), .Y(new_n21382));
  AO21x2_ASAP7_75t_L        g21126(.A1(\a[56] ), .A2(new_n21348), .B(new_n21349), .Y(new_n21383));
  A2O1A1Ixp33_ASAP7_75t_L   g21127(.A1(new_n21381), .A2(new_n21379), .B(new_n21382), .C(new_n21383), .Y(new_n21384));
  INVx1_ASAP7_75t_L         g21128(.A(new_n21212), .Y(new_n21385));
  A2O1A1Ixp33_ASAP7_75t_L   g21129(.A1(new_n21205), .A2(new_n21204), .B(new_n21201), .C(new_n21212), .Y(new_n21386));
  O2A1O1Ixp33_ASAP7_75t_L   g21130(.A1(new_n21212), .A2(new_n21213), .B(new_n21386), .C(new_n21223), .Y(new_n21387));
  O2A1O1Ixp33_ASAP7_75t_L   g21131(.A1(new_n21201), .A2(new_n21207), .B(new_n21385), .C(new_n21387), .Y(new_n21388));
  INVx1_ASAP7_75t_L         g21132(.A(new_n21351), .Y(new_n21389));
  A2O1A1Ixp33_ASAP7_75t_L   g21133(.A1(new_n6389), .A2(new_n11351), .B(new_n21389), .C(new_n11048), .Y(new_n21390));
  O2A1O1Ixp33_ASAP7_75t_L   g21134(.A1(new_n21352), .A2(new_n11048), .B(new_n21390), .C(new_n21375), .Y(new_n21391));
  A2O1A1Ixp33_ASAP7_75t_L   g21135(.A1(new_n21376), .A2(new_n21375), .B(new_n21391), .C(new_n21388), .Y(new_n21392));
  O2A1O1Ixp33_ASAP7_75t_L   g21136(.A1(new_n21388), .A2(new_n21380), .B(new_n21392), .C(new_n21383), .Y(new_n21393));
  A2O1A1O1Ixp25_ASAP7_75t_L g21137(.A1(new_n21348), .A2(\a[56] ), .B(new_n21349), .C(new_n21384), .D(new_n21393), .Y(new_n21394));
  A2O1A1O1Ixp25_ASAP7_75t_L g21138(.A1(new_n21192), .A2(\a[56] ), .B(new_n21193), .C(new_n21229), .D(new_n21225), .Y(new_n21395));
  NAND2xp33_ASAP7_75t_L     g21139(.A(new_n21395), .B(new_n21394), .Y(new_n21396));
  O2A1O1Ixp33_ASAP7_75t_L   g21140(.A1(new_n21232), .A2(new_n21233), .B(new_n21226), .C(new_n21394), .Y(new_n21397));
  INVx1_ASAP7_75t_L         g21141(.A(new_n21397), .Y(new_n21398));
  NAND2xp33_ASAP7_75t_L     g21142(.A(new_n21396), .B(new_n21398), .Y(new_n21399));
  INVx1_ASAP7_75t_L         g21143(.A(new_n21399), .Y(new_n21400));
  A2O1A1Ixp33_ASAP7_75t_L   g21144(.A1(\a[53] ), .A2(new_n21343), .B(new_n21344), .C(new_n21400), .Y(new_n21401));
  AOI211xp5_ASAP7_75t_L     g21145(.A1(new_n21343), .A2(\a[53] ), .B(new_n21344), .C(new_n21399), .Y(new_n21402));
  A2O1A1O1Ixp25_ASAP7_75t_L g21146(.A1(new_n21343), .A2(\a[53] ), .B(new_n21344), .C(new_n21401), .D(new_n21402), .Y(new_n21403));
  O2A1O1Ixp33_ASAP7_75t_L   g21147(.A1(new_n21057), .A2(new_n21068), .B(new_n21235), .C(new_n21249), .Y(new_n21404));
  NAND2xp33_ASAP7_75t_L     g21148(.A(new_n21403), .B(new_n21404), .Y(new_n21405));
  O2A1O1Ixp33_ASAP7_75t_L   g21149(.A1(new_n21240), .A2(new_n21236), .B(new_n21250), .C(new_n21403), .Y(new_n21406));
  INVx1_ASAP7_75t_L         g21150(.A(new_n21406), .Y(new_n21407));
  AND2x2_ASAP7_75t_L        g21151(.A(new_n21405), .B(new_n21407), .Y(new_n21408));
  INVx1_ASAP7_75t_L         g21152(.A(new_n21408), .Y(new_n21409));
  NOR2xp33_ASAP7_75t_L      g21153(.A(new_n8755), .B(new_n10065), .Y(new_n21410));
  AOI221xp5_ASAP7_75t_L     g21154(.A1(new_n8175), .A2(\b[51] ), .B1(new_n8484), .B2(\b[49] ), .C(new_n21410), .Y(new_n21411));
  O2A1O1Ixp33_ASAP7_75t_L   g21155(.A1(new_n8176), .A2(new_n8789), .B(new_n21411), .C(new_n8172), .Y(new_n21412));
  O2A1O1Ixp33_ASAP7_75t_L   g21156(.A1(new_n8176), .A2(new_n8789), .B(new_n21411), .C(\a[50] ), .Y(new_n21413));
  INVx1_ASAP7_75t_L         g21157(.A(new_n21413), .Y(new_n21414));
  OAI211xp5_ASAP7_75t_L     g21158(.A1(new_n8172), .A2(new_n21412), .B(new_n21409), .C(new_n21414), .Y(new_n21415));
  O2A1O1Ixp33_ASAP7_75t_L   g21159(.A1(new_n21412), .A2(new_n8172), .B(new_n21414), .C(new_n21409), .Y(new_n21416));
  INVx1_ASAP7_75t_L         g21160(.A(new_n21416), .Y(new_n21417));
  AND2x2_ASAP7_75t_L        g21161(.A(new_n21415), .B(new_n21417), .Y(new_n21418));
  INVx1_ASAP7_75t_L         g21162(.A(new_n21418), .Y(new_n21419));
  O2A1O1Ixp33_ASAP7_75t_L   g21163(.A1(new_n21252), .A2(new_n21254), .B(new_n21265), .C(new_n21419), .Y(new_n21420));
  A2O1A1O1Ixp25_ASAP7_75t_L g21164(.A1(new_n21262), .A2(\a[50] ), .B(new_n21263), .C(new_n21255), .D(new_n21256), .Y(new_n21421));
  INVx1_ASAP7_75t_L         g21165(.A(new_n21421), .Y(new_n21422));
  NOR2xp33_ASAP7_75t_L      g21166(.A(new_n21422), .B(new_n21418), .Y(new_n21423));
  NOR2xp33_ASAP7_75t_L      g21167(.A(new_n21423), .B(new_n21420), .Y(new_n21424));
  XOR2x2_ASAP7_75t_L        g21168(.A(new_n21339), .B(new_n21424), .Y(new_n21425));
  INVx1_ASAP7_75t_L         g21169(.A(new_n21425), .Y(new_n21426));
  A2O1A1O1Ixp25_ASAP7_75t_L g21170(.A1(new_n21275), .A2(new_n21276), .B(new_n21279), .C(new_n21268), .D(new_n21426), .Y(new_n21427));
  INVx1_ASAP7_75t_L         g21171(.A(new_n21427), .Y(new_n21428));
  NAND3xp33_ASAP7_75t_L     g21172(.A(new_n21426), .B(new_n21278), .C(new_n21268), .Y(new_n21429));
  NAND2xp33_ASAP7_75t_L     g21173(.A(new_n21429), .B(new_n21428), .Y(new_n21430));
  INVx1_ASAP7_75t_L         g21174(.A(new_n21332), .Y(new_n21431));
  O2A1O1Ixp33_ASAP7_75t_L   g21175(.A1(new_n21330), .A2(new_n6439), .B(new_n21431), .C(new_n21430), .Y(new_n21432));
  INVx1_ASAP7_75t_L         g21176(.A(new_n21430), .Y(new_n21433));
  NAND2xp33_ASAP7_75t_L     g21177(.A(new_n21333), .B(new_n21433), .Y(new_n21434));
  A2O1A1O1Ixp25_ASAP7_75t_L g21178(.A1(new_n21184), .A2(\a[44] ), .B(new_n21185), .C(new_n21285), .D(new_n21282), .Y(new_n21435));
  OAI211xp5_ASAP7_75t_L     g21179(.A1(new_n21432), .A2(new_n21333), .B(new_n21434), .C(new_n21435), .Y(new_n21436));
  INVx1_ASAP7_75t_L         g21180(.A(new_n21432), .Y(new_n21437));
  O2A1O1Ixp33_ASAP7_75t_L   g21181(.A1(new_n21330), .A2(new_n6439), .B(new_n21431), .C(new_n21433), .Y(new_n21438));
  INVx1_ASAP7_75t_L         g21182(.A(new_n21435), .Y(new_n21439));
  A2O1A1Ixp33_ASAP7_75t_L   g21183(.A1(new_n21437), .A2(new_n21433), .B(new_n21438), .C(new_n21439), .Y(new_n21440));
  AND2x2_ASAP7_75t_L        g21184(.A(new_n21436), .B(new_n21440), .Y(new_n21441));
  INVx1_ASAP7_75t_L         g21185(.A(new_n21441), .Y(new_n21442));
  NOR2xp33_ASAP7_75t_L      g21186(.A(new_n11626), .B(new_n5641), .Y(new_n21443));
  AOI221xp5_ASAP7_75t_L     g21187(.A1(\b[58] ), .A2(new_n5920), .B1(\b[59] ), .B2(new_n5623), .C(new_n21443), .Y(new_n21444));
  O2A1O1Ixp33_ASAP7_75t_L   g21188(.A1(new_n5630), .A2(new_n11634), .B(new_n21444), .C(new_n5626), .Y(new_n21445));
  O2A1O1Ixp33_ASAP7_75t_L   g21189(.A1(new_n5630), .A2(new_n11634), .B(new_n21444), .C(\a[41] ), .Y(new_n21446));
  INVx1_ASAP7_75t_L         g21190(.A(new_n21446), .Y(new_n21447));
  O2A1O1Ixp33_ASAP7_75t_L   g21191(.A1(new_n21445), .A2(new_n5626), .B(new_n21447), .C(new_n21442), .Y(new_n21448));
  INVx1_ASAP7_75t_L         g21192(.A(new_n21448), .Y(new_n21449));
  O2A1O1Ixp33_ASAP7_75t_L   g21193(.A1(new_n21445), .A2(new_n5626), .B(new_n21447), .C(new_n21441), .Y(new_n21450));
  AOI21xp33_ASAP7_75t_L     g21194(.A1(new_n21449), .A2(new_n21441), .B(new_n21450), .Y(new_n21451));
  A2O1A1O1Ixp25_ASAP7_75t_L g21195(.A1(new_n21179), .A2(new_n21117), .B(new_n21180), .C(new_n21286), .D(new_n21298), .Y(new_n21452));
  NAND2xp33_ASAP7_75t_L     g21196(.A(new_n21452), .B(new_n21451), .Y(new_n21453));
  O2A1O1Ixp33_ASAP7_75t_L   g21197(.A1(new_n21288), .A2(new_n21289), .B(new_n21299), .C(new_n21451), .Y(new_n21454));
  INVx1_ASAP7_75t_L         g21198(.A(new_n21454), .Y(new_n21455));
  AND2x2_ASAP7_75t_L        g21199(.A(new_n21453), .B(new_n21455), .Y(new_n21456));
  INVx1_ASAP7_75t_L         g21200(.A(new_n21456), .Y(new_n21457));
  NOR2xp33_ASAP7_75t_L      g21201(.A(new_n12956), .B(new_n4908), .Y(new_n21458));
  AOI221xp5_ASAP7_75t_L     g21202(.A1(\b[61] ), .A2(new_n5139), .B1(\b[62] ), .B2(new_n4916), .C(new_n21458), .Y(new_n21459));
  O2A1O1Ixp33_ASAP7_75t_L   g21203(.A1(new_n4911), .A2(new_n17815), .B(new_n21459), .C(new_n4906), .Y(new_n21460));
  O2A1O1Ixp33_ASAP7_75t_L   g21204(.A1(new_n4911), .A2(new_n17815), .B(new_n21459), .C(\a[38] ), .Y(new_n21461));
  INVx1_ASAP7_75t_L         g21205(.A(new_n21461), .Y(new_n21462));
  O2A1O1Ixp33_ASAP7_75t_L   g21206(.A1(new_n21460), .A2(new_n4906), .B(new_n21462), .C(new_n21457), .Y(new_n21463));
  INVx1_ASAP7_75t_L         g21207(.A(new_n21463), .Y(new_n21464));
  O2A1O1Ixp33_ASAP7_75t_L   g21208(.A1(new_n21460), .A2(new_n4906), .B(new_n21462), .C(new_n21456), .Y(new_n21465));
  AOI21xp33_ASAP7_75t_L     g21209(.A1(new_n21464), .A2(new_n21456), .B(new_n21465), .Y(new_n21466));
  NAND3xp33_ASAP7_75t_L     g21210(.A(new_n21314), .B(new_n21305), .C(new_n21466), .Y(new_n21467));
  O2A1O1Ixp33_ASAP7_75t_L   g21211(.A1(new_n21301), .A2(new_n21302), .B(new_n21314), .C(new_n21466), .Y(new_n21468));
  INVx1_ASAP7_75t_L         g21212(.A(new_n21468), .Y(new_n21469));
  NAND2xp33_ASAP7_75t_L     g21213(.A(new_n21467), .B(new_n21469), .Y(new_n21470));
  O2A1O1Ixp33_ASAP7_75t_L   g21214(.A1(new_n21320), .A2(new_n21316), .B(new_n21177), .C(new_n21470), .Y(new_n21471));
  A2O1A1Ixp33_ASAP7_75t_L   g21215(.A1(new_n21170), .A2(new_n21318), .B(new_n21316), .C(new_n21177), .Y(new_n21472));
  AOI21xp33_ASAP7_75t_L     g21216(.A1(new_n21469), .A2(new_n21467), .B(new_n21472), .Y(new_n21473));
  NOR2xp33_ASAP7_75t_L      g21217(.A(new_n21473), .B(new_n21471), .Y(new_n21474));
  A2O1A1Ixp33_ASAP7_75t_L   g21218(.A1(new_n21167), .A2(new_n21326), .B(new_n21323), .C(new_n21474), .Y(new_n21475));
  INVx1_ASAP7_75t_L         g21219(.A(new_n21475), .Y(new_n21476));
  A2O1A1Ixp33_ASAP7_75t_L   g21220(.A1(new_n21158), .A2(new_n21160), .B(new_n21163), .C(new_n21326), .Y(new_n21477));
  A2O1A1Ixp33_ASAP7_75t_L   g21221(.A1(new_n21155), .A2(new_n21324), .B(new_n21322), .C(new_n21477), .Y(new_n21478));
  NOR2xp33_ASAP7_75t_L      g21222(.A(new_n21474), .B(new_n21478), .Y(new_n21479));
  NOR2xp33_ASAP7_75t_L      g21223(.A(new_n21476), .B(new_n21479), .Y(\f[99] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21224(.A1(new_n21306), .A2(new_n21314), .B(new_n21315), .C(new_n21319), .Y(new_n21481));
  A2O1A1Ixp33_ASAP7_75t_L   g21225(.A1(new_n21287), .A2(new_n21299), .B(new_n21451), .C(new_n21449), .Y(new_n21482));
  AOI22xp33_ASAP7_75t_L     g21226(.A1(new_n4916), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5139), .Y(new_n21483));
  INVx1_ASAP7_75t_L         g21227(.A(new_n21483), .Y(new_n21484));
  A2O1A1Ixp33_ASAP7_75t_L   g21228(.A1(new_n4905), .A2(new_n4907), .B(new_n4649), .C(new_n21483), .Y(new_n21485));
  O2A1O1Ixp33_ASAP7_75t_L   g21229(.A1(new_n21484), .A2(new_n17329), .B(new_n21485), .C(new_n4906), .Y(new_n21486));
  O2A1O1Ixp33_ASAP7_75t_L   g21230(.A1(new_n4911), .A2(new_n12993), .B(new_n21483), .C(\a[38] ), .Y(new_n21487));
  OAI21xp33_ASAP7_75t_L     g21231(.A1(new_n21486), .A2(new_n21487), .B(new_n21482), .Y(new_n21488));
  NOR2xp33_ASAP7_75t_L      g21232(.A(new_n21487), .B(new_n21486), .Y(new_n21489));
  NAND3xp33_ASAP7_75t_L     g21233(.A(new_n21455), .B(new_n21449), .C(new_n21489), .Y(new_n21490));
  NAND2xp33_ASAP7_75t_L     g21234(.A(new_n21488), .B(new_n21490), .Y(new_n21491));
  NOR2xp33_ASAP7_75t_L      g21235(.A(new_n10309), .B(new_n7318), .Y(new_n21492));
  AOI221xp5_ASAP7_75t_L     g21236(.A1(new_n7333), .A2(\b[54] ), .B1(new_n7609), .B2(\b[53] ), .C(new_n21492), .Y(new_n21493));
  O2A1O1Ixp33_ASAP7_75t_L   g21237(.A1(new_n7321), .A2(new_n15849), .B(new_n21493), .C(new_n7316), .Y(new_n21494));
  INVx1_ASAP7_75t_L         g21238(.A(new_n21494), .Y(new_n21495));
  O2A1O1Ixp33_ASAP7_75t_L   g21239(.A1(new_n7321), .A2(new_n15849), .B(new_n21493), .C(\a[47] ), .Y(new_n21496));
  NOR2xp33_ASAP7_75t_L      g21240(.A(new_n7249), .B(new_n10388), .Y(new_n21497));
  AOI221xp5_ASAP7_75t_L     g21241(.A1(new_n10086), .A2(\b[46] ), .B1(new_n11361), .B2(\b[44] ), .C(new_n21497), .Y(new_n21498));
  O2A1O1Ixp33_ASAP7_75t_L   g21242(.A1(new_n10088), .A2(new_n7279), .B(new_n21498), .C(new_n10083), .Y(new_n21499));
  INVx1_ASAP7_75t_L         g21243(.A(new_n21499), .Y(new_n21500));
  O2A1O1Ixp33_ASAP7_75t_L   g21244(.A1(new_n10088), .A2(new_n7279), .B(new_n21498), .C(\a[56] ), .Y(new_n21501));
  NOR2xp33_ASAP7_75t_L      g21245(.A(new_n4613), .B(new_n13030), .Y(new_n21502));
  O2A1O1Ixp33_ASAP7_75t_L   g21246(.A1(new_n12669), .A2(new_n12671), .B(\b[37] ), .C(new_n21502), .Y(new_n21503));
  INVx1_ASAP7_75t_L         g21247(.A(new_n21503), .Y(new_n21504));
  O2A1O1Ixp33_ASAP7_75t_L   g21248(.A1(new_n4581), .A2(new_n12672), .B(new_n21196), .C(\a[35] ), .Y(new_n21505));
  INVx1_ASAP7_75t_L         g21249(.A(new_n21505), .Y(new_n21506));
  O2A1O1Ixp33_ASAP7_75t_L   g21250(.A1(new_n21361), .A2(new_n21358), .B(new_n21506), .C(new_n21504), .Y(new_n21507));
  NOR2xp33_ASAP7_75t_L      g21251(.A(new_n21504), .B(new_n21507), .Y(new_n21508));
  O2A1O1Ixp33_ASAP7_75t_L   g21252(.A1(new_n21361), .A2(new_n21358), .B(new_n21506), .C(new_n21503), .Y(new_n21509));
  NOR2xp33_ASAP7_75t_L      g21253(.A(new_n5570), .B(new_n12318), .Y(new_n21510));
  AOI221xp5_ASAP7_75t_L     g21254(.A1(new_n11995), .A2(\b[40] ), .B1(new_n13314), .B2(\b[38] ), .C(new_n21510), .Y(new_n21511));
  O2A1O1Ixp33_ASAP7_75t_L   g21255(.A1(new_n11998), .A2(new_n5862), .B(new_n21511), .C(new_n11987), .Y(new_n21512));
  O2A1O1Ixp33_ASAP7_75t_L   g21256(.A1(new_n11998), .A2(new_n5862), .B(new_n21511), .C(\a[62] ), .Y(new_n21513));
  INVx1_ASAP7_75t_L         g21257(.A(new_n21513), .Y(new_n21514));
  INVx1_ASAP7_75t_L         g21258(.A(new_n21360), .Y(new_n21515));
  INVx1_ASAP7_75t_L         g21259(.A(new_n21507), .Y(new_n21516));
  O2A1O1Ixp33_ASAP7_75t_L   g21260(.A1(new_n21505), .A2(new_n21515), .B(new_n21516), .C(new_n21508), .Y(new_n21517));
  O2A1O1Ixp33_ASAP7_75t_L   g21261(.A1(new_n11987), .A2(new_n21512), .B(new_n21514), .C(new_n21517), .Y(new_n21518));
  INVx1_ASAP7_75t_L         g21262(.A(new_n21518), .Y(new_n21519));
  INVx1_ASAP7_75t_L         g21263(.A(new_n21517), .Y(new_n21520));
  O2A1O1Ixp33_ASAP7_75t_L   g21264(.A1(new_n11987), .A2(new_n21512), .B(new_n21514), .C(new_n21520), .Y(new_n21521));
  O2A1O1Ixp33_ASAP7_75t_L   g21265(.A1(new_n21508), .A2(new_n21509), .B(new_n21519), .C(new_n21521), .Y(new_n21522));
  O2A1O1Ixp33_ASAP7_75t_L   g21266(.A1(new_n11998), .A2(new_n5578), .B(new_n21369), .C(\a[62] ), .Y(new_n21523));
  O2A1O1Ixp33_ASAP7_75t_L   g21267(.A1(new_n21373), .A2(new_n21523), .B(new_n21367), .C(new_n21365), .Y(new_n21524));
  NAND2xp33_ASAP7_75t_L     g21268(.A(new_n21522), .B(new_n21524), .Y(new_n21525));
  A2O1A1Ixp33_ASAP7_75t_L   g21269(.A1(\a[62] ), .A2(new_n21372), .B(new_n21523), .C(new_n21367), .Y(new_n21526));
  O2A1O1Ixp33_ASAP7_75t_L   g21270(.A1(new_n21205), .A2(new_n21364), .B(new_n21526), .C(new_n21522), .Y(new_n21527));
  INVx1_ASAP7_75t_L         g21271(.A(new_n21527), .Y(new_n21528));
  AND2x2_ASAP7_75t_L        g21272(.A(new_n21525), .B(new_n21528), .Y(new_n21529));
  NOR2xp33_ASAP7_75t_L      g21273(.A(new_n6110), .B(new_n11354), .Y(new_n21530));
  AOI221xp5_ASAP7_75t_L     g21274(.A1(\b[43] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[42] ), .C(new_n21530), .Y(new_n21531));
  O2A1O1Ixp33_ASAP7_75t_L   g21275(.A1(new_n11053), .A2(new_n6679), .B(new_n21531), .C(new_n11048), .Y(new_n21532));
  INVx1_ASAP7_75t_L         g21276(.A(new_n21532), .Y(new_n21533));
  O2A1O1Ixp33_ASAP7_75t_L   g21277(.A1(new_n11053), .A2(new_n6679), .B(new_n21531), .C(\a[59] ), .Y(new_n21534));
  A2O1A1Ixp33_ASAP7_75t_L   g21278(.A1(\a[59] ), .A2(new_n21533), .B(new_n21534), .C(new_n21529), .Y(new_n21535));
  INVx1_ASAP7_75t_L         g21279(.A(new_n21534), .Y(new_n21536));
  O2A1O1Ixp33_ASAP7_75t_L   g21280(.A1(new_n21532), .A2(new_n11048), .B(new_n21536), .C(new_n21529), .Y(new_n21537));
  AOI21xp33_ASAP7_75t_L     g21281(.A1(new_n21535), .A2(new_n21529), .B(new_n21537), .Y(new_n21538));
  A2O1A1O1Ixp25_ASAP7_75t_L g21282(.A1(new_n21353), .A2(\a[59] ), .B(new_n21354), .C(new_n21375), .D(new_n21380), .Y(new_n21539));
  NAND2xp33_ASAP7_75t_L     g21283(.A(new_n21538), .B(new_n21539), .Y(new_n21540));
  O2A1O1Ixp33_ASAP7_75t_L   g21284(.A1(new_n21378), .A2(new_n21388), .B(new_n21376), .C(new_n21538), .Y(new_n21541));
  INVx1_ASAP7_75t_L         g21285(.A(new_n21541), .Y(new_n21542));
  NAND2xp33_ASAP7_75t_L     g21286(.A(new_n21542), .B(new_n21540), .Y(new_n21543));
  INVx1_ASAP7_75t_L         g21287(.A(new_n21501), .Y(new_n21544));
  O2A1O1Ixp33_ASAP7_75t_L   g21288(.A1(new_n21499), .A2(new_n10083), .B(new_n21544), .C(new_n21543), .Y(new_n21545));
  INVx1_ASAP7_75t_L         g21289(.A(new_n21545), .Y(new_n21546));
  NOR2xp33_ASAP7_75t_L      g21290(.A(new_n21543), .B(new_n21545), .Y(new_n21547));
  A2O1A1O1Ixp25_ASAP7_75t_L g21291(.A1(new_n21500), .A2(\a[56] ), .B(new_n21501), .C(new_n21546), .D(new_n21547), .Y(new_n21548));
  A2O1A1O1Ixp25_ASAP7_75t_L g21292(.A1(new_n21381), .A2(new_n21379), .B(new_n21382), .C(new_n21383), .D(new_n21397), .Y(new_n21549));
  NAND2xp33_ASAP7_75t_L     g21293(.A(new_n21549), .B(new_n21548), .Y(new_n21550));
  INVx1_ASAP7_75t_L         g21294(.A(new_n21543), .Y(new_n21551));
  O2A1O1Ixp33_ASAP7_75t_L   g21295(.A1(new_n21499), .A2(new_n10083), .B(new_n21544), .C(new_n21551), .Y(new_n21552));
  INVx1_ASAP7_75t_L         g21296(.A(new_n21552), .Y(new_n21553));
  O2A1O1Ixp33_ASAP7_75t_L   g21297(.A1(new_n21543), .A2(new_n21545), .B(new_n21553), .C(new_n21549), .Y(new_n21554));
  INVx1_ASAP7_75t_L         g21298(.A(new_n21554), .Y(new_n21555));
  AND2x2_ASAP7_75t_L        g21299(.A(new_n21550), .B(new_n21555), .Y(new_n21556));
  NOR2xp33_ASAP7_75t_L      g21300(.A(new_n7860), .B(new_n10400), .Y(new_n21557));
  AOI221xp5_ASAP7_75t_L     g21301(.A1(new_n9102), .A2(\b[49] ), .B1(new_n10398), .B2(\b[47] ), .C(new_n21557), .Y(new_n21558));
  O2A1O1Ixp33_ASAP7_75t_L   g21302(.A1(new_n9104), .A2(new_n14802), .B(new_n21558), .C(new_n9099), .Y(new_n21559));
  INVx1_ASAP7_75t_L         g21303(.A(new_n21559), .Y(new_n21560));
  O2A1O1Ixp33_ASAP7_75t_L   g21304(.A1(new_n9104), .A2(new_n14802), .B(new_n21558), .C(\a[53] ), .Y(new_n21561));
  A2O1A1Ixp33_ASAP7_75t_L   g21305(.A1(\a[53] ), .A2(new_n21560), .B(new_n21561), .C(new_n21556), .Y(new_n21562));
  INVx1_ASAP7_75t_L         g21306(.A(new_n21561), .Y(new_n21563));
  O2A1O1Ixp33_ASAP7_75t_L   g21307(.A1(new_n21559), .A2(new_n9099), .B(new_n21563), .C(new_n21556), .Y(new_n21564));
  AOI21xp33_ASAP7_75t_L     g21308(.A1(new_n21562), .A2(new_n21556), .B(new_n21564), .Y(new_n21565));
  AND3x1_ASAP7_75t_L        g21309(.A(new_n21407), .B(new_n21565), .C(new_n21401), .Y(new_n21566));
  A2O1A1O1Ixp25_ASAP7_75t_L g21310(.A1(new_n21238), .A2(new_n21250), .B(new_n21403), .C(new_n21401), .D(new_n21565), .Y(new_n21567));
  NOR2xp33_ASAP7_75t_L      g21311(.A(new_n21567), .B(new_n21566), .Y(new_n21568));
  NOR2xp33_ASAP7_75t_L      g21312(.A(new_n8779), .B(new_n10065), .Y(new_n21569));
  AOI221xp5_ASAP7_75t_L     g21313(.A1(new_n8175), .A2(\b[52] ), .B1(new_n8484), .B2(\b[50] ), .C(new_n21569), .Y(new_n21570));
  O2A1O1Ixp33_ASAP7_75t_L   g21314(.A1(new_n8176), .A2(new_n17363), .B(new_n21570), .C(new_n8172), .Y(new_n21571));
  INVx1_ASAP7_75t_L         g21315(.A(new_n21571), .Y(new_n21572));
  O2A1O1Ixp33_ASAP7_75t_L   g21316(.A1(new_n8176), .A2(new_n17363), .B(new_n21570), .C(\a[50] ), .Y(new_n21573));
  A2O1A1Ixp33_ASAP7_75t_L   g21317(.A1(\a[50] ), .A2(new_n21572), .B(new_n21573), .C(new_n21568), .Y(new_n21574));
  A2O1A1Ixp33_ASAP7_75t_L   g21318(.A1(new_n21572), .A2(\a[50] ), .B(new_n21573), .C(new_n21574), .Y(new_n21575));
  INVx1_ASAP7_75t_L         g21319(.A(new_n21575), .Y(new_n21576));
  AOI21xp33_ASAP7_75t_L     g21320(.A1(new_n21574), .A2(new_n21568), .B(new_n21576), .Y(new_n21577));
  O2A1O1Ixp33_ASAP7_75t_L   g21321(.A1(new_n21421), .A2(new_n21419), .B(new_n21417), .C(new_n21577), .Y(new_n21578));
  INVx1_ASAP7_75t_L         g21322(.A(new_n21578), .Y(new_n21579));
  O2A1O1Ixp33_ASAP7_75t_L   g21323(.A1(new_n21421), .A2(new_n21419), .B(new_n21417), .C(new_n21578), .Y(new_n21580));
  A2O1A1O1Ixp25_ASAP7_75t_L g21324(.A1(new_n21574), .A2(new_n21568), .B(new_n21576), .C(new_n21579), .D(new_n21580), .Y(new_n21581));
  INVx1_ASAP7_75t_L         g21325(.A(new_n21496), .Y(new_n21582));
  O2A1O1Ixp33_ASAP7_75t_L   g21326(.A1(new_n21494), .A2(new_n7316), .B(new_n21582), .C(new_n21581), .Y(new_n21583));
  INVx1_ASAP7_75t_L         g21327(.A(new_n21583), .Y(new_n21584));
  O2A1O1Ixp33_ASAP7_75t_L   g21328(.A1(new_n21256), .A2(new_n21266), .B(new_n21415), .C(new_n21416), .Y(new_n21585));
  A2O1A1Ixp33_ASAP7_75t_L   g21329(.A1(new_n21574), .A2(new_n21568), .B(new_n21576), .C(new_n21585), .Y(new_n21586));
  O2A1O1Ixp33_ASAP7_75t_L   g21330(.A1(new_n21585), .A2(new_n21578), .B(new_n21586), .C(new_n21583), .Y(new_n21587));
  A2O1A1O1Ixp25_ASAP7_75t_L g21331(.A1(new_n21495), .A2(\a[47] ), .B(new_n21496), .C(new_n21584), .D(new_n21587), .Y(new_n21588));
  A2O1A1O1Ixp25_ASAP7_75t_L g21332(.A1(new_n21337), .A2(\a[47] ), .B(new_n21338), .C(new_n21424), .D(new_n21427), .Y(new_n21589));
  NAND2xp33_ASAP7_75t_L     g21333(.A(new_n21589), .B(new_n21588), .Y(new_n21590));
  A2O1A1Ixp33_ASAP7_75t_L   g21334(.A1(\a[47] ), .A2(new_n21495), .B(new_n21496), .C(new_n21581), .Y(new_n21591));
  O2A1O1Ixp33_ASAP7_75t_L   g21335(.A1(new_n21581), .A2(new_n21583), .B(new_n21591), .C(new_n21589), .Y(new_n21592));
  INVx1_ASAP7_75t_L         g21336(.A(new_n21592), .Y(new_n21593));
  NAND2xp33_ASAP7_75t_L     g21337(.A(new_n21590), .B(new_n21593), .Y(new_n21594));
  INVx1_ASAP7_75t_L         g21338(.A(new_n21594), .Y(new_n21595));
  NOR2xp33_ASAP7_75t_L      g21339(.A(new_n10978), .B(new_n7304), .Y(new_n21596));
  AOI221xp5_ASAP7_75t_L     g21340(.A1(\b[56] ), .A2(new_n6742), .B1(\b[58] ), .B2(new_n6442), .C(new_n21596), .Y(new_n21597));
  O2A1O1Ixp33_ASAP7_75t_L   g21341(.A1(new_n6443), .A2(new_n20073), .B(new_n21597), .C(new_n6439), .Y(new_n21598));
  O2A1O1Ixp33_ASAP7_75t_L   g21342(.A1(new_n6443), .A2(new_n20073), .B(new_n21597), .C(\a[44] ), .Y(new_n21599));
  INVx1_ASAP7_75t_L         g21343(.A(new_n21599), .Y(new_n21600));
  O2A1O1Ixp33_ASAP7_75t_L   g21344(.A1(new_n21598), .A2(new_n6439), .B(new_n21600), .C(new_n21594), .Y(new_n21601));
  INVx1_ASAP7_75t_L         g21345(.A(new_n21601), .Y(new_n21602));
  NAND2xp33_ASAP7_75t_L     g21346(.A(new_n21595), .B(new_n21602), .Y(new_n21603));
  O2A1O1Ixp33_ASAP7_75t_L   g21347(.A1(new_n21598), .A2(new_n6439), .B(new_n21600), .C(new_n21595), .Y(new_n21604));
  INVx1_ASAP7_75t_L         g21348(.A(new_n21604), .Y(new_n21605));
  O2A1O1Ixp33_ASAP7_75t_L   g21349(.A1(new_n21433), .A2(new_n21438), .B(new_n21439), .C(new_n21432), .Y(new_n21606));
  NAND3xp33_ASAP7_75t_L     g21350(.A(new_n21603), .B(new_n21605), .C(new_n21606), .Y(new_n21607));
  O2A1O1Ixp33_ASAP7_75t_L   g21351(.A1(new_n21594), .A2(new_n21601), .B(new_n21605), .C(new_n21606), .Y(new_n21608));
  INVx1_ASAP7_75t_L         g21352(.A(new_n21608), .Y(new_n21609));
  AND2x2_ASAP7_75t_L        g21353(.A(new_n21607), .B(new_n21609), .Y(new_n21610));
  NOR2xp33_ASAP7_75t_L      g21354(.A(new_n12258), .B(new_n5641), .Y(new_n21611));
  AOI221xp5_ASAP7_75t_L     g21355(.A1(\b[59] ), .A2(new_n5920), .B1(\b[60] ), .B2(new_n5623), .C(new_n21611), .Y(new_n21612));
  O2A1O1Ixp33_ASAP7_75t_L   g21356(.A1(new_n5630), .A2(new_n14764), .B(new_n21612), .C(new_n5626), .Y(new_n21613));
  INVx1_ASAP7_75t_L         g21357(.A(new_n21613), .Y(new_n21614));
  O2A1O1Ixp33_ASAP7_75t_L   g21358(.A1(new_n5630), .A2(new_n14764), .B(new_n21612), .C(\a[41] ), .Y(new_n21615));
  A2O1A1Ixp33_ASAP7_75t_L   g21359(.A1(\a[41] ), .A2(new_n21614), .B(new_n21615), .C(new_n21610), .Y(new_n21616));
  NOR2xp33_ASAP7_75t_L      g21360(.A(new_n5626), .B(new_n21613), .Y(new_n21617));
  OR3x1_ASAP7_75t_L         g21361(.A(new_n21610), .B(new_n21617), .C(new_n21615), .Y(new_n21618));
  AND3x1_ASAP7_75t_L        g21362(.A(new_n21490), .B(new_n21618), .C(new_n21488), .Y(new_n21619));
  NAND3xp33_ASAP7_75t_L     g21363(.A(new_n21491), .B(new_n21616), .C(new_n21618), .Y(new_n21620));
  A2O1A1Ixp33_ASAP7_75t_L   g21364(.A1(new_n21616), .A2(new_n21619), .B(new_n21491), .C(new_n21620), .Y(new_n21621));
  INVx1_ASAP7_75t_L         g21365(.A(new_n21621), .Y(new_n21622));
  A2O1A1Ixp33_ASAP7_75t_L   g21366(.A1(new_n21139), .A2(new_n21127), .B(new_n21301), .C(new_n21314), .Y(new_n21623));
  O2A1O1Ixp33_ASAP7_75t_L   g21367(.A1(new_n21465), .A2(new_n21456), .B(new_n21623), .C(new_n21463), .Y(new_n21624));
  NAND2xp33_ASAP7_75t_L     g21368(.A(new_n21622), .B(new_n21624), .Y(new_n21625));
  A2O1A1O1Ixp25_ASAP7_75t_L g21369(.A1(new_n21305), .A2(new_n21314), .B(new_n21466), .C(new_n21464), .D(new_n21622), .Y(new_n21626));
  INVx1_ASAP7_75t_L         g21370(.A(new_n21626), .Y(new_n21627));
  AND2x2_ASAP7_75t_L        g21371(.A(new_n21625), .B(new_n21627), .Y(new_n21628));
  INVx1_ASAP7_75t_L         g21372(.A(new_n21628), .Y(new_n21629));
  A2O1A1O1Ixp25_ASAP7_75t_L g21373(.A1(new_n21177), .A2(new_n21481), .B(new_n21470), .C(new_n21475), .D(new_n21629), .Y(new_n21630));
  A2O1A1Ixp33_ASAP7_75t_L   g21374(.A1(new_n21481), .A2(new_n21177), .B(new_n21470), .C(new_n21475), .Y(new_n21631));
  NOR2xp33_ASAP7_75t_L      g21375(.A(new_n21628), .B(new_n21631), .Y(new_n21632));
  NOR2xp33_ASAP7_75t_L      g21376(.A(new_n21630), .B(new_n21632), .Y(\f[100] ));
  INVx1_ASAP7_75t_L         g21377(.A(new_n21471), .Y(new_n21634));
  A2O1A1Ixp33_ASAP7_75t_L   g21378(.A1(new_n21475), .A2(new_n21634), .B(new_n21629), .C(new_n21627), .Y(new_n21635));
  INVx1_ASAP7_75t_L         g21379(.A(new_n21491), .Y(new_n21636));
  NAND3xp33_ASAP7_75t_L     g21380(.A(new_n21636), .B(new_n21616), .C(new_n21618), .Y(new_n21637));
  O2A1O1Ixp33_ASAP7_75t_L   g21381(.A1(new_n21617), .A2(new_n21615), .B(new_n21607), .C(new_n21608), .Y(new_n21638));
  INVx1_ASAP7_75t_L         g21382(.A(new_n21638), .Y(new_n21639));
  NOR2xp33_ASAP7_75t_L      g21383(.A(new_n12956), .B(new_n5144), .Y(new_n21640));
  A2O1A1Ixp33_ASAP7_75t_L   g21384(.A1(new_n12986), .A2(new_n4912), .B(new_n21640), .C(\a[38] ), .Y(new_n21641));
  INVx1_ASAP7_75t_L         g21385(.A(new_n21641), .Y(new_n21642));
  A2O1A1Ixp33_ASAP7_75t_L   g21386(.A1(new_n12986), .A2(new_n4912), .B(new_n21640), .C(new_n4906), .Y(new_n21643));
  O2A1O1Ixp33_ASAP7_75t_L   g21387(.A1(new_n21642), .A2(new_n4906), .B(new_n21643), .C(new_n21638), .Y(new_n21644));
  INVx1_ASAP7_75t_L         g21388(.A(new_n21644), .Y(new_n21645));
  O2A1O1Ixp33_ASAP7_75t_L   g21389(.A1(new_n21642), .A2(new_n4906), .B(new_n21643), .C(new_n21639), .Y(new_n21646));
  NOR2xp33_ASAP7_75t_L      g21390(.A(new_n10309), .B(new_n7312), .Y(new_n21647));
  AOI221xp5_ASAP7_75t_L     g21391(.A1(\b[54] ), .A2(new_n7609), .B1(\b[56] ), .B2(new_n7334), .C(new_n21647), .Y(new_n21648));
  INVx1_ASAP7_75t_L         g21392(.A(new_n21648), .Y(new_n21649));
  A2O1A1Ixp33_ASAP7_75t_L   g21393(.A1(new_n11579), .A2(new_n7322), .B(new_n21649), .C(\a[47] ), .Y(new_n21650));
  O2A1O1Ixp33_ASAP7_75t_L   g21394(.A1(new_n7321), .A2(new_n10339), .B(new_n21648), .C(\a[47] ), .Y(new_n21651));
  AO21x2_ASAP7_75t_L        g21395(.A1(\a[47] ), .A2(new_n21650), .B(new_n21651), .Y(new_n21652));
  A2O1A1O1Ixp25_ASAP7_75t_L g21396(.A1(new_n21343), .A2(\a[53] ), .B(new_n21344), .C(new_n21400), .D(new_n21406), .Y(new_n21653));
  A2O1A1O1Ixp25_ASAP7_75t_L g21397(.A1(new_n21560), .A2(\a[53] ), .B(new_n21561), .C(new_n21550), .D(new_n21554), .Y(new_n21654));
  INVx1_ASAP7_75t_L         g21398(.A(new_n21654), .Y(new_n21655));
  NOR2xp33_ASAP7_75t_L      g21399(.A(new_n7270), .B(new_n10388), .Y(new_n21656));
  AOI221xp5_ASAP7_75t_L     g21400(.A1(new_n10086), .A2(\b[47] ), .B1(new_n11361), .B2(\b[45] ), .C(new_n21656), .Y(new_n21657));
  O2A1O1Ixp33_ASAP7_75t_L   g21401(.A1(new_n10088), .A2(new_n7560), .B(new_n21657), .C(new_n10083), .Y(new_n21658));
  INVx1_ASAP7_75t_L         g21402(.A(new_n21658), .Y(new_n21659));
  O2A1O1Ixp33_ASAP7_75t_L   g21403(.A1(new_n10088), .A2(new_n7560), .B(new_n21657), .C(\a[56] ), .Y(new_n21660));
  O2A1O1Ixp33_ASAP7_75t_L   g21404(.A1(new_n21515), .A2(new_n21505), .B(new_n21503), .C(new_n21518), .Y(new_n21661));
  NOR2xp33_ASAP7_75t_L      g21405(.A(new_n5074), .B(new_n13030), .Y(new_n21662));
  INVx1_ASAP7_75t_L         g21406(.A(new_n21662), .Y(new_n21663));
  O2A1O1Ixp33_ASAP7_75t_L   g21407(.A1(new_n12672), .A2(new_n5311), .B(new_n21663), .C(new_n21504), .Y(new_n21664));
  O2A1O1Ixp33_ASAP7_75t_L   g21408(.A1(new_n12672), .A2(new_n5311), .B(new_n21663), .C(new_n21503), .Y(new_n21665));
  INVx1_ASAP7_75t_L         g21409(.A(new_n21665), .Y(new_n21666));
  O2A1O1Ixp33_ASAP7_75t_L   g21410(.A1(new_n21664), .A2(new_n21504), .B(new_n21666), .C(new_n21661), .Y(new_n21667));
  INVx1_ASAP7_75t_L         g21411(.A(new_n21667), .Y(new_n21668));
  O2A1O1Ixp33_ASAP7_75t_L   g21412(.A1(new_n21504), .A2(new_n21664), .B(new_n21666), .C(new_n21667), .Y(new_n21669));
  O2A1O1Ixp33_ASAP7_75t_L   g21413(.A1(new_n21507), .A2(new_n21518), .B(new_n21668), .C(new_n21669), .Y(new_n21670));
  INVx1_ASAP7_75t_L         g21414(.A(new_n21670), .Y(new_n21671));
  NOR2xp33_ASAP7_75t_L      g21415(.A(new_n5855), .B(new_n12318), .Y(new_n21672));
  AOI221xp5_ASAP7_75t_L     g21416(.A1(new_n11995), .A2(\b[41] ), .B1(new_n13314), .B2(\b[39] ), .C(new_n21672), .Y(new_n21673));
  O2A1O1Ixp33_ASAP7_75t_L   g21417(.A1(new_n11998), .A2(new_n6117), .B(new_n21673), .C(new_n11987), .Y(new_n21674));
  OAI21xp33_ASAP7_75t_L     g21418(.A1(new_n11998), .A2(new_n6117), .B(new_n21673), .Y(new_n21675));
  NAND2xp33_ASAP7_75t_L     g21419(.A(new_n11987), .B(new_n21675), .Y(new_n21676));
  O2A1O1Ixp33_ASAP7_75t_L   g21420(.A1(new_n21674), .A2(new_n11987), .B(new_n21676), .C(new_n21670), .Y(new_n21677));
  INVx1_ASAP7_75t_L         g21421(.A(new_n21677), .Y(new_n21678));
  O2A1O1Ixp33_ASAP7_75t_L   g21422(.A1(new_n21674), .A2(new_n11987), .B(new_n21676), .C(new_n21671), .Y(new_n21679));
  NOR2xp33_ASAP7_75t_L      g21423(.A(new_n6378), .B(new_n11354), .Y(new_n21680));
  AOI221xp5_ASAP7_75t_L     g21424(.A1(\b[44] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[43] ), .C(new_n21680), .Y(new_n21681));
  O2A1O1Ixp33_ASAP7_75t_L   g21425(.A1(new_n11053), .A2(new_n6951), .B(new_n21681), .C(new_n11048), .Y(new_n21682));
  INVx1_ASAP7_75t_L         g21426(.A(new_n21682), .Y(new_n21683));
  O2A1O1Ixp33_ASAP7_75t_L   g21427(.A1(new_n11053), .A2(new_n6951), .B(new_n21681), .C(\a[59] ), .Y(new_n21684));
  AOI21xp33_ASAP7_75t_L     g21428(.A1(new_n21683), .A2(\a[59] ), .B(new_n21684), .Y(new_n21685));
  A2O1A1Ixp33_ASAP7_75t_L   g21429(.A1(new_n21678), .A2(new_n21671), .B(new_n21679), .C(new_n21685), .Y(new_n21686));
  A2O1A1O1Ixp25_ASAP7_75t_L g21430(.A1(new_n13028), .A2(\b[36] ), .B(new_n21355), .C(new_n21359), .D(new_n21505), .Y(new_n21687));
  O2A1O1Ixp33_ASAP7_75t_L   g21431(.A1(new_n21504), .A2(new_n21687), .B(new_n21519), .C(new_n21667), .Y(new_n21688));
  O2A1O1Ixp33_ASAP7_75t_L   g21432(.A1(new_n21688), .A2(new_n21669), .B(new_n21678), .C(new_n21679), .Y(new_n21689));
  A2O1A1Ixp33_ASAP7_75t_L   g21433(.A1(\a[59] ), .A2(new_n21683), .B(new_n21684), .C(new_n21689), .Y(new_n21690));
  AND2x2_ASAP7_75t_L        g21434(.A(new_n21686), .B(new_n21690), .Y(new_n21691));
  A2O1A1O1Ixp25_ASAP7_75t_L g21435(.A1(new_n21533), .A2(\a[59] ), .B(new_n21534), .C(new_n21525), .D(new_n21527), .Y(new_n21692));
  NAND2xp33_ASAP7_75t_L     g21436(.A(new_n21692), .B(new_n21691), .Y(new_n21693));
  O2A1O1Ixp33_ASAP7_75t_L   g21437(.A1(new_n21522), .A2(new_n21524), .B(new_n21535), .C(new_n21691), .Y(new_n21694));
  INVx1_ASAP7_75t_L         g21438(.A(new_n21694), .Y(new_n21695));
  AND2x2_ASAP7_75t_L        g21439(.A(new_n21693), .B(new_n21695), .Y(new_n21696));
  A2O1A1Ixp33_ASAP7_75t_L   g21440(.A1(\a[56] ), .A2(new_n21659), .B(new_n21660), .C(new_n21696), .Y(new_n21697));
  AND2x2_ASAP7_75t_L        g21441(.A(new_n21696), .B(new_n21697), .Y(new_n21698));
  A2O1A1O1Ixp25_ASAP7_75t_L g21442(.A1(new_n21659), .A2(\a[56] ), .B(new_n21660), .C(new_n21697), .D(new_n21698), .Y(new_n21699));
  A2O1A1O1Ixp25_ASAP7_75t_L g21443(.A1(new_n21500), .A2(\a[56] ), .B(new_n21501), .C(new_n21540), .D(new_n21541), .Y(new_n21700));
  NAND2xp33_ASAP7_75t_L     g21444(.A(new_n21700), .B(new_n21699), .Y(new_n21701));
  O2A1O1Ixp33_ASAP7_75t_L   g21445(.A1(new_n21538), .A2(new_n21539), .B(new_n21546), .C(new_n21699), .Y(new_n21702));
  INVx1_ASAP7_75t_L         g21446(.A(new_n21702), .Y(new_n21703));
  AND2x2_ASAP7_75t_L        g21447(.A(new_n21701), .B(new_n21703), .Y(new_n21704));
  NOR2xp33_ASAP7_75t_L      g21448(.A(new_n8427), .B(new_n10400), .Y(new_n21705));
  AOI221xp5_ASAP7_75t_L     g21449(.A1(new_n9102), .A2(\b[50] ), .B1(new_n10398), .B2(\b[48] ), .C(new_n21705), .Y(new_n21706));
  O2A1O1Ixp33_ASAP7_75t_L   g21450(.A1(new_n9104), .A2(new_n8764), .B(new_n21706), .C(new_n9099), .Y(new_n21707));
  INVx1_ASAP7_75t_L         g21451(.A(new_n21707), .Y(new_n21708));
  O2A1O1Ixp33_ASAP7_75t_L   g21452(.A1(new_n9104), .A2(new_n8764), .B(new_n21706), .C(\a[53] ), .Y(new_n21709));
  AOI211xp5_ASAP7_75t_L     g21453(.A1(new_n21708), .A2(\a[53] ), .B(new_n21709), .C(new_n21704), .Y(new_n21710));
  A2O1A1Ixp33_ASAP7_75t_L   g21454(.A1(\a[53] ), .A2(new_n21708), .B(new_n21709), .C(new_n21704), .Y(new_n21711));
  INVx1_ASAP7_75t_L         g21455(.A(new_n21711), .Y(new_n21712));
  NOR2xp33_ASAP7_75t_L      g21456(.A(new_n21710), .B(new_n21712), .Y(new_n21713));
  NAND2xp33_ASAP7_75t_L     g21457(.A(new_n21655), .B(new_n21713), .Y(new_n21714));
  NOR2xp33_ASAP7_75t_L      g21458(.A(new_n9355), .B(new_n10065), .Y(new_n21715));
  AOI221xp5_ASAP7_75t_L     g21459(.A1(new_n8175), .A2(\b[53] ), .B1(new_n8484), .B2(\b[51] ), .C(new_n21715), .Y(new_n21716));
  O2A1O1Ixp33_ASAP7_75t_L   g21460(.A1(new_n8176), .A2(new_n9691), .B(new_n21716), .C(new_n8172), .Y(new_n21717));
  INVx1_ASAP7_75t_L         g21461(.A(new_n21717), .Y(new_n21718));
  O2A1O1Ixp33_ASAP7_75t_L   g21462(.A1(new_n8176), .A2(new_n9691), .B(new_n21716), .C(\a[50] ), .Y(new_n21719));
  O2A1O1Ixp33_ASAP7_75t_L   g21463(.A1(new_n21548), .A2(new_n21549), .B(new_n21562), .C(new_n21713), .Y(new_n21720));
  INVx1_ASAP7_75t_L         g21464(.A(new_n21720), .Y(new_n21721));
  NAND2xp33_ASAP7_75t_L     g21465(.A(new_n21654), .B(new_n21713), .Y(new_n21722));
  NAND2xp33_ASAP7_75t_L     g21466(.A(new_n21722), .B(new_n21721), .Y(new_n21723));
  A2O1A1Ixp33_ASAP7_75t_L   g21467(.A1(new_n21718), .A2(\a[50] ), .B(new_n21719), .C(new_n21723), .Y(new_n21724));
  AOI21xp33_ASAP7_75t_L     g21468(.A1(new_n21718), .A2(\a[50] ), .B(new_n21719), .Y(new_n21725));
  NAND2xp33_ASAP7_75t_L     g21469(.A(new_n21725), .B(new_n21722), .Y(new_n21726));
  A2O1A1Ixp33_ASAP7_75t_L   g21470(.A1(new_n21655), .A2(new_n21714), .B(new_n21726), .C(new_n21724), .Y(new_n21727));
  O2A1O1Ixp33_ASAP7_75t_L   g21471(.A1(new_n21565), .A2(new_n21653), .B(new_n21574), .C(new_n21727), .Y(new_n21728));
  A2O1A1Ixp33_ASAP7_75t_L   g21472(.A1(new_n21407), .A2(new_n21401), .B(new_n21565), .C(new_n21574), .Y(new_n21729));
  O2A1O1Ixp33_ASAP7_75t_L   g21473(.A1(new_n21726), .A2(new_n21720), .B(new_n21724), .C(new_n21729), .Y(new_n21730));
  NOR2xp33_ASAP7_75t_L      g21474(.A(new_n21730), .B(new_n21728), .Y(new_n21731));
  XOR2x2_ASAP7_75t_L        g21475(.A(new_n21652), .B(new_n21731), .Y(new_n21732));
  INVx1_ASAP7_75t_L         g21476(.A(new_n21732), .Y(new_n21733));
  O2A1O1Ixp33_ASAP7_75t_L   g21477(.A1(new_n21577), .A2(new_n21585), .B(new_n21584), .C(new_n21733), .Y(new_n21734));
  INVx1_ASAP7_75t_L         g21478(.A(new_n21734), .Y(new_n21735));
  INVx1_ASAP7_75t_L         g21479(.A(new_n21581), .Y(new_n21736));
  A2O1A1O1Ixp25_ASAP7_75t_L g21480(.A1(new_n21495), .A2(\a[47] ), .B(new_n21496), .C(new_n21736), .D(new_n21578), .Y(new_n21737));
  NAND2xp33_ASAP7_75t_L     g21481(.A(new_n21733), .B(new_n21737), .Y(new_n21738));
  AND2x2_ASAP7_75t_L        g21482(.A(new_n21738), .B(new_n21735), .Y(new_n21739));
  INVx1_ASAP7_75t_L         g21483(.A(new_n21739), .Y(new_n21740));
  NOR2xp33_ASAP7_75t_L      g21484(.A(new_n10978), .B(new_n6741), .Y(new_n21741));
  AOI221xp5_ASAP7_75t_L     g21485(.A1(\b[59] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[58] ), .C(new_n21741), .Y(new_n21742));
  O2A1O1Ixp33_ASAP7_75t_L   g21486(.A1(new_n6443), .A2(new_n11597), .B(new_n21742), .C(new_n6439), .Y(new_n21743));
  O2A1O1Ixp33_ASAP7_75t_L   g21487(.A1(new_n6443), .A2(new_n11597), .B(new_n21742), .C(\a[44] ), .Y(new_n21744));
  INVx1_ASAP7_75t_L         g21488(.A(new_n21744), .Y(new_n21745));
  O2A1O1Ixp33_ASAP7_75t_L   g21489(.A1(new_n21743), .A2(new_n6439), .B(new_n21745), .C(new_n21740), .Y(new_n21746));
  INVx1_ASAP7_75t_L         g21490(.A(new_n21746), .Y(new_n21747));
  O2A1O1Ixp33_ASAP7_75t_L   g21491(.A1(new_n21743), .A2(new_n6439), .B(new_n21745), .C(new_n21739), .Y(new_n21748));
  AOI21xp33_ASAP7_75t_L     g21492(.A1(new_n21747), .A2(new_n21739), .B(new_n21748), .Y(new_n21749));
  INVx1_ASAP7_75t_L         g21493(.A(new_n21598), .Y(new_n21750));
  A2O1A1O1Ixp25_ASAP7_75t_L g21494(.A1(new_n21750), .A2(\a[44] ), .B(new_n21599), .C(new_n21590), .D(new_n21592), .Y(new_n21751));
  NAND2xp33_ASAP7_75t_L     g21495(.A(new_n21751), .B(new_n21749), .Y(new_n21752));
  INVx1_ASAP7_75t_L         g21496(.A(new_n21751), .Y(new_n21753));
  A2O1A1Ixp33_ASAP7_75t_L   g21497(.A1(new_n21747), .A2(new_n21739), .B(new_n21748), .C(new_n21753), .Y(new_n21754));
  AND2x2_ASAP7_75t_L        g21498(.A(new_n21754), .B(new_n21752), .Y(new_n21755));
  INVx1_ASAP7_75t_L         g21499(.A(new_n21755), .Y(new_n21756));
  NOR2xp33_ASAP7_75t_L      g21500(.A(new_n12603), .B(new_n5641), .Y(new_n21757));
  AOI221xp5_ASAP7_75t_L     g21501(.A1(\b[60] ), .A2(new_n5920), .B1(\b[61] ), .B2(new_n5623), .C(new_n21757), .Y(new_n21758));
  O2A1O1Ixp33_ASAP7_75t_L   g21502(.A1(new_n5630), .A2(new_n12610), .B(new_n21758), .C(new_n5626), .Y(new_n21759));
  O2A1O1Ixp33_ASAP7_75t_L   g21503(.A1(new_n5630), .A2(new_n12610), .B(new_n21758), .C(\a[41] ), .Y(new_n21760));
  INVx1_ASAP7_75t_L         g21504(.A(new_n21760), .Y(new_n21761));
  O2A1O1Ixp33_ASAP7_75t_L   g21505(.A1(new_n21759), .A2(new_n5626), .B(new_n21761), .C(new_n21756), .Y(new_n21762));
  INVx1_ASAP7_75t_L         g21506(.A(new_n21762), .Y(new_n21763));
  O2A1O1Ixp33_ASAP7_75t_L   g21507(.A1(new_n21759), .A2(new_n5626), .B(new_n21761), .C(new_n21755), .Y(new_n21764));
  AOI21xp33_ASAP7_75t_L     g21508(.A1(new_n21763), .A2(new_n21755), .B(new_n21764), .Y(new_n21765));
  A2O1A1Ixp33_ASAP7_75t_L   g21509(.A1(new_n21645), .A2(new_n21639), .B(new_n21646), .C(new_n21765), .Y(new_n21766));
  A2O1A1O1Ixp25_ASAP7_75t_L g21510(.A1(new_n12603), .A2(new_n14444), .B(new_n4911), .C(new_n5144), .D(new_n12956), .Y(new_n21767));
  A2O1A1O1Ixp25_ASAP7_75t_L g21511(.A1(new_n4912), .A2(new_n14172), .B(new_n5139), .C(\b[63] ), .D(new_n4906), .Y(new_n21768));
  A2O1A1O1Ixp25_ASAP7_75t_L g21512(.A1(new_n21605), .A2(new_n21603), .B(new_n21606), .C(new_n21616), .D(new_n21644), .Y(new_n21769));
  A2O1A1O1Ixp25_ASAP7_75t_L g21513(.A1(new_n21641), .A2(new_n21767), .B(new_n21768), .C(new_n21645), .D(new_n21769), .Y(new_n21770));
  A2O1A1Ixp33_ASAP7_75t_L   g21514(.A1(new_n21755), .A2(new_n21763), .B(new_n21764), .C(new_n21770), .Y(new_n21771));
  AND2x2_ASAP7_75t_L        g21515(.A(new_n21766), .B(new_n21771), .Y(new_n21772));
  A2O1A1O1Ixp25_ASAP7_75t_L g21516(.A1(new_n21455), .A2(new_n21449), .B(new_n21489), .C(new_n21637), .D(new_n21772), .Y(new_n21773));
  AND3x1_ASAP7_75t_L        g21517(.A(new_n21772), .B(new_n21637), .C(new_n21488), .Y(new_n21774));
  NOR2xp33_ASAP7_75t_L      g21518(.A(new_n21773), .B(new_n21774), .Y(new_n21775));
  XOR2x2_ASAP7_75t_L        g21519(.A(new_n21775), .B(new_n21635), .Y(\f[101] ));
  NOR2xp33_ASAP7_75t_L      g21520(.A(new_n9683), .B(new_n10065), .Y(new_n21777));
  AOI221xp5_ASAP7_75t_L     g21521(.A1(new_n8175), .A2(\b[54] ), .B1(new_n8484), .B2(\b[52] ), .C(new_n21777), .Y(new_n21778));
  O2A1O1Ixp33_ASAP7_75t_L   g21522(.A1(new_n8176), .A2(new_n9718), .B(new_n21778), .C(new_n8172), .Y(new_n21779));
  INVx1_ASAP7_75t_L         g21523(.A(new_n21779), .Y(new_n21780));
  O2A1O1Ixp33_ASAP7_75t_L   g21524(.A1(new_n8176), .A2(new_n9718), .B(new_n21778), .C(\a[50] ), .Y(new_n21781));
  NOR2xp33_ASAP7_75t_L      g21525(.A(new_n7552), .B(new_n10388), .Y(new_n21782));
  AOI221xp5_ASAP7_75t_L     g21526(.A1(new_n10086), .A2(\b[48] ), .B1(new_n11361), .B2(\b[46] ), .C(new_n21782), .Y(new_n21783));
  INVx1_ASAP7_75t_L         g21527(.A(new_n21783), .Y(new_n21784));
  A2O1A1Ixp33_ASAP7_75t_L   g21528(.A1(new_n11656), .A2(new_n10386), .B(new_n21784), .C(\a[56] ), .Y(new_n21785));
  O2A1O1Ixp33_ASAP7_75t_L   g21529(.A1(new_n10088), .A2(new_n7868), .B(new_n21783), .C(\a[56] ), .Y(new_n21786));
  INVx1_ASAP7_75t_L         g21530(.A(new_n21689), .Y(new_n21787));
  A2O1A1Ixp33_ASAP7_75t_L   g21531(.A1(\a[59] ), .A2(new_n21683), .B(new_n21684), .C(new_n21787), .Y(new_n21788));
  O2A1O1Ixp33_ASAP7_75t_L   g21532(.A1(new_n12669), .A2(new_n12671), .B(\b[38] ), .C(new_n21662), .Y(new_n21789));
  NOR2xp33_ASAP7_75t_L      g21533(.A(new_n5311), .B(new_n13030), .Y(new_n21790));
  INVx1_ASAP7_75t_L         g21534(.A(new_n21790), .Y(new_n21791));
  A2O1A1Ixp33_ASAP7_75t_L   g21535(.A1(new_n13028), .A2(\b[37] ), .B(new_n21502), .C(\a[38] ), .Y(new_n21792));
  NOR2xp33_ASAP7_75t_L      g21536(.A(\a[38] ), .B(new_n21504), .Y(new_n21793));
  INVx1_ASAP7_75t_L         g21537(.A(new_n21793), .Y(new_n21794));
  AND2x2_ASAP7_75t_L        g21538(.A(new_n21792), .B(new_n21794), .Y(new_n21795));
  O2A1O1Ixp33_ASAP7_75t_L   g21539(.A1(new_n5570), .A2(new_n12672), .B(new_n21791), .C(new_n21795), .Y(new_n21796));
  INVx1_ASAP7_75t_L         g21540(.A(new_n21796), .Y(new_n21797));
  O2A1O1Ixp33_ASAP7_75t_L   g21541(.A1(new_n12669), .A2(new_n12671), .B(\b[39] ), .C(new_n21790), .Y(new_n21798));
  NAND2xp33_ASAP7_75t_L     g21542(.A(new_n21798), .B(new_n21795), .Y(new_n21799));
  AND2x2_ASAP7_75t_L        g21543(.A(new_n21799), .B(new_n21797), .Y(new_n21800));
  INVx1_ASAP7_75t_L         g21544(.A(new_n21800), .Y(new_n21801));
  O2A1O1Ixp33_ASAP7_75t_L   g21545(.A1(new_n21504), .A2(new_n21789), .B(new_n21668), .C(new_n21801), .Y(new_n21802));
  NOR3xp33_ASAP7_75t_L      g21546(.A(new_n21667), .B(new_n21800), .C(new_n21664), .Y(new_n21803));
  NOR2xp33_ASAP7_75t_L      g21547(.A(new_n21803), .B(new_n21802), .Y(new_n21804));
  NAND2xp33_ASAP7_75t_L     g21548(.A(\b[42] ), .B(new_n11995), .Y(new_n21805));
  OAI221xp5_ASAP7_75t_L     g21549(.A1(new_n12318), .A2(new_n6110), .B1(new_n5855), .B2(new_n12320), .C(new_n21805), .Y(new_n21806));
  A2O1A1Ixp33_ASAP7_75t_L   g21550(.A1(new_n6389), .A2(new_n11997), .B(new_n21806), .C(\a[62] ), .Y(new_n21807));
  NAND2xp33_ASAP7_75t_L     g21551(.A(\a[62] ), .B(new_n21807), .Y(new_n21808));
  A2O1A1Ixp33_ASAP7_75t_L   g21552(.A1(new_n6389), .A2(new_n11997), .B(new_n21806), .C(new_n11987), .Y(new_n21809));
  NAND2xp33_ASAP7_75t_L     g21553(.A(new_n21809), .B(new_n21808), .Y(new_n21810));
  NAND2xp33_ASAP7_75t_L     g21554(.A(new_n21810), .B(new_n21804), .Y(new_n21811));
  NAND2xp33_ASAP7_75t_L     g21555(.A(new_n21804), .B(new_n21811), .Y(new_n21812));
  NAND2xp33_ASAP7_75t_L     g21556(.A(new_n21810), .B(new_n21811), .Y(new_n21813));
  AND2x2_ASAP7_75t_L        g21557(.A(new_n21812), .B(new_n21813), .Y(new_n21814));
  NOR2xp33_ASAP7_75t_L      g21558(.A(new_n6671), .B(new_n11354), .Y(new_n21815));
  AOI221xp5_ASAP7_75t_L     g21559(.A1(\b[45] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[44] ), .C(new_n21815), .Y(new_n21816));
  O2A1O1Ixp33_ASAP7_75t_L   g21560(.A1(new_n11053), .A2(new_n7255), .B(new_n21816), .C(new_n11048), .Y(new_n21817));
  O2A1O1Ixp33_ASAP7_75t_L   g21561(.A1(new_n11053), .A2(new_n7255), .B(new_n21816), .C(\a[59] ), .Y(new_n21818));
  INVx1_ASAP7_75t_L         g21562(.A(new_n21818), .Y(new_n21819));
  O2A1O1Ixp33_ASAP7_75t_L   g21563(.A1(new_n21817), .A2(new_n11048), .B(new_n21819), .C(new_n21814), .Y(new_n21820));
  INVx1_ASAP7_75t_L         g21564(.A(new_n21814), .Y(new_n21821));
  O2A1O1Ixp33_ASAP7_75t_L   g21565(.A1(new_n21817), .A2(new_n11048), .B(new_n21819), .C(new_n21821), .Y(new_n21822));
  INVx1_ASAP7_75t_L         g21566(.A(new_n21822), .Y(new_n21823));
  A2O1A1O1Ixp25_ASAP7_75t_L g21567(.A1(new_n21683), .A2(\a[59] ), .B(new_n21684), .C(new_n21787), .D(new_n21677), .Y(new_n21824));
  O2A1O1Ixp33_ASAP7_75t_L   g21568(.A1(new_n21814), .A2(new_n21820), .B(new_n21823), .C(new_n21824), .Y(new_n21825));
  O2A1O1Ixp33_ASAP7_75t_L   g21569(.A1(new_n21814), .A2(new_n21820), .B(new_n21823), .C(new_n21825), .Y(new_n21826));
  INVx1_ASAP7_75t_L         g21570(.A(new_n21826), .Y(new_n21827));
  A2O1A1Ixp33_ASAP7_75t_L   g21571(.A1(new_n21788), .A2(new_n21678), .B(new_n21825), .C(new_n21827), .Y(new_n21828));
  A2O1A1Ixp33_ASAP7_75t_L   g21572(.A1(\a[56] ), .A2(new_n21785), .B(new_n21786), .C(new_n21828), .Y(new_n21829));
  AO21x2_ASAP7_75t_L        g21573(.A1(\a[56] ), .A2(new_n21785), .B(new_n21786), .Y(new_n21830));
  O2A1O1Ixp33_ASAP7_75t_L   g21574(.A1(new_n21824), .A2(new_n21825), .B(new_n21827), .C(new_n21830), .Y(new_n21831));
  A2O1A1O1Ixp25_ASAP7_75t_L g21575(.A1(new_n21785), .A2(\a[56] ), .B(new_n21786), .C(new_n21829), .D(new_n21831), .Y(new_n21832));
  A2O1A1O1Ixp25_ASAP7_75t_L g21576(.A1(new_n21659), .A2(\a[56] ), .B(new_n21660), .C(new_n21693), .D(new_n21694), .Y(new_n21833));
  XOR2x2_ASAP7_75t_L        g21577(.A(new_n21833), .B(new_n21832), .Y(new_n21834));
  INVx1_ASAP7_75t_L         g21578(.A(new_n21834), .Y(new_n21835));
  NOR2xp33_ASAP7_75t_L      g21579(.A(new_n8755), .B(new_n10400), .Y(new_n21836));
  AOI221xp5_ASAP7_75t_L     g21580(.A1(new_n9102), .A2(\b[51] ), .B1(new_n10398), .B2(\b[49] ), .C(new_n21836), .Y(new_n21837));
  O2A1O1Ixp33_ASAP7_75t_L   g21581(.A1(new_n9104), .A2(new_n8789), .B(new_n21837), .C(new_n9099), .Y(new_n21838));
  O2A1O1Ixp33_ASAP7_75t_L   g21582(.A1(new_n9104), .A2(new_n8789), .B(new_n21837), .C(\a[53] ), .Y(new_n21839));
  INVx1_ASAP7_75t_L         g21583(.A(new_n21839), .Y(new_n21840));
  OAI211xp5_ASAP7_75t_L     g21584(.A1(new_n9099), .A2(new_n21838), .B(new_n21835), .C(new_n21840), .Y(new_n21841));
  O2A1O1Ixp33_ASAP7_75t_L   g21585(.A1(new_n21838), .A2(new_n9099), .B(new_n21840), .C(new_n21835), .Y(new_n21842));
  INVx1_ASAP7_75t_L         g21586(.A(new_n21842), .Y(new_n21843));
  AND2x2_ASAP7_75t_L        g21587(.A(new_n21841), .B(new_n21843), .Y(new_n21844));
  INVx1_ASAP7_75t_L         g21588(.A(new_n21844), .Y(new_n21845));
  O2A1O1Ixp33_ASAP7_75t_L   g21589(.A1(new_n21699), .A2(new_n21700), .B(new_n21711), .C(new_n21845), .Y(new_n21846));
  INVx1_ASAP7_75t_L         g21590(.A(new_n21846), .Y(new_n21847));
  A2O1A1O1Ixp25_ASAP7_75t_L g21591(.A1(new_n21708), .A2(\a[53] ), .B(new_n21709), .C(new_n21701), .D(new_n21702), .Y(new_n21848));
  NAND2xp33_ASAP7_75t_L     g21592(.A(new_n21848), .B(new_n21845), .Y(new_n21849));
  AND2x2_ASAP7_75t_L        g21593(.A(new_n21849), .B(new_n21847), .Y(new_n21850));
  A2O1A1Ixp33_ASAP7_75t_L   g21594(.A1(new_n21780), .A2(\a[50] ), .B(new_n21781), .C(new_n21850), .Y(new_n21851));
  NOR2xp33_ASAP7_75t_L      g21595(.A(new_n8172), .B(new_n21779), .Y(new_n21852));
  OR3x1_ASAP7_75t_L         g21596(.A(new_n21850), .B(new_n21852), .C(new_n21781), .Y(new_n21853));
  AND2x2_ASAP7_75t_L        g21597(.A(new_n21851), .B(new_n21853), .Y(new_n21854));
  INVx1_ASAP7_75t_L         g21598(.A(new_n21854), .Y(new_n21855));
  A2O1A1O1Ixp25_ASAP7_75t_L g21599(.A1(new_n21721), .A2(new_n21722), .B(new_n21725), .C(new_n21714), .D(new_n21855), .Y(new_n21856));
  INVx1_ASAP7_75t_L         g21600(.A(new_n21856), .Y(new_n21857));
  NAND3xp33_ASAP7_75t_L     g21601(.A(new_n21855), .B(new_n21724), .C(new_n21714), .Y(new_n21858));
  NAND2xp33_ASAP7_75t_L     g21602(.A(new_n21858), .B(new_n21857), .Y(new_n21859));
  INVx1_ASAP7_75t_L         g21603(.A(new_n21859), .Y(new_n21860));
  NOR2xp33_ASAP7_75t_L      g21604(.A(new_n10332), .B(new_n7312), .Y(new_n21861));
  AOI221xp5_ASAP7_75t_L     g21605(.A1(\b[55] ), .A2(new_n7609), .B1(\b[57] ), .B2(new_n7334), .C(new_n21861), .Y(new_n21862));
  O2A1O1Ixp33_ASAP7_75t_L   g21606(.A1(new_n7321), .A2(new_n17096), .B(new_n21862), .C(new_n7316), .Y(new_n21863));
  O2A1O1Ixp33_ASAP7_75t_L   g21607(.A1(new_n7321), .A2(new_n17096), .B(new_n21862), .C(\a[47] ), .Y(new_n21864));
  INVx1_ASAP7_75t_L         g21608(.A(new_n21864), .Y(new_n21865));
  O2A1O1Ixp33_ASAP7_75t_L   g21609(.A1(new_n21863), .A2(new_n7316), .B(new_n21865), .C(new_n21859), .Y(new_n21866));
  INVx1_ASAP7_75t_L         g21610(.A(new_n21866), .Y(new_n21867));
  O2A1O1Ixp33_ASAP7_75t_L   g21611(.A1(new_n21863), .A2(new_n7316), .B(new_n21865), .C(new_n21860), .Y(new_n21868));
  AOI21xp33_ASAP7_75t_L     g21612(.A1(new_n21867), .A2(new_n21860), .B(new_n21868), .Y(new_n21869));
  A2O1A1O1Ixp25_ASAP7_75t_L g21613(.A1(new_n21650), .A2(\a[47] ), .B(new_n21651), .C(new_n21731), .D(new_n21728), .Y(new_n21870));
  NAND2xp33_ASAP7_75t_L     g21614(.A(new_n21870), .B(new_n21869), .Y(new_n21871));
  INVx1_ASAP7_75t_L         g21615(.A(new_n21870), .Y(new_n21872));
  A2O1A1Ixp33_ASAP7_75t_L   g21616(.A1(new_n21867), .A2(new_n21860), .B(new_n21868), .C(new_n21872), .Y(new_n21873));
  AND2x2_ASAP7_75t_L        g21617(.A(new_n21873), .B(new_n21871), .Y(new_n21874));
  INVx1_ASAP7_75t_L         g21618(.A(new_n21874), .Y(new_n21875));
  NOR2xp33_ASAP7_75t_L      g21619(.A(new_n11303), .B(new_n6741), .Y(new_n21876));
  AOI221xp5_ASAP7_75t_L     g21620(.A1(\b[60] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[59] ), .C(new_n21876), .Y(new_n21877));
  O2A1O1Ixp33_ASAP7_75t_L   g21621(.A1(new_n6443), .A2(new_n11634), .B(new_n21877), .C(new_n6439), .Y(new_n21878));
  O2A1O1Ixp33_ASAP7_75t_L   g21622(.A1(new_n6443), .A2(new_n11634), .B(new_n21877), .C(\a[44] ), .Y(new_n21879));
  INVx1_ASAP7_75t_L         g21623(.A(new_n21879), .Y(new_n21880));
  O2A1O1Ixp33_ASAP7_75t_L   g21624(.A1(new_n21878), .A2(new_n6439), .B(new_n21880), .C(new_n21875), .Y(new_n21881));
  INVx1_ASAP7_75t_L         g21625(.A(new_n21881), .Y(new_n21882));
  O2A1O1Ixp33_ASAP7_75t_L   g21626(.A1(new_n21878), .A2(new_n6439), .B(new_n21880), .C(new_n21874), .Y(new_n21883));
  AOI21xp33_ASAP7_75t_L     g21627(.A1(new_n21882), .A2(new_n21874), .B(new_n21883), .Y(new_n21884));
  O2A1O1Ixp33_ASAP7_75t_L   g21628(.A1(new_n21578), .A2(new_n21583), .B(new_n21732), .C(new_n21746), .Y(new_n21885));
  NAND2xp33_ASAP7_75t_L     g21629(.A(new_n21885), .B(new_n21884), .Y(new_n21886));
  O2A1O1Ixp33_ASAP7_75t_L   g21630(.A1(new_n21737), .A2(new_n21733), .B(new_n21747), .C(new_n21884), .Y(new_n21887));
  INVx1_ASAP7_75t_L         g21631(.A(new_n21887), .Y(new_n21888));
  AND2x2_ASAP7_75t_L        g21632(.A(new_n21886), .B(new_n21888), .Y(new_n21889));
  INVx1_ASAP7_75t_L         g21633(.A(new_n21889), .Y(new_n21890));
  NOR2xp33_ASAP7_75t_L      g21634(.A(new_n12956), .B(new_n5641), .Y(new_n21891));
  AOI221xp5_ASAP7_75t_L     g21635(.A1(\b[61] ), .A2(new_n5920), .B1(\b[62] ), .B2(new_n5623), .C(new_n21891), .Y(new_n21892));
  O2A1O1Ixp33_ASAP7_75t_L   g21636(.A1(new_n5630), .A2(new_n17815), .B(new_n21892), .C(new_n5626), .Y(new_n21893));
  O2A1O1Ixp33_ASAP7_75t_L   g21637(.A1(new_n5630), .A2(new_n17815), .B(new_n21892), .C(\a[41] ), .Y(new_n21894));
  INVx1_ASAP7_75t_L         g21638(.A(new_n21894), .Y(new_n21895));
  O2A1O1Ixp33_ASAP7_75t_L   g21639(.A1(new_n21893), .A2(new_n5626), .B(new_n21895), .C(new_n21890), .Y(new_n21896));
  INVx1_ASAP7_75t_L         g21640(.A(new_n21896), .Y(new_n21897));
  O2A1O1Ixp33_ASAP7_75t_L   g21641(.A1(new_n21893), .A2(new_n5626), .B(new_n21895), .C(new_n21889), .Y(new_n21898));
  AOI21xp33_ASAP7_75t_L     g21642(.A1(new_n21897), .A2(new_n21889), .B(new_n21898), .Y(new_n21899));
  A2O1A1O1Ixp25_ASAP7_75t_L g21643(.A1(new_n21747), .A2(new_n21739), .B(new_n21748), .C(new_n21753), .D(new_n21762), .Y(new_n21900));
  NAND2xp33_ASAP7_75t_L     g21644(.A(new_n21900), .B(new_n21899), .Y(new_n21901));
  O2A1O1Ixp33_ASAP7_75t_L   g21645(.A1(new_n21749), .A2(new_n21751), .B(new_n21763), .C(new_n21899), .Y(new_n21902));
  INVx1_ASAP7_75t_L         g21646(.A(new_n21902), .Y(new_n21903));
  AND2x2_ASAP7_75t_L        g21647(.A(new_n21901), .B(new_n21903), .Y(new_n21904));
  INVx1_ASAP7_75t_L         g21648(.A(new_n21904), .Y(new_n21905));
  O2A1O1Ixp33_ASAP7_75t_L   g21649(.A1(new_n21770), .A2(new_n21765), .B(new_n21645), .C(new_n21905), .Y(new_n21906));
  INVx1_ASAP7_75t_L         g21650(.A(new_n21646), .Y(new_n21907));
  O2A1O1Ixp33_ASAP7_75t_L   g21651(.A1(new_n21638), .A2(new_n21644), .B(new_n21907), .C(new_n21765), .Y(new_n21908));
  NOR3xp33_ASAP7_75t_L      g21652(.A(new_n21904), .B(new_n21908), .C(new_n21644), .Y(new_n21909));
  NOR2xp33_ASAP7_75t_L      g21653(.A(new_n21909), .B(new_n21906), .Y(new_n21910));
  A2O1A1Ixp33_ASAP7_75t_L   g21654(.A1(new_n21635), .A2(new_n21775), .B(new_n21773), .C(new_n21910), .Y(new_n21911));
  INVx1_ASAP7_75t_L         g21655(.A(new_n21911), .Y(new_n21912));
  A2O1A1Ixp33_ASAP7_75t_L   g21656(.A1(new_n21631), .A2(new_n21628), .B(new_n21626), .C(new_n21775), .Y(new_n21913));
  A2O1A1Ixp33_ASAP7_75t_L   g21657(.A1(new_n21637), .A2(new_n21488), .B(new_n21772), .C(new_n21913), .Y(new_n21914));
  NOR2xp33_ASAP7_75t_L      g21658(.A(new_n21910), .B(new_n21914), .Y(new_n21915));
  NOR2xp33_ASAP7_75t_L      g21659(.A(new_n21912), .B(new_n21915), .Y(\f[102] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21660(.A1(new_n21641), .A2(new_n21767), .B(new_n21768), .C(new_n21639), .D(new_n21908), .Y(new_n21917));
  A2O1A1Ixp33_ASAP7_75t_L   g21661(.A1(new_n21735), .A2(new_n21747), .B(new_n21884), .C(new_n21882), .Y(new_n21918));
  AOI22xp33_ASAP7_75t_L     g21662(.A1(new_n5623), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5920), .Y(new_n21919));
  INVx1_ASAP7_75t_L         g21663(.A(new_n21919), .Y(new_n21920));
  A2O1A1Ixp33_ASAP7_75t_L   g21664(.A1(new_n5625), .A2(new_n5627), .B(new_n5348), .C(new_n21919), .Y(new_n21921));
  O2A1O1Ixp33_ASAP7_75t_L   g21665(.A1(new_n21920), .A2(new_n17329), .B(new_n21921), .C(new_n5626), .Y(new_n21922));
  O2A1O1Ixp33_ASAP7_75t_L   g21666(.A1(new_n5630), .A2(new_n12993), .B(new_n21919), .C(\a[41] ), .Y(new_n21923));
  OAI21xp33_ASAP7_75t_L     g21667(.A1(new_n21922), .A2(new_n21923), .B(new_n21918), .Y(new_n21924));
  NOR2xp33_ASAP7_75t_L      g21668(.A(new_n21923), .B(new_n21922), .Y(new_n21925));
  NAND3xp33_ASAP7_75t_L     g21669(.A(new_n21888), .B(new_n21882), .C(new_n21925), .Y(new_n21926));
  NAND2xp33_ASAP7_75t_L     g21670(.A(new_n21924), .B(new_n21926), .Y(new_n21927));
  INVx1_ASAP7_75t_L         g21671(.A(new_n21927), .Y(new_n21928));
  NOR2xp33_ASAP7_75t_L      g21672(.A(new_n7860), .B(new_n10388), .Y(new_n21929));
  AOI221xp5_ASAP7_75t_L     g21673(.A1(new_n10086), .A2(\b[49] ), .B1(new_n11361), .B2(\b[47] ), .C(new_n21929), .Y(new_n21930));
  O2A1O1Ixp33_ASAP7_75t_L   g21674(.A1(new_n10088), .A2(new_n14802), .B(new_n21930), .C(new_n10083), .Y(new_n21931));
  INVx1_ASAP7_75t_L         g21675(.A(new_n21931), .Y(new_n21932));
  O2A1O1Ixp33_ASAP7_75t_L   g21676(.A1(new_n10088), .A2(new_n14802), .B(new_n21930), .C(\a[56] ), .Y(new_n21933));
  INVx1_ASAP7_75t_L         g21677(.A(new_n21802), .Y(new_n21934));
  NOR2xp33_ASAP7_75t_L      g21678(.A(new_n5570), .B(new_n13030), .Y(new_n21935));
  O2A1O1Ixp33_ASAP7_75t_L   g21679(.A1(new_n12669), .A2(new_n12671), .B(\b[40] ), .C(new_n21935), .Y(new_n21936));
  A2O1A1Ixp33_ASAP7_75t_L   g21680(.A1(new_n21504), .A2(new_n4906), .B(new_n21796), .C(new_n21936), .Y(new_n21937));
  A2O1A1O1Ixp25_ASAP7_75t_L g21681(.A1(new_n13028), .A2(\b[37] ), .B(new_n21502), .C(new_n4906), .D(new_n21796), .Y(new_n21938));
  A2O1A1Ixp33_ASAP7_75t_L   g21682(.A1(new_n13028), .A2(\b[40] ), .B(new_n21935), .C(new_n21938), .Y(new_n21939));
  NAND2xp33_ASAP7_75t_L     g21683(.A(new_n21937), .B(new_n21939), .Y(new_n21940));
  NAND2xp33_ASAP7_75t_L     g21684(.A(\b[43] ), .B(new_n11995), .Y(new_n21941));
  OAI221xp5_ASAP7_75t_L     g21685(.A1(new_n12318), .A2(new_n6378), .B1(new_n6110), .B2(new_n12320), .C(new_n21941), .Y(new_n21942));
  AOI21xp33_ASAP7_75t_L     g21686(.A1(new_n6682), .A2(new_n11997), .B(new_n21942), .Y(new_n21943));
  NAND2xp33_ASAP7_75t_L     g21687(.A(\a[62] ), .B(new_n21943), .Y(new_n21944));
  A2O1A1Ixp33_ASAP7_75t_L   g21688(.A1(new_n6682), .A2(new_n11997), .B(new_n21942), .C(new_n11987), .Y(new_n21945));
  AOI21xp33_ASAP7_75t_L     g21689(.A1(new_n21944), .A2(new_n21945), .B(new_n21940), .Y(new_n21946));
  AND3x1_ASAP7_75t_L        g21690(.A(new_n21944), .B(new_n21945), .C(new_n21940), .Y(new_n21947));
  NOR2xp33_ASAP7_75t_L      g21691(.A(new_n21946), .B(new_n21947), .Y(new_n21948));
  INVx1_ASAP7_75t_L         g21692(.A(new_n21948), .Y(new_n21949));
  A2O1A1O1Ixp25_ASAP7_75t_L g21693(.A1(new_n21809), .A2(new_n21808), .B(new_n21803), .C(new_n21934), .D(new_n21949), .Y(new_n21950));
  INVx1_ASAP7_75t_L         g21694(.A(new_n21950), .Y(new_n21951));
  NAND3xp33_ASAP7_75t_L     g21695(.A(new_n21811), .B(new_n21934), .C(new_n21949), .Y(new_n21952));
  AND2x2_ASAP7_75t_L        g21696(.A(new_n21952), .B(new_n21951), .Y(new_n21953));
  INVx1_ASAP7_75t_L         g21697(.A(new_n21953), .Y(new_n21954));
  NOR2xp33_ASAP7_75t_L      g21698(.A(new_n6944), .B(new_n11354), .Y(new_n21955));
  AOI221xp5_ASAP7_75t_L     g21699(.A1(\b[46] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[45] ), .C(new_n21955), .Y(new_n21956));
  O2A1O1Ixp33_ASAP7_75t_L   g21700(.A1(new_n11053), .A2(new_n7279), .B(new_n21956), .C(new_n11048), .Y(new_n21957));
  O2A1O1Ixp33_ASAP7_75t_L   g21701(.A1(new_n11053), .A2(new_n7279), .B(new_n21956), .C(\a[59] ), .Y(new_n21958));
  INVx1_ASAP7_75t_L         g21702(.A(new_n21958), .Y(new_n21959));
  O2A1O1Ixp33_ASAP7_75t_L   g21703(.A1(new_n21957), .A2(new_n11048), .B(new_n21959), .C(new_n21954), .Y(new_n21960));
  INVx1_ASAP7_75t_L         g21704(.A(new_n21960), .Y(new_n21961));
  O2A1O1Ixp33_ASAP7_75t_L   g21705(.A1(new_n21957), .A2(new_n11048), .B(new_n21959), .C(new_n21953), .Y(new_n21962));
  AO21x2_ASAP7_75t_L        g21706(.A1(new_n21953), .A2(new_n21961), .B(new_n21962), .Y(new_n21963));
  OR3x1_ASAP7_75t_L         g21707(.A(new_n21963), .B(new_n21820), .C(new_n21825), .Y(new_n21964));
  INVx1_ASAP7_75t_L         g21708(.A(new_n21820), .Y(new_n21965));
  A2O1A1Ixp33_ASAP7_75t_L   g21709(.A1(new_n21823), .A2(new_n21814), .B(new_n21824), .C(new_n21965), .Y(new_n21966));
  A2O1A1Ixp33_ASAP7_75t_L   g21710(.A1(new_n21961), .A2(new_n21953), .B(new_n21962), .C(new_n21966), .Y(new_n21967));
  NAND2xp33_ASAP7_75t_L     g21711(.A(new_n21967), .B(new_n21964), .Y(new_n21968));
  INVx1_ASAP7_75t_L         g21712(.A(new_n21968), .Y(new_n21969));
  A2O1A1Ixp33_ASAP7_75t_L   g21713(.A1(\a[56] ), .A2(new_n21932), .B(new_n21933), .C(new_n21969), .Y(new_n21970));
  INVx1_ASAP7_75t_L         g21714(.A(new_n21970), .Y(new_n21971));
  NOR2xp33_ASAP7_75t_L      g21715(.A(new_n21968), .B(new_n21971), .Y(new_n21972));
  A2O1A1O1Ixp25_ASAP7_75t_L g21716(.A1(new_n21932), .A2(\a[56] ), .B(new_n21933), .C(new_n21970), .D(new_n21972), .Y(new_n21973));
  A2O1A1Ixp33_ASAP7_75t_L   g21717(.A1(new_n21813), .A2(new_n21812), .B(new_n21820), .C(new_n21823), .Y(new_n21974));
  O2A1O1Ixp33_ASAP7_75t_L   g21718(.A1(new_n21689), .A2(new_n21685), .B(new_n21678), .C(new_n21974), .Y(new_n21975));
  O2A1O1Ixp33_ASAP7_75t_L   g21719(.A1(new_n21691), .A2(new_n21692), .B(new_n21697), .C(new_n21832), .Y(new_n21976));
  O2A1O1Ixp33_ASAP7_75t_L   g21720(.A1(new_n21826), .A2(new_n21975), .B(new_n21830), .C(new_n21976), .Y(new_n21977));
  NAND2xp33_ASAP7_75t_L     g21721(.A(new_n21977), .B(new_n21973), .Y(new_n21978));
  A2O1A1Ixp33_ASAP7_75t_L   g21722(.A1(\a[56] ), .A2(new_n21932), .B(new_n21933), .C(new_n21968), .Y(new_n21979));
  O2A1O1Ixp33_ASAP7_75t_L   g21723(.A1(new_n21968), .A2(new_n21971), .B(new_n21979), .C(new_n21977), .Y(new_n21980));
  INVx1_ASAP7_75t_L         g21724(.A(new_n21980), .Y(new_n21981));
  AND2x2_ASAP7_75t_L        g21725(.A(new_n21978), .B(new_n21981), .Y(new_n21982));
  NOR2xp33_ASAP7_75t_L      g21726(.A(new_n8779), .B(new_n10400), .Y(new_n21983));
  AOI221xp5_ASAP7_75t_L     g21727(.A1(new_n9102), .A2(\b[52] ), .B1(new_n10398), .B2(\b[50] ), .C(new_n21983), .Y(new_n21984));
  O2A1O1Ixp33_ASAP7_75t_L   g21728(.A1(new_n9104), .A2(new_n17363), .B(new_n21984), .C(new_n9099), .Y(new_n21985));
  INVx1_ASAP7_75t_L         g21729(.A(new_n21985), .Y(new_n21986));
  O2A1O1Ixp33_ASAP7_75t_L   g21730(.A1(new_n9104), .A2(new_n17363), .B(new_n21984), .C(\a[53] ), .Y(new_n21987));
  A2O1A1Ixp33_ASAP7_75t_L   g21731(.A1(\a[53] ), .A2(new_n21986), .B(new_n21987), .C(new_n21982), .Y(new_n21988));
  A2O1A1Ixp33_ASAP7_75t_L   g21732(.A1(new_n21986), .A2(\a[53] ), .B(new_n21987), .C(new_n21988), .Y(new_n21989));
  INVx1_ASAP7_75t_L         g21733(.A(new_n21989), .Y(new_n21990));
  AOI21xp33_ASAP7_75t_L     g21734(.A1(new_n21988), .A2(new_n21982), .B(new_n21990), .Y(new_n21991));
  INVx1_ASAP7_75t_L         g21735(.A(new_n21991), .Y(new_n21992));
  O2A1O1Ixp33_ASAP7_75t_L   g21736(.A1(new_n21848), .A2(new_n21845), .B(new_n21843), .C(new_n21991), .Y(new_n21993));
  INVx1_ASAP7_75t_L         g21737(.A(new_n21993), .Y(new_n21994));
  O2A1O1Ixp33_ASAP7_75t_L   g21738(.A1(new_n21848), .A2(new_n21845), .B(new_n21843), .C(new_n21992), .Y(new_n21995));
  A2O1A1O1Ixp25_ASAP7_75t_L g21739(.A1(new_n21988), .A2(new_n21982), .B(new_n21990), .C(new_n21994), .D(new_n21995), .Y(new_n21996));
  NOR2xp33_ASAP7_75t_L      g21740(.A(new_n9709), .B(new_n10065), .Y(new_n21997));
  AOI221xp5_ASAP7_75t_L     g21741(.A1(new_n8175), .A2(\b[55] ), .B1(new_n8484), .B2(\b[53] ), .C(new_n21997), .Y(new_n21998));
  O2A1O1Ixp33_ASAP7_75t_L   g21742(.A1(new_n8176), .A2(new_n15849), .B(new_n21998), .C(new_n8172), .Y(new_n21999));
  O2A1O1Ixp33_ASAP7_75t_L   g21743(.A1(new_n8176), .A2(new_n15849), .B(new_n21998), .C(\a[50] ), .Y(new_n22000));
  INVx1_ASAP7_75t_L         g21744(.A(new_n22000), .Y(new_n22001));
  O2A1O1Ixp33_ASAP7_75t_L   g21745(.A1(new_n21999), .A2(new_n8172), .B(new_n22001), .C(new_n21996), .Y(new_n22002));
  INVx1_ASAP7_75t_L         g21746(.A(new_n22002), .Y(new_n22003));
  O2A1O1Ixp33_ASAP7_75t_L   g21747(.A1(new_n8172), .A2(new_n21999), .B(new_n22001), .C(new_n22002), .Y(new_n22004));
  A2O1A1O1Ixp25_ASAP7_75t_L g21748(.A1(new_n21994), .A2(new_n21992), .B(new_n21995), .C(new_n22003), .D(new_n22004), .Y(new_n22005));
  O2A1O1Ixp33_ASAP7_75t_L   g21749(.A1(new_n21852), .A2(new_n21781), .B(new_n21850), .C(new_n21856), .Y(new_n22006));
  NAND2xp33_ASAP7_75t_L     g21750(.A(new_n22006), .B(new_n22005), .Y(new_n22007));
  A2O1A1O1Ixp25_ASAP7_75t_L g21751(.A1(new_n21724), .A2(new_n21714), .B(new_n21855), .C(new_n21851), .D(new_n22005), .Y(new_n22008));
  INVx1_ASAP7_75t_L         g21752(.A(new_n22008), .Y(new_n22009));
  AND2x2_ASAP7_75t_L        g21753(.A(new_n22007), .B(new_n22009), .Y(new_n22010));
  INVx1_ASAP7_75t_L         g21754(.A(new_n22010), .Y(new_n22011));
  NOR2xp33_ASAP7_75t_L      g21755(.A(new_n11303), .B(new_n7318), .Y(new_n22012));
  AOI221xp5_ASAP7_75t_L     g21756(.A1(new_n7333), .A2(\b[57] ), .B1(new_n7609), .B2(\b[56] ), .C(new_n22012), .Y(new_n22013));
  O2A1O1Ixp33_ASAP7_75t_L   g21757(.A1(new_n7321), .A2(new_n20073), .B(new_n22013), .C(new_n7316), .Y(new_n22014));
  O2A1O1Ixp33_ASAP7_75t_L   g21758(.A1(new_n7321), .A2(new_n20073), .B(new_n22013), .C(\a[47] ), .Y(new_n22015));
  INVx1_ASAP7_75t_L         g21759(.A(new_n22015), .Y(new_n22016));
  O2A1O1Ixp33_ASAP7_75t_L   g21760(.A1(new_n22014), .A2(new_n7316), .B(new_n22016), .C(new_n22011), .Y(new_n22017));
  INVx1_ASAP7_75t_L         g21761(.A(new_n22017), .Y(new_n22018));
  O2A1O1Ixp33_ASAP7_75t_L   g21762(.A1(new_n22014), .A2(new_n7316), .B(new_n22016), .C(new_n22010), .Y(new_n22019));
  AOI21xp33_ASAP7_75t_L     g21763(.A1(new_n22018), .A2(new_n22010), .B(new_n22019), .Y(new_n22020));
  O2A1O1Ixp33_ASAP7_75t_L   g21764(.A1(new_n21860), .A2(new_n21868), .B(new_n21872), .C(new_n21866), .Y(new_n22021));
  NAND2xp33_ASAP7_75t_L     g21765(.A(new_n22021), .B(new_n22020), .Y(new_n22022));
  O2A1O1Ixp33_ASAP7_75t_L   g21766(.A1(new_n21869), .A2(new_n21870), .B(new_n21867), .C(new_n22020), .Y(new_n22023));
  INVx1_ASAP7_75t_L         g21767(.A(new_n22023), .Y(new_n22024));
  AND2x2_ASAP7_75t_L        g21768(.A(new_n22022), .B(new_n22024), .Y(new_n22025));
  NOR2xp33_ASAP7_75t_L      g21769(.A(new_n11591), .B(new_n6741), .Y(new_n22026));
  AOI221xp5_ASAP7_75t_L     g21770(.A1(\b[61] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[60] ), .C(new_n22026), .Y(new_n22027));
  O2A1O1Ixp33_ASAP7_75t_L   g21771(.A1(new_n6443), .A2(new_n14764), .B(new_n22027), .C(new_n6439), .Y(new_n22028));
  INVx1_ASAP7_75t_L         g21772(.A(new_n22028), .Y(new_n22029));
  O2A1O1Ixp33_ASAP7_75t_L   g21773(.A1(new_n6443), .A2(new_n14764), .B(new_n22027), .C(\a[44] ), .Y(new_n22030));
  A2O1A1Ixp33_ASAP7_75t_L   g21774(.A1(\a[44] ), .A2(new_n22029), .B(new_n22030), .C(new_n22025), .Y(new_n22031));
  NOR2xp33_ASAP7_75t_L      g21775(.A(new_n6439), .B(new_n22028), .Y(new_n22032));
  OR3x1_ASAP7_75t_L         g21776(.A(new_n22025), .B(new_n22032), .C(new_n22030), .Y(new_n22033));
  NAND3xp33_ASAP7_75t_L     g21777(.A(new_n21928), .B(new_n22031), .C(new_n22033), .Y(new_n22034));
  NAND2xp33_ASAP7_75t_L     g21778(.A(new_n21928), .B(new_n22034), .Y(new_n22035));
  NAND3xp33_ASAP7_75t_L     g21779(.A(new_n21927), .B(new_n22031), .C(new_n22033), .Y(new_n22036));
  NAND2xp33_ASAP7_75t_L     g21780(.A(new_n22036), .B(new_n22035), .Y(new_n22037));
  INVx1_ASAP7_75t_L         g21781(.A(new_n22037), .Y(new_n22038));
  NAND3xp33_ASAP7_75t_L     g21782(.A(new_n21903), .B(new_n22038), .C(new_n21897), .Y(new_n22039));
  O2A1O1Ixp33_ASAP7_75t_L   g21783(.A1(new_n21899), .A2(new_n21900), .B(new_n21897), .C(new_n22038), .Y(new_n22040));
  INVx1_ASAP7_75t_L         g21784(.A(new_n22040), .Y(new_n22041));
  AND2x2_ASAP7_75t_L        g21785(.A(new_n22039), .B(new_n22041), .Y(new_n22042));
  INVx1_ASAP7_75t_L         g21786(.A(new_n22042), .Y(new_n22043));
  O2A1O1Ixp33_ASAP7_75t_L   g21787(.A1(new_n21905), .A2(new_n21917), .B(new_n21911), .C(new_n22043), .Y(new_n22044));
  NOR3xp33_ASAP7_75t_L      g21788(.A(new_n21912), .B(new_n22042), .C(new_n21906), .Y(new_n22045));
  NOR2xp33_ASAP7_75t_L      g21789(.A(new_n22044), .B(new_n22045), .Y(\f[103] ));
  INVx1_ASAP7_75t_L         g21790(.A(new_n21906), .Y(new_n22047));
  A2O1A1Ixp33_ASAP7_75t_L   g21791(.A1(new_n21911), .A2(new_n22047), .B(new_n22043), .C(new_n22041), .Y(new_n22048));
  O2A1O1Ixp33_ASAP7_75t_L   g21792(.A1(new_n22032), .A2(new_n22030), .B(new_n22022), .C(new_n22023), .Y(new_n22049));
  INVx1_ASAP7_75t_L         g21793(.A(new_n22049), .Y(new_n22050));
  NOR2xp33_ASAP7_75t_L      g21794(.A(new_n12956), .B(new_n5925), .Y(new_n22051));
  A2O1A1Ixp33_ASAP7_75t_L   g21795(.A1(new_n12986), .A2(new_n5637), .B(new_n22051), .C(\a[41] ), .Y(new_n22052));
  INVx1_ASAP7_75t_L         g21796(.A(new_n22052), .Y(new_n22053));
  A2O1A1Ixp33_ASAP7_75t_L   g21797(.A1(new_n12986), .A2(new_n5637), .B(new_n22051), .C(new_n5626), .Y(new_n22054));
  O2A1O1Ixp33_ASAP7_75t_L   g21798(.A1(new_n22053), .A2(new_n5626), .B(new_n22054), .C(new_n22049), .Y(new_n22055));
  INVx1_ASAP7_75t_L         g21799(.A(new_n22055), .Y(new_n22056));
  O2A1O1Ixp33_ASAP7_75t_L   g21800(.A1(new_n22053), .A2(new_n5626), .B(new_n22054), .C(new_n22050), .Y(new_n22057));
  O2A1O1Ixp33_ASAP7_75t_L   g21801(.A1(new_n21702), .A2(new_n21712), .B(new_n21841), .C(new_n21842), .Y(new_n22058));
  NOR2xp33_ASAP7_75t_L      g21802(.A(new_n10309), .B(new_n10065), .Y(new_n22059));
  AOI221xp5_ASAP7_75t_L     g21803(.A1(new_n8175), .A2(\b[56] ), .B1(new_n8484), .B2(\b[54] ), .C(new_n22059), .Y(new_n22060));
  O2A1O1Ixp33_ASAP7_75t_L   g21804(.A1(new_n8176), .A2(new_n10339), .B(new_n22060), .C(new_n8172), .Y(new_n22061));
  INVx1_ASAP7_75t_L         g21805(.A(new_n22061), .Y(new_n22062));
  O2A1O1Ixp33_ASAP7_75t_L   g21806(.A1(new_n8176), .A2(new_n10339), .B(new_n22060), .C(\a[50] ), .Y(new_n22063));
  NOR2xp33_ASAP7_75t_L      g21807(.A(new_n9355), .B(new_n10400), .Y(new_n22064));
  AOI221xp5_ASAP7_75t_L     g21808(.A1(new_n9102), .A2(\b[53] ), .B1(new_n10398), .B2(\b[51] ), .C(new_n22064), .Y(new_n22065));
  O2A1O1Ixp33_ASAP7_75t_L   g21809(.A1(new_n9104), .A2(new_n9691), .B(new_n22065), .C(new_n9099), .Y(new_n22066));
  INVx1_ASAP7_75t_L         g21810(.A(new_n22066), .Y(new_n22067));
  O2A1O1Ixp33_ASAP7_75t_L   g21811(.A1(new_n9104), .A2(new_n9691), .B(new_n22065), .C(\a[53] ), .Y(new_n22068));
  A2O1A1O1Ixp25_ASAP7_75t_L g21812(.A1(new_n21804), .A2(new_n21810), .B(new_n21802), .C(new_n21948), .D(new_n21960), .Y(new_n22069));
  A2O1A1O1Ixp25_ASAP7_75t_L g21813(.A1(new_n21504), .A2(new_n4906), .B(new_n21796), .C(new_n21936), .D(new_n21946), .Y(new_n22070));
  INVx1_ASAP7_75t_L         g21814(.A(new_n22070), .Y(new_n22071));
  INVx1_ASAP7_75t_L         g21815(.A(new_n21936), .Y(new_n22072));
  NOR2xp33_ASAP7_75t_L      g21816(.A(new_n5855), .B(new_n13030), .Y(new_n22073));
  INVx1_ASAP7_75t_L         g21817(.A(new_n22073), .Y(new_n22074));
  O2A1O1Ixp33_ASAP7_75t_L   g21818(.A1(new_n12672), .A2(new_n6110), .B(new_n22074), .C(new_n22072), .Y(new_n22075));
  INVx1_ASAP7_75t_L         g21819(.A(new_n22075), .Y(new_n22076));
  O2A1O1Ixp33_ASAP7_75t_L   g21820(.A1(new_n12672), .A2(new_n6110), .B(new_n22074), .C(new_n21936), .Y(new_n22077));
  A2O1A1Ixp33_ASAP7_75t_L   g21821(.A1(new_n21936), .A2(new_n22076), .B(new_n22077), .C(new_n22071), .Y(new_n22078));
  INVx1_ASAP7_75t_L         g21822(.A(new_n22077), .Y(new_n22079));
  O2A1O1Ixp33_ASAP7_75t_L   g21823(.A1(new_n22075), .A2(new_n22072), .B(new_n22079), .C(new_n22071), .Y(new_n22080));
  NOR2xp33_ASAP7_75t_L      g21824(.A(new_n6671), .B(new_n12318), .Y(new_n22081));
  AOI221xp5_ASAP7_75t_L     g21825(.A1(new_n11995), .A2(\b[44] ), .B1(new_n13314), .B2(\b[42] ), .C(new_n22081), .Y(new_n22082));
  OAI21xp33_ASAP7_75t_L     g21826(.A1(new_n11998), .A2(new_n6951), .B(new_n22082), .Y(new_n22083));
  NOR2xp33_ASAP7_75t_L      g21827(.A(new_n11987), .B(new_n22083), .Y(new_n22084));
  O2A1O1Ixp33_ASAP7_75t_L   g21828(.A1(new_n11998), .A2(new_n6951), .B(new_n22082), .C(\a[62] ), .Y(new_n22085));
  NOR2xp33_ASAP7_75t_L      g21829(.A(new_n22085), .B(new_n22084), .Y(new_n22086));
  A2O1A1Ixp33_ASAP7_75t_L   g21830(.A1(new_n22078), .A2(new_n22071), .B(new_n22080), .C(new_n22086), .Y(new_n22087));
  A2O1A1Ixp33_ASAP7_75t_L   g21831(.A1(new_n13028), .A2(\b[37] ), .B(new_n21502), .C(new_n4906), .Y(new_n22088));
  A2O1A1O1Ixp25_ASAP7_75t_L g21832(.A1(new_n21792), .A2(new_n21794), .B(new_n21798), .C(new_n22088), .D(new_n22072), .Y(new_n22089));
  O2A1O1Ixp33_ASAP7_75t_L   g21833(.A1(new_n22089), .A2(new_n21946), .B(new_n22078), .C(new_n22080), .Y(new_n22090));
  NAND2xp33_ASAP7_75t_L     g21834(.A(\a[62] ), .B(new_n22083), .Y(new_n22091));
  A2O1A1Ixp33_ASAP7_75t_L   g21835(.A1(new_n22083), .A2(new_n22091), .B(new_n22084), .C(new_n22090), .Y(new_n22092));
  AND2x2_ASAP7_75t_L        g21836(.A(new_n22087), .B(new_n22092), .Y(new_n22093));
  NOR2xp33_ASAP7_75t_L      g21837(.A(new_n7249), .B(new_n11354), .Y(new_n22094));
  AOI221xp5_ASAP7_75t_L     g21838(.A1(\b[47] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[46] ), .C(new_n22094), .Y(new_n22095));
  O2A1O1Ixp33_ASAP7_75t_L   g21839(.A1(new_n11053), .A2(new_n7560), .B(new_n22095), .C(new_n11048), .Y(new_n22096));
  NOR2xp33_ASAP7_75t_L      g21840(.A(new_n11048), .B(new_n22096), .Y(new_n22097));
  O2A1O1Ixp33_ASAP7_75t_L   g21841(.A1(new_n11053), .A2(new_n7560), .B(new_n22095), .C(\a[59] ), .Y(new_n22098));
  NOR2xp33_ASAP7_75t_L      g21842(.A(new_n22098), .B(new_n22097), .Y(new_n22099));
  XOR2x2_ASAP7_75t_L        g21843(.A(new_n22099), .B(new_n22093), .Y(new_n22100));
  INVx1_ASAP7_75t_L         g21844(.A(new_n22100), .Y(new_n22101));
  NAND2xp33_ASAP7_75t_L     g21845(.A(new_n22069), .B(new_n22101), .Y(new_n22102));
  A2O1A1O1Ixp25_ASAP7_75t_L g21846(.A1(new_n21811), .A2(new_n21934), .B(new_n21949), .C(new_n21961), .D(new_n22101), .Y(new_n22103));
  INVx1_ASAP7_75t_L         g21847(.A(new_n22103), .Y(new_n22104));
  AND2x2_ASAP7_75t_L        g21848(.A(new_n22102), .B(new_n22104), .Y(new_n22105));
  NOR2xp33_ASAP7_75t_L      g21849(.A(new_n8427), .B(new_n10388), .Y(new_n22106));
  AOI221xp5_ASAP7_75t_L     g21850(.A1(new_n10086), .A2(\b[50] ), .B1(new_n11361), .B2(\b[48] ), .C(new_n22106), .Y(new_n22107));
  O2A1O1Ixp33_ASAP7_75t_L   g21851(.A1(new_n10088), .A2(new_n8764), .B(new_n22107), .C(new_n10083), .Y(new_n22108));
  INVx1_ASAP7_75t_L         g21852(.A(new_n22108), .Y(new_n22109));
  O2A1O1Ixp33_ASAP7_75t_L   g21853(.A1(new_n10088), .A2(new_n8764), .B(new_n22107), .C(\a[56] ), .Y(new_n22110));
  AOI211xp5_ASAP7_75t_L     g21854(.A1(new_n22109), .A2(\a[56] ), .B(new_n22110), .C(new_n22105), .Y(new_n22111));
  A2O1A1Ixp33_ASAP7_75t_L   g21855(.A1(\a[56] ), .A2(new_n22109), .B(new_n22110), .C(new_n22105), .Y(new_n22112));
  INVx1_ASAP7_75t_L         g21856(.A(new_n22112), .Y(new_n22113));
  NOR2xp33_ASAP7_75t_L      g21857(.A(new_n22111), .B(new_n22113), .Y(new_n22114));
  A2O1A1Ixp33_ASAP7_75t_L   g21858(.A1(new_n21966), .A2(new_n21963), .B(new_n21971), .C(new_n22114), .Y(new_n22115));
  INVx1_ASAP7_75t_L         g21859(.A(new_n22115), .Y(new_n22116));
  O2A1O1Ixp33_ASAP7_75t_L   g21860(.A1(new_n21820), .A2(new_n21825), .B(new_n21963), .C(new_n21971), .Y(new_n22117));
  NAND2xp33_ASAP7_75t_L     g21861(.A(new_n22117), .B(new_n22114), .Y(new_n22118));
  A2O1A1Ixp33_ASAP7_75t_L   g21862(.A1(new_n21970), .A2(new_n21967), .B(new_n22116), .C(new_n22118), .Y(new_n22119));
  NAND2xp33_ASAP7_75t_L     g21863(.A(new_n21967), .B(new_n21970), .Y(new_n22120));
  AOI21xp33_ASAP7_75t_L     g21864(.A1(new_n22067), .A2(\a[53] ), .B(new_n22068), .Y(new_n22121));
  NAND2xp33_ASAP7_75t_L     g21865(.A(new_n22121), .B(new_n22118), .Y(new_n22122));
  O2A1O1Ixp33_ASAP7_75t_L   g21866(.A1(new_n22111), .A2(new_n22113), .B(new_n22120), .C(new_n22122), .Y(new_n22123));
  A2O1A1O1Ixp25_ASAP7_75t_L g21867(.A1(new_n22067), .A2(\a[53] ), .B(new_n22068), .C(new_n22119), .D(new_n22123), .Y(new_n22124));
  INVx1_ASAP7_75t_L         g21868(.A(new_n22124), .Y(new_n22125));
  O2A1O1Ixp33_ASAP7_75t_L   g21869(.A1(new_n21973), .A2(new_n21977), .B(new_n21988), .C(new_n22125), .Y(new_n22126));
  A2O1A1O1Ixp25_ASAP7_75t_L g21870(.A1(new_n21986), .A2(\a[53] ), .B(new_n21987), .C(new_n21978), .D(new_n21980), .Y(new_n22127));
  NAND2xp33_ASAP7_75t_L     g21871(.A(new_n22127), .B(new_n22124), .Y(new_n22128));
  A2O1A1Ixp33_ASAP7_75t_L   g21872(.A1(new_n21988), .A2(new_n21981), .B(new_n22126), .C(new_n22128), .Y(new_n22129));
  INVx1_ASAP7_75t_L         g21873(.A(new_n22127), .Y(new_n22130));
  O2A1O1Ixp33_ASAP7_75t_L   g21874(.A1(new_n22117), .A2(new_n22116), .B(new_n22118), .C(new_n22121), .Y(new_n22131));
  AOI21xp33_ASAP7_75t_L     g21875(.A1(new_n22062), .A2(\a[50] ), .B(new_n22063), .Y(new_n22132));
  NAND2xp33_ASAP7_75t_L     g21876(.A(new_n22132), .B(new_n22128), .Y(new_n22133));
  O2A1O1Ixp33_ASAP7_75t_L   g21877(.A1(new_n22131), .A2(new_n22123), .B(new_n22130), .C(new_n22133), .Y(new_n22134));
  A2O1A1O1Ixp25_ASAP7_75t_L g21878(.A1(new_n22062), .A2(\a[50] ), .B(new_n22063), .C(new_n22129), .D(new_n22134), .Y(new_n22135));
  INVx1_ASAP7_75t_L         g21879(.A(new_n22135), .Y(new_n22136));
  O2A1O1Ixp33_ASAP7_75t_L   g21880(.A1(new_n21991), .A2(new_n22058), .B(new_n22003), .C(new_n22136), .Y(new_n22137));
  INVx1_ASAP7_75t_L         g21881(.A(new_n22137), .Y(new_n22138));
  O2A1O1Ixp33_ASAP7_75t_L   g21882(.A1(new_n21842), .A2(new_n21846), .B(new_n21992), .C(new_n22002), .Y(new_n22139));
  NAND2xp33_ASAP7_75t_L     g21883(.A(new_n22136), .B(new_n22139), .Y(new_n22140));
  AND2x2_ASAP7_75t_L        g21884(.A(new_n22140), .B(new_n22138), .Y(new_n22141));
  INVx1_ASAP7_75t_L         g21885(.A(new_n22141), .Y(new_n22142));
  NOR2xp33_ASAP7_75t_L      g21886(.A(new_n11591), .B(new_n7318), .Y(new_n22143));
  AOI221xp5_ASAP7_75t_L     g21887(.A1(new_n7333), .A2(\b[58] ), .B1(new_n7609), .B2(\b[57] ), .C(new_n22143), .Y(new_n22144));
  O2A1O1Ixp33_ASAP7_75t_L   g21888(.A1(new_n7321), .A2(new_n11597), .B(new_n22144), .C(new_n7316), .Y(new_n22145));
  O2A1O1Ixp33_ASAP7_75t_L   g21889(.A1(new_n7321), .A2(new_n11597), .B(new_n22144), .C(\a[47] ), .Y(new_n22146));
  INVx1_ASAP7_75t_L         g21890(.A(new_n22146), .Y(new_n22147));
  O2A1O1Ixp33_ASAP7_75t_L   g21891(.A1(new_n22145), .A2(new_n7316), .B(new_n22147), .C(new_n22142), .Y(new_n22148));
  INVx1_ASAP7_75t_L         g21892(.A(new_n22148), .Y(new_n22149));
  O2A1O1Ixp33_ASAP7_75t_L   g21893(.A1(new_n22145), .A2(new_n7316), .B(new_n22147), .C(new_n22141), .Y(new_n22150));
  AOI21xp33_ASAP7_75t_L     g21894(.A1(new_n22149), .A2(new_n22141), .B(new_n22150), .Y(new_n22151));
  A2O1A1Ixp33_ASAP7_75t_L   g21895(.A1(new_n21857), .A2(new_n21851), .B(new_n22005), .C(new_n22018), .Y(new_n22152));
  INVx1_ASAP7_75t_L         g21896(.A(new_n22152), .Y(new_n22153));
  NAND2xp33_ASAP7_75t_L     g21897(.A(new_n22151), .B(new_n22153), .Y(new_n22154));
  O2A1O1Ixp33_ASAP7_75t_L   g21898(.A1(new_n22005), .A2(new_n22006), .B(new_n22018), .C(new_n22151), .Y(new_n22155));
  INVx1_ASAP7_75t_L         g21899(.A(new_n22155), .Y(new_n22156));
  AND2x2_ASAP7_75t_L        g21900(.A(new_n22156), .B(new_n22154), .Y(new_n22157));
  INVx1_ASAP7_75t_L         g21901(.A(new_n22157), .Y(new_n22158));
  NOR2xp33_ASAP7_75t_L      g21902(.A(new_n11626), .B(new_n6741), .Y(new_n22159));
  AOI221xp5_ASAP7_75t_L     g21903(.A1(\b[62] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[61] ), .C(new_n22159), .Y(new_n22160));
  O2A1O1Ixp33_ASAP7_75t_L   g21904(.A1(new_n6443), .A2(new_n12610), .B(new_n22160), .C(new_n6439), .Y(new_n22161));
  O2A1O1Ixp33_ASAP7_75t_L   g21905(.A1(new_n6443), .A2(new_n12610), .B(new_n22160), .C(\a[44] ), .Y(new_n22162));
  INVx1_ASAP7_75t_L         g21906(.A(new_n22162), .Y(new_n22163));
  O2A1O1Ixp33_ASAP7_75t_L   g21907(.A1(new_n22161), .A2(new_n6439), .B(new_n22163), .C(new_n22158), .Y(new_n22164));
  INVx1_ASAP7_75t_L         g21908(.A(new_n22164), .Y(new_n22165));
  O2A1O1Ixp33_ASAP7_75t_L   g21909(.A1(new_n22161), .A2(new_n6439), .B(new_n22163), .C(new_n22157), .Y(new_n22166));
  AOI21xp33_ASAP7_75t_L     g21910(.A1(new_n22165), .A2(new_n22157), .B(new_n22166), .Y(new_n22167));
  A2O1A1Ixp33_ASAP7_75t_L   g21911(.A1(new_n22056), .A2(new_n22050), .B(new_n22057), .C(new_n22167), .Y(new_n22168));
  A2O1A1O1Ixp25_ASAP7_75t_L g21912(.A1(new_n12603), .A2(new_n14444), .B(new_n5630), .C(new_n5925), .D(new_n12956), .Y(new_n22169));
  A2O1A1O1Ixp25_ASAP7_75t_L g21913(.A1(new_n5637), .A2(new_n14172), .B(new_n5920), .C(\b[63] ), .D(new_n5626), .Y(new_n22170));
  O2A1O1Ixp33_ASAP7_75t_L   g21914(.A1(new_n22020), .A2(new_n22021), .B(new_n22031), .C(new_n22055), .Y(new_n22171));
  A2O1A1O1Ixp25_ASAP7_75t_L g21915(.A1(new_n22052), .A2(new_n22169), .B(new_n22170), .C(new_n22056), .D(new_n22171), .Y(new_n22172));
  A2O1A1Ixp33_ASAP7_75t_L   g21916(.A1(new_n22157), .A2(new_n22165), .B(new_n22166), .C(new_n22172), .Y(new_n22173));
  AND2x2_ASAP7_75t_L        g21917(.A(new_n22168), .B(new_n22173), .Y(new_n22174));
  A2O1A1O1Ixp25_ASAP7_75t_L g21918(.A1(new_n21888), .A2(new_n21882), .B(new_n21925), .C(new_n22034), .D(new_n22174), .Y(new_n22175));
  AND3x1_ASAP7_75t_L        g21919(.A(new_n22174), .B(new_n22034), .C(new_n21924), .Y(new_n22176));
  NOR2xp33_ASAP7_75t_L      g21920(.A(new_n22175), .B(new_n22176), .Y(new_n22177));
  XOR2x2_ASAP7_75t_L        g21921(.A(new_n22177), .B(new_n22048), .Y(\f[104] ));
  O2A1O1Ixp33_ASAP7_75t_L   g21922(.A1(new_n22127), .A2(new_n22126), .B(new_n22128), .C(new_n22132), .Y(new_n22179));
  NOR2xp33_ASAP7_75t_L      g21923(.A(new_n10332), .B(new_n10065), .Y(new_n22180));
  AOI221xp5_ASAP7_75t_L     g21924(.A1(new_n8175), .A2(\b[57] ), .B1(new_n8484), .B2(\b[55] ), .C(new_n22180), .Y(new_n22181));
  O2A1O1Ixp33_ASAP7_75t_L   g21925(.A1(new_n8176), .A2(new_n17096), .B(new_n22181), .C(new_n8172), .Y(new_n22182));
  INVx1_ASAP7_75t_L         g21926(.A(new_n22182), .Y(new_n22183));
  O2A1O1Ixp33_ASAP7_75t_L   g21927(.A1(new_n8176), .A2(new_n17096), .B(new_n22181), .C(\a[50] ), .Y(new_n22184));
  AO21x2_ASAP7_75t_L        g21928(.A1(\a[50] ), .A2(new_n22183), .B(new_n22184), .Y(new_n22185));
  A2O1A1Ixp33_ASAP7_75t_L   g21929(.A1(new_n21966), .A2(new_n21963), .B(new_n21971), .C(new_n22115), .Y(new_n22186));
  INVx1_ASAP7_75t_L         g21930(.A(new_n21935), .Y(new_n22187));
  O2A1O1Ixp33_ASAP7_75t_L   g21931(.A1(new_n5855), .A2(new_n12672), .B(new_n22187), .C(new_n5626), .Y(new_n22188));
  NOR2xp33_ASAP7_75t_L      g21932(.A(\a[41] ), .B(new_n22072), .Y(new_n22189));
  NOR2xp33_ASAP7_75t_L      g21933(.A(new_n22188), .B(new_n22189), .Y(new_n22190));
  NOR2xp33_ASAP7_75t_L      g21934(.A(new_n6110), .B(new_n13030), .Y(new_n22191));
  O2A1O1Ixp33_ASAP7_75t_L   g21935(.A1(new_n12669), .A2(new_n12671), .B(\b[42] ), .C(new_n22191), .Y(new_n22192));
  NAND2xp33_ASAP7_75t_L     g21936(.A(new_n22192), .B(new_n22190), .Y(new_n22193));
  INVx1_ASAP7_75t_L         g21937(.A(new_n22190), .Y(new_n22194));
  A2O1A1Ixp33_ASAP7_75t_L   g21938(.A1(\b[42] ), .A2(new_n13028), .B(new_n22191), .C(new_n22194), .Y(new_n22195));
  AND2x2_ASAP7_75t_L        g21939(.A(new_n22193), .B(new_n22195), .Y(new_n22196));
  INVx1_ASAP7_75t_L         g21940(.A(new_n22196), .Y(new_n22197));
  NOR2xp33_ASAP7_75t_L      g21941(.A(new_n6944), .B(new_n12318), .Y(new_n22198));
  AOI221xp5_ASAP7_75t_L     g21942(.A1(new_n11995), .A2(\b[45] ), .B1(new_n13314), .B2(\b[43] ), .C(new_n22198), .Y(new_n22199));
  O2A1O1Ixp33_ASAP7_75t_L   g21943(.A1(new_n11998), .A2(new_n7255), .B(new_n22199), .C(new_n11987), .Y(new_n22200));
  O2A1O1Ixp33_ASAP7_75t_L   g21944(.A1(new_n11998), .A2(new_n7255), .B(new_n22199), .C(\a[62] ), .Y(new_n22201));
  INVx1_ASAP7_75t_L         g21945(.A(new_n22201), .Y(new_n22202));
  O2A1O1Ixp33_ASAP7_75t_L   g21946(.A1(new_n22200), .A2(new_n11987), .B(new_n22202), .C(new_n22197), .Y(new_n22203));
  INVx1_ASAP7_75t_L         g21947(.A(new_n22203), .Y(new_n22204));
  O2A1O1Ixp33_ASAP7_75t_L   g21948(.A1(new_n22200), .A2(new_n11987), .B(new_n22202), .C(new_n22196), .Y(new_n22205));
  AOI21xp33_ASAP7_75t_L     g21949(.A1(new_n22204), .A2(new_n22196), .B(new_n22205), .Y(new_n22206));
  O2A1O1Ixp33_ASAP7_75t_L   g21950(.A1(new_n21936), .A2(new_n22077), .B(new_n22071), .C(new_n22075), .Y(new_n22207));
  AND2x2_ASAP7_75t_L        g21951(.A(new_n22206), .B(new_n22207), .Y(new_n22208));
  O2A1O1Ixp33_ASAP7_75t_L   g21952(.A1(new_n12669), .A2(new_n12671), .B(\b[41] ), .C(new_n22073), .Y(new_n22209));
  O2A1O1Ixp33_ASAP7_75t_L   g21953(.A1(new_n22072), .A2(new_n22209), .B(new_n22078), .C(new_n22206), .Y(new_n22210));
  NOR2xp33_ASAP7_75t_L      g21954(.A(new_n22210), .B(new_n22208), .Y(new_n22211));
  NOR2xp33_ASAP7_75t_L      g21955(.A(new_n7270), .B(new_n11354), .Y(new_n22212));
  AOI221xp5_ASAP7_75t_L     g21956(.A1(\b[48] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[47] ), .C(new_n22212), .Y(new_n22213));
  O2A1O1Ixp33_ASAP7_75t_L   g21957(.A1(new_n11053), .A2(new_n7868), .B(new_n22213), .C(new_n11048), .Y(new_n22214));
  INVx1_ASAP7_75t_L         g21958(.A(new_n22214), .Y(new_n22215));
  O2A1O1Ixp33_ASAP7_75t_L   g21959(.A1(new_n11053), .A2(new_n7868), .B(new_n22213), .C(\a[59] ), .Y(new_n22216));
  A2O1A1Ixp33_ASAP7_75t_L   g21960(.A1(\a[59] ), .A2(new_n22215), .B(new_n22216), .C(new_n22211), .Y(new_n22217));
  INVx1_ASAP7_75t_L         g21961(.A(new_n22216), .Y(new_n22218));
  O2A1O1Ixp33_ASAP7_75t_L   g21962(.A1(new_n22214), .A2(new_n11048), .B(new_n22218), .C(new_n22211), .Y(new_n22219));
  AO21x2_ASAP7_75t_L        g21963(.A1(new_n22211), .A2(new_n22217), .B(new_n22219), .Y(new_n22220));
  INVx1_ASAP7_75t_L         g21964(.A(new_n22086), .Y(new_n22221));
  A2O1A1Ixp33_ASAP7_75t_L   g21965(.A1(new_n22078), .A2(new_n22071), .B(new_n22080), .C(new_n22221), .Y(new_n22222));
  A2O1A1Ixp33_ASAP7_75t_L   g21966(.A1(new_n22092), .A2(new_n22087), .B(new_n22099), .C(new_n22222), .Y(new_n22223));
  XOR2x2_ASAP7_75t_L        g21967(.A(new_n22223), .B(new_n22220), .Y(new_n22224));
  NOR2xp33_ASAP7_75t_L      g21968(.A(new_n8755), .B(new_n10388), .Y(new_n22225));
  AOI221xp5_ASAP7_75t_L     g21969(.A1(new_n10086), .A2(\b[51] ), .B1(new_n11361), .B2(\b[49] ), .C(new_n22225), .Y(new_n22226));
  O2A1O1Ixp33_ASAP7_75t_L   g21970(.A1(new_n10088), .A2(new_n8789), .B(new_n22226), .C(new_n10083), .Y(new_n22227));
  O2A1O1Ixp33_ASAP7_75t_L   g21971(.A1(new_n10088), .A2(new_n8789), .B(new_n22226), .C(\a[56] ), .Y(new_n22228));
  INVx1_ASAP7_75t_L         g21972(.A(new_n22228), .Y(new_n22229));
  INVx1_ASAP7_75t_L         g21973(.A(new_n22224), .Y(new_n22230));
  O2A1O1Ixp33_ASAP7_75t_L   g21974(.A1(new_n10083), .A2(new_n22227), .B(new_n22229), .C(new_n22230), .Y(new_n22231));
  INVx1_ASAP7_75t_L         g21975(.A(new_n22231), .Y(new_n22232));
  O2A1O1Ixp33_ASAP7_75t_L   g21976(.A1(new_n10083), .A2(new_n22227), .B(new_n22229), .C(new_n22224), .Y(new_n22233));
  AOI21xp33_ASAP7_75t_L     g21977(.A1(new_n22232), .A2(new_n22224), .B(new_n22233), .Y(new_n22234));
  O2A1O1Ixp33_ASAP7_75t_L   g21978(.A1(new_n22069), .A2(new_n22101), .B(new_n22112), .C(new_n22234), .Y(new_n22235));
  A2O1A1O1Ixp25_ASAP7_75t_L g21979(.A1(new_n22109), .A2(\a[56] ), .B(new_n22110), .C(new_n22102), .D(new_n22103), .Y(new_n22236));
  A2O1A1Ixp33_ASAP7_75t_L   g21980(.A1(new_n22232), .A2(new_n22224), .B(new_n22233), .C(new_n22236), .Y(new_n22237));
  A2O1A1Ixp33_ASAP7_75t_L   g21981(.A1(new_n22112), .A2(new_n22104), .B(new_n22235), .C(new_n22237), .Y(new_n22238));
  INVx1_ASAP7_75t_L         g21982(.A(new_n22238), .Y(new_n22239));
  NOR2xp33_ASAP7_75t_L      g21983(.A(new_n9683), .B(new_n10400), .Y(new_n22240));
  AOI221xp5_ASAP7_75t_L     g21984(.A1(new_n9102), .A2(\b[54] ), .B1(new_n10398), .B2(\b[52] ), .C(new_n22240), .Y(new_n22241));
  O2A1O1Ixp33_ASAP7_75t_L   g21985(.A1(new_n9104), .A2(new_n9718), .B(new_n22241), .C(new_n9099), .Y(new_n22242));
  O2A1O1Ixp33_ASAP7_75t_L   g21986(.A1(new_n9104), .A2(new_n9718), .B(new_n22241), .C(\a[53] ), .Y(new_n22243));
  INVx1_ASAP7_75t_L         g21987(.A(new_n22243), .Y(new_n22244));
  OAI211xp5_ASAP7_75t_L     g21988(.A1(new_n9099), .A2(new_n22242), .B(new_n22239), .C(new_n22244), .Y(new_n22245));
  O2A1O1Ixp33_ASAP7_75t_L   g21989(.A1(new_n22242), .A2(new_n9099), .B(new_n22244), .C(new_n22239), .Y(new_n22246));
  INVx1_ASAP7_75t_L         g21990(.A(new_n22246), .Y(new_n22247));
  AND2x2_ASAP7_75t_L        g21991(.A(new_n22245), .B(new_n22247), .Y(new_n22248));
  INVx1_ASAP7_75t_L         g21992(.A(new_n22248), .Y(new_n22249));
  A2O1A1O1Ixp25_ASAP7_75t_L g21993(.A1(new_n22186), .A2(new_n22118), .B(new_n22121), .C(new_n22115), .D(new_n22249), .Y(new_n22250));
  INVx1_ASAP7_75t_L         g21994(.A(new_n22250), .Y(new_n22251));
  A2O1A1O1Ixp25_ASAP7_75t_L g21995(.A1(new_n22067), .A2(\a[53] ), .B(new_n22068), .C(new_n22119), .D(new_n22116), .Y(new_n22252));
  NAND2xp33_ASAP7_75t_L     g21996(.A(new_n22252), .B(new_n22249), .Y(new_n22253));
  AO21x2_ASAP7_75t_L        g21997(.A1(new_n22253), .A2(new_n22251), .B(new_n22185), .Y(new_n22254));
  AND2x2_ASAP7_75t_L        g21998(.A(new_n22253), .B(new_n22251), .Y(new_n22255));
  A2O1A1Ixp33_ASAP7_75t_L   g21999(.A1(new_n22183), .A2(\a[50] ), .B(new_n22184), .C(new_n22255), .Y(new_n22256));
  AND2x2_ASAP7_75t_L        g22000(.A(new_n22254), .B(new_n22256), .Y(new_n22257));
  A2O1A1Ixp33_ASAP7_75t_L   g22001(.A1(new_n22124), .A2(new_n22130), .B(new_n22179), .C(new_n22257), .Y(new_n22258));
  A2O1A1O1Ixp25_ASAP7_75t_L g22002(.A1(new_n22062), .A2(\a[50] ), .B(new_n22063), .C(new_n22129), .D(new_n22126), .Y(new_n22259));
  INVx1_ASAP7_75t_L         g22003(.A(new_n22257), .Y(new_n22260));
  NAND2xp33_ASAP7_75t_L     g22004(.A(new_n22259), .B(new_n22260), .Y(new_n22261));
  AND2x2_ASAP7_75t_L        g22005(.A(new_n22258), .B(new_n22261), .Y(new_n22262));
  INVx1_ASAP7_75t_L         g22006(.A(new_n22262), .Y(new_n22263));
  NOR2xp33_ASAP7_75t_L      g22007(.A(new_n11626), .B(new_n7318), .Y(new_n22264));
  AOI221xp5_ASAP7_75t_L     g22008(.A1(new_n7333), .A2(\b[59] ), .B1(new_n7609), .B2(\b[58] ), .C(new_n22264), .Y(new_n22265));
  O2A1O1Ixp33_ASAP7_75t_L   g22009(.A1(new_n7321), .A2(new_n11634), .B(new_n22265), .C(new_n7316), .Y(new_n22266));
  O2A1O1Ixp33_ASAP7_75t_L   g22010(.A1(new_n7321), .A2(new_n11634), .B(new_n22265), .C(\a[47] ), .Y(new_n22267));
  INVx1_ASAP7_75t_L         g22011(.A(new_n22267), .Y(new_n22268));
  O2A1O1Ixp33_ASAP7_75t_L   g22012(.A1(new_n22266), .A2(new_n7316), .B(new_n22268), .C(new_n22263), .Y(new_n22269));
  INVx1_ASAP7_75t_L         g22013(.A(new_n22269), .Y(new_n22270));
  O2A1O1Ixp33_ASAP7_75t_L   g22014(.A1(new_n22266), .A2(new_n7316), .B(new_n22268), .C(new_n22262), .Y(new_n22271));
  AOI21xp33_ASAP7_75t_L     g22015(.A1(new_n22270), .A2(new_n22262), .B(new_n22271), .Y(new_n22272));
  O2A1O1Ixp33_ASAP7_75t_L   g22016(.A1(new_n21993), .A2(new_n22002), .B(new_n22135), .C(new_n22148), .Y(new_n22273));
  NAND2xp33_ASAP7_75t_L     g22017(.A(new_n22272), .B(new_n22273), .Y(new_n22274));
  O2A1O1Ixp33_ASAP7_75t_L   g22018(.A1(new_n22139), .A2(new_n22136), .B(new_n22149), .C(new_n22272), .Y(new_n22275));
  INVx1_ASAP7_75t_L         g22019(.A(new_n22275), .Y(new_n22276));
  AND2x2_ASAP7_75t_L        g22020(.A(new_n22274), .B(new_n22276), .Y(new_n22277));
  INVx1_ASAP7_75t_L         g22021(.A(new_n22277), .Y(new_n22278));
  NOR2xp33_ASAP7_75t_L      g22022(.A(new_n12258), .B(new_n6741), .Y(new_n22279));
  AOI221xp5_ASAP7_75t_L     g22023(.A1(\b[63] ), .A2(new_n6442), .B1(new_n6436), .B2(\b[62] ), .C(new_n22279), .Y(new_n22280));
  O2A1O1Ixp33_ASAP7_75t_L   g22024(.A1(new_n6443), .A2(new_n17815), .B(new_n22280), .C(new_n6439), .Y(new_n22281));
  O2A1O1Ixp33_ASAP7_75t_L   g22025(.A1(new_n6443), .A2(new_n17815), .B(new_n22280), .C(\a[44] ), .Y(new_n22282));
  INVx1_ASAP7_75t_L         g22026(.A(new_n22282), .Y(new_n22283));
  O2A1O1Ixp33_ASAP7_75t_L   g22027(.A1(new_n22281), .A2(new_n6439), .B(new_n22283), .C(new_n22278), .Y(new_n22284));
  INVx1_ASAP7_75t_L         g22028(.A(new_n22284), .Y(new_n22285));
  O2A1O1Ixp33_ASAP7_75t_L   g22029(.A1(new_n22281), .A2(new_n6439), .B(new_n22283), .C(new_n22277), .Y(new_n22286));
  AOI21xp33_ASAP7_75t_L     g22030(.A1(new_n22285), .A2(new_n22277), .B(new_n22286), .Y(new_n22287));
  A2O1A1O1Ixp25_ASAP7_75t_L g22031(.A1(new_n22149), .A2(new_n22141), .B(new_n22150), .C(new_n22152), .D(new_n22164), .Y(new_n22288));
  NAND2xp33_ASAP7_75t_L     g22032(.A(new_n22287), .B(new_n22288), .Y(new_n22289));
  O2A1O1Ixp33_ASAP7_75t_L   g22033(.A1(new_n22151), .A2(new_n22153), .B(new_n22165), .C(new_n22287), .Y(new_n22290));
  INVx1_ASAP7_75t_L         g22034(.A(new_n22290), .Y(new_n22291));
  AND2x2_ASAP7_75t_L        g22035(.A(new_n22289), .B(new_n22291), .Y(new_n22292));
  INVx1_ASAP7_75t_L         g22036(.A(new_n22292), .Y(new_n22293));
  O2A1O1Ixp33_ASAP7_75t_L   g22037(.A1(new_n22172), .A2(new_n22167), .B(new_n22056), .C(new_n22293), .Y(new_n22294));
  INVx1_ASAP7_75t_L         g22038(.A(new_n22057), .Y(new_n22295));
  O2A1O1Ixp33_ASAP7_75t_L   g22039(.A1(new_n22049), .A2(new_n22055), .B(new_n22295), .C(new_n22167), .Y(new_n22296));
  NOR3xp33_ASAP7_75t_L      g22040(.A(new_n22292), .B(new_n22296), .C(new_n22055), .Y(new_n22297));
  NOR2xp33_ASAP7_75t_L      g22041(.A(new_n22297), .B(new_n22294), .Y(new_n22298));
  A2O1A1Ixp33_ASAP7_75t_L   g22042(.A1(new_n22048), .A2(new_n22177), .B(new_n22175), .C(new_n22298), .Y(new_n22299));
  INVx1_ASAP7_75t_L         g22043(.A(new_n22299), .Y(new_n22300));
  A2O1A1Ixp33_ASAP7_75t_L   g22044(.A1(new_n21754), .A2(new_n21763), .B(new_n21899), .C(new_n21897), .Y(new_n22301));
  A2O1A1Ixp33_ASAP7_75t_L   g22045(.A1(new_n22301), .A2(new_n22037), .B(new_n22044), .C(new_n22177), .Y(new_n22302));
  A2O1A1Ixp33_ASAP7_75t_L   g22046(.A1(new_n22034), .A2(new_n21924), .B(new_n22174), .C(new_n22302), .Y(new_n22303));
  NOR2xp33_ASAP7_75t_L      g22047(.A(new_n22298), .B(new_n22303), .Y(new_n22304));
  NOR2xp33_ASAP7_75t_L      g22048(.A(new_n22300), .B(new_n22304), .Y(\f[105] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g22049(.A1(new_n22052), .A2(new_n22169), .B(new_n22170), .C(new_n22050), .D(new_n22296), .Y(new_n22306));
  NAND2xp33_ASAP7_75t_L     g22050(.A(\b[60] ), .B(new_n7333), .Y(new_n22307));
  OAI221xp5_ASAP7_75t_L     g22051(.A1(new_n7318), .A2(new_n12258), .B1(new_n11591), .B2(new_n7614), .C(new_n22307), .Y(new_n22308));
  A2O1A1Ixp33_ASAP7_75t_L   g22052(.A1(new_n12269), .A2(new_n7322), .B(new_n22308), .C(\a[47] ), .Y(new_n22309));
  NAND2xp33_ASAP7_75t_L     g22053(.A(\a[47] ), .B(new_n22309), .Y(new_n22310));
  A2O1A1Ixp33_ASAP7_75t_L   g22054(.A1(new_n12269), .A2(new_n7322), .B(new_n22308), .C(new_n7316), .Y(new_n22311));
  NAND2xp33_ASAP7_75t_L     g22055(.A(new_n22311), .B(new_n22310), .Y(new_n22312));
  INVx1_ASAP7_75t_L         g22056(.A(new_n22252), .Y(new_n22313));
  A2O1A1Ixp33_ASAP7_75t_L   g22057(.A1(new_n22217), .A2(new_n22211), .B(new_n22219), .C(new_n22223), .Y(new_n22314));
  O2A1O1Ixp33_ASAP7_75t_L   g22058(.A1(new_n5855), .A2(new_n12672), .B(new_n22187), .C(\a[41] ), .Y(new_n22315));
  A2O1A1O1Ixp25_ASAP7_75t_L g22059(.A1(new_n13028), .A2(\b[42] ), .B(new_n22191), .C(new_n22194), .D(new_n22315), .Y(new_n22316));
  NOR2xp33_ASAP7_75t_L      g22060(.A(new_n6378), .B(new_n13030), .Y(new_n22317));
  O2A1O1Ixp33_ASAP7_75t_L   g22061(.A1(new_n12669), .A2(new_n12671), .B(\b[43] ), .C(new_n22317), .Y(new_n22318));
  INVx1_ASAP7_75t_L         g22062(.A(new_n22318), .Y(new_n22319));
  INVx1_ASAP7_75t_L         g22063(.A(new_n22315), .Y(new_n22320));
  O2A1O1Ixp33_ASAP7_75t_L   g22064(.A1(new_n22192), .A2(new_n22190), .B(new_n22320), .C(new_n22319), .Y(new_n22321));
  NAND2xp33_ASAP7_75t_L     g22065(.A(new_n22318), .B(new_n22316), .Y(new_n22322));
  NOR2xp33_ASAP7_75t_L      g22066(.A(new_n7249), .B(new_n12318), .Y(new_n22323));
  AOI221xp5_ASAP7_75t_L     g22067(.A1(new_n11995), .A2(\b[46] ), .B1(new_n13314), .B2(\b[44] ), .C(new_n22323), .Y(new_n22324));
  INVx1_ASAP7_75t_L         g22068(.A(new_n22324), .Y(new_n22325));
  A2O1A1Ixp33_ASAP7_75t_L   g22069(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n22324), .Y(new_n22326));
  O2A1O1Ixp33_ASAP7_75t_L   g22070(.A1(new_n22325), .A2(new_n7278), .B(new_n22326), .C(new_n11987), .Y(new_n22327));
  O2A1O1Ixp33_ASAP7_75t_L   g22071(.A1(new_n11998), .A2(new_n7279), .B(new_n22324), .C(\a[62] ), .Y(new_n22328));
  NOR2xp33_ASAP7_75t_L      g22072(.A(new_n22327), .B(new_n22328), .Y(new_n22329));
  O2A1O1Ixp33_ASAP7_75t_L   g22073(.A1(new_n22316), .A2(new_n22321), .B(new_n22322), .C(new_n22329), .Y(new_n22330));
  INVx1_ASAP7_75t_L         g22074(.A(new_n22330), .Y(new_n22331));
  A2O1A1Ixp33_ASAP7_75t_L   g22075(.A1(new_n22320), .A2(new_n22195), .B(new_n22321), .C(new_n22322), .Y(new_n22332));
  OR3x1_ASAP7_75t_L         g22076(.A(new_n22328), .B(new_n22332), .C(new_n22327), .Y(new_n22333));
  AND2x2_ASAP7_75t_L        g22077(.A(new_n22333), .B(new_n22331), .Y(new_n22334));
  INVx1_ASAP7_75t_L         g22078(.A(new_n22334), .Y(new_n22335));
  O2A1O1Ixp33_ASAP7_75t_L   g22079(.A1(new_n22206), .A2(new_n22207), .B(new_n22204), .C(new_n22335), .Y(new_n22336));
  INVx1_ASAP7_75t_L         g22080(.A(new_n22336), .Y(new_n22337));
  INVx1_ASAP7_75t_L         g22081(.A(new_n22207), .Y(new_n22338));
  O2A1O1Ixp33_ASAP7_75t_L   g22082(.A1(new_n22205), .A2(new_n22196), .B(new_n22338), .C(new_n22203), .Y(new_n22339));
  NAND2xp33_ASAP7_75t_L     g22083(.A(new_n22339), .B(new_n22335), .Y(new_n22340));
  AND2x2_ASAP7_75t_L        g22084(.A(new_n22340), .B(new_n22337), .Y(new_n22341));
  NOR2xp33_ASAP7_75t_L      g22085(.A(new_n7552), .B(new_n11354), .Y(new_n22342));
  AOI221xp5_ASAP7_75t_L     g22086(.A1(\b[49] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[48] ), .C(new_n22342), .Y(new_n22343));
  O2A1O1Ixp33_ASAP7_75t_L   g22087(.A1(new_n11053), .A2(new_n14802), .B(new_n22343), .C(new_n11048), .Y(new_n22344));
  INVx1_ASAP7_75t_L         g22088(.A(new_n22344), .Y(new_n22345));
  O2A1O1Ixp33_ASAP7_75t_L   g22089(.A1(new_n11053), .A2(new_n14802), .B(new_n22343), .C(\a[59] ), .Y(new_n22346));
  A2O1A1Ixp33_ASAP7_75t_L   g22090(.A1(\a[59] ), .A2(new_n22345), .B(new_n22346), .C(new_n22341), .Y(new_n22347));
  INVx1_ASAP7_75t_L         g22091(.A(new_n22346), .Y(new_n22348));
  O2A1O1Ixp33_ASAP7_75t_L   g22092(.A1(new_n22344), .A2(new_n11048), .B(new_n22348), .C(new_n22341), .Y(new_n22349));
  AOI21xp33_ASAP7_75t_L     g22093(.A1(new_n22347), .A2(new_n22341), .B(new_n22349), .Y(new_n22350));
  NAND3xp33_ASAP7_75t_L     g22094(.A(new_n22350), .B(new_n22314), .C(new_n22217), .Y(new_n22351));
  NAND2xp33_ASAP7_75t_L     g22095(.A(new_n22217), .B(new_n22314), .Y(new_n22352));
  A2O1A1Ixp33_ASAP7_75t_L   g22096(.A1(new_n22347), .A2(new_n22341), .B(new_n22349), .C(new_n22352), .Y(new_n22353));
  NAND2xp33_ASAP7_75t_L     g22097(.A(new_n22353), .B(new_n22351), .Y(new_n22354));
  INVx1_ASAP7_75t_L         g22098(.A(new_n22354), .Y(new_n22355));
  NOR2xp33_ASAP7_75t_L      g22099(.A(new_n8779), .B(new_n10388), .Y(new_n22356));
  AOI221xp5_ASAP7_75t_L     g22100(.A1(new_n10086), .A2(\b[52] ), .B1(new_n11361), .B2(\b[50] ), .C(new_n22356), .Y(new_n22357));
  INVx1_ASAP7_75t_L         g22101(.A(new_n22357), .Y(new_n22358));
  A2O1A1Ixp33_ASAP7_75t_L   g22102(.A1(new_n9367), .A2(new_n10386), .B(new_n22358), .C(\a[56] ), .Y(new_n22359));
  O2A1O1Ixp33_ASAP7_75t_L   g22103(.A1(new_n10088), .A2(new_n17363), .B(new_n22357), .C(\a[56] ), .Y(new_n22360));
  A2O1A1Ixp33_ASAP7_75t_L   g22104(.A1(\a[56] ), .A2(new_n22359), .B(new_n22360), .C(new_n22355), .Y(new_n22361));
  NAND2xp33_ASAP7_75t_L     g22105(.A(new_n22355), .B(new_n22361), .Y(new_n22362));
  A2O1A1Ixp33_ASAP7_75t_L   g22106(.A1(\a[56] ), .A2(new_n22359), .B(new_n22360), .C(new_n22354), .Y(new_n22363));
  A2O1A1Ixp33_ASAP7_75t_L   g22107(.A1(new_n22112), .A2(new_n22104), .B(new_n22234), .C(new_n22232), .Y(new_n22364));
  INVx1_ASAP7_75t_L         g22108(.A(new_n22364), .Y(new_n22365));
  AND3x1_ASAP7_75t_L        g22109(.A(new_n22365), .B(new_n22363), .C(new_n22362), .Y(new_n22366));
  AOI211xp5_ASAP7_75t_L     g22110(.A1(new_n22359), .A2(\a[56] ), .B(new_n22360), .C(new_n22354), .Y(new_n22367));
  A2O1A1O1Ixp25_ASAP7_75t_L g22111(.A1(new_n22359), .A2(\a[56] ), .B(new_n22360), .C(new_n22361), .D(new_n22367), .Y(new_n22368));
  O2A1O1Ixp33_ASAP7_75t_L   g22112(.A1(new_n22236), .A2(new_n22234), .B(new_n22232), .C(new_n22368), .Y(new_n22369));
  NOR2xp33_ASAP7_75t_L      g22113(.A(new_n22366), .B(new_n22369), .Y(new_n22370));
  NOR2xp33_ASAP7_75t_L      g22114(.A(new_n9709), .B(new_n10400), .Y(new_n22371));
  AOI221xp5_ASAP7_75t_L     g22115(.A1(new_n9102), .A2(\b[55] ), .B1(new_n10398), .B2(\b[53] ), .C(new_n22371), .Y(new_n22372));
  O2A1O1Ixp33_ASAP7_75t_L   g22116(.A1(new_n9104), .A2(new_n15849), .B(new_n22372), .C(new_n9099), .Y(new_n22373));
  INVx1_ASAP7_75t_L         g22117(.A(new_n22373), .Y(new_n22374));
  O2A1O1Ixp33_ASAP7_75t_L   g22118(.A1(new_n9104), .A2(new_n15849), .B(new_n22372), .C(\a[53] ), .Y(new_n22375));
  A2O1A1Ixp33_ASAP7_75t_L   g22119(.A1(\a[53] ), .A2(new_n22374), .B(new_n22375), .C(new_n22370), .Y(new_n22376));
  INVx1_ASAP7_75t_L         g22120(.A(new_n22375), .Y(new_n22377));
  O2A1O1Ixp33_ASAP7_75t_L   g22121(.A1(new_n22373), .A2(new_n9099), .B(new_n22377), .C(new_n22370), .Y(new_n22378));
  AOI21xp33_ASAP7_75t_L     g22122(.A1(new_n22376), .A2(new_n22370), .B(new_n22378), .Y(new_n22379));
  A2O1A1Ixp33_ASAP7_75t_L   g22123(.A1(new_n22245), .A2(new_n22313), .B(new_n22246), .C(new_n22379), .Y(new_n22380));
  O2A1O1Ixp33_ASAP7_75t_L   g22124(.A1(new_n22116), .A2(new_n22131), .B(new_n22245), .C(new_n22246), .Y(new_n22381));
  A2O1A1Ixp33_ASAP7_75t_L   g22125(.A1(new_n22376), .A2(new_n22370), .B(new_n22378), .C(new_n22381), .Y(new_n22382));
  AND2x2_ASAP7_75t_L        g22126(.A(new_n22382), .B(new_n22380), .Y(new_n22383));
  INVx1_ASAP7_75t_L         g22127(.A(new_n22383), .Y(new_n22384));
  NOR2xp33_ASAP7_75t_L      g22128(.A(new_n10978), .B(new_n10065), .Y(new_n22385));
  AOI221xp5_ASAP7_75t_L     g22129(.A1(new_n8175), .A2(\b[58] ), .B1(new_n8484), .B2(\b[56] ), .C(new_n22385), .Y(new_n22386));
  O2A1O1Ixp33_ASAP7_75t_L   g22130(.A1(new_n8176), .A2(new_n20073), .B(new_n22386), .C(new_n8172), .Y(new_n22387));
  INVx1_ASAP7_75t_L         g22131(.A(new_n22387), .Y(new_n22388));
  O2A1O1Ixp33_ASAP7_75t_L   g22132(.A1(new_n8176), .A2(new_n20073), .B(new_n22386), .C(\a[50] ), .Y(new_n22389));
  AOI21xp33_ASAP7_75t_L     g22133(.A1(new_n22388), .A2(\a[50] ), .B(new_n22389), .Y(new_n22390));
  INVx1_ASAP7_75t_L         g22134(.A(new_n22390), .Y(new_n22391));
  NOR2xp33_ASAP7_75t_L      g22135(.A(new_n22391), .B(new_n22384), .Y(new_n22392));
  INVx1_ASAP7_75t_L         g22136(.A(new_n22392), .Y(new_n22393));
  A2O1A1Ixp33_ASAP7_75t_L   g22137(.A1(\a[50] ), .A2(new_n22388), .B(new_n22389), .C(new_n22384), .Y(new_n22394));
  AND2x2_ASAP7_75t_L        g22138(.A(new_n22394), .B(new_n22393), .Y(new_n22395));
  INVx1_ASAP7_75t_L         g22139(.A(new_n22395), .Y(new_n22396));
  O2A1O1Ixp33_ASAP7_75t_L   g22140(.A1(new_n22259), .A2(new_n22260), .B(new_n22256), .C(new_n22396), .Y(new_n22397));
  INVx1_ASAP7_75t_L         g22141(.A(new_n22397), .Y(new_n22398));
  O2A1O1Ixp33_ASAP7_75t_L   g22142(.A1(new_n22259), .A2(new_n22260), .B(new_n22256), .C(new_n22395), .Y(new_n22399));
  A2O1A1Ixp33_ASAP7_75t_L   g22143(.A1(new_n22398), .A2(new_n22395), .B(new_n22399), .C(new_n22312), .Y(new_n22400));
  A2O1A1Ixp33_ASAP7_75t_L   g22144(.A1(new_n22398), .A2(new_n22395), .B(new_n22399), .C(new_n22400), .Y(new_n22401));
  INVx1_ASAP7_75t_L         g22145(.A(new_n22401), .Y(new_n22402));
  A2O1A1Ixp33_ASAP7_75t_L   g22146(.A1(new_n22149), .A2(new_n22138), .B(new_n22272), .C(new_n22270), .Y(new_n22403));
  AOI22xp33_ASAP7_75t_L     g22147(.A1(new_n6436), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n6742), .Y(new_n22404));
  INVx1_ASAP7_75t_L         g22148(.A(new_n22404), .Y(new_n22405));
  A2O1A1Ixp33_ASAP7_75t_L   g22149(.A1(new_n6438), .A2(new_n6440), .B(new_n6152), .C(new_n22404), .Y(new_n22406));
  O2A1O1Ixp33_ASAP7_75t_L   g22150(.A1(new_n22405), .A2(new_n17329), .B(new_n22406), .C(new_n6439), .Y(new_n22407));
  O2A1O1Ixp33_ASAP7_75t_L   g22151(.A1(new_n6443), .A2(new_n12993), .B(new_n22404), .C(\a[44] ), .Y(new_n22408));
  OAI21xp33_ASAP7_75t_L     g22152(.A1(new_n22407), .A2(new_n22408), .B(new_n22403), .Y(new_n22409));
  NOR2xp33_ASAP7_75t_L      g22153(.A(new_n22408), .B(new_n22407), .Y(new_n22410));
  NAND3xp33_ASAP7_75t_L     g22154(.A(new_n22276), .B(new_n22270), .C(new_n22410), .Y(new_n22411));
  NAND2xp33_ASAP7_75t_L     g22155(.A(new_n22409), .B(new_n22411), .Y(new_n22412));
  INVx1_ASAP7_75t_L         g22156(.A(new_n22412), .Y(new_n22413));
  A2O1A1Ixp33_ASAP7_75t_L   g22157(.A1(new_n22312), .A2(new_n22400), .B(new_n22402), .C(new_n22413), .Y(new_n22414));
  AOI211xp5_ASAP7_75t_L     g22158(.A1(new_n22312), .A2(new_n22400), .B(new_n22402), .C(new_n22412), .Y(new_n22415));
  A2O1A1O1Ixp25_ASAP7_75t_L g22159(.A1(new_n22400), .A2(new_n22312), .B(new_n22402), .C(new_n22414), .D(new_n22415), .Y(new_n22416));
  NAND3xp33_ASAP7_75t_L     g22160(.A(new_n22291), .B(new_n22285), .C(new_n22416), .Y(new_n22417));
  A2O1A1O1Ixp25_ASAP7_75t_L g22161(.A1(new_n22156), .A2(new_n22165), .B(new_n22287), .C(new_n22285), .D(new_n22416), .Y(new_n22418));
  INVx1_ASAP7_75t_L         g22162(.A(new_n22418), .Y(new_n22419));
  AND2x2_ASAP7_75t_L        g22163(.A(new_n22419), .B(new_n22417), .Y(new_n22420));
  INVx1_ASAP7_75t_L         g22164(.A(new_n22420), .Y(new_n22421));
  O2A1O1Ixp33_ASAP7_75t_L   g22165(.A1(new_n22293), .A2(new_n22306), .B(new_n22299), .C(new_n22421), .Y(new_n22422));
  NOR3xp33_ASAP7_75t_L      g22166(.A(new_n22300), .B(new_n22420), .C(new_n22294), .Y(new_n22423));
  NOR2xp33_ASAP7_75t_L      g22167(.A(new_n22422), .B(new_n22423), .Y(\f[106] ));
  INVx1_ASAP7_75t_L         g22168(.A(new_n22294), .Y(new_n22425));
  A2O1A1Ixp33_ASAP7_75t_L   g22169(.A1(new_n22299), .A2(new_n22425), .B(new_n22421), .C(new_n22419), .Y(new_n22426));
  A2O1A1O1Ixp25_ASAP7_75t_L g22170(.A1(new_n12603), .A2(new_n14444), .B(new_n6443), .C(new_n6741), .D(new_n12956), .Y(new_n22427));
  NOR2xp33_ASAP7_75t_L      g22171(.A(new_n12956), .B(new_n6741), .Y(new_n22428));
  A2O1A1Ixp33_ASAP7_75t_L   g22172(.A1(new_n12986), .A2(new_n6450), .B(new_n22428), .C(\a[44] ), .Y(new_n22429));
  A2O1A1O1Ixp25_ASAP7_75t_L g22173(.A1(new_n6450), .A2(new_n14172), .B(new_n6742), .C(\b[63] ), .D(new_n6439), .Y(new_n22430));
  INVx1_ASAP7_75t_L         g22174(.A(new_n22258), .Y(new_n22431));
  A2O1A1O1Ixp25_ASAP7_75t_L g22175(.A1(new_n22183), .A2(\a[50] ), .B(new_n22184), .C(new_n22255), .D(new_n22431), .Y(new_n22432));
  A2O1A1O1Ixp25_ASAP7_75t_L g22176(.A1(new_n12986), .A2(new_n6450), .B(new_n22428), .C(new_n22429), .D(new_n22430), .Y(new_n22433));
  O2A1O1Ixp33_ASAP7_75t_L   g22177(.A1(new_n22432), .A2(new_n22396), .B(new_n22400), .C(new_n22433), .Y(new_n22434));
  INVx1_ASAP7_75t_L         g22178(.A(new_n22434), .Y(new_n22435));
  O2A1O1Ixp33_ASAP7_75t_L   g22179(.A1(new_n22432), .A2(new_n22396), .B(new_n22400), .C(new_n22434), .Y(new_n22436));
  A2O1A1O1Ixp25_ASAP7_75t_L g22180(.A1(new_n22429), .A2(new_n22427), .B(new_n22430), .C(new_n22435), .D(new_n22436), .Y(new_n22437));
  INVx1_ASAP7_75t_L         g22181(.A(new_n22437), .Y(new_n22438));
  NOR2xp33_ASAP7_75t_L      g22182(.A(new_n10309), .B(new_n10400), .Y(new_n22439));
  AOI221xp5_ASAP7_75t_L     g22183(.A1(new_n9102), .A2(\b[56] ), .B1(new_n10398), .B2(\b[54] ), .C(new_n22439), .Y(new_n22440));
  O2A1O1Ixp33_ASAP7_75t_L   g22184(.A1(new_n9104), .A2(new_n10339), .B(new_n22440), .C(new_n9099), .Y(new_n22441));
  INVx1_ASAP7_75t_L         g22185(.A(new_n22441), .Y(new_n22442));
  O2A1O1Ixp33_ASAP7_75t_L   g22186(.A1(new_n9104), .A2(new_n10339), .B(new_n22440), .C(\a[53] ), .Y(new_n22443));
  NOR2xp33_ASAP7_75t_L      g22187(.A(new_n9355), .B(new_n10388), .Y(new_n22444));
  AOI221xp5_ASAP7_75t_L     g22188(.A1(new_n10086), .A2(\b[53] ), .B1(new_n11361), .B2(\b[51] ), .C(new_n22444), .Y(new_n22445));
  O2A1O1Ixp33_ASAP7_75t_L   g22189(.A1(new_n10088), .A2(new_n9691), .B(new_n22445), .C(new_n10083), .Y(new_n22446));
  INVx1_ASAP7_75t_L         g22190(.A(new_n22446), .Y(new_n22447));
  O2A1O1Ixp33_ASAP7_75t_L   g22191(.A1(new_n10088), .A2(new_n9691), .B(new_n22445), .C(\a[56] ), .Y(new_n22448));
  INVx1_ASAP7_75t_L         g22192(.A(new_n22339), .Y(new_n22449));
  INVx1_ASAP7_75t_L         g22193(.A(new_n22347), .Y(new_n22450));
  O2A1O1Ixp33_ASAP7_75t_L   g22194(.A1(new_n22327), .A2(new_n22328), .B(new_n22332), .C(new_n22321), .Y(new_n22451));
  NAND2xp33_ASAP7_75t_L     g22195(.A(\b[43] ), .B(new_n13029), .Y(new_n22452));
  O2A1O1Ixp33_ASAP7_75t_L   g22196(.A1(new_n12672), .A2(new_n6944), .B(new_n22452), .C(new_n22319), .Y(new_n22453));
  INVx1_ASAP7_75t_L         g22197(.A(new_n22317), .Y(new_n22454));
  A2O1A1Ixp33_ASAP7_75t_L   g22198(.A1(new_n12685), .A2(new_n12686), .B(new_n6944), .C(new_n22452), .Y(new_n22455));
  O2A1O1Ixp33_ASAP7_75t_L   g22199(.A1(new_n6671), .A2(new_n12672), .B(new_n22454), .C(new_n22455), .Y(new_n22456));
  NOR2xp33_ASAP7_75t_L      g22200(.A(new_n22456), .B(new_n22453), .Y(new_n22457));
  INVx1_ASAP7_75t_L         g22201(.A(new_n22457), .Y(new_n22458));
  NAND2xp33_ASAP7_75t_L     g22202(.A(\b[47] ), .B(new_n11995), .Y(new_n22459));
  OAI221xp5_ASAP7_75t_L     g22203(.A1(new_n12318), .A2(new_n7270), .B1(new_n7249), .B2(new_n12320), .C(new_n22459), .Y(new_n22460));
  AOI21xp33_ASAP7_75t_L     g22204(.A1(new_n8726), .A2(new_n11997), .B(new_n22460), .Y(new_n22461));
  NAND2xp33_ASAP7_75t_L     g22205(.A(\a[62] ), .B(new_n22461), .Y(new_n22462));
  A2O1A1Ixp33_ASAP7_75t_L   g22206(.A1(new_n8726), .A2(new_n11997), .B(new_n22460), .C(new_n11987), .Y(new_n22463));
  AOI21xp33_ASAP7_75t_L     g22207(.A1(new_n22462), .A2(new_n22463), .B(new_n22458), .Y(new_n22464));
  NAND2xp33_ASAP7_75t_L     g22208(.A(new_n22463), .B(new_n22462), .Y(new_n22465));
  NOR2xp33_ASAP7_75t_L      g22209(.A(new_n22457), .B(new_n22465), .Y(new_n22466));
  NOR2xp33_ASAP7_75t_L      g22210(.A(new_n22464), .B(new_n22466), .Y(new_n22467));
  INVx1_ASAP7_75t_L         g22211(.A(new_n22467), .Y(new_n22468));
  O2A1O1Ixp33_ASAP7_75t_L   g22212(.A1(new_n22319), .A2(new_n22316), .B(new_n22331), .C(new_n22468), .Y(new_n22469));
  NOR2xp33_ASAP7_75t_L      g22213(.A(new_n7860), .B(new_n11354), .Y(new_n22470));
  AOI221xp5_ASAP7_75t_L     g22214(.A1(\b[50] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[49] ), .C(new_n22470), .Y(new_n22471));
  O2A1O1Ixp33_ASAP7_75t_L   g22215(.A1(new_n11053), .A2(new_n8764), .B(new_n22471), .C(new_n11048), .Y(new_n22472));
  NOR2xp33_ASAP7_75t_L      g22216(.A(new_n11048), .B(new_n22472), .Y(new_n22473));
  O2A1O1Ixp33_ASAP7_75t_L   g22217(.A1(new_n11053), .A2(new_n8764), .B(new_n22471), .C(\a[59] ), .Y(new_n22474));
  NOR2xp33_ASAP7_75t_L      g22218(.A(new_n22474), .B(new_n22473), .Y(new_n22475));
  INVx1_ASAP7_75t_L         g22219(.A(new_n22475), .Y(new_n22476));
  INVx1_ASAP7_75t_L         g22220(.A(new_n22469), .Y(new_n22477));
  O2A1O1Ixp33_ASAP7_75t_L   g22221(.A1(new_n22319), .A2(new_n22316), .B(new_n22331), .C(new_n22467), .Y(new_n22478));
  A2O1A1Ixp33_ASAP7_75t_L   g22222(.A1(new_n22477), .A2(new_n22467), .B(new_n22478), .C(new_n22476), .Y(new_n22479));
  INVx1_ASAP7_75t_L         g22223(.A(new_n22479), .Y(new_n22480));
  AOI21xp33_ASAP7_75t_L     g22224(.A1(new_n22467), .A2(new_n22451), .B(new_n22476), .Y(new_n22481));
  O2A1O1Ixp33_ASAP7_75t_L   g22225(.A1(new_n22469), .A2(new_n22451), .B(new_n22481), .C(new_n22480), .Y(new_n22482));
  A2O1A1Ixp33_ASAP7_75t_L   g22226(.A1(new_n22334), .A2(new_n22449), .B(new_n22450), .C(new_n22482), .Y(new_n22483));
  INVx1_ASAP7_75t_L         g22227(.A(new_n22483), .Y(new_n22484));
  A2O1A1O1Ixp25_ASAP7_75t_L g22228(.A1(new_n22345), .A2(\a[59] ), .B(new_n22346), .C(new_n22340), .D(new_n22336), .Y(new_n22485));
  NAND2xp33_ASAP7_75t_L     g22229(.A(new_n22485), .B(new_n22482), .Y(new_n22486));
  A2O1A1Ixp33_ASAP7_75t_L   g22230(.A1(new_n22347), .A2(new_n22337), .B(new_n22484), .C(new_n22486), .Y(new_n22487));
  AOI21xp33_ASAP7_75t_L     g22231(.A1(new_n22447), .A2(\a[56] ), .B(new_n22448), .Y(new_n22488));
  NAND2xp33_ASAP7_75t_L     g22232(.A(new_n22488), .B(new_n22486), .Y(new_n22489));
  O2A1O1Ixp33_ASAP7_75t_L   g22233(.A1(new_n22336), .A2(new_n22450), .B(new_n22483), .C(new_n22489), .Y(new_n22490));
  A2O1A1O1Ixp25_ASAP7_75t_L g22234(.A1(new_n22447), .A2(\a[56] ), .B(new_n22448), .C(new_n22487), .D(new_n22490), .Y(new_n22491));
  INVx1_ASAP7_75t_L         g22235(.A(new_n22491), .Y(new_n22492));
  A2O1A1O1Ixp25_ASAP7_75t_L g22236(.A1(new_n22314), .A2(new_n22217), .B(new_n22350), .C(new_n22361), .D(new_n22492), .Y(new_n22493));
  INVx1_ASAP7_75t_L         g22237(.A(new_n22493), .Y(new_n22494));
  NAND2xp33_ASAP7_75t_L     g22238(.A(new_n22491), .B(new_n22494), .Y(new_n22495));
  A2O1A1Ixp33_ASAP7_75t_L   g22239(.A1(new_n22361), .A2(new_n22353), .B(new_n22493), .C(new_n22495), .Y(new_n22496));
  A2O1A1Ixp33_ASAP7_75t_L   g22240(.A1(new_n22314), .A2(new_n22217), .B(new_n22350), .C(new_n22361), .Y(new_n22497));
  O2A1O1Ixp33_ASAP7_75t_L   g22241(.A1(new_n22485), .A2(new_n22484), .B(new_n22486), .C(new_n22488), .Y(new_n22498));
  AOI21xp33_ASAP7_75t_L     g22242(.A1(new_n22442), .A2(\a[53] ), .B(new_n22443), .Y(new_n22499));
  NAND2xp33_ASAP7_75t_L     g22243(.A(new_n22499), .B(new_n22495), .Y(new_n22500));
  O2A1O1Ixp33_ASAP7_75t_L   g22244(.A1(new_n22498), .A2(new_n22490), .B(new_n22497), .C(new_n22500), .Y(new_n22501));
  A2O1A1O1Ixp25_ASAP7_75t_L g22245(.A1(new_n22442), .A2(\a[53] ), .B(new_n22443), .C(new_n22496), .D(new_n22501), .Y(new_n22502));
  INVx1_ASAP7_75t_L         g22246(.A(new_n22502), .Y(new_n22503));
  O2A1O1Ixp33_ASAP7_75t_L   g22247(.A1(new_n22368), .A2(new_n22365), .B(new_n22376), .C(new_n22503), .Y(new_n22504));
  A2O1A1O1Ixp25_ASAP7_75t_L g22248(.A1(new_n22374), .A2(\a[53] ), .B(new_n22375), .C(new_n22370), .D(new_n22369), .Y(new_n22505));
  INVx1_ASAP7_75t_L         g22249(.A(new_n22505), .Y(new_n22506));
  A2O1A1O1Ixp25_ASAP7_75t_L g22250(.A1(new_n22314), .A2(new_n22217), .B(new_n22350), .C(new_n22361), .D(new_n22491), .Y(new_n22507));
  INVx1_ASAP7_75t_L         g22251(.A(new_n22507), .Y(new_n22508));
  O2A1O1Ixp33_ASAP7_75t_L   g22252(.A1(new_n22492), .A2(new_n22493), .B(new_n22508), .C(new_n22499), .Y(new_n22509));
  INVx1_ASAP7_75t_L         g22253(.A(new_n22509), .Y(new_n22510));
  O2A1O1Ixp33_ASAP7_75t_L   g22254(.A1(new_n22500), .A2(new_n22507), .B(new_n22510), .C(new_n22506), .Y(new_n22511));
  NOR2xp33_ASAP7_75t_L      g22255(.A(new_n22511), .B(new_n22504), .Y(new_n22512));
  NOR2xp33_ASAP7_75t_L      g22256(.A(new_n11303), .B(new_n10065), .Y(new_n22513));
  AOI221xp5_ASAP7_75t_L     g22257(.A1(new_n8175), .A2(\b[59] ), .B1(new_n8484), .B2(\b[57] ), .C(new_n22513), .Y(new_n22514));
  INVx1_ASAP7_75t_L         g22258(.A(new_n22514), .Y(new_n22515));
  A2O1A1Ixp33_ASAP7_75t_L   g22259(.A1(new_n12577), .A2(new_n8490), .B(new_n22515), .C(\a[50] ), .Y(new_n22516));
  O2A1O1Ixp33_ASAP7_75t_L   g22260(.A1(new_n8176), .A2(new_n11597), .B(new_n22514), .C(\a[50] ), .Y(new_n22517));
  A2O1A1Ixp33_ASAP7_75t_L   g22261(.A1(\a[50] ), .A2(new_n22516), .B(new_n22517), .C(new_n22512), .Y(new_n22518));
  NAND2xp33_ASAP7_75t_L     g22262(.A(new_n22512), .B(new_n22518), .Y(new_n22519));
  A2O1A1Ixp33_ASAP7_75t_L   g22263(.A1(new_n22516), .A2(\a[50] ), .B(new_n22517), .C(new_n22518), .Y(new_n22520));
  AND2x2_ASAP7_75t_L        g22264(.A(new_n22519), .B(new_n22520), .Y(new_n22521));
  INVx1_ASAP7_75t_L         g22265(.A(new_n22521), .Y(new_n22522));
  O2A1O1Ixp33_ASAP7_75t_L   g22266(.A1(new_n22381), .A2(new_n22379), .B(new_n22394), .C(new_n22521), .Y(new_n22523));
  INVx1_ASAP7_75t_L         g22267(.A(new_n22523), .Y(new_n22524));
  O2A1O1Ixp33_ASAP7_75t_L   g22268(.A1(new_n22381), .A2(new_n22379), .B(new_n22394), .C(new_n22522), .Y(new_n22525));
  INVx1_ASAP7_75t_L         g22269(.A(new_n22525), .Y(new_n22526));
  A2O1A1Ixp33_ASAP7_75t_L   g22270(.A1(new_n22520), .A2(new_n22519), .B(new_n22523), .C(new_n22526), .Y(new_n22527));
  NOR2xp33_ASAP7_75t_L      g22271(.A(new_n12258), .B(new_n7312), .Y(new_n22528));
  AOI221xp5_ASAP7_75t_L     g22272(.A1(\b[60] ), .A2(new_n7609), .B1(\b[62] ), .B2(new_n7334), .C(new_n22528), .Y(new_n22529));
  O2A1O1Ixp33_ASAP7_75t_L   g22273(.A1(new_n7321), .A2(new_n12610), .B(new_n22529), .C(new_n7316), .Y(new_n22530));
  INVx1_ASAP7_75t_L         g22274(.A(new_n22530), .Y(new_n22531));
  O2A1O1Ixp33_ASAP7_75t_L   g22275(.A1(new_n7321), .A2(new_n12610), .B(new_n22529), .C(\a[47] ), .Y(new_n22532));
  A2O1A1Ixp33_ASAP7_75t_L   g22276(.A1(\a[47] ), .A2(new_n22531), .B(new_n22532), .C(new_n22527), .Y(new_n22533));
  INVx1_ASAP7_75t_L         g22277(.A(new_n22532), .Y(new_n22534));
  O2A1O1Ixp33_ASAP7_75t_L   g22278(.A1(new_n22530), .A2(new_n7316), .B(new_n22534), .C(new_n22527), .Y(new_n22535));
  A2O1A1O1Ixp25_ASAP7_75t_L g22279(.A1(new_n22524), .A2(new_n22522), .B(new_n22525), .C(new_n22533), .D(new_n22535), .Y(new_n22536));
  NAND2xp33_ASAP7_75t_L     g22280(.A(new_n22536), .B(new_n22438), .Y(new_n22537));
  A2O1A1Ixp33_ASAP7_75t_L   g22281(.A1(new_n22527), .A2(new_n22533), .B(new_n22535), .C(new_n22437), .Y(new_n22538));
  AND2x2_ASAP7_75t_L        g22282(.A(new_n22538), .B(new_n22537), .Y(new_n22539));
  A2O1A1O1Ixp25_ASAP7_75t_L g22283(.A1(new_n22276), .A2(new_n22270), .B(new_n22410), .C(new_n22414), .D(new_n22539), .Y(new_n22540));
  A2O1A1O1Ixp25_ASAP7_75t_L g22284(.A1(new_n22138), .A2(new_n22149), .B(new_n22272), .C(new_n22270), .D(new_n22410), .Y(new_n22541));
  A2O1A1O1Ixp25_ASAP7_75t_L g22285(.A1(new_n22400), .A2(new_n22312), .B(new_n22402), .C(new_n22411), .D(new_n22541), .Y(new_n22542));
  AND2x2_ASAP7_75t_L        g22286(.A(new_n22539), .B(new_n22542), .Y(new_n22543));
  NOR2xp33_ASAP7_75t_L      g22287(.A(new_n22543), .B(new_n22540), .Y(new_n22544));
  XOR2x2_ASAP7_75t_L        g22288(.A(new_n22544), .B(new_n22426), .Y(\f[107] ));
  O2A1O1Ixp33_ASAP7_75t_L   g22289(.A1(new_n22418), .A2(new_n22422), .B(new_n22544), .C(new_n22540), .Y(new_n22546));
  O2A1O1Ixp33_ASAP7_75t_L   g22290(.A1(new_n22399), .A2(new_n22395), .B(new_n22312), .C(new_n22397), .Y(new_n22547));
  NOR2xp33_ASAP7_75t_L      g22291(.A(new_n11591), .B(new_n10065), .Y(new_n22548));
  AOI221xp5_ASAP7_75t_L     g22292(.A1(new_n8175), .A2(\b[60] ), .B1(new_n8484), .B2(\b[58] ), .C(new_n22548), .Y(new_n22549));
  O2A1O1Ixp33_ASAP7_75t_L   g22293(.A1(new_n8176), .A2(new_n11634), .B(new_n22549), .C(new_n8172), .Y(new_n22550));
  INVx1_ASAP7_75t_L         g22294(.A(new_n22550), .Y(new_n22551));
  O2A1O1Ixp33_ASAP7_75t_L   g22295(.A1(new_n8176), .A2(new_n11634), .B(new_n22549), .C(\a[50] ), .Y(new_n22552));
  AO21x2_ASAP7_75t_L        g22296(.A1(\a[50] ), .A2(new_n22551), .B(new_n22552), .Y(new_n22553));
  NOR2xp33_ASAP7_75t_L      g22297(.A(new_n10332), .B(new_n10400), .Y(new_n22554));
  AOI221xp5_ASAP7_75t_L     g22298(.A1(new_n9102), .A2(\b[57] ), .B1(new_n10398), .B2(\b[55] ), .C(new_n22554), .Y(new_n22555));
  O2A1O1Ixp33_ASAP7_75t_L   g22299(.A1(new_n9104), .A2(new_n17096), .B(new_n22555), .C(new_n9099), .Y(new_n22556));
  INVx1_ASAP7_75t_L         g22300(.A(new_n22556), .Y(new_n22557));
  O2A1O1Ixp33_ASAP7_75t_L   g22301(.A1(new_n9104), .A2(new_n17096), .B(new_n22555), .C(\a[53] ), .Y(new_n22558));
  AOI21xp33_ASAP7_75t_L     g22302(.A1(new_n22557), .A2(\a[53] ), .B(new_n22558), .Y(new_n22559));
  INVx1_ASAP7_75t_L         g22303(.A(new_n22559), .Y(new_n22560));
  NOR2xp33_ASAP7_75t_L      g22304(.A(new_n9683), .B(new_n10388), .Y(new_n22561));
  AOI221xp5_ASAP7_75t_L     g22305(.A1(new_n10086), .A2(\b[54] ), .B1(new_n11361), .B2(\b[52] ), .C(new_n22561), .Y(new_n22562));
  O2A1O1Ixp33_ASAP7_75t_L   g22306(.A1(new_n10088), .A2(new_n9718), .B(new_n22562), .C(new_n10083), .Y(new_n22563));
  O2A1O1Ixp33_ASAP7_75t_L   g22307(.A1(new_n10088), .A2(new_n9718), .B(new_n22562), .C(\a[56] ), .Y(new_n22564));
  INVx1_ASAP7_75t_L         g22308(.A(new_n22564), .Y(new_n22565));
  INVx1_ASAP7_75t_L         g22309(.A(new_n22453), .Y(new_n22566));
  NOR2xp33_ASAP7_75t_L      g22310(.A(new_n6944), .B(new_n13030), .Y(new_n22567));
  A2O1A1Ixp33_ASAP7_75t_L   g22311(.A1(new_n13028), .A2(\b[45] ), .B(new_n22567), .C(new_n6439), .Y(new_n22568));
  INVx1_ASAP7_75t_L         g22312(.A(new_n22568), .Y(new_n22569));
  O2A1O1Ixp33_ASAP7_75t_L   g22313(.A1(new_n12669), .A2(new_n12671), .B(\b[45] ), .C(new_n22567), .Y(new_n22570));
  NAND2xp33_ASAP7_75t_L     g22314(.A(\a[44] ), .B(new_n22570), .Y(new_n22571));
  INVx1_ASAP7_75t_L         g22315(.A(new_n22571), .Y(new_n22572));
  NOR2xp33_ASAP7_75t_L      g22316(.A(new_n22569), .B(new_n22572), .Y(new_n22573));
  INVx1_ASAP7_75t_L         g22317(.A(new_n22573), .Y(new_n22574));
  O2A1O1Ixp33_ASAP7_75t_L   g22318(.A1(new_n6671), .A2(new_n12672), .B(new_n22454), .C(new_n22574), .Y(new_n22575));
  INVx1_ASAP7_75t_L         g22319(.A(new_n22575), .Y(new_n22576));
  NOR2xp33_ASAP7_75t_L      g22320(.A(new_n22319), .B(new_n22574), .Y(new_n22577));
  A2O1A1O1Ixp25_ASAP7_75t_L g22321(.A1(new_n13028), .A2(\b[43] ), .B(new_n22317), .C(new_n22576), .D(new_n22577), .Y(new_n22578));
  INVx1_ASAP7_75t_L         g22322(.A(new_n22578), .Y(new_n22579));
  A2O1A1O1Ixp25_ASAP7_75t_L g22323(.A1(new_n22463), .A2(new_n22462), .B(new_n22458), .C(new_n22566), .D(new_n22579), .Y(new_n22580));
  A2O1A1Ixp33_ASAP7_75t_L   g22324(.A1(new_n22462), .A2(new_n22463), .B(new_n22458), .C(new_n22566), .Y(new_n22581));
  A2O1A1Ixp33_ASAP7_75t_L   g22325(.A1(new_n13028), .A2(\b[43] ), .B(new_n22317), .C(new_n22574), .Y(new_n22582));
  O2A1O1Ixp33_ASAP7_75t_L   g22326(.A1(new_n22574), .A2(new_n22575), .B(new_n22582), .C(new_n22581), .Y(new_n22583));
  A2O1A1O1Ixp25_ASAP7_75t_L g22327(.A1(new_n22463), .A2(new_n22462), .B(new_n22456), .C(new_n22566), .D(new_n22578), .Y(new_n22584));
  A2O1A1Ixp33_ASAP7_75t_L   g22328(.A1(new_n22465), .A2(new_n22457), .B(new_n22453), .C(new_n22578), .Y(new_n22585));
  OAI22xp33_ASAP7_75t_L     g22329(.A1(new_n12320), .A2(new_n7270), .B1(new_n7552), .B2(new_n12318), .Y(new_n22586));
  AOI221xp5_ASAP7_75t_L     g22330(.A1(new_n11995), .A2(\b[48] ), .B1(new_n11997), .B2(new_n11656), .C(new_n22586), .Y(new_n22587));
  XNOR2x2_ASAP7_75t_L       g22331(.A(new_n11987), .B(new_n22587), .Y(new_n22588));
  O2A1O1Ixp33_ASAP7_75t_L   g22332(.A1(new_n22578), .A2(new_n22584), .B(new_n22585), .C(new_n22588), .Y(new_n22589));
  INVx1_ASAP7_75t_L         g22333(.A(new_n22589), .Y(new_n22590));
  NOR2xp33_ASAP7_75t_L      g22334(.A(new_n22588), .B(new_n22589), .Y(new_n22591));
  O2A1O1Ixp33_ASAP7_75t_L   g22335(.A1(new_n22580), .A2(new_n22583), .B(new_n22590), .C(new_n22591), .Y(new_n22592));
  NOR2xp33_ASAP7_75t_L      g22336(.A(new_n8427), .B(new_n11354), .Y(new_n22593));
  AOI221xp5_ASAP7_75t_L     g22337(.A1(\b[51] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[50] ), .C(new_n22593), .Y(new_n22594));
  O2A1O1Ixp33_ASAP7_75t_L   g22338(.A1(new_n11053), .A2(new_n8789), .B(new_n22594), .C(new_n11048), .Y(new_n22595));
  O2A1O1Ixp33_ASAP7_75t_L   g22339(.A1(new_n11053), .A2(new_n8789), .B(new_n22594), .C(\a[59] ), .Y(new_n22596));
  INVx1_ASAP7_75t_L         g22340(.A(new_n22596), .Y(new_n22597));
  OAI211xp5_ASAP7_75t_L     g22341(.A1(new_n11048), .A2(new_n22595), .B(new_n22592), .C(new_n22597), .Y(new_n22598));
  O2A1O1Ixp33_ASAP7_75t_L   g22342(.A1(new_n22595), .A2(new_n11048), .B(new_n22597), .C(new_n22592), .Y(new_n22599));
  INVx1_ASAP7_75t_L         g22343(.A(new_n22599), .Y(new_n22600));
  NAND2xp33_ASAP7_75t_L     g22344(.A(new_n22598), .B(new_n22600), .Y(new_n22601));
  O2A1O1Ixp33_ASAP7_75t_L   g22345(.A1(new_n22451), .A2(new_n22468), .B(new_n22479), .C(new_n22601), .Y(new_n22602));
  AOI211xp5_ASAP7_75t_L     g22346(.A1(new_n22600), .A2(new_n22598), .B(new_n22469), .C(new_n22480), .Y(new_n22603));
  NOR2xp33_ASAP7_75t_L      g22347(.A(new_n22603), .B(new_n22602), .Y(new_n22604));
  INVx1_ASAP7_75t_L         g22348(.A(new_n22604), .Y(new_n22605));
  OAI211xp5_ASAP7_75t_L     g22349(.A1(new_n10083), .A2(new_n22563), .B(new_n22605), .C(new_n22565), .Y(new_n22606));
  O2A1O1Ixp33_ASAP7_75t_L   g22350(.A1(new_n10083), .A2(new_n22563), .B(new_n22565), .C(new_n22605), .Y(new_n22607));
  INVx1_ASAP7_75t_L         g22351(.A(new_n22607), .Y(new_n22608));
  NAND2xp33_ASAP7_75t_L     g22352(.A(new_n22606), .B(new_n22608), .Y(new_n22609));
  A2O1A1O1Ixp25_ASAP7_75t_L g22353(.A1(new_n22486), .A2(new_n22485), .B(new_n22488), .C(new_n22483), .D(new_n22609), .Y(new_n22610));
  INVx1_ASAP7_75t_L         g22354(.A(new_n22610), .Y(new_n22611));
  A2O1A1O1Ixp25_ASAP7_75t_L g22355(.A1(new_n22447), .A2(\a[56] ), .B(new_n22448), .C(new_n22487), .D(new_n22484), .Y(new_n22612));
  NAND2xp33_ASAP7_75t_L     g22356(.A(new_n22612), .B(new_n22609), .Y(new_n22613));
  AO21x2_ASAP7_75t_L        g22357(.A1(new_n22613), .A2(new_n22611), .B(new_n22560), .Y(new_n22614));
  AND2x2_ASAP7_75t_L        g22358(.A(new_n22613), .B(new_n22611), .Y(new_n22615));
  A2O1A1Ixp33_ASAP7_75t_L   g22359(.A1(new_n22557), .A2(\a[53] ), .B(new_n22558), .C(new_n22615), .Y(new_n22616));
  AND2x2_ASAP7_75t_L        g22360(.A(new_n22614), .B(new_n22616), .Y(new_n22617));
  INVx1_ASAP7_75t_L         g22361(.A(new_n22617), .Y(new_n22618));
  A2O1A1O1Ixp25_ASAP7_75t_L g22362(.A1(new_n22508), .A2(new_n22492), .B(new_n22499), .C(new_n22494), .D(new_n22618), .Y(new_n22619));
  NOR3xp33_ASAP7_75t_L      g22363(.A(new_n22617), .B(new_n22509), .C(new_n22493), .Y(new_n22620));
  NOR2xp33_ASAP7_75t_L      g22364(.A(new_n22620), .B(new_n22619), .Y(new_n22621));
  XOR2x2_ASAP7_75t_L        g22365(.A(new_n22553), .B(new_n22621), .Y(new_n22622));
  INVx1_ASAP7_75t_L         g22366(.A(new_n22622), .Y(new_n22623));
  O2A1O1Ixp33_ASAP7_75t_L   g22367(.A1(new_n22505), .A2(new_n22503), .B(new_n22518), .C(new_n22623), .Y(new_n22624));
  INVx1_ASAP7_75t_L         g22368(.A(new_n22624), .Y(new_n22625));
  A2O1A1O1Ixp25_ASAP7_75t_L g22369(.A1(new_n22516), .A2(\a[50] ), .B(new_n22517), .C(new_n22512), .D(new_n22504), .Y(new_n22626));
  NAND2xp33_ASAP7_75t_L     g22370(.A(new_n22626), .B(new_n22623), .Y(new_n22627));
  AND2x2_ASAP7_75t_L        g22371(.A(new_n22627), .B(new_n22625), .Y(new_n22628));
  NOR2xp33_ASAP7_75t_L      g22372(.A(new_n12603), .B(new_n7312), .Y(new_n22629));
  AOI221xp5_ASAP7_75t_L     g22373(.A1(\b[61] ), .A2(new_n7609), .B1(\b[63] ), .B2(new_n7334), .C(new_n22629), .Y(new_n22630));
  O2A1O1Ixp33_ASAP7_75t_L   g22374(.A1(new_n7321), .A2(new_n17815), .B(new_n22630), .C(new_n7316), .Y(new_n22631));
  INVx1_ASAP7_75t_L         g22375(.A(new_n22631), .Y(new_n22632));
  O2A1O1Ixp33_ASAP7_75t_L   g22376(.A1(new_n7321), .A2(new_n17815), .B(new_n22630), .C(\a[47] ), .Y(new_n22633));
  A2O1A1Ixp33_ASAP7_75t_L   g22377(.A1(\a[47] ), .A2(new_n22632), .B(new_n22633), .C(new_n22628), .Y(new_n22634));
  INVx1_ASAP7_75t_L         g22378(.A(new_n22633), .Y(new_n22635));
  O2A1O1Ixp33_ASAP7_75t_L   g22379(.A1(new_n22631), .A2(new_n7316), .B(new_n22635), .C(new_n22628), .Y(new_n22636));
  AOI21xp33_ASAP7_75t_L     g22380(.A1(new_n22634), .A2(new_n22628), .B(new_n22636), .Y(new_n22637));
  AND3x1_ASAP7_75t_L        g22381(.A(new_n22533), .B(new_n22637), .C(new_n22524), .Y(new_n22638));
  O2A1O1Ixp33_ASAP7_75t_L   g22382(.A1(new_n22252), .A2(new_n22249), .B(new_n22247), .C(new_n22379), .Y(new_n22639));
  A2O1A1O1Ixp25_ASAP7_75t_L g22383(.A1(new_n22388), .A2(\a[50] ), .B(new_n22389), .C(new_n22384), .D(new_n22639), .Y(new_n22640));
  O2A1O1Ixp33_ASAP7_75t_L   g22384(.A1(new_n22521), .A2(new_n22640), .B(new_n22533), .C(new_n22637), .Y(new_n22641));
  NOR2xp33_ASAP7_75t_L      g22385(.A(new_n22641), .B(new_n22638), .Y(new_n22642));
  INVx1_ASAP7_75t_L         g22386(.A(new_n22642), .Y(new_n22643));
  A2O1A1Ixp33_ASAP7_75t_L   g22387(.A1(new_n22527), .A2(new_n22533), .B(new_n22535), .C(new_n22438), .Y(new_n22644));
  O2A1O1Ixp33_ASAP7_75t_L   g22388(.A1(new_n22433), .A2(new_n22547), .B(new_n22644), .C(new_n22643), .Y(new_n22645));
  A2O1A1Ixp33_ASAP7_75t_L   g22389(.A1(new_n22427), .A2(new_n22429), .B(new_n22430), .C(new_n22547), .Y(new_n22646));
  O2A1O1Ixp33_ASAP7_75t_L   g22390(.A1(new_n22547), .A2(new_n22434), .B(new_n22646), .C(new_n22536), .Y(new_n22647));
  NOR3xp33_ASAP7_75t_L      g22391(.A(new_n22647), .B(new_n22642), .C(new_n22434), .Y(new_n22648));
  NOR2xp33_ASAP7_75t_L      g22392(.A(new_n22648), .B(new_n22645), .Y(new_n22649));
  XNOR2x2_ASAP7_75t_L       g22393(.A(new_n22649), .B(new_n22546), .Y(\f[108] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g22394(.A1(new_n22533), .A2(new_n22527), .B(new_n22535), .C(new_n22438), .D(new_n22434), .Y(new_n22651));
  A2O1A1Ixp33_ASAP7_75t_L   g22395(.A1(new_n22426), .A2(new_n22544), .B(new_n22540), .C(new_n22649), .Y(new_n22652));
  NOR2xp33_ASAP7_75t_L      g22396(.A(new_n11626), .B(new_n10065), .Y(new_n22653));
  AOI221xp5_ASAP7_75t_L     g22397(.A1(new_n8175), .A2(\b[61] ), .B1(new_n8484), .B2(\b[59] ), .C(new_n22653), .Y(new_n22654));
  O2A1O1Ixp33_ASAP7_75t_L   g22398(.A1(new_n8176), .A2(new_n14764), .B(new_n22654), .C(new_n8172), .Y(new_n22655));
  INVx1_ASAP7_75t_L         g22399(.A(new_n22655), .Y(new_n22656));
  O2A1O1Ixp33_ASAP7_75t_L   g22400(.A1(new_n8176), .A2(new_n14764), .B(new_n22654), .C(\a[50] ), .Y(new_n22657));
  AOI21xp33_ASAP7_75t_L     g22401(.A1(new_n22656), .A2(\a[50] ), .B(new_n22657), .Y(new_n22658));
  O2A1O1Ixp33_ASAP7_75t_L   g22402(.A1(new_n22484), .A2(new_n22498), .B(new_n22606), .C(new_n22607), .Y(new_n22659));
  O2A1O1Ixp33_ASAP7_75t_L   g22403(.A1(new_n22478), .A2(new_n22467), .B(new_n22476), .C(new_n22469), .Y(new_n22660));
  NOR2xp33_ASAP7_75t_L      g22404(.A(new_n8755), .B(new_n11354), .Y(new_n22661));
  AOI221xp5_ASAP7_75t_L     g22405(.A1(\b[52] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[51] ), .C(new_n22661), .Y(new_n22662));
  O2A1O1Ixp33_ASAP7_75t_L   g22406(.A1(new_n11053), .A2(new_n17363), .B(new_n22662), .C(new_n11048), .Y(new_n22663));
  INVx1_ASAP7_75t_L         g22407(.A(new_n22663), .Y(new_n22664));
  O2A1O1Ixp33_ASAP7_75t_L   g22408(.A1(new_n11053), .A2(new_n17363), .B(new_n22662), .C(\a[59] ), .Y(new_n22665));
  NOR2xp33_ASAP7_75t_L      g22409(.A(new_n7249), .B(new_n13030), .Y(new_n22666));
  A2O1A1O1Ixp25_ASAP7_75t_L g22410(.A1(new_n13028), .A2(\b[43] ), .B(new_n22317), .C(new_n22571), .D(new_n22569), .Y(new_n22667));
  A2O1A1Ixp33_ASAP7_75t_L   g22411(.A1(new_n13028), .A2(\b[46] ), .B(new_n22666), .C(new_n22667), .Y(new_n22668));
  O2A1O1Ixp33_ASAP7_75t_L   g22412(.A1(new_n12669), .A2(new_n12671), .B(\b[46] ), .C(new_n22666), .Y(new_n22669));
  INVx1_ASAP7_75t_L         g22413(.A(new_n22669), .Y(new_n22670));
  O2A1O1Ixp33_ASAP7_75t_L   g22414(.A1(new_n22318), .A2(new_n22572), .B(new_n22568), .C(new_n22670), .Y(new_n22671));
  INVx1_ASAP7_75t_L         g22415(.A(new_n22671), .Y(new_n22672));
  NAND2xp33_ASAP7_75t_L     g22416(.A(new_n22668), .B(new_n22672), .Y(new_n22673));
  INVx1_ASAP7_75t_L         g22417(.A(new_n22673), .Y(new_n22674));
  NOR2xp33_ASAP7_75t_L      g22418(.A(new_n7860), .B(new_n12318), .Y(new_n22675));
  AOI221xp5_ASAP7_75t_L     g22419(.A1(new_n11995), .A2(\b[49] ), .B1(new_n13314), .B2(\b[47] ), .C(new_n22675), .Y(new_n22676));
  O2A1O1Ixp33_ASAP7_75t_L   g22420(.A1(new_n11998), .A2(new_n14802), .B(new_n22676), .C(new_n11987), .Y(new_n22677));
  INVx1_ASAP7_75t_L         g22421(.A(new_n22677), .Y(new_n22678));
  O2A1O1Ixp33_ASAP7_75t_L   g22422(.A1(new_n11998), .A2(new_n14802), .B(new_n22676), .C(\a[62] ), .Y(new_n22679));
  AOI211xp5_ASAP7_75t_L     g22423(.A1(new_n22678), .A2(\a[62] ), .B(new_n22679), .C(new_n22674), .Y(new_n22680));
  A2O1A1Ixp33_ASAP7_75t_L   g22424(.A1(new_n22678), .A2(\a[62] ), .B(new_n22679), .C(new_n22674), .Y(new_n22681));
  INVx1_ASAP7_75t_L         g22425(.A(new_n22681), .Y(new_n22682));
  NOR2xp33_ASAP7_75t_L      g22426(.A(new_n22680), .B(new_n22682), .Y(new_n22683));
  A2O1A1Ixp33_ASAP7_75t_L   g22427(.A1(new_n22579), .A2(new_n22581), .B(new_n22589), .C(new_n22683), .Y(new_n22684));
  A2O1A1Ixp33_ASAP7_75t_L   g22428(.A1(new_n22579), .A2(new_n22581), .B(new_n22589), .C(new_n22684), .Y(new_n22685));
  O2A1O1Ixp33_ASAP7_75t_L   g22429(.A1(new_n22453), .A2(new_n22464), .B(new_n22579), .C(new_n22589), .Y(new_n22686));
  NAND2xp33_ASAP7_75t_L     g22430(.A(new_n22686), .B(new_n22683), .Y(new_n22687));
  NAND2xp33_ASAP7_75t_L     g22431(.A(new_n22687), .B(new_n22685), .Y(new_n22688));
  AOI21xp33_ASAP7_75t_L     g22432(.A1(new_n22664), .A2(\a[59] ), .B(new_n22665), .Y(new_n22689));
  NAND2xp33_ASAP7_75t_L     g22433(.A(new_n22689), .B(new_n22687), .Y(new_n22690));
  O2A1O1Ixp33_ASAP7_75t_L   g22434(.A1(new_n22584), .A2(new_n22589), .B(new_n22684), .C(new_n22690), .Y(new_n22691));
  A2O1A1O1Ixp25_ASAP7_75t_L g22435(.A1(new_n22664), .A2(\a[59] ), .B(new_n22665), .C(new_n22688), .D(new_n22691), .Y(new_n22692));
  INVx1_ASAP7_75t_L         g22436(.A(new_n22692), .Y(new_n22693));
  O2A1O1Ixp33_ASAP7_75t_L   g22437(.A1(new_n22660), .A2(new_n22601), .B(new_n22600), .C(new_n22693), .Y(new_n22694));
  NOR3xp33_ASAP7_75t_L      g22438(.A(new_n22692), .B(new_n22602), .C(new_n22599), .Y(new_n22695));
  NOR2xp33_ASAP7_75t_L      g22439(.A(new_n22695), .B(new_n22694), .Y(new_n22696));
  INVx1_ASAP7_75t_L         g22440(.A(new_n22696), .Y(new_n22697));
  NOR2xp33_ASAP7_75t_L      g22441(.A(new_n9709), .B(new_n10388), .Y(new_n22698));
  AOI221xp5_ASAP7_75t_L     g22442(.A1(new_n10086), .A2(\b[55] ), .B1(new_n11361), .B2(\b[53] ), .C(new_n22698), .Y(new_n22699));
  O2A1O1Ixp33_ASAP7_75t_L   g22443(.A1(new_n10088), .A2(new_n15849), .B(new_n22699), .C(new_n10083), .Y(new_n22700));
  O2A1O1Ixp33_ASAP7_75t_L   g22444(.A1(new_n10088), .A2(new_n15849), .B(new_n22699), .C(\a[56] ), .Y(new_n22701));
  INVx1_ASAP7_75t_L         g22445(.A(new_n22701), .Y(new_n22702));
  O2A1O1Ixp33_ASAP7_75t_L   g22446(.A1(new_n22700), .A2(new_n10083), .B(new_n22702), .C(new_n22697), .Y(new_n22703));
  INVx1_ASAP7_75t_L         g22447(.A(new_n22703), .Y(new_n22704));
  O2A1O1Ixp33_ASAP7_75t_L   g22448(.A1(new_n22700), .A2(new_n10083), .B(new_n22702), .C(new_n22696), .Y(new_n22705));
  AOI211xp5_ASAP7_75t_L     g22449(.A1(new_n22704), .A2(new_n22696), .B(new_n22705), .C(new_n22659), .Y(new_n22706));
  INVx1_ASAP7_75t_L         g22450(.A(new_n22659), .Y(new_n22707));
  INVx1_ASAP7_75t_L         g22451(.A(new_n22705), .Y(new_n22708));
  O2A1O1Ixp33_ASAP7_75t_L   g22452(.A1(new_n22697), .A2(new_n22703), .B(new_n22708), .C(new_n22707), .Y(new_n22709));
  NOR2xp33_ASAP7_75t_L      g22453(.A(new_n22709), .B(new_n22706), .Y(new_n22710));
  NAND2xp33_ASAP7_75t_L     g22454(.A(\b[57] ), .B(new_n9096), .Y(new_n22711));
  OAI221xp5_ASAP7_75t_L     g22455(.A1(new_n9440), .A2(new_n10332), .B1(new_n11303), .B2(new_n9439), .C(new_n22711), .Y(new_n22712));
  A2O1A1Ixp33_ASAP7_75t_L   g22456(.A1(new_n11314), .A2(new_n9437), .B(new_n22712), .C(\a[53] ), .Y(new_n22713));
  NAND2xp33_ASAP7_75t_L     g22457(.A(\a[53] ), .B(new_n22713), .Y(new_n22714));
  A2O1A1Ixp33_ASAP7_75t_L   g22458(.A1(new_n11314), .A2(new_n9437), .B(new_n22712), .C(new_n9099), .Y(new_n22715));
  NAND2xp33_ASAP7_75t_L     g22459(.A(new_n22715), .B(new_n22714), .Y(new_n22716));
  XNOR2x2_ASAP7_75t_L       g22460(.A(new_n22716), .B(new_n22710), .Y(new_n22717));
  INVx1_ASAP7_75t_L         g22461(.A(new_n22717), .Y(new_n22718));
  A2O1A1O1Ixp25_ASAP7_75t_L g22462(.A1(new_n22442), .A2(\a[53] ), .B(new_n22443), .C(new_n22496), .D(new_n22493), .Y(new_n22719));
  O2A1O1Ixp33_ASAP7_75t_L   g22463(.A1(new_n22719), .A2(new_n22618), .B(new_n22616), .C(new_n22718), .Y(new_n22720));
  A2O1A1Ixp33_ASAP7_75t_L   g22464(.A1(new_n22615), .A2(new_n22560), .B(new_n22619), .C(new_n22718), .Y(new_n22721));
  O2A1O1Ixp33_ASAP7_75t_L   g22465(.A1(new_n22718), .A2(new_n22720), .B(new_n22721), .C(new_n22658), .Y(new_n22722));
  INVx1_ASAP7_75t_L         g22466(.A(new_n22722), .Y(new_n22723));
  O2A1O1Ixp33_ASAP7_75t_L   g22467(.A1(new_n22718), .A2(new_n22720), .B(new_n22721), .C(new_n22722), .Y(new_n22724));
  A2O1A1O1Ixp25_ASAP7_75t_L g22468(.A1(new_n22656), .A2(\a[50] ), .B(new_n22657), .C(new_n22723), .D(new_n22724), .Y(new_n22725));
  AOI22xp33_ASAP7_75t_L     g22469(.A1(new_n7333), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n7609), .Y(new_n22726));
  INVx1_ASAP7_75t_L         g22470(.A(new_n22726), .Y(new_n22727));
  A2O1A1Ixp33_ASAP7_75t_L   g22471(.A1(new_n7315), .A2(new_n7317), .B(new_n7000), .C(new_n22726), .Y(new_n22728));
  O2A1O1Ixp33_ASAP7_75t_L   g22472(.A1(new_n22727), .A2(new_n17329), .B(new_n22728), .C(new_n7316), .Y(new_n22729));
  O2A1O1Ixp33_ASAP7_75t_L   g22473(.A1(new_n7321), .A2(new_n12993), .B(new_n22726), .C(\a[47] ), .Y(new_n22730));
  NOR2xp33_ASAP7_75t_L      g22474(.A(new_n22730), .B(new_n22729), .Y(new_n22731));
  INVx1_ASAP7_75t_L         g22475(.A(new_n22731), .Y(new_n22732));
  A2O1A1Ixp33_ASAP7_75t_L   g22476(.A1(new_n22621), .A2(new_n22553), .B(new_n22624), .C(new_n22732), .Y(new_n22733));
  A2O1A1O1Ixp25_ASAP7_75t_L g22477(.A1(new_n22551), .A2(\a[50] ), .B(new_n22552), .C(new_n22621), .D(new_n22624), .Y(new_n22734));
  NAND2xp33_ASAP7_75t_L     g22478(.A(new_n22731), .B(new_n22734), .Y(new_n22735));
  NAND2xp33_ASAP7_75t_L     g22479(.A(new_n22733), .B(new_n22735), .Y(new_n22736));
  INVx1_ASAP7_75t_L         g22480(.A(new_n22724), .Y(new_n22737));
  O2A1O1Ixp33_ASAP7_75t_L   g22481(.A1(new_n22658), .A2(new_n22722), .B(new_n22737), .C(new_n22736), .Y(new_n22738));
  NAND3xp33_ASAP7_75t_L     g22482(.A(new_n22735), .B(new_n22733), .C(new_n22725), .Y(new_n22739));
  A2O1A1O1Ixp25_ASAP7_75t_L g22483(.A1(new_n22632), .A2(\a[47] ), .B(new_n22633), .C(new_n22628), .D(new_n22641), .Y(new_n22740));
  OAI211xp5_ASAP7_75t_L     g22484(.A1(new_n22725), .A2(new_n22738), .B(new_n22740), .C(new_n22739), .Y(new_n22741));
  O2A1O1Ixp33_ASAP7_75t_L   g22485(.A1(new_n22725), .A2(new_n22738), .B(new_n22739), .C(new_n22740), .Y(new_n22742));
  INVx1_ASAP7_75t_L         g22486(.A(new_n22742), .Y(new_n22743));
  AND2x2_ASAP7_75t_L        g22487(.A(new_n22741), .B(new_n22743), .Y(new_n22744));
  INVx1_ASAP7_75t_L         g22488(.A(new_n22744), .Y(new_n22745));
  O2A1O1Ixp33_ASAP7_75t_L   g22489(.A1(new_n22643), .A2(new_n22651), .B(new_n22652), .C(new_n22745), .Y(new_n22746));
  A2O1A1Ixp33_ASAP7_75t_L   g22490(.A1(new_n22644), .A2(new_n22435), .B(new_n22643), .C(new_n22652), .Y(new_n22747));
  NOR2xp33_ASAP7_75t_L      g22491(.A(new_n22744), .B(new_n22747), .Y(new_n22748));
  NOR2xp33_ASAP7_75t_L      g22492(.A(new_n22746), .B(new_n22748), .Y(\f[109] ));
  O2A1O1Ixp33_ASAP7_75t_L   g22493(.A1(new_n22469), .A2(new_n22480), .B(new_n22598), .C(new_n22599), .Y(new_n22750));
  NOR2xp33_ASAP7_75t_L      g22494(.A(new_n10309), .B(new_n10388), .Y(new_n22751));
  AOI221xp5_ASAP7_75t_L     g22495(.A1(new_n10086), .A2(\b[56] ), .B1(new_n11361), .B2(\b[54] ), .C(new_n22751), .Y(new_n22752));
  O2A1O1Ixp33_ASAP7_75t_L   g22496(.A1(new_n10088), .A2(new_n10339), .B(new_n22752), .C(new_n10083), .Y(new_n22753));
  INVx1_ASAP7_75t_L         g22497(.A(new_n22753), .Y(new_n22754));
  O2A1O1Ixp33_ASAP7_75t_L   g22498(.A1(new_n10088), .A2(new_n10339), .B(new_n22752), .C(\a[56] ), .Y(new_n22755));
  A2O1A1Ixp33_ASAP7_75t_L   g22499(.A1(new_n22687), .A2(new_n22686), .B(new_n22689), .C(new_n22684), .Y(new_n22756));
  NOR2xp33_ASAP7_75t_L      g22500(.A(new_n8779), .B(new_n11354), .Y(new_n22757));
  AOI221xp5_ASAP7_75t_L     g22501(.A1(\b[53] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[52] ), .C(new_n22757), .Y(new_n22758));
  O2A1O1Ixp33_ASAP7_75t_L   g22502(.A1(new_n11053), .A2(new_n9691), .B(new_n22758), .C(new_n11048), .Y(new_n22759));
  NOR2xp33_ASAP7_75t_L      g22503(.A(new_n11048), .B(new_n22759), .Y(new_n22760));
  O2A1O1Ixp33_ASAP7_75t_L   g22504(.A1(new_n11053), .A2(new_n9691), .B(new_n22758), .C(\a[59] ), .Y(new_n22761));
  NOR2xp33_ASAP7_75t_L      g22505(.A(new_n22761), .B(new_n22760), .Y(new_n22762));
  NOR2xp33_ASAP7_75t_L      g22506(.A(new_n7270), .B(new_n13030), .Y(new_n22763));
  INVx1_ASAP7_75t_L         g22507(.A(new_n22763), .Y(new_n22764));
  O2A1O1Ixp33_ASAP7_75t_L   g22508(.A1(new_n12672), .A2(new_n7552), .B(new_n22764), .C(new_n22670), .Y(new_n22765));
  INVx1_ASAP7_75t_L         g22509(.A(new_n22667), .Y(new_n22766));
  O2A1O1Ixp33_ASAP7_75t_L   g22510(.A1(new_n12669), .A2(new_n12671), .B(\b[47] ), .C(new_n22763), .Y(new_n22767));
  A2O1A1Ixp33_ASAP7_75t_L   g22511(.A1(new_n13028), .A2(\b[46] ), .B(new_n22666), .C(new_n22767), .Y(new_n22768));
  A2O1A1Ixp33_ASAP7_75t_L   g22512(.A1(new_n22766), .A2(new_n22669), .B(new_n22682), .C(new_n22768), .Y(new_n22769));
  A2O1A1O1Ixp25_ASAP7_75t_L g22513(.A1(new_n13028), .A2(\b[47] ), .B(new_n22763), .C(new_n22669), .D(new_n22769), .Y(new_n22770));
  O2A1O1Ixp33_ASAP7_75t_L   g22514(.A1(new_n22670), .A2(new_n22667), .B(new_n22681), .C(new_n22770), .Y(new_n22771));
  INVx1_ASAP7_75t_L         g22515(.A(new_n22771), .Y(new_n22772));
  A2O1A1O1Ixp25_ASAP7_75t_L g22516(.A1(new_n13028), .A2(\b[46] ), .B(new_n22666), .C(new_n22767), .D(new_n22770), .Y(new_n22773));
  INVx1_ASAP7_75t_L         g22517(.A(new_n22773), .Y(new_n22774));
  OAI22xp33_ASAP7_75t_L     g22518(.A1(new_n12320), .A2(new_n7860), .B1(new_n8427), .B2(new_n12318), .Y(new_n22775));
  AOI221xp5_ASAP7_75t_L     g22519(.A1(new_n11995), .A2(\b[50] ), .B1(new_n11997), .B2(new_n8763), .C(new_n22775), .Y(new_n22776));
  XNOR2x2_ASAP7_75t_L       g22520(.A(new_n11987), .B(new_n22776), .Y(new_n22777));
  INVx1_ASAP7_75t_L         g22521(.A(new_n22777), .Y(new_n22778));
  O2A1O1Ixp33_ASAP7_75t_L   g22522(.A1(new_n22765), .A2(new_n22774), .B(new_n22772), .C(new_n22778), .Y(new_n22779));
  A2O1A1O1Ixp25_ASAP7_75t_L g22523(.A1(new_n13028), .A2(\b[47] ), .B(new_n22763), .C(new_n22669), .D(new_n22774), .Y(new_n22780));
  NOR3xp33_ASAP7_75t_L      g22524(.A(new_n22780), .B(new_n22777), .C(new_n22771), .Y(new_n22781));
  NOR2xp33_ASAP7_75t_L      g22525(.A(new_n22779), .B(new_n22781), .Y(new_n22782));
  NOR2xp33_ASAP7_75t_L      g22526(.A(new_n22762), .B(new_n22782), .Y(new_n22783));
  NOR4xp25_ASAP7_75t_L      g22527(.A(new_n22781), .B(new_n22760), .C(new_n22761), .D(new_n22779), .Y(new_n22784));
  NOR2xp33_ASAP7_75t_L      g22528(.A(new_n22784), .B(new_n22783), .Y(new_n22785));
  NAND2xp33_ASAP7_75t_L     g22529(.A(new_n22756), .B(new_n22785), .Y(new_n22786));
  NAND2xp33_ASAP7_75t_L     g22530(.A(new_n22756), .B(new_n22786), .Y(new_n22787));
  NAND2xp33_ASAP7_75t_L     g22531(.A(new_n22785), .B(new_n22786), .Y(new_n22788));
  NAND2xp33_ASAP7_75t_L     g22532(.A(new_n22788), .B(new_n22787), .Y(new_n22789));
  AOI21xp33_ASAP7_75t_L     g22533(.A1(new_n22754), .A2(\a[56] ), .B(new_n22755), .Y(new_n22790));
  NAND2xp33_ASAP7_75t_L     g22534(.A(new_n22790), .B(new_n22788), .Y(new_n22791));
  O2A1O1Ixp33_ASAP7_75t_L   g22535(.A1(new_n22783), .A2(new_n22784), .B(new_n22756), .C(new_n22791), .Y(new_n22792));
  A2O1A1O1Ixp25_ASAP7_75t_L g22536(.A1(new_n22754), .A2(\a[56] ), .B(new_n22755), .C(new_n22789), .D(new_n22792), .Y(new_n22793));
  INVx1_ASAP7_75t_L         g22537(.A(new_n22793), .Y(new_n22794));
  O2A1O1Ixp33_ASAP7_75t_L   g22538(.A1(new_n22750), .A2(new_n22693), .B(new_n22704), .C(new_n22794), .Y(new_n22795));
  INVx1_ASAP7_75t_L         g22539(.A(new_n22700), .Y(new_n22796));
  A2O1A1O1Ixp25_ASAP7_75t_L g22540(.A1(new_n22796), .A2(\a[56] ), .B(new_n22701), .C(new_n22696), .D(new_n22694), .Y(new_n22797));
  INVx1_ASAP7_75t_L         g22541(.A(new_n22797), .Y(new_n22798));
  A2O1A1O1Ixp25_ASAP7_75t_L g22542(.A1(new_n22687), .A2(new_n22686), .B(new_n22689), .C(new_n22684), .D(new_n22785), .Y(new_n22799));
  A2O1A1Ixp33_ASAP7_75t_L   g22543(.A1(new_n22754), .A2(\a[56] ), .B(new_n22755), .C(new_n22789), .Y(new_n22800));
  O2A1O1Ixp33_ASAP7_75t_L   g22544(.A1(new_n22791), .A2(new_n22799), .B(new_n22800), .C(new_n22798), .Y(new_n22801));
  NOR2xp33_ASAP7_75t_L      g22545(.A(new_n22801), .B(new_n22795), .Y(new_n22802));
  INVx1_ASAP7_75t_L         g22546(.A(new_n22802), .Y(new_n22803));
  NOR2xp33_ASAP7_75t_L      g22547(.A(new_n11303), .B(new_n10400), .Y(new_n22804));
  AOI221xp5_ASAP7_75t_L     g22548(.A1(new_n9102), .A2(\b[59] ), .B1(new_n10398), .B2(\b[57] ), .C(new_n22804), .Y(new_n22805));
  O2A1O1Ixp33_ASAP7_75t_L   g22549(.A1(new_n9104), .A2(new_n11597), .B(new_n22805), .C(new_n9099), .Y(new_n22806));
  O2A1O1Ixp33_ASAP7_75t_L   g22550(.A1(new_n9104), .A2(new_n11597), .B(new_n22805), .C(\a[53] ), .Y(new_n22807));
  INVx1_ASAP7_75t_L         g22551(.A(new_n22807), .Y(new_n22808));
  O2A1O1Ixp33_ASAP7_75t_L   g22552(.A1(new_n22806), .A2(new_n9099), .B(new_n22808), .C(new_n22803), .Y(new_n22809));
  INVx1_ASAP7_75t_L         g22553(.A(new_n22809), .Y(new_n22810));
  O2A1O1Ixp33_ASAP7_75t_L   g22554(.A1(new_n22806), .A2(new_n9099), .B(new_n22808), .C(new_n22802), .Y(new_n22811));
  AOI21xp33_ASAP7_75t_L     g22555(.A1(new_n22810), .A2(new_n22802), .B(new_n22811), .Y(new_n22812));
  O2A1O1Ixp33_ASAP7_75t_L   g22556(.A1(new_n22697), .A2(new_n22703), .B(new_n22708), .C(new_n22659), .Y(new_n22813));
  INVx1_ASAP7_75t_L         g22557(.A(new_n22813), .Y(new_n22814));
  A2O1A1O1Ixp25_ASAP7_75t_L g22558(.A1(new_n22714), .A2(new_n22715), .B(new_n22710), .C(new_n22814), .D(new_n22812), .Y(new_n22815));
  INVx1_ASAP7_75t_L         g22559(.A(new_n22815), .Y(new_n22816));
  INVx1_ASAP7_75t_L         g22560(.A(new_n22812), .Y(new_n22817));
  A2O1A1O1Ixp25_ASAP7_75t_L g22561(.A1(new_n22714), .A2(new_n22715), .B(new_n22710), .C(new_n22814), .D(new_n22817), .Y(new_n22818));
  A2O1A1O1Ixp25_ASAP7_75t_L g22562(.A1(new_n22810), .A2(new_n22802), .B(new_n22811), .C(new_n22816), .D(new_n22818), .Y(new_n22819));
  INVx1_ASAP7_75t_L         g22563(.A(new_n22819), .Y(new_n22820));
  NOR2xp33_ASAP7_75t_L      g22564(.A(new_n12258), .B(new_n10065), .Y(new_n22821));
  AOI221xp5_ASAP7_75t_L     g22565(.A1(new_n8175), .A2(\b[62] ), .B1(new_n8484), .B2(\b[60] ), .C(new_n22821), .Y(new_n22822));
  O2A1O1Ixp33_ASAP7_75t_L   g22566(.A1(new_n8176), .A2(new_n12610), .B(new_n22822), .C(new_n8172), .Y(new_n22823));
  O2A1O1Ixp33_ASAP7_75t_L   g22567(.A1(new_n8176), .A2(new_n12610), .B(new_n22822), .C(\a[50] ), .Y(new_n22824));
  INVx1_ASAP7_75t_L         g22568(.A(new_n22824), .Y(new_n22825));
  O2A1O1Ixp33_ASAP7_75t_L   g22569(.A1(new_n22823), .A2(new_n8172), .B(new_n22825), .C(new_n22819), .Y(new_n22826));
  INVx1_ASAP7_75t_L         g22570(.A(new_n22826), .Y(new_n22827));
  O2A1O1Ixp33_ASAP7_75t_L   g22571(.A1(new_n22823), .A2(new_n8172), .B(new_n22825), .C(new_n22820), .Y(new_n22828));
  INVx1_ASAP7_75t_L         g22572(.A(new_n22720), .Y(new_n22829));
  NOR2xp33_ASAP7_75t_L      g22573(.A(new_n12956), .B(new_n7614), .Y(new_n22830));
  INVx1_ASAP7_75t_L         g22574(.A(new_n22830), .Y(new_n22831));
  A2O1A1Ixp33_ASAP7_75t_L   g22575(.A1(new_n14444), .A2(new_n12603), .B(new_n12956), .C(new_n22831), .Y(new_n22832));
  O2A1O1Ixp33_ASAP7_75t_L   g22576(.A1(new_n7322), .A2(new_n22830), .B(new_n22832), .C(new_n7316), .Y(new_n22833));
  O2A1O1Ixp33_ASAP7_75t_L   g22577(.A1(new_n7321), .A2(new_n13573), .B(new_n22831), .C(\a[47] ), .Y(new_n22834));
  NOR2xp33_ASAP7_75t_L      g22578(.A(new_n22834), .B(new_n22833), .Y(new_n22835));
  A2O1A1O1Ixp25_ASAP7_75t_L g22579(.A1(new_n22718), .A2(new_n22721), .B(new_n22658), .C(new_n22829), .D(new_n22835), .Y(new_n22836));
  NOR4xp25_ASAP7_75t_L      g22580(.A(new_n22722), .B(new_n22834), .C(new_n22720), .D(new_n22833), .Y(new_n22837));
  NOR2xp33_ASAP7_75t_L      g22581(.A(new_n22836), .B(new_n22837), .Y(new_n22838));
  A2O1A1Ixp33_ASAP7_75t_L   g22582(.A1(new_n22827), .A2(new_n22820), .B(new_n22828), .C(new_n22838), .Y(new_n22839));
  A2O1A1Ixp33_ASAP7_75t_L   g22583(.A1(new_n22827), .A2(new_n22820), .B(new_n22828), .C(new_n22839), .Y(new_n22840));
  A2O1A1O1Ixp25_ASAP7_75t_L g22584(.A1(new_n22816), .A2(new_n22817), .B(new_n22818), .C(new_n22827), .D(new_n22828), .Y(new_n22841));
  NAND2xp33_ASAP7_75t_L     g22585(.A(new_n22838), .B(new_n22841), .Y(new_n22842));
  A2O1A1O1Ixp25_ASAP7_75t_L g22586(.A1(new_n22621), .A2(new_n22553), .B(new_n22624), .C(new_n22732), .D(new_n22738), .Y(new_n22843));
  AND3x1_ASAP7_75t_L        g22587(.A(new_n22840), .B(new_n22843), .C(new_n22842), .Y(new_n22844));
  INVx1_ASAP7_75t_L         g22588(.A(new_n22840), .Y(new_n22845));
  INVx1_ASAP7_75t_L         g22589(.A(new_n22843), .Y(new_n22846));
  A2O1A1Ixp33_ASAP7_75t_L   g22590(.A1(new_n22839), .A2(new_n22838), .B(new_n22845), .C(new_n22846), .Y(new_n22847));
  INVx1_ASAP7_75t_L         g22591(.A(new_n22847), .Y(new_n22848));
  NOR2xp33_ASAP7_75t_L      g22592(.A(new_n22844), .B(new_n22848), .Y(new_n22849));
  INVx1_ASAP7_75t_L         g22593(.A(new_n22645), .Y(new_n22850));
  A2O1A1Ixp33_ASAP7_75t_L   g22594(.A1(new_n22652), .A2(new_n22850), .B(new_n22745), .C(new_n22743), .Y(new_n22851));
  XOR2x2_ASAP7_75t_L        g22595(.A(new_n22849), .B(new_n22851), .Y(\f[110] ));
  NOR2xp33_ASAP7_75t_L      g22596(.A(new_n12603), .B(new_n10065), .Y(new_n22853));
  AOI221xp5_ASAP7_75t_L     g22597(.A1(new_n8175), .A2(\b[63] ), .B1(new_n8484), .B2(\b[61] ), .C(new_n22853), .Y(new_n22854));
  O2A1O1Ixp33_ASAP7_75t_L   g22598(.A1(new_n8176), .A2(new_n17815), .B(new_n22854), .C(new_n8172), .Y(new_n22855));
  INVx1_ASAP7_75t_L         g22599(.A(new_n22855), .Y(new_n22856));
  O2A1O1Ixp33_ASAP7_75t_L   g22600(.A1(new_n8176), .A2(new_n17815), .B(new_n22854), .C(\a[50] ), .Y(new_n22857));
  NOR2xp33_ASAP7_75t_L      g22601(.A(new_n11591), .B(new_n10400), .Y(new_n22858));
  AOI221xp5_ASAP7_75t_L     g22602(.A1(new_n9102), .A2(\b[60] ), .B1(new_n10398), .B2(\b[58] ), .C(new_n22858), .Y(new_n22859));
  O2A1O1Ixp33_ASAP7_75t_L   g22603(.A1(new_n9104), .A2(new_n11634), .B(new_n22859), .C(new_n9099), .Y(new_n22860));
  INVx1_ASAP7_75t_L         g22604(.A(new_n22860), .Y(new_n22861));
  O2A1O1Ixp33_ASAP7_75t_L   g22605(.A1(new_n9104), .A2(new_n11634), .B(new_n22859), .C(\a[53] ), .Y(new_n22862));
  AO21x2_ASAP7_75t_L        g22606(.A1(\a[53] ), .A2(new_n22861), .B(new_n22862), .Y(new_n22863));
  NOR2xp33_ASAP7_75t_L      g22607(.A(new_n10332), .B(new_n10388), .Y(new_n22864));
  AOI221xp5_ASAP7_75t_L     g22608(.A1(new_n10086), .A2(\b[57] ), .B1(new_n11361), .B2(\b[55] ), .C(new_n22864), .Y(new_n22865));
  O2A1O1Ixp33_ASAP7_75t_L   g22609(.A1(new_n10088), .A2(new_n17096), .B(new_n22865), .C(new_n10083), .Y(new_n22866));
  INVx1_ASAP7_75t_L         g22610(.A(new_n22866), .Y(new_n22867));
  O2A1O1Ixp33_ASAP7_75t_L   g22611(.A1(new_n10088), .A2(new_n17096), .B(new_n22865), .C(\a[56] ), .Y(new_n22868));
  AOI21xp33_ASAP7_75t_L     g22612(.A1(new_n22867), .A2(\a[56] ), .B(new_n22868), .Y(new_n22869));
  INVx1_ASAP7_75t_L         g22613(.A(new_n22869), .Y(new_n22870));
  O2A1O1Ixp33_ASAP7_75t_L   g22614(.A1(new_n22765), .A2(new_n22774), .B(new_n22772), .C(new_n22777), .Y(new_n22871));
  INVx1_ASAP7_75t_L         g22615(.A(new_n22871), .Y(new_n22872));
  NOR2xp33_ASAP7_75t_L      g22616(.A(new_n7552), .B(new_n13030), .Y(new_n22873));
  O2A1O1Ixp33_ASAP7_75t_L   g22617(.A1(new_n7552), .A2(new_n12672), .B(new_n22764), .C(new_n7316), .Y(new_n22874));
  AOI211xp5_ASAP7_75t_L     g22618(.A1(new_n13028), .A2(\b[47] ), .B(new_n22763), .C(\a[47] ), .Y(new_n22875));
  NOR2xp33_ASAP7_75t_L      g22619(.A(new_n22875), .B(new_n22874), .Y(new_n22876));
  INVx1_ASAP7_75t_L         g22620(.A(new_n22876), .Y(new_n22877));
  A2O1A1Ixp33_ASAP7_75t_L   g22621(.A1(new_n13028), .A2(\b[48] ), .B(new_n22873), .C(new_n22877), .Y(new_n22878));
  O2A1O1Ixp33_ASAP7_75t_L   g22622(.A1(new_n12669), .A2(new_n12671), .B(\b[48] ), .C(new_n22873), .Y(new_n22879));
  NAND2xp33_ASAP7_75t_L     g22623(.A(new_n22879), .B(new_n22876), .Y(new_n22880));
  AND2x2_ASAP7_75t_L        g22624(.A(new_n22880), .B(new_n22878), .Y(new_n22881));
  NOR2xp33_ASAP7_75t_L      g22625(.A(new_n8755), .B(new_n12318), .Y(new_n22882));
  AOI221xp5_ASAP7_75t_L     g22626(.A1(new_n11995), .A2(\b[51] ), .B1(new_n13314), .B2(\b[49] ), .C(new_n22882), .Y(new_n22883));
  O2A1O1Ixp33_ASAP7_75t_L   g22627(.A1(new_n11998), .A2(new_n8789), .B(new_n22883), .C(new_n11987), .Y(new_n22884));
  O2A1O1Ixp33_ASAP7_75t_L   g22628(.A1(new_n11998), .A2(new_n8789), .B(new_n22883), .C(\a[62] ), .Y(new_n22885));
  INVx1_ASAP7_75t_L         g22629(.A(new_n22885), .Y(new_n22886));
  INVx1_ASAP7_75t_L         g22630(.A(new_n22881), .Y(new_n22887));
  O2A1O1Ixp33_ASAP7_75t_L   g22631(.A1(new_n11987), .A2(new_n22884), .B(new_n22886), .C(new_n22887), .Y(new_n22888));
  INVx1_ASAP7_75t_L         g22632(.A(new_n22888), .Y(new_n22889));
  O2A1O1Ixp33_ASAP7_75t_L   g22633(.A1(new_n11987), .A2(new_n22884), .B(new_n22886), .C(new_n22881), .Y(new_n22890));
  AOI21xp33_ASAP7_75t_L     g22634(.A1(new_n22889), .A2(new_n22881), .B(new_n22890), .Y(new_n22891));
  O2A1O1Ixp33_ASAP7_75t_L   g22635(.A1(new_n22765), .A2(new_n22769), .B(new_n22768), .C(new_n22891), .Y(new_n22892));
  INVx1_ASAP7_75t_L         g22636(.A(new_n22892), .Y(new_n22893));
  INVx1_ASAP7_75t_L         g22637(.A(new_n22891), .Y(new_n22894));
  O2A1O1Ixp33_ASAP7_75t_L   g22638(.A1(new_n22765), .A2(new_n22769), .B(new_n22768), .C(new_n22894), .Y(new_n22895));
  A2O1A1O1Ixp25_ASAP7_75t_L g22639(.A1(new_n22889), .A2(new_n22881), .B(new_n22890), .C(new_n22893), .D(new_n22895), .Y(new_n22896));
  NOR2xp33_ASAP7_75t_L      g22640(.A(new_n9355), .B(new_n11354), .Y(new_n22897));
  AOI221xp5_ASAP7_75t_L     g22641(.A1(\b[54] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[53] ), .C(new_n22897), .Y(new_n22898));
  O2A1O1Ixp33_ASAP7_75t_L   g22642(.A1(new_n11053), .A2(new_n9718), .B(new_n22898), .C(new_n11048), .Y(new_n22899));
  O2A1O1Ixp33_ASAP7_75t_L   g22643(.A1(new_n11053), .A2(new_n9718), .B(new_n22898), .C(\a[59] ), .Y(new_n22900));
  INVx1_ASAP7_75t_L         g22644(.A(new_n22900), .Y(new_n22901));
  OAI211xp5_ASAP7_75t_L     g22645(.A1(new_n11048), .A2(new_n22899), .B(new_n22896), .C(new_n22901), .Y(new_n22902));
  O2A1O1Ixp33_ASAP7_75t_L   g22646(.A1(new_n22899), .A2(new_n11048), .B(new_n22901), .C(new_n22896), .Y(new_n22903));
  INVx1_ASAP7_75t_L         g22647(.A(new_n22903), .Y(new_n22904));
  NAND2xp33_ASAP7_75t_L     g22648(.A(new_n22902), .B(new_n22904), .Y(new_n22905));
  O2A1O1Ixp33_ASAP7_75t_L   g22649(.A1(new_n22762), .A2(new_n22782), .B(new_n22872), .C(new_n22905), .Y(new_n22906));
  INVx1_ASAP7_75t_L         g22650(.A(new_n22906), .Y(new_n22907));
  O2A1O1Ixp33_ASAP7_75t_L   g22651(.A1(new_n22771), .A2(new_n22780), .B(new_n22778), .C(new_n22783), .Y(new_n22908));
  NAND2xp33_ASAP7_75t_L     g22652(.A(new_n22905), .B(new_n22908), .Y(new_n22909));
  AO21x2_ASAP7_75t_L        g22653(.A1(new_n22907), .A2(new_n22909), .B(new_n22870), .Y(new_n22910));
  AND2x2_ASAP7_75t_L        g22654(.A(new_n22907), .B(new_n22909), .Y(new_n22911));
  A2O1A1Ixp33_ASAP7_75t_L   g22655(.A1(new_n22867), .A2(\a[56] ), .B(new_n22868), .C(new_n22911), .Y(new_n22912));
  AND2x2_ASAP7_75t_L        g22656(.A(new_n22910), .B(new_n22912), .Y(new_n22913));
  INVx1_ASAP7_75t_L         g22657(.A(new_n22913), .Y(new_n22914));
  A2O1A1O1Ixp25_ASAP7_75t_L g22658(.A1(new_n22787), .A2(new_n22788), .B(new_n22790), .C(new_n22786), .D(new_n22914), .Y(new_n22915));
  A2O1A1Ixp33_ASAP7_75t_L   g22659(.A1(new_n22787), .A2(new_n22788), .B(new_n22790), .C(new_n22786), .Y(new_n22916));
  NOR2xp33_ASAP7_75t_L      g22660(.A(new_n22916), .B(new_n22913), .Y(new_n22917));
  NOR2xp33_ASAP7_75t_L      g22661(.A(new_n22917), .B(new_n22915), .Y(new_n22918));
  XOR2x2_ASAP7_75t_L        g22662(.A(new_n22863), .B(new_n22918), .Y(new_n22919));
  INVx1_ASAP7_75t_L         g22663(.A(new_n22919), .Y(new_n22920));
  O2A1O1Ixp33_ASAP7_75t_L   g22664(.A1(new_n22797), .A2(new_n22794), .B(new_n22810), .C(new_n22920), .Y(new_n22921));
  INVx1_ASAP7_75t_L         g22665(.A(new_n22921), .Y(new_n22922));
  O2A1O1Ixp33_ASAP7_75t_L   g22666(.A1(new_n22694), .A2(new_n22703), .B(new_n22793), .C(new_n22809), .Y(new_n22923));
  NAND2xp33_ASAP7_75t_L     g22667(.A(new_n22920), .B(new_n22923), .Y(new_n22924));
  AND2x2_ASAP7_75t_L        g22668(.A(new_n22924), .B(new_n22922), .Y(new_n22925));
  A2O1A1Ixp33_ASAP7_75t_L   g22669(.A1(\a[50] ), .A2(new_n22856), .B(new_n22857), .C(new_n22925), .Y(new_n22926));
  AND2x2_ASAP7_75t_L        g22670(.A(new_n22925), .B(new_n22926), .Y(new_n22927));
  A2O1A1O1Ixp25_ASAP7_75t_L g22671(.A1(new_n22856), .A2(\a[50] ), .B(new_n22857), .C(new_n22926), .D(new_n22927), .Y(new_n22928));
  INVx1_ASAP7_75t_L         g22672(.A(new_n22928), .Y(new_n22929));
  NOR3xp33_ASAP7_75t_L      g22673(.A(new_n22929), .B(new_n22826), .C(new_n22815), .Y(new_n22930));
  O2A1O1Ixp33_ASAP7_75t_L   g22674(.A1(new_n22709), .A2(new_n22706), .B(new_n22716), .C(new_n22813), .Y(new_n22931));
  O2A1O1Ixp33_ASAP7_75t_L   g22675(.A1(new_n22812), .A2(new_n22931), .B(new_n22827), .C(new_n22928), .Y(new_n22932));
  NOR2xp33_ASAP7_75t_L      g22676(.A(new_n22932), .B(new_n22930), .Y(new_n22933));
  INVx1_ASAP7_75t_L         g22677(.A(new_n22933), .Y(new_n22934));
  A2O1A1O1Ixp25_ASAP7_75t_L g22678(.A1(new_n22820), .A2(new_n22827), .B(new_n22828), .C(new_n22838), .D(new_n22836), .Y(new_n22935));
  AND2x2_ASAP7_75t_L        g22679(.A(new_n22935), .B(new_n22934), .Y(new_n22936));
  A2O1A1O1Ixp25_ASAP7_75t_L g22680(.A1(new_n22615), .A2(new_n22560), .B(new_n22619), .C(new_n22717), .D(new_n22722), .Y(new_n22937));
  O2A1O1Ixp33_ASAP7_75t_L   g22681(.A1(new_n22937), .A2(new_n22835), .B(new_n22839), .C(new_n22934), .Y(new_n22938));
  NOR2xp33_ASAP7_75t_L      g22682(.A(new_n22938), .B(new_n22936), .Y(new_n22939));
  A2O1A1Ixp33_ASAP7_75t_L   g22683(.A1(new_n22851), .A2(new_n22849), .B(new_n22848), .C(new_n22939), .Y(new_n22940));
  INVx1_ASAP7_75t_L         g22684(.A(new_n22940), .Y(new_n22941));
  A2O1A1Ixp33_ASAP7_75t_L   g22685(.A1(new_n22747), .A2(new_n22744), .B(new_n22742), .C(new_n22849), .Y(new_n22942));
  A2O1A1Ixp33_ASAP7_75t_L   g22686(.A1(new_n22842), .A2(new_n22840), .B(new_n22843), .C(new_n22942), .Y(new_n22943));
  NOR2xp33_ASAP7_75t_L      g22687(.A(new_n22939), .B(new_n22943), .Y(new_n22944));
  NOR2xp33_ASAP7_75t_L      g22688(.A(new_n22941), .B(new_n22944), .Y(\f[111] ));
  A2O1A1Ixp33_ASAP7_75t_L   g22689(.A1(new_n22861), .A2(\a[53] ), .B(new_n22862), .C(new_n22918), .Y(new_n22946));
  A2O1A1O1Ixp25_ASAP7_75t_L g22690(.A1(new_n22867), .A2(\a[56] ), .B(new_n22868), .C(new_n22911), .D(new_n22915), .Y(new_n22947));
  INVx1_ASAP7_75t_L         g22691(.A(new_n22947), .Y(new_n22948));
  NOR2xp33_ASAP7_75t_L      g22692(.A(new_n10978), .B(new_n10388), .Y(new_n22949));
  AOI221xp5_ASAP7_75t_L     g22693(.A1(new_n10086), .A2(\b[58] ), .B1(new_n11361), .B2(\b[56] ), .C(new_n22949), .Y(new_n22950));
  O2A1O1Ixp33_ASAP7_75t_L   g22694(.A1(new_n10088), .A2(new_n20073), .B(new_n22950), .C(new_n10083), .Y(new_n22951));
  O2A1O1Ixp33_ASAP7_75t_L   g22695(.A1(new_n10088), .A2(new_n20073), .B(new_n22950), .C(\a[56] ), .Y(new_n22952));
  INVx1_ASAP7_75t_L         g22696(.A(new_n22952), .Y(new_n22953));
  NOR2xp33_ASAP7_75t_L      g22697(.A(new_n9683), .B(new_n11354), .Y(new_n22954));
  AOI221xp5_ASAP7_75t_L     g22698(.A1(\b[55] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[54] ), .C(new_n22954), .Y(new_n22955));
  O2A1O1Ixp33_ASAP7_75t_L   g22699(.A1(new_n11053), .A2(new_n15849), .B(new_n22955), .C(new_n11048), .Y(new_n22956));
  INVx1_ASAP7_75t_L         g22700(.A(new_n22956), .Y(new_n22957));
  O2A1O1Ixp33_ASAP7_75t_L   g22701(.A1(new_n11053), .A2(new_n15849), .B(new_n22955), .C(\a[59] ), .Y(new_n22958));
  NOR2xp33_ASAP7_75t_L      g22702(.A(new_n7860), .B(new_n13030), .Y(new_n22959));
  O2A1O1Ixp33_ASAP7_75t_L   g22703(.A1(new_n12669), .A2(new_n12671), .B(\b[49] ), .C(new_n22959), .Y(new_n22960));
  INVx1_ASAP7_75t_L         g22704(.A(new_n22960), .Y(new_n22961));
  O2A1O1Ixp33_ASAP7_75t_L   g22705(.A1(\a[47] ), .A2(new_n22767), .B(new_n22878), .C(new_n22961), .Y(new_n22962));
  INVx1_ASAP7_75t_L         g22706(.A(new_n22962), .Y(new_n22963));
  INVx1_ASAP7_75t_L         g22707(.A(new_n22879), .Y(new_n22964));
  O2A1O1Ixp33_ASAP7_75t_L   g22708(.A1(new_n7552), .A2(new_n12672), .B(new_n22764), .C(\a[47] ), .Y(new_n22965));
  O2A1O1Ixp33_ASAP7_75t_L   g22709(.A1(new_n22875), .A2(new_n22874), .B(new_n22964), .C(new_n22965), .Y(new_n22966));
  A2O1A1Ixp33_ASAP7_75t_L   g22710(.A1(new_n13028), .A2(\b[49] ), .B(new_n22959), .C(new_n22966), .Y(new_n22967));
  NAND2xp33_ASAP7_75t_L     g22711(.A(new_n22967), .B(new_n22963), .Y(new_n22968));
  NOR2xp33_ASAP7_75t_L      g22712(.A(new_n8779), .B(new_n12318), .Y(new_n22969));
  AOI221xp5_ASAP7_75t_L     g22713(.A1(new_n11995), .A2(\b[52] ), .B1(new_n13314), .B2(\b[50] ), .C(new_n22969), .Y(new_n22970));
  INVx1_ASAP7_75t_L         g22714(.A(new_n22970), .Y(new_n22971));
  A2O1A1Ixp33_ASAP7_75t_L   g22715(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n22970), .Y(new_n22972));
  O2A1O1Ixp33_ASAP7_75t_L   g22716(.A1(new_n22971), .A2(new_n9367), .B(new_n22972), .C(new_n11987), .Y(new_n22973));
  O2A1O1Ixp33_ASAP7_75t_L   g22717(.A1(new_n11998), .A2(new_n17363), .B(new_n22970), .C(\a[62] ), .Y(new_n22974));
  NOR2xp33_ASAP7_75t_L      g22718(.A(new_n22973), .B(new_n22974), .Y(new_n22975));
  NOR2xp33_ASAP7_75t_L      g22719(.A(new_n22968), .B(new_n22975), .Y(new_n22976));
  INVx1_ASAP7_75t_L         g22720(.A(new_n22976), .Y(new_n22977));
  NAND2xp33_ASAP7_75t_L     g22721(.A(new_n22968), .B(new_n22975), .Y(new_n22978));
  NAND2xp33_ASAP7_75t_L     g22722(.A(new_n22978), .B(new_n22977), .Y(new_n22979));
  O2A1O1Ixp33_ASAP7_75t_L   g22723(.A1(new_n22891), .A2(new_n22773), .B(new_n22889), .C(new_n22979), .Y(new_n22980));
  A2O1A1O1Ixp25_ASAP7_75t_L g22724(.A1(new_n22767), .A2(new_n22670), .B(new_n22770), .C(new_n22894), .D(new_n22888), .Y(new_n22981));
  NAND3xp33_ASAP7_75t_L     g22725(.A(new_n22981), .B(new_n22977), .C(new_n22978), .Y(new_n22982));
  A2O1A1Ixp33_ASAP7_75t_L   g22726(.A1(new_n22893), .A2(new_n22889), .B(new_n22980), .C(new_n22982), .Y(new_n22983));
  AOI21xp33_ASAP7_75t_L     g22727(.A1(new_n22957), .A2(\a[59] ), .B(new_n22958), .Y(new_n22984));
  NAND2xp33_ASAP7_75t_L     g22728(.A(new_n22984), .B(new_n22982), .Y(new_n22985));
  O2A1O1Ixp33_ASAP7_75t_L   g22729(.A1(new_n22888), .A2(new_n22892), .B(new_n22979), .C(new_n22985), .Y(new_n22986));
  A2O1A1O1Ixp25_ASAP7_75t_L g22730(.A1(new_n22957), .A2(\a[59] ), .B(new_n22958), .C(new_n22983), .D(new_n22986), .Y(new_n22987));
  INVx1_ASAP7_75t_L         g22731(.A(new_n22987), .Y(new_n22988));
  O2A1O1Ixp33_ASAP7_75t_L   g22732(.A1(new_n22905), .A2(new_n22908), .B(new_n22904), .C(new_n22988), .Y(new_n22989));
  O2A1O1Ixp33_ASAP7_75t_L   g22733(.A1(new_n22871), .A2(new_n22783), .B(new_n22902), .C(new_n22903), .Y(new_n22990));
  INVx1_ASAP7_75t_L         g22734(.A(new_n22990), .Y(new_n22991));
  O2A1O1Ixp33_ASAP7_75t_L   g22735(.A1(new_n22773), .A2(new_n22891), .B(new_n22889), .C(new_n22980), .Y(new_n22992));
  O2A1O1Ixp33_ASAP7_75t_L   g22736(.A1(new_n22981), .A2(new_n22980), .B(new_n22982), .C(new_n22984), .Y(new_n22993));
  INVx1_ASAP7_75t_L         g22737(.A(new_n22993), .Y(new_n22994));
  O2A1O1Ixp33_ASAP7_75t_L   g22738(.A1(new_n22985), .A2(new_n22992), .B(new_n22994), .C(new_n22991), .Y(new_n22995));
  NOR2xp33_ASAP7_75t_L      g22739(.A(new_n22989), .B(new_n22995), .Y(new_n22996));
  INVx1_ASAP7_75t_L         g22740(.A(new_n22996), .Y(new_n22997));
  O2A1O1Ixp33_ASAP7_75t_L   g22741(.A1(new_n10083), .A2(new_n22951), .B(new_n22953), .C(new_n22997), .Y(new_n22998));
  OA211x2_ASAP7_75t_L       g22742(.A1(new_n22951), .A2(new_n10083), .B(new_n22997), .C(new_n22953), .Y(new_n22999));
  NOR2xp33_ASAP7_75t_L      g22743(.A(new_n22998), .B(new_n22999), .Y(new_n23000));
  A2O1A1Ixp33_ASAP7_75t_L   g22744(.A1(new_n22911), .A2(new_n22870), .B(new_n22915), .C(new_n23000), .Y(new_n23001));
  NAND2xp33_ASAP7_75t_L     g22745(.A(\b[60] ), .B(new_n9096), .Y(new_n23002));
  OAI221xp5_ASAP7_75t_L     g22746(.A1(new_n9440), .A2(new_n11591), .B1(new_n12258), .B2(new_n9439), .C(new_n23002), .Y(new_n23003));
  A2O1A1Ixp33_ASAP7_75t_L   g22747(.A1(new_n12269), .A2(new_n9437), .B(new_n23003), .C(\a[53] ), .Y(new_n23004));
  AOI211xp5_ASAP7_75t_L     g22748(.A1(new_n12269), .A2(new_n9437), .B(new_n23003), .C(new_n9099), .Y(new_n23005));
  A2O1A1O1Ixp25_ASAP7_75t_L g22749(.A1(new_n12269), .A2(new_n9437), .B(new_n23003), .C(new_n23004), .D(new_n23005), .Y(new_n23006));
  INVx1_ASAP7_75t_L         g22750(.A(new_n23001), .Y(new_n23007));
  NAND2xp33_ASAP7_75t_L     g22751(.A(new_n23000), .B(new_n23001), .Y(new_n23008));
  O2A1O1Ixp33_ASAP7_75t_L   g22752(.A1(new_n22947), .A2(new_n23007), .B(new_n23008), .C(new_n23006), .Y(new_n23009));
  INVx1_ASAP7_75t_L         g22753(.A(new_n23009), .Y(new_n23010));
  NAND2xp33_ASAP7_75t_L     g22754(.A(new_n23006), .B(new_n23008), .Y(new_n23011));
  A2O1A1Ixp33_ASAP7_75t_L   g22755(.A1(new_n22948), .A2(new_n23001), .B(new_n23011), .C(new_n23010), .Y(new_n23012));
  O2A1O1Ixp33_ASAP7_75t_L   g22756(.A1(new_n22923), .A2(new_n22920), .B(new_n22946), .C(new_n23012), .Y(new_n23013));
  INVx1_ASAP7_75t_L         g22757(.A(new_n23013), .Y(new_n23014));
  A2O1A1O1Ixp25_ASAP7_75t_L g22758(.A1(new_n22861), .A2(\a[53] ), .B(new_n22862), .C(new_n22918), .D(new_n22921), .Y(new_n23015));
  NAND2xp33_ASAP7_75t_L     g22759(.A(new_n23012), .B(new_n23015), .Y(new_n23016));
  AND2x2_ASAP7_75t_L        g22760(.A(new_n23014), .B(new_n23016), .Y(new_n23017));
  INVx1_ASAP7_75t_L         g22761(.A(new_n23017), .Y(new_n23018));
  AOI22xp33_ASAP7_75t_L     g22762(.A1(new_n8169), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n8484), .Y(new_n23019));
  O2A1O1Ixp33_ASAP7_75t_L   g22763(.A1(new_n8176), .A2(new_n12993), .B(new_n23019), .C(new_n8172), .Y(new_n23020));
  O2A1O1Ixp33_ASAP7_75t_L   g22764(.A1(new_n8176), .A2(new_n12993), .B(new_n23019), .C(\a[50] ), .Y(new_n23021));
  INVx1_ASAP7_75t_L         g22765(.A(new_n23021), .Y(new_n23022));
  O2A1O1Ixp33_ASAP7_75t_L   g22766(.A1(new_n23020), .A2(new_n8172), .B(new_n23022), .C(new_n23018), .Y(new_n23023));
  INVx1_ASAP7_75t_L         g22767(.A(new_n23023), .Y(new_n23024));
  O2A1O1Ixp33_ASAP7_75t_L   g22768(.A1(new_n23020), .A2(new_n8172), .B(new_n23022), .C(new_n23017), .Y(new_n23025));
  AOI21xp33_ASAP7_75t_L     g22769(.A1(new_n23024), .A2(new_n23017), .B(new_n23025), .Y(new_n23026));
  A2O1A1O1Ixp25_ASAP7_75t_L g22770(.A1(new_n22856), .A2(\a[50] ), .B(new_n22857), .C(new_n22925), .D(new_n22932), .Y(new_n23027));
  NAND2xp33_ASAP7_75t_L     g22771(.A(new_n23026), .B(new_n23027), .Y(new_n23028));
  A2O1A1O1Ixp25_ASAP7_75t_L g22772(.A1(new_n22827), .A2(new_n22816), .B(new_n22928), .C(new_n22926), .D(new_n23026), .Y(new_n23029));
  INVx1_ASAP7_75t_L         g22773(.A(new_n23029), .Y(new_n23030));
  AND2x2_ASAP7_75t_L        g22774(.A(new_n23028), .B(new_n23030), .Y(new_n23031));
  INVx1_ASAP7_75t_L         g22775(.A(new_n23031), .Y(new_n23032));
  O2A1O1Ixp33_ASAP7_75t_L   g22776(.A1(new_n22934), .A2(new_n22935), .B(new_n22940), .C(new_n23032), .Y(new_n23033));
  INVx1_ASAP7_75t_L         g22777(.A(new_n22938), .Y(new_n23034));
  A2O1A1Ixp33_ASAP7_75t_L   g22778(.A1(new_n22942), .A2(new_n22847), .B(new_n22936), .C(new_n23034), .Y(new_n23035));
  NOR2xp33_ASAP7_75t_L      g22779(.A(new_n23031), .B(new_n23035), .Y(new_n23036));
  NOR2xp33_ASAP7_75t_L      g22780(.A(new_n23033), .B(new_n23036), .Y(\f[112] ));
  NOR2xp33_ASAP7_75t_L      g22781(.A(new_n9355), .B(new_n12318), .Y(new_n23038));
  AOI221xp5_ASAP7_75t_L     g22782(.A1(new_n11995), .A2(\b[53] ), .B1(new_n13314), .B2(\b[51] ), .C(new_n23038), .Y(new_n23039));
  O2A1O1Ixp33_ASAP7_75t_L   g22783(.A1(new_n11998), .A2(new_n9691), .B(new_n23039), .C(new_n11987), .Y(new_n23040));
  INVx1_ASAP7_75t_L         g22784(.A(new_n23039), .Y(new_n23041));
  A2O1A1Ixp33_ASAP7_75t_L   g22785(.A1(new_n9690), .A2(new_n11997), .B(new_n23041), .C(new_n11987), .Y(new_n23042));
  NOR2xp33_ASAP7_75t_L      g22786(.A(new_n8427), .B(new_n13030), .Y(new_n23043));
  INVx1_ASAP7_75t_L         g22787(.A(new_n23043), .Y(new_n23044));
  O2A1O1Ixp33_ASAP7_75t_L   g22788(.A1(new_n12672), .A2(new_n8755), .B(new_n23044), .C(new_n22961), .Y(new_n23045));
  INVx1_ASAP7_75t_L         g22789(.A(new_n23045), .Y(new_n23046));
  NOR2xp33_ASAP7_75t_L      g22790(.A(new_n22961), .B(new_n23045), .Y(new_n23047));
  A2O1A1O1Ixp25_ASAP7_75t_L g22791(.A1(new_n13028), .A2(\b[50] ), .B(new_n23043), .C(new_n23046), .D(new_n23047), .Y(new_n23048));
  O2A1O1Ixp33_ASAP7_75t_L   g22792(.A1(new_n11987), .A2(new_n23040), .B(new_n23042), .C(new_n23048), .Y(new_n23049));
  O2A1O1Ixp33_ASAP7_75t_L   g22793(.A1(new_n11987), .A2(new_n23040), .B(new_n23042), .C(new_n23049), .Y(new_n23050));
  OAI21xp33_ASAP7_75t_L     g22794(.A1(new_n11987), .A2(new_n23040), .B(new_n23042), .Y(new_n23051));
  A2O1A1Ixp33_ASAP7_75t_L   g22795(.A1(\b[50] ), .A2(new_n13028), .B(new_n23043), .C(new_n22961), .Y(new_n23052));
  O2A1O1Ixp33_ASAP7_75t_L   g22796(.A1(new_n23045), .A2(new_n22961), .B(new_n23052), .C(new_n23051), .Y(new_n23053));
  NOR4xp25_ASAP7_75t_L      g22797(.A(new_n23050), .B(new_n22962), .C(new_n23053), .D(new_n22976), .Y(new_n23054));
  O2A1O1Ixp33_ASAP7_75t_L   g22798(.A1(new_n12672), .A2(new_n8755), .B(new_n23044), .C(new_n22960), .Y(new_n23055));
  INVx1_ASAP7_75t_L         g22799(.A(new_n23049), .Y(new_n23056));
  O2A1O1Ixp33_ASAP7_75t_L   g22800(.A1(new_n23047), .A2(new_n23055), .B(new_n23056), .C(new_n23050), .Y(new_n23057));
  O2A1O1Ixp33_ASAP7_75t_L   g22801(.A1(new_n22961), .A2(new_n22966), .B(new_n22977), .C(new_n23057), .Y(new_n23058));
  NOR2xp33_ASAP7_75t_L      g22802(.A(new_n23054), .B(new_n23058), .Y(new_n23059));
  INVx1_ASAP7_75t_L         g22803(.A(new_n23059), .Y(new_n23060));
  NOR2xp33_ASAP7_75t_L      g22804(.A(new_n9709), .B(new_n11354), .Y(new_n23061));
  AOI221xp5_ASAP7_75t_L     g22805(.A1(\b[56] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[55] ), .C(new_n23061), .Y(new_n23062));
  O2A1O1Ixp33_ASAP7_75t_L   g22806(.A1(new_n11053), .A2(new_n10339), .B(new_n23062), .C(new_n11048), .Y(new_n23063));
  O2A1O1Ixp33_ASAP7_75t_L   g22807(.A1(new_n11053), .A2(new_n10339), .B(new_n23062), .C(\a[59] ), .Y(new_n23064));
  INVx1_ASAP7_75t_L         g22808(.A(new_n23064), .Y(new_n23065));
  OAI211xp5_ASAP7_75t_L     g22809(.A1(new_n11048), .A2(new_n23063), .B(new_n23060), .C(new_n23065), .Y(new_n23066));
  O2A1O1Ixp33_ASAP7_75t_L   g22810(.A1(new_n23063), .A2(new_n11048), .B(new_n23065), .C(new_n23060), .Y(new_n23067));
  INVx1_ASAP7_75t_L         g22811(.A(new_n23067), .Y(new_n23068));
  AND2x2_ASAP7_75t_L        g22812(.A(new_n23066), .B(new_n23068), .Y(new_n23069));
  INVx1_ASAP7_75t_L         g22813(.A(new_n23069), .Y(new_n23070));
  O2A1O1Ixp33_ASAP7_75t_L   g22814(.A1(new_n22981), .A2(new_n22979), .B(new_n22994), .C(new_n23070), .Y(new_n23071));
  INVx1_ASAP7_75t_L         g22815(.A(new_n23071), .Y(new_n23072));
  A2O1A1O1Ixp25_ASAP7_75t_L g22816(.A1(new_n22957), .A2(\a[59] ), .B(new_n22958), .C(new_n22983), .D(new_n22980), .Y(new_n23073));
  NAND2xp33_ASAP7_75t_L     g22817(.A(new_n23073), .B(new_n23070), .Y(new_n23074));
  AND2x2_ASAP7_75t_L        g22818(.A(new_n23074), .B(new_n23072), .Y(new_n23075));
  INVx1_ASAP7_75t_L         g22819(.A(new_n23075), .Y(new_n23076));
  NOR2xp33_ASAP7_75t_L      g22820(.A(new_n11303), .B(new_n10388), .Y(new_n23077));
  AOI221xp5_ASAP7_75t_L     g22821(.A1(new_n10086), .A2(\b[59] ), .B1(new_n11361), .B2(\b[57] ), .C(new_n23077), .Y(new_n23078));
  O2A1O1Ixp33_ASAP7_75t_L   g22822(.A1(new_n10088), .A2(new_n11597), .B(new_n23078), .C(new_n10083), .Y(new_n23079));
  O2A1O1Ixp33_ASAP7_75t_L   g22823(.A1(new_n10088), .A2(new_n11597), .B(new_n23078), .C(\a[56] ), .Y(new_n23080));
  INVx1_ASAP7_75t_L         g22824(.A(new_n23080), .Y(new_n23081));
  O2A1O1Ixp33_ASAP7_75t_L   g22825(.A1(new_n23079), .A2(new_n10083), .B(new_n23081), .C(new_n23076), .Y(new_n23082));
  INVx1_ASAP7_75t_L         g22826(.A(new_n23082), .Y(new_n23083));
  O2A1O1Ixp33_ASAP7_75t_L   g22827(.A1(new_n23079), .A2(new_n10083), .B(new_n23081), .C(new_n23075), .Y(new_n23084));
  AOI21xp33_ASAP7_75t_L     g22828(.A1(new_n23083), .A2(new_n23075), .B(new_n23084), .Y(new_n23085));
  O2A1O1Ixp33_ASAP7_75t_L   g22829(.A1(new_n22903), .A2(new_n22906), .B(new_n22987), .C(new_n22998), .Y(new_n23086));
  NAND2xp33_ASAP7_75t_L     g22830(.A(new_n23086), .B(new_n23085), .Y(new_n23087));
  INVx1_ASAP7_75t_L         g22831(.A(new_n22998), .Y(new_n23088));
  O2A1O1Ixp33_ASAP7_75t_L   g22832(.A1(new_n22990), .A2(new_n22988), .B(new_n23088), .C(new_n23085), .Y(new_n23089));
  INVx1_ASAP7_75t_L         g22833(.A(new_n23089), .Y(new_n23090));
  AND2x2_ASAP7_75t_L        g22834(.A(new_n23087), .B(new_n23090), .Y(new_n23091));
  INVx1_ASAP7_75t_L         g22835(.A(new_n23091), .Y(new_n23092));
  NOR2xp33_ASAP7_75t_L      g22836(.A(new_n12258), .B(new_n10400), .Y(new_n23093));
  AOI221xp5_ASAP7_75t_L     g22837(.A1(new_n9102), .A2(\b[62] ), .B1(new_n10398), .B2(\b[60] ), .C(new_n23093), .Y(new_n23094));
  O2A1O1Ixp33_ASAP7_75t_L   g22838(.A1(new_n9104), .A2(new_n12610), .B(new_n23094), .C(new_n9099), .Y(new_n23095));
  O2A1O1Ixp33_ASAP7_75t_L   g22839(.A1(new_n9104), .A2(new_n12610), .B(new_n23094), .C(\a[53] ), .Y(new_n23096));
  INVx1_ASAP7_75t_L         g22840(.A(new_n23096), .Y(new_n23097));
  O2A1O1Ixp33_ASAP7_75t_L   g22841(.A1(new_n23095), .A2(new_n9099), .B(new_n23097), .C(new_n23092), .Y(new_n23098));
  INVx1_ASAP7_75t_L         g22842(.A(new_n23098), .Y(new_n23099));
  O2A1O1Ixp33_ASAP7_75t_L   g22843(.A1(new_n23095), .A2(new_n9099), .B(new_n23097), .C(new_n23091), .Y(new_n23100));
  NOR2xp33_ASAP7_75t_L      g22844(.A(new_n12956), .B(new_n8483), .Y(new_n23101));
  INVx1_ASAP7_75t_L         g22845(.A(new_n23101), .Y(new_n23102));
  A2O1A1Ixp33_ASAP7_75t_L   g22846(.A1(new_n14444), .A2(new_n12603), .B(new_n12956), .C(new_n23102), .Y(new_n23103));
  O2A1O1Ixp33_ASAP7_75t_L   g22847(.A1(new_n8490), .A2(new_n23101), .B(new_n23103), .C(new_n8172), .Y(new_n23104));
  O2A1O1Ixp33_ASAP7_75t_L   g22848(.A1(new_n8176), .A2(new_n13573), .B(new_n23102), .C(\a[50] ), .Y(new_n23105));
  NOR2xp33_ASAP7_75t_L      g22849(.A(new_n23105), .B(new_n23104), .Y(new_n23106));
  A2O1A1O1Ixp25_ASAP7_75t_L g22850(.A1(new_n22947), .A2(new_n23008), .B(new_n23006), .C(new_n23001), .D(new_n23106), .Y(new_n23107));
  NOR4xp25_ASAP7_75t_L      g22851(.A(new_n23009), .B(new_n23105), .C(new_n23007), .D(new_n23104), .Y(new_n23108));
  NOR2xp33_ASAP7_75t_L      g22852(.A(new_n23107), .B(new_n23108), .Y(new_n23109));
  A2O1A1Ixp33_ASAP7_75t_L   g22853(.A1(new_n23099), .A2(new_n23091), .B(new_n23100), .C(new_n23109), .Y(new_n23110));
  AND2x2_ASAP7_75t_L        g22854(.A(new_n23109), .B(new_n23110), .Y(new_n23111));
  A2O1A1O1Ixp25_ASAP7_75t_L g22855(.A1(new_n23099), .A2(new_n23091), .B(new_n23100), .C(new_n23110), .D(new_n23111), .Y(new_n23112));
  INVx1_ASAP7_75t_L         g22856(.A(new_n23112), .Y(new_n23113));
  A2O1A1Ixp33_ASAP7_75t_L   g22857(.A1(new_n22922), .A2(new_n22946), .B(new_n23012), .C(new_n23024), .Y(new_n23114));
  NOR2xp33_ASAP7_75t_L      g22858(.A(new_n23113), .B(new_n23114), .Y(new_n23115));
  O2A1O1Ixp33_ASAP7_75t_L   g22859(.A1(new_n23015), .A2(new_n23012), .B(new_n23024), .C(new_n23112), .Y(new_n23116));
  NOR2xp33_ASAP7_75t_L      g22860(.A(new_n23116), .B(new_n23115), .Y(new_n23117));
  A2O1A1Ixp33_ASAP7_75t_L   g22861(.A1(new_n22940), .A2(new_n23034), .B(new_n23032), .C(new_n23030), .Y(new_n23118));
  XOR2x2_ASAP7_75t_L        g22862(.A(new_n23117), .B(new_n23118), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g22863(.A(new_n11591), .B(new_n10388), .Y(new_n23120));
  AOI221xp5_ASAP7_75t_L     g22864(.A1(new_n10086), .A2(\b[60] ), .B1(new_n11361), .B2(\b[58] ), .C(new_n23120), .Y(new_n23121));
  INVx1_ASAP7_75t_L         g22865(.A(new_n23121), .Y(new_n23122));
  A2O1A1Ixp33_ASAP7_75t_L   g22866(.A1(new_n13839), .A2(new_n10386), .B(new_n23122), .C(\a[56] ), .Y(new_n23123));
  O2A1O1Ixp33_ASAP7_75t_L   g22867(.A1(new_n10088), .A2(new_n11634), .B(new_n23121), .C(\a[56] ), .Y(new_n23124));
  A2O1A1Ixp33_ASAP7_75t_L   g22868(.A1(new_n22977), .A2(new_n22963), .B(new_n23057), .C(new_n23068), .Y(new_n23125));
  O2A1O1Ixp33_ASAP7_75t_L   g22869(.A1(new_n22960), .A2(new_n23055), .B(new_n23051), .C(new_n23045), .Y(new_n23126));
  NOR2xp33_ASAP7_75t_L      g22870(.A(new_n8755), .B(new_n13030), .Y(new_n23127));
  A2O1A1Ixp33_ASAP7_75t_L   g22871(.A1(new_n13028), .A2(\b[51] ), .B(new_n23127), .C(new_n8172), .Y(new_n23128));
  INVx1_ASAP7_75t_L         g22872(.A(new_n23128), .Y(new_n23129));
  O2A1O1Ixp33_ASAP7_75t_L   g22873(.A1(new_n12669), .A2(new_n12671), .B(\b[51] ), .C(new_n23127), .Y(new_n23130));
  NAND2xp33_ASAP7_75t_L     g22874(.A(\a[50] ), .B(new_n23130), .Y(new_n23131));
  INVx1_ASAP7_75t_L         g22875(.A(new_n23131), .Y(new_n23132));
  NOR2xp33_ASAP7_75t_L      g22876(.A(new_n23129), .B(new_n23132), .Y(new_n23133));
  A2O1A1Ixp33_ASAP7_75t_L   g22877(.A1(new_n13028), .A2(\b[49] ), .B(new_n22959), .C(new_n23133), .Y(new_n23134));
  OAI21xp33_ASAP7_75t_L     g22878(.A1(new_n23129), .A2(new_n23132), .B(new_n22960), .Y(new_n23135));
  AND2x2_ASAP7_75t_L        g22879(.A(new_n23135), .B(new_n23134), .Y(new_n23136));
  NOR2xp33_ASAP7_75t_L      g22880(.A(new_n9683), .B(new_n12318), .Y(new_n23137));
  AOI221xp5_ASAP7_75t_L     g22881(.A1(new_n11995), .A2(\b[54] ), .B1(new_n13314), .B2(\b[52] ), .C(new_n23137), .Y(new_n23138));
  O2A1O1Ixp33_ASAP7_75t_L   g22882(.A1(new_n11998), .A2(new_n9718), .B(new_n23138), .C(new_n11987), .Y(new_n23139));
  NOR2xp33_ASAP7_75t_L      g22883(.A(new_n11987), .B(new_n23139), .Y(new_n23140));
  O2A1O1Ixp33_ASAP7_75t_L   g22884(.A1(new_n11998), .A2(new_n9718), .B(new_n23138), .C(\a[62] ), .Y(new_n23141));
  NOR2xp33_ASAP7_75t_L      g22885(.A(new_n23141), .B(new_n23140), .Y(new_n23142));
  INVx1_ASAP7_75t_L         g22886(.A(new_n23136), .Y(new_n23143));
  O2A1O1Ixp33_ASAP7_75t_L   g22887(.A1(new_n12669), .A2(new_n12671), .B(\b[50] ), .C(new_n23043), .Y(new_n23144));
  O2A1O1Ixp33_ASAP7_75t_L   g22888(.A1(new_n22961), .A2(new_n23144), .B(new_n23056), .C(new_n23143), .Y(new_n23145));
  O2A1O1Ixp33_ASAP7_75t_L   g22889(.A1(new_n22961), .A2(new_n23144), .B(new_n23056), .C(new_n23136), .Y(new_n23146));
  INVx1_ASAP7_75t_L         g22890(.A(new_n23146), .Y(new_n23147));
  O2A1O1Ixp33_ASAP7_75t_L   g22891(.A1(new_n23143), .A2(new_n23145), .B(new_n23147), .C(new_n23142), .Y(new_n23148));
  NOR2xp33_ASAP7_75t_L      g22892(.A(new_n23143), .B(new_n23145), .Y(new_n23149));
  NOR3xp33_ASAP7_75t_L      g22893(.A(new_n23149), .B(new_n23141), .C(new_n23140), .Y(new_n23150));
  O2A1O1Ixp33_ASAP7_75t_L   g22894(.A1(new_n23136), .A2(new_n23126), .B(new_n23150), .C(new_n23148), .Y(new_n23151));
  NOR2xp33_ASAP7_75t_L      g22895(.A(new_n10309), .B(new_n11354), .Y(new_n23152));
  AOI221xp5_ASAP7_75t_L     g22896(.A1(\b[57] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[56] ), .C(new_n23152), .Y(new_n23153));
  O2A1O1Ixp33_ASAP7_75t_L   g22897(.A1(new_n11053), .A2(new_n17096), .B(new_n23153), .C(new_n11048), .Y(new_n23154));
  INVx1_ASAP7_75t_L         g22898(.A(new_n23154), .Y(new_n23155));
  O2A1O1Ixp33_ASAP7_75t_L   g22899(.A1(new_n11053), .A2(new_n17096), .B(new_n23153), .C(\a[59] ), .Y(new_n23156));
  A2O1A1Ixp33_ASAP7_75t_L   g22900(.A1(new_n23155), .A2(\a[59] ), .B(new_n23156), .C(new_n23151), .Y(new_n23157));
  A2O1A1Ixp33_ASAP7_75t_L   g22901(.A1(new_n23155), .A2(\a[59] ), .B(new_n23156), .C(new_n23157), .Y(new_n23158));
  INVx1_ASAP7_75t_L         g22902(.A(new_n23158), .Y(new_n23159));
  A2O1A1Ixp33_ASAP7_75t_L   g22903(.A1(new_n23151), .A2(new_n23157), .B(new_n23159), .C(new_n23125), .Y(new_n23160));
  AOI21xp33_ASAP7_75t_L     g22904(.A1(new_n23157), .A2(new_n23151), .B(new_n23125), .Y(new_n23161));
  NAND2xp33_ASAP7_75t_L     g22905(.A(new_n23158), .B(new_n23161), .Y(new_n23162));
  NAND2xp33_ASAP7_75t_L     g22906(.A(new_n23160), .B(new_n23162), .Y(new_n23163));
  INVx1_ASAP7_75t_L         g22907(.A(new_n23163), .Y(new_n23164));
  A2O1A1Ixp33_ASAP7_75t_L   g22908(.A1(new_n23123), .A2(\a[56] ), .B(new_n23124), .C(new_n23164), .Y(new_n23165));
  AO21x2_ASAP7_75t_L        g22909(.A1(\a[56] ), .A2(new_n23123), .B(new_n23124), .Y(new_n23166));
  AO21x2_ASAP7_75t_L        g22910(.A1(new_n23160), .A2(new_n23162), .B(new_n23166), .Y(new_n23167));
  AND2x2_ASAP7_75t_L        g22911(.A(new_n23167), .B(new_n23165), .Y(new_n23168));
  INVx1_ASAP7_75t_L         g22912(.A(new_n23168), .Y(new_n23169));
  O2A1O1Ixp33_ASAP7_75t_L   g22913(.A1(new_n23073), .A2(new_n23070), .B(new_n23083), .C(new_n23169), .Y(new_n23170));
  INVx1_ASAP7_75t_L         g22914(.A(new_n23170), .Y(new_n23171));
  O2A1O1Ixp33_ASAP7_75t_L   g22915(.A1(new_n22980), .A2(new_n22993), .B(new_n23069), .C(new_n23082), .Y(new_n23172));
  NAND2xp33_ASAP7_75t_L     g22916(.A(new_n23169), .B(new_n23172), .Y(new_n23173));
  NAND2xp33_ASAP7_75t_L     g22917(.A(new_n23173), .B(new_n23171), .Y(new_n23174));
  INVx1_ASAP7_75t_L         g22918(.A(new_n23174), .Y(new_n23175));
  NOR2xp33_ASAP7_75t_L      g22919(.A(new_n12603), .B(new_n10400), .Y(new_n23176));
  AOI221xp5_ASAP7_75t_L     g22920(.A1(new_n9102), .A2(\b[63] ), .B1(new_n10398), .B2(\b[61] ), .C(new_n23176), .Y(new_n23177));
  O2A1O1Ixp33_ASAP7_75t_L   g22921(.A1(new_n9104), .A2(new_n17815), .B(new_n23177), .C(new_n9099), .Y(new_n23178));
  O2A1O1Ixp33_ASAP7_75t_L   g22922(.A1(new_n9104), .A2(new_n17815), .B(new_n23177), .C(\a[53] ), .Y(new_n23179));
  INVx1_ASAP7_75t_L         g22923(.A(new_n23179), .Y(new_n23180));
  O2A1O1Ixp33_ASAP7_75t_L   g22924(.A1(new_n23178), .A2(new_n9099), .B(new_n23180), .C(new_n23174), .Y(new_n23181));
  INVx1_ASAP7_75t_L         g22925(.A(new_n23181), .Y(new_n23182));
  O2A1O1Ixp33_ASAP7_75t_L   g22926(.A1(new_n23178), .A2(new_n9099), .B(new_n23180), .C(new_n23175), .Y(new_n23183));
  INVx1_ASAP7_75t_L         g22927(.A(new_n22989), .Y(new_n23184));
  A2O1A1Ixp33_ASAP7_75t_L   g22928(.A1(new_n23088), .A2(new_n23184), .B(new_n23085), .C(new_n23099), .Y(new_n23185));
  AOI211xp5_ASAP7_75t_L     g22929(.A1(new_n23175), .A2(new_n23182), .B(new_n23183), .C(new_n23185), .Y(new_n23186));
  AOI21xp33_ASAP7_75t_L     g22930(.A1(new_n23182), .A2(new_n23175), .B(new_n23183), .Y(new_n23187));
  O2A1O1Ixp33_ASAP7_75t_L   g22931(.A1(new_n23085), .A2(new_n23086), .B(new_n23099), .C(new_n23187), .Y(new_n23188));
  NOR2xp33_ASAP7_75t_L      g22932(.A(new_n23188), .B(new_n23186), .Y(new_n23189));
  INVx1_ASAP7_75t_L         g22933(.A(new_n23189), .Y(new_n23190));
  A2O1A1O1Ixp25_ASAP7_75t_L g22934(.A1(new_n23091), .A2(new_n23099), .B(new_n23100), .C(new_n23109), .D(new_n23107), .Y(new_n23191));
  AND2x2_ASAP7_75t_L        g22935(.A(new_n23191), .B(new_n23190), .Y(new_n23192));
  A2O1A1O1Ixp25_ASAP7_75t_L g22936(.A1(new_n22911), .A2(new_n22870), .B(new_n22915), .C(new_n23000), .D(new_n23009), .Y(new_n23193));
  O2A1O1Ixp33_ASAP7_75t_L   g22937(.A1(new_n23193), .A2(new_n23106), .B(new_n23110), .C(new_n23190), .Y(new_n23194));
  NOR2xp33_ASAP7_75t_L      g22938(.A(new_n23194), .B(new_n23192), .Y(new_n23195));
  A2O1A1Ixp33_ASAP7_75t_L   g22939(.A1(new_n23118), .A2(new_n23117), .B(new_n23116), .C(new_n23195), .Y(new_n23196));
  INVx1_ASAP7_75t_L         g22940(.A(new_n23196), .Y(new_n23197));
  A2O1A1Ixp33_ASAP7_75t_L   g22941(.A1(new_n23035), .A2(new_n23031), .B(new_n23029), .C(new_n23117), .Y(new_n23198));
  A2O1A1Ixp33_ASAP7_75t_L   g22942(.A1(new_n23024), .A2(new_n23014), .B(new_n23112), .C(new_n23198), .Y(new_n23199));
  NOR2xp33_ASAP7_75t_L      g22943(.A(new_n23195), .B(new_n23199), .Y(new_n23200));
  NOR2xp33_ASAP7_75t_L      g22944(.A(new_n23197), .B(new_n23200), .Y(\f[114] ));
  NAND2xp33_ASAP7_75t_L     g22945(.A(new_n23157), .B(new_n23160), .Y(new_n23202));
  INVx1_ASAP7_75t_L         g22946(.A(new_n23202), .Y(new_n23203));
  NOR2xp33_ASAP7_75t_L      g22947(.A(new_n10332), .B(new_n11354), .Y(new_n23204));
  AOI221xp5_ASAP7_75t_L     g22948(.A1(\b[58] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[57] ), .C(new_n23204), .Y(new_n23205));
  O2A1O1Ixp33_ASAP7_75t_L   g22949(.A1(new_n11053), .A2(new_n20073), .B(new_n23205), .C(new_n11048), .Y(new_n23206));
  O2A1O1Ixp33_ASAP7_75t_L   g22950(.A1(new_n11053), .A2(new_n20073), .B(new_n23205), .C(\a[59] ), .Y(new_n23207));
  INVx1_ASAP7_75t_L         g22951(.A(new_n23207), .Y(new_n23208));
  INVx1_ASAP7_75t_L         g22952(.A(new_n23145), .Y(new_n23209));
  O2A1O1Ixp33_ASAP7_75t_L   g22953(.A1(new_n23045), .A2(new_n23049), .B(new_n23209), .C(new_n23149), .Y(new_n23210));
  NOR2xp33_ASAP7_75t_L      g22954(.A(new_n8779), .B(new_n13030), .Y(new_n23211));
  A2O1A1O1Ixp25_ASAP7_75t_L g22955(.A1(new_n13028), .A2(\b[49] ), .B(new_n22959), .C(new_n23131), .D(new_n23129), .Y(new_n23212));
  A2O1A1Ixp33_ASAP7_75t_L   g22956(.A1(new_n13028), .A2(\b[52] ), .B(new_n23211), .C(new_n23212), .Y(new_n23213));
  O2A1O1Ixp33_ASAP7_75t_L   g22957(.A1(new_n12669), .A2(new_n12671), .B(\b[52] ), .C(new_n23211), .Y(new_n23214));
  INVx1_ASAP7_75t_L         g22958(.A(new_n23214), .Y(new_n23215));
  O2A1O1Ixp33_ASAP7_75t_L   g22959(.A1(new_n22960), .A2(new_n23132), .B(new_n23128), .C(new_n23215), .Y(new_n23216));
  INVx1_ASAP7_75t_L         g22960(.A(new_n23216), .Y(new_n23217));
  NAND2xp33_ASAP7_75t_L     g22961(.A(new_n23213), .B(new_n23217), .Y(new_n23218));
  NOR2xp33_ASAP7_75t_L      g22962(.A(new_n9709), .B(new_n12318), .Y(new_n23219));
  AOI221xp5_ASAP7_75t_L     g22963(.A1(new_n11995), .A2(\b[55] ), .B1(new_n13314), .B2(\b[53] ), .C(new_n23219), .Y(new_n23220));
  O2A1O1Ixp33_ASAP7_75t_L   g22964(.A1(new_n11998), .A2(new_n15849), .B(new_n23220), .C(new_n11987), .Y(new_n23221));
  O2A1O1Ixp33_ASAP7_75t_L   g22965(.A1(new_n11998), .A2(new_n15849), .B(new_n23220), .C(\a[62] ), .Y(new_n23222));
  INVx1_ASAP7_75t_L         g22966(.A(new_n23222), .Y(new_n23223));
  OAI211xp5_ASAP7_75t_L     g22967(.A1(new_n11987), .A2(new_n23221), .B(new_n23223), .C(new_n23218), .Y(new_n23224));
  O2A1O1Ixp33_ASAP7_75t_L   g22968(.A1(new_n11987), .A2(new_n23221), .B(new_n23223), .C(new_n23218), .Y(new_n23225));
  INVx1_ASAP7_75t_L         g22969(.A(new_n23225), .Y(new_n23226));
  AND2x2_ASAP7_75t_L        g22970(.A(new_n23224), .B(new_n23226), .Y(new_n23227));
  INVx1_ASAP7_75t_L         g22971(.A(new_n23227), .Y(new_n23228));
  O2A1O1Ixp33_ASAP7_75t_L   g22972(.A1(new_n23142), .A2(new_n23210), .B(new_n23209), .C(new_n23228), .Y(new_n23229));
  NOR3xp33_ASAP7_75t_L      g22973(.A(new_n23227), .B(new_n23148), .C(new_n23145), .Y(new_n23230));
  NOR2xp33_ASAP7_75t_L      g22974(.A(new_n23230), .B(new_n23229), .Y(new_n23231));
  INVx1_ASAP7_75t_L         g22975(.A(new_n23231), .Y(new_n23232));
  O2A1O1Ixp33_ASAP7_75t_L   g22976(.A1(new_n11048), .A2(new_n23206), .B(new_n23208), .C(new_n23232), .Y(new_n23233));
  INVx1_ASAP7_75t_L         g22977(.A(new_n23233), .Y(new_n23234));
  OAI211xp5_ASAP7_75t_L     g22978(.A1(new_n11048), .A2(new_n23206), .B(new_n23232), .C(new_n23208), .Y(new_n23235));
  AND2x2_ASAP7_75t_L        g22979(.A(new_n23235), .B(new_n23234), .Y(new_n23236));
  INVx1_ASAP7_75t_L         g22980(.A(new_n23236), .Y(new_n23237));
  NOR2xp33_ASAP7_75t_L      g22981(.A(new_n23203), .B(new_n23237), .Y(new_n23238));
  NOR2xp33_ASAP7_75t_L      g22982(.A(new_n11626), .B(new_n10388), .Y(new_n23239));
  AOI221xp5_ASAP7_75t_L     g22983(.A1(new_n10086), .A2(\b[61] ), .B1(new_n11361), .B2(\b[59] ), .C(new_n23239), .Y(new_n23240));
  O2A1O1Ixp33_ASAP7_75t_L   g22984(.A1(new_n10088), .A2(new_n14764), .B(new_n23240), .C(new_n10083), .Y(new_n23241));
  INVx1_ASAP7_75t_L         g22985(.A(new_n23241), .Y(new_n23242));
  O2A1O1Ixp33_ASAP7_75t_L   g22986(.A1(new_n10088), .A2(new_n14764), .B(new_n23240), .C(\a[56] ), .Y(new_n23243));
  AOI21xp33_ASAP7_75t_L     g22987(.A1(new_n23242), .A2(\a[56] ), .B(new_n23243), .Y(new_n23244));
  NOR2xp33_ASAP7_75t_L      g22988(.A(new_n23203), .B(new_n23236), .Y(new_n23245));
  INVx1_ASAP7_75t_L         g22989(.A(new_n23245), .Y(new_n23246));
  O2A1O1Ixp33_ASAP7_75t_L   g22990(.A1(new_n23237), .A2(new_n23238), .B(new_n23246), .C(new_n23244), .Y(new_n23247));
  INVx1_ASAP7_75t_L         g22991(.A(new_n23244), .Y(new_n23248));
  AOI21xp33_ASAP7_75t_L     g22992(.A1(new_n23236), .A2(new_n23203), .B(new_n23248), .Y(new_n23249));
  O2A1O1Ixp33_ASAP7_75t_L   g22993(.A1(new_n23238), .A2(new_n23203), .B(new_n23249), .C(new_n23247), .Y(new_n23250));
  INVx1_ASAP7_75t_L         g22994(.A(new_n23250), .Y(new_n23251));
  O2A1O1Ixp33_ASAP7_75t_L   g22995(.A1(new_n23172), .A2(new_n23169), .B(new_n23165), .C(new_n23251), .Y(new_n23252));
  INVx1_ASAP7_75t_L         g22996(.A(new_n23252), .Y(new_n23253));
  A2O1A1O1Ixp25_ASAP7_75t_L g22997(.A1(new_n23123), .A2(\a[56] ), .B(new_n23124), .C(new_n23164), .D(new_n23170), .Y(new_n23254));
  A2O1A1Ixp33_ASAP7_75t_L   g22998(.A1(new_n23249), .A2(new_n23246), .B(new_n23247), .C(new_n23254), .Y(new_n23255));
  NAND2xp33_ASAP7_75t_L     g22999(.A(new_n23253), .B(new_n23255), .Y(new_n23256));
  INVx1_ASAP7_75t_L         g23000(.A(new_n23256), .Y(new_n23257));
  AOI22xp33_ASAP7_75t_L     g23001(.A1(new_n9096), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n10398), .Y(new_n23258));
  O2A1O1Ixp33_ASAP7_75t_L   g23002(.A1(new_n9104), .A2(new_n12993), .B(new_n23258), .C(new_n9099), .Y(new_n23259));
  O2A1O1Ixp33_ASAP7_75t_L   g23003(.A1(new_n9104), .A2(new_n12993), .B(new_n23258), .C(\a[53] ), .Y(new_n23260));
  INVx1_ASAP7_75t_L         g23004(.A(new_n23260), .Y(new_n23261));
  O2A1O1Ixp33_ASAP7_75t_L   g23005(.A1(new_n23259), .A2(new_n9099), .B(new_n23261), .C(new_n23256), .Y(new_n23262));
  INVx1_ASAP7_75t_L         g23006(.A(new_n23262), .Y(new_n23263));
  O2A1O1Ixp33_ASAP7_75t_L   g23007(.A1(new_n23259), .A2(new_n9099), .B(new_n23261), .C(new_n23257), .Y(new_n23264));
  AOI21xp33_ASAP7_75t_L     g23008(.A1(new_n23263), .A2(new_n23257), .B(new_n23264), .Y(new_n23265));
  O2A1O1Ixp33_ASAP7_75t_L   g23009(.A1(new_n23183), .A2(new_n23175), .B(new_n23185), .C(new_n23181), .Y(new_n23266));
  NAND2xp33_ASAP7_75t_L     g23010(.A(new_n23265), .B(new_n23266), .Y(new_n23267));
  A2O1A1O1Ixp25_ASAP7_75t_L g23011(.A1(new_n23099), .A2(new_n23090), .B(new_n23187), .C(new_n23182), .D(new_n23265), .Y(new_n23268));
  INVx1_ASAP7_75t_L         g23012(.A(new_n23268), .Y(new_n23269));
  AND2x2_ASAP7_75t_L        g23013(.A(new_n23269), .B(new_n23267), .Y(new_n23270));
  INVx1_ASAP7_75t_L         g23014(.A(new_n23270), .Y(new_n23271));
  O2A1O1Ixp33_ASAP7_75t_L   g23015(.A1(new_n23190), .A2(new_n23191), .B(new_n23196), .C(new_n23271), .Y(new_n23272));
  NOR3xp33_ASAP7_75t_L      g23016(.A(new_n23197), .B(new_n23270), .C(new_n23194), .Y(new_n23273));
  NOR2xp33_ASAP7_75t_L      g23017(.A(new_n23272), .B(new_n23273), .Y(\f[115] ));
  NOR2xp33_ASAP7_75t_L      g23018(.A(new_n9355), .B(new_n13030), .Y(new_n23275));
  INVx1_ASAP7_75t_L         g23019(.A(new_n23275), .Y(new_n23276));
  O2A1O1Ixp33_ASAP7_75t_L   g23020(.A1(new_n12672), .A2(new_n9683), .B(new_n23276), .C(new_n23215), .Y(new_n23277));
  INVx1_ASAP7_75t_L         g23021(.A(new_n23277), .Y(new_n23278));
  INVx1_ASAP7_75t_L         g23022(.A(new_n23212), .Y(new_n23279));
  O2A1O1Ixp33_ASAP7_75t_L   g23023(.A1(new_n12669), .A2(new_n12671), .B(\b[53] ), .C(new_n23275), .Y(new_n23280));
  A2O1A1Ixp33_ASAP7_75t_L   g23024(.A1(new_n13028), .A2(\b[52] ), .B(new_n23211), .C(new_n23280), .Y(new_n23281));
  A2O1A1Ixp33_ASAP7_75t_L   g23025(.A1(new_n23279), .A2(new_n23214), .B(new_n23225), .C(new_n23281), .Y(new_n23282));
  A2O1A1O1Ixp25_ASAP7_75t_L g23026(.A1(new_n13028), .A2(\b[53] ), .B(new_n23275), .C(new_n23214), .D(new_n23282), .Y(new_n23283));
  O2A1O1Ixp33_ASAP7_75t_L   g23027(.A1(new_n23215), .A2(new_n23212), .B(new_n23226), .C(new_n23283), .Y(new_n23284));
  A2O1A1O1Ixp25_ASAP7_75t_L g23028(.A1(new_n13028), .A2(\b[52] ), .B(new_n23211), .C(new_n23280), .D(new_n23283), .Y(new_n23285));
  OAI22xp33_ASAP7_75t_L     g23029(.A1(new_n12320), .A2(new_n9709), .B1(new_n10309), .B2(new_n12318), .Y(new_n23286));
  AOI221xp5_ASAP7_75t_L     g23030(.A1(new_n11995), .A2(\b[56] ), .B1(new_n11997), .B2(new_n11579), .C(new_n23286), .Y(new_n23287));
  XNOR2x2_ASAP7_75t_L       g23031(.A(new_n11987), .B(new_n23287), .Y(new_n23288));
  A2O1A1Ixp33_ASAP7_75t_L   g23032(.A1(new_n23285), .A2(new_n23278), .B(new_n23284), .C(new_n23288), .Y(new_n23289));
  O2A1O1Ixp33_ASAP7_75t_L   g23033(.A1(new_n23280), .A2(new_n23215), .B(new_n23285), .C(new_n23284), .Y(new_n23290));
  INVx1_ASAP7_75t_L         g23034(.A(new_n23288), .Y(new_n23291));
  NAND2xp33_ASAP7_75t_L     g23035(.A(new_n23291), .B(new_n23290), .Y(new_n23292));
  AND2x2_ASAP7_75t_L        g23036(.A(new_n23289), .B(new_n23292), .Y(new_n23293));
  NOR2xp33_ASAP7_75t_L      g23037(.A(new_n10978), .B(new_n11354), .Y(new_n23294));
  AOI221xp5_ASAP7_75t_L     g23038(.A1(\b[59] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[58] ), .C(new_n23294), .Y(new_n23295));
  O2A1O1Ixp33_ASAP7_75t_L   g23039(.A1(new_n11053), .A2(new_n11597), .B(new_n23295), .C(new_n11048), .Y(new_n23296));
  NOR2xp33_ASAP7_75t_L      g23040(.A(new_n11048), .B(new_n23296), .Y(new_n23297));
  O2A1O1Ixp33_ASAP7_75t_L   g23041(.A1(new_n11053), .A2(new_n11597), .B(new_n23295), .C(\a[59] ), .Y(new_n23298));
  NOR2xp33_ASAP7_75t_L      g23042(.A(new_n23298), .B(new_n23297), .Y(new_n23299));
  XOR2x2_ASAP7_75t_L        g23043(.A(new_n23299), .B(new_n23293), .Y(new_n23300));
  NOR3xp33_ASAP7_75t_L      g23044(.A(new_n23300), .B(new_n23233), .C(new_n23229), .Y(new_n23301));
  O2A1O1Ixp33_ASAP7_75t_L   g23045(.A1(new_n23045), .A2(new_n23049), .B(new_n23136), .C(new_n23148), .Y(new_n23302));
  INVx1_ASAP7_75t_L         g23046(.A(new_n23300), .Y(new_n23303));
  O2A1O1Ixp33_ASAP7_75t_L   g23047(.A1(new_n23302), .A2(new_n23228), .B(new_n23234), .C(new_n23303), .Y(new_n23304));
  NOR2xp33_ASAP7_75t_L      g23048(.A(new_n23301), .B(new_n23304), .Y(new_n23305));
  NOR2xp33_ASAP7_75t_L      g23049(.A(new_n12258), .B(new_n10388), .Y(new_n23306));
  AOI221xp5_ASAP7_75t_L     g23050(.A1(new_n10086), .A2(\b[62] ), .B1(new_n11361), .B2(\b[60] ), .C(new_n23306), .Y(new_n23307));
  O2A1O1Ixp33_ASAP7_75t_L   g23051(.A1(new_n10088), .A2(new_n12610), .B(new_n23307), .C(new_n10083), .Y(new_n23308));
  INVx1_ASAP7_75t_L         g23052(.A(new_n23308), .Y(new_n23309));
  O2A1O1Ixp33_ASAP7_75t_L   g23053(.A1(new_n10088), .A2(new_n12610), .B(new_n23307), .C(\a[56] ), .Y(new_n23310));
  A2O1A1Ixp33_ASAP7_75t_L   g23054(.A1(\a[56] ), .A2(new_n23309), .B(new_n23310), .C(new_n23305), .Y(new_n23311));
  INVx1_ASAP7_75t_L         g23055(.A(new_n23310), .Y(new_n23312));
  O2A1O1Ixp33_ASAP7_75t_L   g23056(.A1(new_n23308), .A2(new_n10083), .B(new_n23312), .C(new_n23305), .Y(new_n23313));
  O2A1O1Ixp33_ASAP7_75t_L   g23057(.A1(new_n23245), .A2(new_n23236), .B(new_n23248), .C(new_n23238), .Y(new_n23314));
  NOR2xp33_ASAP7_75t_L      g23058(.A(new_n12956), .B(new_n9440), .Y(new_n23315));
  INVx1_ASAP7_75t_L         g23059(.A(new_n23315), .Y(new_n23316));
  A2O1A1Ixp33_ASAP7_75t_L   g23060(.A1(new_n14444), .A2(new_n12603), .B(new_n12956), .C(new_n23316), .Y(new_n23317));
  O2A1O1Ixp33_ASAP7_75t_L   g23061(.A1(new_n9437), .A2(new_n23315), .B(new_n23317), .C(new_n9099), .Y(new_n23318));
  INVx1_ASAP7_75t_L         g23062(.A(new_n23318), .Y(new_n23319));
  O2A1O1Ixp33_ASAP7_75t_L   g23063(.A1(new_n9104), .A2(new_n13573), .B(new_n23316), .C(\a[53] ), .Y(new_n23320));
  INVx1_ASAP7_75t_L         g23064(.A(new_n23320), .Y(new_n23321));
  NAND2xp33_ASAP7_75t_L     g23065(.A(new_n23321), .B(new_n23319), .Y(new_n23322));
  XNOR2x2_ASAP7_75t_L       g23066(.A(new_n23322), .B(new_n23314), .Y(new_n23323));
  A2O1A1Ixp33_ASAP7_75t_L   g23067(.A1(new_n23311), .A2(new_n23305), .B(new_n23313), .C(new_n23323), .Y(new_n23324));
  AND2x2_ASAP7_75t_L        g23068(.A(new_n23323), .B(new_n23324), .Y(new_n23325));
  A2O1A1O1Ixp25_ASAP7_75t_L g23069(.A1(new_n23311), .A2(new_n23305), .B(new_n23313), .C(new_n23324), .D(new_n23325), .Y(new_n23326));
  A2O1A1O1Ixp25_ASAP7_75t_L g23070(.A1(new_n23164), .A2(new_n23166), .B(new_n23170), .C(new_n23250), .D(new_n23262), .Y(new_n23327));
  AND2x2_ASAP7_75t_L        g23071(.A(new_n23326), .B(new_n23327), .Y(new_n23328));
  O2A1O1Ixp33_ASAP7_75t_L   g23072(.A1(new_n23254), .A2(new_n23251), .B(new_n23263), .C(new_n23326), .Y(new_n23329));
  NOR2xp33_ASAP7_75t_L      g23073(.A(new_n23329), .B(new_n23328), .Y(new_n23330));
  INVx1_ASAP7_75t_L         g23074(.A(new_n23194), .Y(new_n23331));
  A2O1A1Ixp33_ASAP7_75t_L   g23075(.A1(new_n23196), .A2(new_n23331), .B(new_n23271), .C(new_n23269), .Y(new_n23332));
  XOR2x2_ASAP7_75t_L        g23076(.A(new_n23330), .B(new_n23332), .Y(\f[116] ));
  NOR2xp33_ASAP7_75t_L      g23077(.A(new_n12603), .B(new_n10388), .Y(new_n23334));
  AOI221xp5_ASAP7_75t_L     g23078(.A1(new_n10086), .A2(\b[63] ), .B1(new_n11361), .B2(\b[61] ), .C(new_n23334), .Y(new_n23335));
  O2A1O1Ixp33_ASAP7_75t_L   g23079(.A1(new_n10088), .A2(new_n17815), .B(new_n23335), .C(new_n10083), .Y(new_n23336));
  INVx1_ASAP7_75t_L         g23080(.A(new_n23336), .Y(new_n23337));
  O2A1O1Ixp33_ASAP7_75t_L   g23081(.A1(new_n10088), .A2(new_n17815), .B(new_n23335), .C(\a[56] ), .Y(new_n23338));
  AOI21xp33_ASAP7_75t_L     g23082(.A1(new_n23337), .A2(\a[56] ), .B(new_n23338), .Y(new_n23339));
  INVx1_ASAP7_75t_L         g23083(.A(new_n23339), .Y(new_n23340));
  A2O1A1O1Ixp25_ASAP7_75t_L g23084(.A1(new_n23309), .A2(\a[56] ), .B(new_n23310), .C(new_n23305), .D(new_n23304), .Y(new_n23341));
  INVx1_ASAP7_75t_L         g23085(.A(new_n23341), .Y(new_n23342));
  A2O1A1Ixp33_ASAP7_75t_L   g23086(.A1(\a[56] ), .A2(new_n23337), .B(new_n23338), .C(new_n23342), .Y(new_n23343));
  O2A1O1Ixp33_ASAP7_75t_L   g23087(.A1(new_n23145), .A2(new_n23148), .B(new_n23227), .C(new_n23233), .Y(new_n23344));
  O2A1O1Ixp33_ASAP7_75t_L   g23088(.A1(new_n23344), .A2(new_n23303), .B(new_n23311), .C(new_n23340), .Y(new_n23345));
  O2A1O1Ixp33_ASAP7_75t_L   g23089(.A1(new_n9683), .A2(new_n12672), .B(new_n23276), .C(new_n9099), .Y(new_n23346));
  AOI211xp5_ASAP7_75t_L     g23090(.A1(new_n13028), .A2(\b[53] ), .B(new_n23275), .C(\a[53] ), .Y(new_n23347));
  NOR2xp33_ASAP7_75t_L      g23091(.A(new_n23347), .B(new_n23346), .Y(new_n23348));
  NOR2xp33_ASAP7_75t_L      g23092(.A(new_n9683), .B(new_n13030), .Y(new_n23349));
  O2A1O1Ixp33_ASAP7_75t_L   g23093(.A1(new_n12669), .A2(new_n12671), .B(\b[54] ), .C(new_n23349), .Y(new_n23350));
  NAND2xp33_ASAP7_75t_L     g23094(.A(new_n23350), .B(new_n23348), .Y(new_n23351));
  INVx1_ASAP7_75t_L         g23095(.A(new_n23348), .Y(new_n23352));
  A2O1A1Ixp33_ASAP7_75t_L   g23096(.A1(\b[54] ), .A2(new_n13028), .B(new_n23349), .C(new_n23352), .Y(new_n23353));
  AND2x2_ASAP7_75t_L        g23097(.A(new_n23351), .B(new_n23353), .Y(new_n23354));
  INVx1_ASAP7_75t_L         g23098(.A(new_n23354), .Y(new_n23355));
  NOR2xp33_ASAP7_75t_L      g23099(.A(new_n10332), .B(new_n12318), .Y(new_n23356));
  AOI221xp5_ASAP7_75t_L     g23100(.A1(new_n11995), .A2(\b[57] ), .B1(new_n13314), .B2(\b[55] ), .C(new_n23356), .Y(new_n23357));
  O2A1O1Ixp33_ASAP7_75t_L   g23101(.A1(new_n11998), .A2(new_n17096), .B(new_n23357), .C(new_n11987), .Y(new_n23358));
  O2A1O1Ixp33_ASAP7_75t_L   g23102(.A1(new_n11998), .A2(new_n17096), .B(new_n23357), .C(\a[62] ), .Y(new_n23359));
  INVx1_ASAP7_75t_L         g23103(.A(new_n23359), .Y(new_n23360));
  O2A1O1Ixp33_ASAP7_75t_L   g23104(.A1(new_n23358), .A2(new_n11987), .B(new_n23360), .C(new_n23355), .Y(new_n23361));
  INVx1_ASAP7_75t_L         g23105(.A(new_n23361), .Y(new_n23362));
  O2A1O1Ixp33_ASAP7_75t_L   g23106(.A1(new_n23358), .A2(new_n11987), .B(new_n23360), .C(new_n23354), .Y(new_n23363));
  AOI21xp33_ASAP7_75t_L     g23107(.A1(new_n23362), .A2(new_n23354), .B(new_n23363), .Y(new_n23364));
  O2A1O1Ixp33_ASAP7_75t_L   g23108(.A1(new_n23277), .A2(new_n23282), .B(new_n23281), .C(new_n23364), .Y(new_n23365));
  AND2x2_ASAP7_75t_L        g23109(.A(new_n23364), .B(new_n23285), .Y(new_n23366));
  NOR2xp33_ASAP7_75t_L      g23110(.A(new_n23365), .B(new_n23366), .Y(new_n23367));
  NOR2xp33_ASAP7_75t_L      g23111(.A(new_n11303), .B(new_n11354), .Y(new_n23368));
  AOI221xp5_ASAP7_75t_L     g23112(.A1(\b[60] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[59] ), .C(new_n23368), .Y(new_n23369));
  O2A1O1Ixp33_ASAP7_75t_L   g23113(.A1(new_n11053), .A2(new_n11634), .B(new_n23369), .C(new_n11048), .Y(new_n23370));
  INVx1_ASAP7_75t_L         g23114(.A(new_n23370), .Y(new_n23371));
  O2A1O1Ixp33_ASAP7_75t_L   g23115(.A1(new_n11053), .A2(new_n11634), .B(new_n23369), .C(\a[59] ), .Y(new_n23372));
  A2O1A1Ixp33_ASAP7_75t_L   g23116(.A1(new_n23371), .A2(\a[59] ), .B(new_n23372), .C(new_n23367), .Y(new_n23373));
  INVx1_ASAP7_75t_L         g23117(.A(new_n23372), .Y(new_n23374));
  O2A1O1Ixp33_ASAP7_75t_L   g23118(.A1(new_n11048), .A2(new_n23370), .B(new_n23374), .C(new_n23367), .Y(new_n23375));
  A2O1A1Ixp33_ASAP7_75t_L   g23119(.A1(new_n23285), .A2(new_n23278), .B(new_n23284), .C(new_n23291), .Y(new_n23376));
  A2O1A1Ixp33_ASAP7_75t_L   g23120(.A1(new_n23292), .A2(new_n23289), .B(new_n23299), .C(new_n23376), .Y(new_n23377));
  A2O1A1Ixp33_ASAP7_75t_L   g23121(.A1(new_n23373), .A2(new_n23367), .B(new_n23375), .C(new_n23377), .Y(new_n23378));
  AO21x2_ASAP7_75t_L        g23122(.A1(new_n23367), .A2(new_n23373), .B(new_n23375), .Y(new_n23379));
  O2A1O1Ixp33_ASAP7_75t_L   g23123(.A1(new_n23293), .A2(new_n23299), .B(new_n23376), .C(new_n23379), .Y(new_n23380));
  A2O1A1O1Ixp25_ASAP7_75t_L g23124(.A1(new_n23373), .A2(new_n23367), .B(new_n23375), .C(new_n23378), .D(new_n23380), .Y(new_n23381));
  A2O1A1Ixp33_ASAP7_75t_L   g23125(.A1(new_n23343), .A2(new_n23340), .B(new_n23345), .C(new_n23381), .Y(new_n23382));
  A2O1A1O1Ixp25_ASAP7_75t_L g23126(.A1(new_n23337), .A2(\a[56] ), .B(new_n23338), .C(new_n23343), .D(new_n23345), .Y(new_n23383));
  A2O1A1Ixp33_ASAP7_75t_L   g23127(.A1(new_n23379), .A2(new_n23378), .B(new_n23380), .C(new_n23383), .Y(new_n23384));
  NAND2xp33_ASAP7_75t_L     g23128(.A(new_n23382), .B(new_n23384), .Y(new_n23385));
  INVx1_ASAP7_75t_L         g23129(.A(new_n23385), .Y(new_n23386));
  A2O1A1O1Ixp25_ASAP7_75t_L g23130(.A1(new_n23319), .A2(new_n23321), .B(new_n23314), .C(new_n23324), .D(new_n23386), .Y(new_n23387));
  A2O1A1Ixp33_ASAP7_75t_L   g23131(.A1(new_n23319), .A2(new_n23321), .B(new_n23314), .C(new_n23324), .Y(new_n23388));
  NOR2xp33_ASAP7_75t_L      g23132(.A(new_n23388), .B(new_n23385), .Y(new_n23389));
  NOR2xp33_ASAP7_75t_L      g23133(.A(new_n23389), .B(new_n23387), .Y(new_n23390));
  A2O1A1Ixp33_ASAP7_75t_L   g23134(.A1(new_n23332), .A2(new_n23330), .B(new_n23329), .C(new_n23390), .Y(new_n23391));
  INVx1_ASAP7_75t_L         g23135(.A(new_n23391), .Y(new_n23392));
  INVx1_ASAP7_75t_L         g23136(.A(new_n23107), .Y(new_n23393));
  A2O1A1Ixp33_ASAP7_75t_L   g23137(.A1(new_n23110), .A2(new_n23393), .B(new_n23190), .C(new_n23196), .Y(new_n23394));
  A2O1A1Ixp33_ASAP7_75t_L   g23138(.A1(new_n23394), .A2(new_n23270), .B(new_n23268), .C(new_n23330), .Y(new_n23395));
  A2O1A1Ixp33_ASAP7_75t_L   g23139(.A1(new_n23263), .A2(new_n23253), .B(new_n23326), .C(new_n23395), .Y(new_n23396));
  NOR2xp33_ASAP7_75t_L      g23140(.A(new_n23390), .B(new_n23396), .Y(new_n23397));
  NOR2xp33_ASAP7_75t_L      g23141(.A(new_n23392), .B(new_n23397), .Y(\f[117] ));
  A2O1A1Ixp33_ASAP7_75t_L   g23142(.A1(new_n23236), .A2(new_n23202), .B(new_n23247), .C(new_n23322), .Y(new_n23399));
  NOR2xp33_ASAP7_75t_L      g23143(.A(new_n11591), .B(new_n11354), .Y(new_n23400));
  AOI221xp5_ASAP7_75t_L     g23144(.A1(\b[61] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[60] ), .C(new_n23400), .Y(new_n23401));
  O2A1O1Ixp33_ASAP7_75t_L   g23145(.A1(new_n11053), .A2(new_n14764), .B(new_n23401), .C(new_n11048), .Y(new_n23402));
  O2A1O1Ixp33_ASAP7_75t_L   g23146(.A1(new_n11053), .A2(new_n14764), .B(new_n23401), .C(\a[59] ), .Y(new_n23403));
  INVx1_ASAP7_75t_L         g23147(.A(new_n23403), .Y(new_n23404));
  OA21x2_ASAP7_75t_L        g23148(.A1(new_n11048), .A2(new_n23402), .B(new_n23404), .Y(new_n23405));
  NOR2xp33_ASAP7_75t_L      g23149(.A(new_n9709), .B(new_n13030), .Y(new_n23406));
  O2A1O1Ixp33_ASAP7_75t_L   g23150(.A1(new_n12669), .A2(new_n12671), .B(\b[55] ), .C(new_n23406), .Y(new_n23407));
  INVx1_ASAP7_75t_L         g23151(.A(new_n23407), .Y(new_n23408));
  O2A1O1Ixp33_ASAP7_75t_L   g23152(.A1(\a[53] ), .A2(new_n23280), .B(new_n23353), .C(new_n23408), .Y(new_n23409));
  INVx1_ASAP7_75t_L         g23153(.A(new_n23409), .Y(new_n23410));
  INVx1_ASAP7_75t_L         g23154(.A(new_n23350), .Y(new_n23411));
  O2A1O1Ixp33_ASAP7_75t_L   g23155(.A1(new_n9683), .A2(new_n12672), .B(new_n23276), .C(\a[53] ), .Y(new_n23412));
  O2A1O1Ixp33_ASAP7_75t_L   g23156(.A1(new_n23347), .A2(new_n23346), .B(new_n23411), .C(new_n23412), .Y(new_n23413));
  A2O1A1Ixp33_ASAP7_75t_L   g23157(.A1(new_n13028), .A2(\b[55] ), .B(new_n23406), .C(new_n23413), .Y(new_n23414));
  NAND2xp33_ASAP7_75t_L     g23158(.A(new_n23414), .B(new_n23410), .Y(new_n23415));
  NOR2xp33_ASAP7_75t_L      g23159(.A(new_n10978), .B(new_n12318), .Y(new_n23416));
  AOI221xp5_ASAP7_75t_L     g23160(.A1(new_n11995), .A2(\b[58] ), .B1(new_n13314), .B2(\b[56] ), .C(new_n23416), .Y(new_n23417));
  INVx1_ASAP7_75t_L         g23161(.A(new_n23417), .Y(new_n23418));
  A2O1A1Ixp33_ASAP7_75t_L   g23162(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n23417), .Y(new_n23419));
  O2A1O1Ixp33_ASAP7_75t_L   g23163(.A1(new_n23418), .A2(new_n11314), .B(new_n23419), .C(new_n11987), .Y(new_n23420));
  O2A1O1Ixp33_ASAP7_75t_L   g23164(.A1(new_n11998), .A2(new_n20073), .B(new_n23417), .C(\a[62] ), .Y(new_n23421));
  NOR2xp33_ASAP7_75t_L      g23165(.A(new_n23420), .B(new_n23421), .Y(new_n23422));
  NOR2xp33_ASAP7_75t_L      g23166(.A(new_n23415), .B(new_n23422), .Y(new_n23423));
  INVx1_ASAP7_75t_L         g23167(.A(new_n23423), .Y(new_n23424));
  NAND2xp33_ASAP7_75t_L     g23168(.A(new_n23415), .B(new_n23422), .Y(new_n23425));
  NAND2xp33_ASAP7_75t_L     g23169(.A(new_n23425), .B(new_n23424), .Y(new_n23426));
  O2A1O1Ixp33_ASAP7_75t_L   g23170(.A1(new_n23285), .A2(new_n23364), .B(new_n23362), .C(new_n23426), .Y(new_n23427));
  INVx1_ASAP7_75t_L         g23171(.A(new_n23426), .Y(new_n23428));
  O2A1O1Ixp33_ASAP7_75t_L   g23172(.A1(new_n23285), .A2(new_n23364), .B(new_n23362), .C(new_n23428), .Y(new_n23429));
  INVx1_ASAP7_75t_L         g23173(.A(new_n23429), .Y(new_n23430));
  O2A1O1Ixp33_ASAP7_75t_L   g23174(.A1(new_n23426), .A2(new_n23427), .B(new_n23430), .C(new_n23405), .Y(new_n23431));
  OAI21xp33_ASAP7_75t_L     g23175(.A1(new_n23426), .A2(new_n23427), .B(new_n23405), .Y(new_n23432));
  O2A1O1Ixp33_ASAP7_75t_L   g23176(.A1(new_n23361), .A2(new_n23365), .B(new_n23426), .C(new_n23432), .Y(new_n23433));
  NOR2xp33_ASAP7_75t_L      g23177(.A(new_n23433), .B(new_n23431), .Y(new_n23434));
  INVx1_ASAP7_75t_L         g23178(.A(new_n23434), .Y(new_n23435));
  AO21x2_ASAP7_75t_L        g23179(.A1(new_n23373), .A2(new_n23378), .B(new_n23435), .Y(new_n23436));
  NAND3xp33_ASAP7_75t_L     g23180(.A(new_n23435), .B(new_n23378), .C(new_n23373), .Y(new_n23437));
  AND2x2_ASAP7_75t_L        g23181(.A(new_n23437), .B(new_n23436), .Y(new_n23438));
  INVx1_ASAP7_75t_L         g23182(.A(new_n23438), .Y(new_n23439));
  AOI22xp33_ASAP7_75t_L     g23183(.A1(new_n10080), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n11361), .Y(new_n23440));
  O2A1O1Ixp33_ASAP7_75t_L   g23184(.A1(new_n10088), .A2(new_n12993), .B(new_n23440), .C(new_n10083), .Y(new_n23441));
  O2A1O1Ixp33_ASAP7_75t_L   g23185(.A1(new_n10088), .A2(new_n12993), .B(new_n23440), .C(\a[56] ), .Y(new_n23442));
  INVx1_ASAP7_75t_L         g23186(.A(new_n23442), .Y(new_n23443));
  O2A1O1Ixp33_ASAP7_75t_L   g23187(.A1(new_n23441), .A2(new_n10083), .B(new_n23443), .C(new_n23439), .Y(new_n23444));
  INVx1_ASAP7_75t_L         g23188(.A(new_n23444), .Y(new_n23445));
  O2A1O1Ixp33_ASAP7_75t_L   g23189(.A1(new_n23441), .A2(new_n10083), .B(new_n23443), .C(new_n23438), .Y(new_n23446));
  A2O1A1Ixp33_ASAP7_75t_L   g23190(.A1(\a[56] ), .A2(new_n23337), .B(new_n23338), .C(new_n23341), .Y(new_n23447));
  AOI21xp33_ASAP7_75t_L     g23191(.A1(new_n23445), .A2(new_n23438), .B(new_n23446), .Y(new_n23448));
  A2O1A1O1Ixp25_ASAP7_75t_L g23192(.A1(new_n23447), .A2(new_n23341), .B(new_n23381), .C(new_n23343), .D(new_n23448), .Y(new_n23449));
  INVx1_ASAP7_75t_L         g23193(.A(new_n23449), .Y(new_n23450));
  O2A1O1Ixp33_ASAP7_75t_L   g23194(.A1(new_n23383), .A2(new_n23381), .B(new_n23343), .C(new_n23449), .Y(new_n23451));
  A2O1A1O1Ixp25_ASAP7_75t_L g23195(.A1(new_n23445), .A2(new_n23438), .B(new_n23446), .C(new_n23450), .D(new_n23451), .Y(new_n23452));
  A2O1A1O1Ixp25_ASAP7_75t_L g23196(.A1(new_n23324), .A2(new_n23399), .B(new_n23386), .C(new_n23391), .D(new_n23452), .Y(new_n23453));
  INVx1_ASAP7_75t_L         g23197(.A(new_n23452), .Y(new_n23454));
  A2O1A1Ixp33_ASAP7_75t_L   g23198(.A1(new_n23324), .A2(new_n23399), .B(new_n23386), .C(new_n23391), .Y(new_n23455));
  NOR2xp33_ASAP7_75t_L      g23199(.A(new_n23454), .B(new_n23455), .Y(new_n23456));
  NOR2xp33_ASAP7_75t_L      g23200(.A(new_n23453), .B(new_n23456), .Y(\f[118] ));
  NOR2xp33_ASAP7_75t_L      g23201(.A(new_n10309), .B(new_n13030), .Y(new_n23458));
  INVx1_ASAP7_75t_L         g23202(.A(new_n23458), .Y(new_n23459));
  O2A1O1Ixp33_ASAP7_75t_L   g23203(.A1(new_n12672), .A2(new_n10332), .B(new_n23459), .C(new_n23408), .Y(new_n23460));
  NOR2xp33_ASAP7_75t_L      g23204(.A(new_n23408), .B(new_n23460), .Y(new_n23461));
  O2A1O1Ixp33_ASAP7_75t_L   g23205(.A1(new_n12672), .A2(new_n10332), .B(new_n23459), .C(new_n23407), .Y(new_n23462));
  NOR2xp33_ASAP7_75t_L      g23206(.A(new_n11303), .B(new_n12318), .Y(new_n23463));
  AOI221xp5_ASAP7_75t_L     g23207(.A1(new_n11995), .A2(\b[59] ), .B1(new_n13314), .B2(\b[57] ), .C(new_n23463), .Y(new_n23464));
  O2A1O1Ixp33_ASAP7_75t_L   g23208(.A1(new_n11998), .A2(new_n11597), .B(new_n23464), .C(new_n11987), .Y(new_n23465));
  O2A1O1Ixp33_ASAP7_75t_L   g23209(.A1(new_n11998), .A2(new_n11597), .B(new_n23464), .C(\a[62] ), .Y(new_n23466));
  INVx1_ASAP7_75t_L         g23210(.A(new_n23466), .Y(new_n23467));
  INVx1_ASAP7_75t_L         g23211(.A(new_n23460), .Y(new_n23468));
  A2O1A1O1Ixp25_ASAP7_75t_L g23212(.A1(new_n13028), .A2(\b[56] ), .B(new_n23458), .C(new_n23468), .D(new_n23461), .Y(new_n23469));
  O2A1O1Ixp33_ASAP7_75t_L   g23213(.A1(new_n11987), .A2(new_n23465), .B(new_n23467), .C(new_n23469), .Y(new_n23470));
  INVx1_ASAP7_75t_L         g23214(.A(new_n23470), .Y(new_n23471));
  O2A1O1Ixp33_ASAP7_75t_L   g23215(.A1(new_n11987), .A2(new_n23465), .B(new_n23467), .C(new_n23470), .Y(new_n23472));
  O2A1O1Ixp33_ASAP7_75t_L   g23216(.A1(new_n23461), .A2(new_n23462), .B(new_n23471), .C(new_n23472), .Y(new_n23473));
  O2A1O1Ixp33_ASAP7_75t_L   g23217(.A1(new_n23420), .A2(new_n23421), .B(new_n23414), .C(new_n23409), .Y(new_n23474));
  NAND2xp33_ASAP7_75t_L     g23218(.A(new_n23474), .B(new_n23473), .Y(new_n23475));
  O2A1O1Ixp33_ASAP7_75t_L   g23219(.A1(new_n23408), .A2(new_n23413), .B(new_n23424), .C(new_n23473), .Y(new_n23476));
  INVx1_ASAP7_75t_L         g23220(.A(new_n23476), .Y(new_n23477));
  AND2x2_ASAP7_75t_L        g23221(.A(new_n23475), .B(new_n23477), .Y(new_n23478));
  NOR2xp33_ASAP7_75t_L      g23222(.A(new_n11626), .B(new_n11354), .Y(new_n23479));
  AOI221xp5_ASAP7_75t_L     g23223(.A1(\b[62] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[61] ), .C(new_n23479), .Y(new_n23480));
  O2A1O1Ixp33_ASAP7_75t_L   g23224(.A1(new_n11053), .A2(new_n12610), .B(new_n23480), .C(new_n11048), .Y(new_n23481));
  INVx1_ASAP7_75t_L         g23225(.A(new_n23481), .Y(new_n23482));
  O2A1O1Ixp33_ASAP7_75t_L   g23226(.A1(new_n11053), .A2(new_n12610), .B(new_n23480), .C(\a[59] ), .Y(new_n23483));
  A2O1A1Ixp33_ASAP7_75t_L   g23227(.A1(\a[59] ), .A2(new_n23482), .B(new_n23483), .C(new_n23478), .Y(new_n23484));
  NAND2xp33_ASAP7_75t_L     g23228(.A(new_n23478), .B(new_n23484), .Y(new_n23485));
  A2O1A1Ixp33_ASAP7_75t_L   g23229(.A1(new_n23482), .A2(\a[59] ), .B(new_n23483), .C(new_n23484), .Y(new_n23486));
  INVx1_ASAP7_75t_L         g23230(.A(new_n23486), .Y(new_n23487));
  INVx1_ASAP7_75t_L         g23231(.A(new_n23427), .Y(new_n23488));
  NOR2xp33_ASAP7_75t_L      g23232(.A(new_n12956), .B(new_n10390), .Y(new_n23489));
  INVx1_ASAP7_75t_L         g23233(.A(new_n23489), .Y(new_n23490));
  A2O1A1Ixp33_ASAP7_75t_L   g23234(.A1(new_n14444), .A2(new_n12603), .B(new_n12956), .C(new_n23490), .Y(new_n23491));
  O2A1O1Ixp33_ASAP7_75t_L   g23235(.A1(new_n10386), .A2(new_n23489), .B(new_n23491), .C(new_n10083), .Y(new_n23492));
  O2A1O1Ixp33_ASAP7_75t_L   g23236(.A1(new_n10088), .A2(new_n13573), .B(new_n23490), .C(\a[56] ), .Y(new_n23493));
  NOR2xp33_ASAP7_75t_L      g23237(.A(new_n23493), .B(new_n23492), .Y(new_n23494));
  A2O1A1O1Ixp25_ASAP7_75t_L g23238(.A1(new_n23426), .A2(new_n23430), .B(new_n23405), .C(new_n23488), .D(new_n23494), .Y(new_n23495));
  INVx1_ASAP7_75t_L         g23239(.A(new_n23495), .Y(new_n23496));
  O2A1O1Ixp33_ASAP7_75t_L   g23240(.A1(new_n23361), .A2(new_n23365), .B(new_n23428), .C(new_n23431), .Y(new_n23497));
  NAND2xp33_ASAP7_75t_L     g23241(.A(new_n23494), .B(new_n23497), .Y(new_n23498));
  AND2x2_ASAP7_75t_L        g23242(.A(new_n23496), .B(new_n23498), .Y(new_n23499));
  A2O1A1Ixp33_ASAP7_75t_L   g23243(.A1(new_n23484), .A2(new_n23478), .B(new_n23487), .C(new_n23499), .Y(new_n23500));
  INVx1_ASAP7_75t_L         g23244(.A(new_n23500), .Y(new_n23501));
  NAND2xp33_ASAP7_75t_L     g23245(.A(new_n23499), .B(new_n23500), .Y(new_n23502));
  A2O1A1Ixp33_ASAP7_75t_L   g23246(.A1(new_n23486), .A2(new_n23485), .B(new_n23501), .C(new_n23502), .Y(new_n23503));
  A2O1A1Ixp33_ASAP7_75t_L   g23247(.A1(new_n23378), .A2(new_n23373), .B(new_n23435), .C(new_n23445), .Y(new_n23504));
  NOR2xp33_ASAP7_75t_L      g23248(.A(new_n23503), .B(new_n23504), .Y(new_n23505));
  INVx1_ASAP7_75t_L         g23249(.A(new_n23503), .Y(new_n23506));
  A2O1A1O1Ixp25_ASAP7_75t_L g23250(.A1(new_n23378), .A2(new_n23373), .B(new_n23435), .C(new_n23445), .D(new_n23506), .Y(new_n23507));
  NOR2xp33_ASAP7_75t_L      g23251(.A(new_n23507), .B(new_n23505), .Y(new_n23508));
  INVx1_ASAP7_75t_L         g23252(.A(new_n23387), .Y(new_n23509));
  A2O1A1Ixp33_ASAP7_75t_L   g23253(.A1(new_n23391), .A2(new_n23509), .B(new_n23452), .C(new_n23450), .Y(new_n23510));
  XOR2x2_ASAP7_75t_L        g23254(.A(new_n23508), .B(new_n23510), .Y(\f[119] ));
  NOR2xp33_ASAP7_75t_L      g23255(.A(new_n10332), .B(new_n13030), .Y(new_n23512));
  INVx1_ASAP7_75t_L         g23256(.A(new_n23512), .Y(new_n23513));
  O2A1O1Ixp33_ASAP7_75t_L   g23257(.A1(new_n10978), .A2(new_n12672), .B(new_n23513), .C(\a[56] ), .Y(new_n23514));
  O2A1O1Ixp33_ASAP7_75t_L   g23258(.A1(new_n10978), .A2(new_n12672), .B(new_n23513), .C(new_n10083), .Y(new_n23515));
  INVx1_ASAP7_75t_L         g23259(.A(new_n23515), .Y(new_n23516));
  O2A1O1Ixp33_ASAP7_75t_L   g23260(.A1(\a[56] ), .A2(new_n23514), .B(new_n23516), .C(new_n23407), .Y(new_n23517));
  INVx1_ASAP7_75t_L         g23261(.A(new_n23517), .Y(new_n23518));
  O2A1O1Ixp33_ASAP7_75t_L   g23262(.A1(\a[56] ), .A2(new_n23514), .B(new_n23516), .C(new_n23408), .Y(new_n23519));
  A2O1A1O1Ixp25_ASAP7_75t_L g23263(.A1(new_n13028), .A2(\b[55] ), .B(new_n23406), .C(new_n23518), .D(new_n23519), .Y(new_n23520));
  A2O1A1O1Ixp25_ASAP7_75t_L g23264(.A1(new_n13028), .A2(\b[56] ), .B(new_n23458), .C(new_n23407), .D(new_n23470), .Y(new_n23521));
  NAND2xp33_ASAP7_75t_L     g23265(.A(new_n23520), .B(new_n23521), .Y(new_n23522));
  O2A1O1Ixp33_ASAP7_75t_L   g23266(.A1(new_n12669), .A2(new_n12671), .B(\b[56] ), .C(new_n23458), .Y(new_n23523));
  O2A1O1Ixp33_ASAP7_75t_L   g23267(.A1(new_n23408), .A2(new_n23523), .B(new_n23471), .C(new_n23520), .Y(new_n23524));
  INVx1_ASAP7_75t_L         g23268(.A(new_n23524), .Y(new_n23525));
  AND2x2_ASAP7_75t_L        g23269(.A(new_n23522), .B(new_n23525), .Y(new_n23526));
  OAI22xp33_ASAP7_75t_L     g23270(.A1(new_n12320), .A2(new_n11303), .B1(new_n11591), .B2(new_n12318), .Y(new_n23527));
  AOI221xp5_ASAP7_75t_L     g23271(.A1(new_n11995), .A2(\b[60] ), .B1(new_n11997), .B2(new_n13839), .C(new_n23527), .Y(new_n23528));
  XNOR2x2_ASAP7_75t_L       g23272(.A(new_n11987), .B(new_n23528), .Y(new_n23529));
  INVx1_ASAP7_75t_L         g23273(.A(new_n23529), .Y(new_n23530));
  A2O1A1O1Ixp25_ASAP7_75t_L g23274(.A1(new_n23482), .A2(\a[59] ), .B(new_n23483), .C(new_n23475), .D(new_n23476), .Y(new_n23531));
  INVx1_ASAP7_75t_L         g23275(.A(new_n23531), .Y(new_n23532));
  NOR2xp33_ASAP7_75t_L      g23276(.A(new_n12258), .B(new_n11354), .Y(new_n23533));
  AOI221xp5_ASAP7_75t_L     g23277(.A1(\b[63] ), .A2(new_n11051), .B1(new_n11045), .B2(\b[62] ), .C(new_n23533), .Y(new_n23534));
  O2A1O1Ixp33_ASAP7_75t_L   g23278(.A1(new_n11053), .A2(new_n17815), .B(new_n23534), .C(new_n11048), .Y(new_n23535));
  O2A1O1Ixp33_ASAP7_75t_L   g23279(.A1(new_n11053), .A2(new_n17815), .B(new_n23534), .C(\a[59] ), .Y(new_n23536));
  INVx1_ASAP7_75t_L         g23280(.A(new_n23536), .Y(new_n23537));
  O2A1O1Ixp33_ASAP7_75t_L   g23281(.A1(new_n23535), .A2(new_n11048), .B(new_n23537), .C(new_n23531), .Y(new_n23538));
  INVx1_ASAP7_75t_L         g23282(.A(new_n23538), .Y(new_n23539));
  O2A1O1Ixp33_ASAP7_75t_L   g23283(.A1(new_n23535), .A2(new_n11048), .B(new_n23537), .C(new_n23532), .Y(new_n23540));
  O2A1O1Ixp33_ASAP7_75t_L   g23284(.A1(new_n23473), .A2(new_n23474), .B(new_n23484), .C(new_n23538), .Y(new_n23541));
  INVx1_ASAP7_75t_L         g23285(.A(new_n23526), .Y(new_n23542));
  NOR2xp33_ASAP7_75t_L      g23286(.A(new_n23529), .B(new_n23542), .Y(new_n23543));
  INVx1_ASAP7_75t_L         g23287(.A(new_n23543), .Y(new_n23544));
  NAND2xp33_ASAP7_75t_L     g23288(.A(new_n23529), .B(new_n23542), .Y(new_n23545));
  OAI211xp5_ASAP7_75t_L     g23289(.A1(new_n23540), .A2(new_n23541), .B(new_n23544), .C(new_n23545), .Y(new_n23546));
  A2O1A1Ixp33_ASAP7_75t_L   g23290(.A1(new_n23539), .A2(new_n23532), .B(new_n23540), .C(new_n23546), .Y(new_n23547));
  A2O1A1Ixp33_ASAP7_75t_L   g23291(.A1(new_n23525), .A2(new_n23522), .B(new_n23530), .C(new_n23546), .Y(new_n23548));
  A2O1A1Ixp33_ASAP7_75t_L   g23292(.A1(new_n23526), .A2(new_n23530), .B(new_n23548), .C(new_n23547), .Y(new_n23549));
  NOR3xp33_ASAP7_75t_L      g23293(.A(new_n23549), .B(new_n23501), .C(new_n23495), .Y(new_n23550));
  A2O1A1O1Ixp25_ASAP7_75t_L g23294(.A1(new_n23478), .A2(new_n23484), .B(new_n23487), .C(new_n23498), .D(new_n23495), .Y(new_n23551));
  O2A1O1Ixp33_ASAP7_75t_L   g23295(.A1(new_n23543), .A2(new_n23548), .B(new_n23547), .C(new_n23551), .Y(new_n23552));
  NOR2xp33_ASAP7_75t_L      g23296(.A(new_n23552), .B(new_n23550), .Y(new_n23553));
  A2O1A1Ixp33_ASAP7_75t_L   g23297(.A1(new_n23510), .A2(new_n23508), .B(new_n23507), .C(new_n23553), .Y(new_n23554));
  INVx1_ASAP7_75t_L         g23298(.A(new_n23554), .Y(new_n23555));
  AOI211xp5_ASAP7_75t_L     g23299(.A1(new_n23510), .A2(new_n23508), .B(new_n23553), .C(new_n23507), .Y(new_n23556));
  NOR2xp33_ASAP7_75t_L      g23300(.A(new_n23556), .B(new_n23555), .Y(\f[120] ));
  INVx1_ASAP7_75t_L         g23301(.A(new_n23552), .Y(new_n23558));
  O2A1O1Ixp33_ASAP7_75t_L   g23302(.A1(new_n23449), .A2(new_n23453), .B(new_n23508), .C(new_n23507), .Y(new_n23559));
  NOR2xp33_ASAP7_75t_L      g23303(.A(new_n10978), .B(new_n13030), .Y(new_n23560));
  O2A1O1Ixp33_ASAP7_75t_L   g23304(.A1(new_n10083), .A2(new_n23515), .B(new_n23408), .C(new_n23514), .Y(new_n23561));
  A2O1A1Ixp33_ASAP7_75t_L   g23305(.A1(new_n13028), .A2(\b[58] ), .B(new_n23560), .C(new_n23561), .Y(new_n23562));
  INVx1_ASAP7_75t_L         g23306(.A(new_n23514), .Y(new_n23563));
  O2A1O1Ixp33_ASAP7_75t_L   g23307(.A1(new_n12669), .A2(new_n12671), .B(\b[58] ), .C(new_n23560), .Y(new_n23564));
  INVx1_ASAP7_75t_L         g23308(.A(new_n23564), .Y(new_n23565));
  A2O1A1O1Ixp25_ASAP7_75t_L g23309(.A1(\a[56] ), .A2(new_n23516), .B(new_n23407), .C(new_n23563), .D(new_n23565), .Y(new_n23566));
  INVx1_ASAP7_75t_L         g23310(.A(new_n23566), .Y(new_n23567));
  NAND2xp33_ASAP7_75t_L     g23311(.A(\b[61] ), .B(new_n11995), .Y(new_n23568));
  OAI221xp5_ASAP7_75t_L     g23312(.A1(new_n12318), .A2(new_n11626), .B1(new_n11591), .B2(new_n12320), .C(new_n23568), .Y(new_n23569));
  AOI21xp33_ASAP7_75t_L     g23313(.A1(new_n12269), .A2(new_n11997), .B(new_n23569), .Y(new_n23570));
  NAND2xp33_ASAP7_75t_L     g23314(.A(\a[62] ), .B(new_n23570), .Y(new_n23571));
  A2O1A1Ixp33_ASAP7_75t_L   g23315(.A1(new_n12269), .A2(new_n11997), .B(new_n23569), .C(new_n11987), .Y(new_n23572));
  NAND2xp33_ASAP7_75t_L     g23316(.A(new_n23572), .B(new_n23571), .Y(new_n23573));
  NAND3xp33_ASAP7_75t_L     g23317(.A(new_n23573), .B(new_n23567), .C(new_n23562), .Y(new_n23574));
  AO21x2_ASAP7_75t_L        g23318(.A1(new_n23562), .A2(new_n23567), .B(new_n23573), .Y(new_n23575));
  AND2x2_ASAP7_75t_L        g23319(.A(new_n23574), .B(new_n23575), .Y(new_n23576));
  INVx1_ASAP7_75t_L         g23320(.A(new_n23576), .Y(new_n23577));
  O2A1O1Ixp33_ASAP7_75t_L   g23321(.A1(new_n23542), .A2(new_n23529), .B(new_n23525), .C(new_n23577), .Y(new_n23578));
  A2O1A1Ixp33_ASAP7_75t_L   g23322(.A1(new_n23471), .A2(new_n23468), .B(new_n23520), .C(new_n23544), .Y(new_n23579));
  NOR2xp33_ASAP7_75t_L      g23323(.A(new_n23576), .B(new_n23579), .Y(new_n23580));
  NOR2xp33_ASAP7_75t_L      g23324(.A(new_n23578), .B(new_n23580), .Y(new_n23581));
  OAI22xp33_ASAP7_75t_L     g23325(.A1(new_n11352), .A2(new_n12956), .B1(new_n12603), .B2(new_n11354), .Y(new_n23582));
  INVx1_ASAP7_75t_L         g23326(.A(new_n23582), .Y(new_n23583));
  O2A1O1Ixp33_ASAP7_75t_L   g23327(.A1(new_n11053), .A2(new_n12993), .B(new_n23583), .C(new_n11048), .Y(new_n23584));
  INVx1_ASAP7_75t_L         g23328(.A(new_n23584), .Y(new_n23585));
  O2A1O1Ixp33_ASAP7_75t_L   g23329(.A1(new_n11053), .A2(new_n12993), .B(new_n23583), .C(\a[59] ), .Y(new_n23586));
  A2O1A1Ixp33_ASAP7_75t_L   g23330(.A1(\a[59] ), .A2(new_n23585), .B(new_n23586), .C(new_n23581), .Y(new_n23587));
  INVx1_ASAP7_75t_L         g23331(.A(new_n12990), .Y(new_n23588));
  O2A1O1Ixp33_ASAP7_75t_L   g23332(.A1(new_n12987), .A2(new_n23588), .B(new_n11351), .C(new_n23582), .Y(new_n23589));
  NAND2xp33_ASAP7_75t_L     g23333(.A(\a[59] ), .B(new_n23589), .Y(new_n23590));
  O2A1O1Ixp33_ASAP7_75t_L   g23334(.A1(new_n23589), .A2(new_n23584), .B(new_n23590), .C(new_n23581), .Y(new_n23591));
  AOI21xp33_ASAP7_75t_L     g23335(.A1(new_n23587), .A2(new_n23581), .B(new_n23591), .Y(new_n23592));
  NAND3xp33_ASAP7_75t_L     g23336(.A(new_n23592), .B(new_n23546), .C(new_n23539), .Y(new_n23593));
  A2O1A1Ixp33_ASAP7_75t_L   g23337(.A1(new_n23539), .A2(new_n23532), .B(new_n23540), .C(new_n23545), .Y(new_n23594));
  O2A1O1Ixp33_ASAP7_75t_L   g23338(.A1(new_n23543), .A2(new_n23594), .B(new_n23539), .C(new_n23592), .Y(new_n23595));
  INVx1_ASAP7_75t_L         g23339(.A(new_n23595), .Y(new_n23596));
  AND2x2_ASAP7_75t_L        g23340(.A(new_n23593), .B(new_n23596), .Y(new_n23597));
  INVx1_ASAP7_75t_L         g23341(.A(new_n23597), .Y(new_n23598));
  O2A1O1Ixp33_ASAP7_75t_L   g23342(.A1(new_n23550), .A2(new_n23559), .B(new_n23558), .C(new_n23598), .Y(new_n23599));
  NOR3xp33_ASAP7_75t_L      g23343(.A(new_n23555), .B(new_n23597), .C(new_n23552), .Y(new_n23600));
  NOR2xp33_ASAP7_75t_L      g23344(.A(new_n23599), .B(new_n23600), .Y(\f[121] ));
  NOR2xp33_ASAP7_75t_L      g23345(.A(new_n11303), .B(new_n13030), .Y(new_n23602));
  INVx1_ASAP7_75t_L         g23346(.A(new_n23602), .Y(new_n23603));
  O2A1O1Ixp33_ASAP7_75t_L   g23347(.A1(new_n12672), .A2(new_n11591), .B(new_n23603), .C(new_n23565), .Y(new_n23604));
  INVx1_ASAP7_75t_L         g23348(.A(new_n23604), .Y(new_n23605));
  O2A1O1Ixp33_ASAP7_75t_L   g23349(.A1(new_n12669), .A2(new_n12671), .B(\b[59] ), .C(new_n23602), .Y(new_n23606));
  A2O1A1Ixp33_ASAP7_75t_L   g23350(.A1(new_n13028), .A2(\b[58] ), .B(new_n23560), .C(new_n23606), .Y(new_n23607));
  A2O1A1Ixp33_ASAP7_75t_L   g23351(.A1(new_n23573), .A2(new_n23562), .B(new_n23566), .C(new_n23607), .Y(new_n23608));
  A2O1A1O1Ixp25_ASAP7_75t_L g23352(.A1(new_n13028), .A2(\b[59] ), .B(new_n23602), .C(new_n23564), .D(new_n23608), .Y(new_n23609));
  O2A1O1Ixp33_ASAP7_75t_L   g23353(.A1(new_n23565), .A2(new_n23561), .B(new_n23574), .C(new_n23609), .Y(new_n23610));
  A2O1A1O1Ixp25_ASAP7_75t_L g23354(.A1(new_n13028), .A2(\b[58] ), .B(new_n23560), .C(new_n23606), .D(new_n23609), .Y(new_n23611));
  NOR2xp33_ASAP7_75t_L      g23355(.A(new_n12956), .B(new_n11354), .Y(new_n23612));
  A2O1A1Ixp33_ASAP7_75t_L   g23356(.A1(new_n12986), .A2(new_n11351), .B(new_n23612), .C(\a[59] ), .Y(new_n23613));
  A2O1A1Ixp33_ASAP7_75t_L   g23357(.A1(new_n12986), .A2(new_n11351), .B(new_n23612), .C(new_n11048), .Y(new_n23614));
  INVx1_ASAP7_75t_L         g23358(.A(new_n23614), .Y(new_n23615));
  NOR2xp33_ASAP7_75t_L      g23359(.A(new_n12258), .B(new_n12318), .Y(new_n23616));
  AOI221xp5_ASAP7_75t_L     g23360(.A1(new_n11995), .A2(\b[62] ), .B1(new_n13314), .B2(\b[60] ), .C(new_n23616), .Y(new_n23617));
  O2A1O1Ixp33_ASAP7_75t_L   g23361(.A1(new_n11998), .A2(new_n12610), .B(new_n23617), .C(new_n11987), .Y(new_n23618));
  O2A1O1Ixp33_ASAP7_75t_L   g23362(.A1(new_n11998), .A2(new_n12610), .B(new_n23617), .C(\a[62] ), .Y(new_n23619));
  INVx1_ASAP7_75t_L         g23363(.A(new_n23619), .Y(new_n23620));
  OAI21xp33_ASAP7_75t_L     g23364(.A1(new_n11987), .A2(new_n23618), .B(new_n23620), .Y(new_n23621));
  A2O1A1Ixp33_ASAP7_75t_L   g23365(.A1(\a[59] ), .A2(new_n23613), .B(new_n23615), .C(new_n23621), .Y(new_n23622));
  INVx1_ASAP7_75t_L         g23366(.A(new_n23622), .Y(new_n23623));
  O2A1O1Ixp33_ASAP7_75t_L   g23367(.A1(new_n11987), .A2(new_n23618), .B(new_n23620), .C(new_n23623), .Y(new_n23624));
  A2O1A1O1Ixp25_ASAP7_75t_L g23368(.A1(new_n23613), .A2(\a[59] ), .B(new_n23615), .C(new_n23622), .D(new_n23624), .Y(new_n23625));
  A2O1A1Ixp33_ASAP7_75t_L   g23369(.A1(new_n23611), .A2(new_n23605), .B(new_n23610), .C(new_n23625), .Y(new_n23626));
  O2A1O1Ixp33_ASAP7_75t_L   g23370(.A1(new_n23606), .A2(new_n23565), .B(new_n23611), .C(new_n23610), .Y(new_n23627));
  INVx1_ASAP7_75t_L         g23371(.A(new_n23613), .Y(new_n23628));
  O2A1O1Ixp33_ASAP7_75t_L   g23372(.A1(new_n23628), .A2(new_n11048), .B(new_n23614), .C(new_n23621), .Y(new_n23629));
  A2O1A1Ixp33_ASAP7_75t_L   g23373(.A1(new_n23621), .A2(new_n23622), .B(new_n23629), .C(new_n23627), .Y(new_n23630));
  AND2x2_ASAP7_75t_L        g23374(.A(new_n23626), .B(new_n23630), .Y(new_n23631));
  A2O1A1O1Ixp25_ASAP7_75t_L g23375(.A1(new_n23544), .A2(new_n23525), .B(new_n23577), .C(new_n23587), .D(new_n23631), .Y(new_n23632));
  A2O1A1Ixp33_ASAP7_75t_L   g23376(.A1(new_n13573), .A2(\b[63] ), .B(new_n23588), .C(new_n11351), .Y(new_n23633));
  A2O1A1Ixp33_ASAP7_75t_L   g23377(.A1(new_n23633), .A2(new_n23583), .B(new_n23584), .C(new_n23590), .Y(new_n23634));
  A2O1A1Ixp33_ASAP7_75t_L   g23378(.A1(new_n23581), .A2(new_n23634), .B(new_n23578), .C(new_n23631), .Y(new_n23635));
  A2O1A1Ixp33_ASAP7_75t_L   g23379(.A1(new_n23630), .A2(new_n23626), .B(new_n23632), .C(new_n23635), .Y(new_n23636));
  A2O1A1Ixp33_ASAP7_75t_L   g23380(.A1(new_n23554), .A2(new_n23558), .B(new_n23598), .C(new_n23596), .Y(new_n23637));
  INVx1_ASAP7_75t_L         g23381(.A(new_n23637), .Y(new_n23638));
  A2O1A1Ixp33_ASAP7_75t_L   g23382(.A1(new_n23626), .A2(new_n23630), .B(new_n23632), .C(new_n23638), .Y(new_n23639));
  A2O1A1O1Ixp25_ASAP7_75t_L g23383(.A1(new_n23581), .A2(new_n23634), .B(new_n23578), .C(new_n23631), .D(new_n23639), .Y(new_n23640));
  O2A1O1Ixp33_ASAP7_75t_L   g23384(.A1(new_n23595), .A2(new_n23599), .B(new_n23636), .C(new_n23640), .Y(\f[122] ));
  INVx1_ASAP7_75t_L         g23385(.A(new_n23627), .Y(new_n23642));
  A2O1A1Ixp33_ASAP7_75t_L   g23386(.A1(new_n23621), .A2(new_n23622), .B(new_n23629), .C(new_n23642), .Y(new_n23643));
  O2A1O1Ixp33_ASAP7_75t_L   g23387(.A1(new_n23629), .A2(new_n23621), .B(new_n23642), .C(new_n23623), .Y(new_n23644));
  INVx1_ASAP7_75t_L         g23388(.A(new_n23644), .Y(new_n23645));
  O2A1O1Ixp33_ASAP7_75t_L   g23389(.A1(new_n11591), .A2(new_n12672), .B(new_n23603), .C(new_n11048), .Y(new_n23646));
  AOI211xp5_ASAP7_75t_L     g23390(.A1(new_n13028), .A2(\b[59] ), .B(new_n23602), .C(\a[59] ), .Y(new_n23647));
  NOR2xp33_ASAP7_75t_L      g23391(.A(new_n23647), .B(new_n23646), .Y(new_n23648));
  NOR2xp33_ASAP7_75t_L      g23392(.A(new_n11591), .B(new_n13030), .Y(new_n23649));
  O2A1O1Ixp33_ASAP7_75t_L   g23393(.A1(new_n12669), .A2(new_n12671), .B(\b[60] ), .C(new_n23649), .Y(new_n23650));
  NAND2xp33_ASAP7_75t_L     g23394(.A(new_n23650), .B(new_n23648), .Y(new_n23651));
  INVx1_ASAP7_75t_L         g23395(.A(new_n23648), .Y(new_n23652));
  A2O1A1Ixp33_ASAP7_75t_L   g23396(.A1(\b[60] ), .A2(new_n13028), .B(new_n23649), .C(new_n23652), .Y(new_n23653));
  AND2x2_ASAP7_75t_L        g23397(.A(new_n23651), .B(new_n23653), .Y(new_n23654));
  INVx1_ASAP7_75t_L         g23398(.A(new_n23654), .Y(new_n23655));
  NOR2xp33_ASAP7_75t_L      g23399(.A(new_n12603), .B(new_n12318), .Y(new_n23656));
  AOI221xp5_ASAP7_75t_L     g23400(.A1(new_n11995), .A2(\b[63] ), .B1(new_n13314), .B2(\b[61] ), .C(new_n23656), .Y(new_n23657));
  O2A1O1Ixp33_ASAP7_75t_L   g23401(.A1(new_n11998), .A2(new_n17815), .B(new_n23657), .C(new_n11987), .Y(new_n23658));
  O2A1O1Ixp33_ASAP7_75t_L   g23402(.A1(new_n11998), .A2(new_n17815), .B(new_n23657), .C(\a[62] ), .Y(new_n23659));
  INVx1_ASAP7_75t_L         g23403(.A(new_n23659), .Y(new_n23660));
  O2A1O1Ixp33_ASAP7_75t_L   g23404(.A1(new_n11987), .A2(new_n23658), .B(new_n23660), .C(new_n23655), .Y(new_n23661));
  INVx1_ASAP7_75t_L         g23405(.A(new_n23658), .Y(new_n23662));
  A2O1A1Ixp33_ASAP7_75t_L   g23406(.A1(new_n23662), .A2(\a[62] ), .B(new_n23659), .C(new_n23655), .Y(new_n23663));
  O2A1O1Ixp33_ASAP7_75t_L   g23407(.A1(new_n23655), .A2(new_n23661), .B(new_n23663), .C(new_n23611), .Y(new_n23664));
  A2O1A1Ixp33_ASAP7_75t_L   g23408(.A1(new_n23662), .A2(\a[62] ), .B(new_n23659), .C(new_n23654), .Y(new_n23665));
  NOR2xp33_ASAP7_75t_L      g23409(.A(new_n23655), .B(new_n23661), .Y(new_n23666));
  A2O1A1O1Ixp25_ASAP7_75t_L g23410(.A1(new_n23662), .A2(\a[62] ), .B(new_n23659), .C(new_n23665), .D(new_n23666), .Y(new_n23667));
  AND2x2_ASAP7_75t_L        g23411(.A(new_n23611), .B(new_n23667), .Y(new_n23668));
  NOR2xp33_ASAP7_75t_L      g23412(.A(new_n23664), .B(new_n23668), .Y(new_n23669));
  NAND2xp33_ASAP7_75t_L     g23413(.A(new_n23669), .B(new_n23645), .Y(new_n23670));
  INVx1_ASAP7_75t_L         g23414(.A(new_n23670), .Y(new_n23671));
  NAND2xp33_ASAP7_75t_L     g23415(.A(new_n23644), .B(new_n23669), .Y(new_n23672));
  A2O1A1Ixp33_ASAP7_75t_L   g23416(.A1(new_n23643), .A2(new_n23622), .B(new_n23671), .C(new_n23672), .Y(new_n23673));
  O2A1O1Ixp33_ASAP7_75t_L   g23417(.A1(new_n23595), .A2(new_n23599), .B(new_n23636), .C(new_n23632), .Y(new_n23674));
  NAND2xp33_ASAP7_75t_L     g23418(.A(new_n23672), .B(new_n23674), .Y(new_n23675));
  O2A1O1Ixp33_ASAP7_75t_L   g23419(.A1(new_n23664), .A2(new_n23668), .B(new_n23645), .C(new_n23675), .Y(new_n23676));
  A2O1A1O1Ixp25_ASAP7_75t_L g23420(.A1(new_n23637), .A2(new_n23636), .B(new_n23632), .C(new_n23673), .D(new_n23676), .Y(\f[123] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g23421(.A1(new_n23662), .A2(\a[62] ), .B(new_n23659), .C(new_n23654), .D(new_n23664), .Y(new_n23678));
  NOR2xp33_ASAP7_75t_L      g23422(.A(new_n11626), .B(new_n13030), .Y(new_n23679));
  O2A1O1Ixp33_ASAP7_75t_L   g23423(.A1(new_n12669), .A2(new_n12671), .B(\b[61] ), .C(new_n23679), .Y(new_n23680));
  INVx1_ASAP7_75t_L         g23424(.A(new_n23680), .Y(new_n23681));
  O2A1O1Ixp33_ASAP7_75t_L   g23425(.A1(new_n11591), .A2(new_n12672), .B(new_n23603), .C(\a[59] ), .Y(new_n23682));
  INVx1_ASAP7_75t_L         g23426(.A(new_n23682), .Y(new_n23683));
  O2A1O1Ixp33_ASAP7_75t_L   g23427(.A1(new_n23650), .A2(new_n23648), .B(new_n23683), .C(new_n23681), .Y(new_n23684));
  INVx1_ASAP7_75t_L         g23428(.A(new_n23679), .Y(new_n23685));
  NAND2xp33_ASAP7_75t_L     g23429(.A(new_n23683), .B(new_n23653), .Y(new_n23686));
  O2A1O1Ixp33_ASAP7_75t_L   g23430(.A1(new_n12258), .A2(new_n12672), .B(new_n23685), .C(new_n23686), .Y(new_n23687));
  NOR2xp33_ASAP7_75t_L      g23431(.A(new_n23684), .B(new_n23687), .Y(new_n23688));
  NOR2xp33_ASAP7_75t_L      g23432(.A(new_n12956), .B(new_n12318), .Y(new_n23689));
  AOI21xp33_ASAP7_75t_L     g23433(.A1(new_n13314), .A2(\b[62] ), .B(new_n23689), .Y(new_n23690));
  INVx1_ASAP7_75t_L         g23434(.A(new_n23690), .Y(new_n23691));
  A2O1A1Ixp33_ASAP7_75t_L   g23435(.A1(new_n11992), .A2(new_n11993), .B(new_n11720), .C(new_n23690), .Y(new_n23692));
  O2A1O1Ixp33_ASAP7_75t_L   g23436(.A1(new_n23691), .A2(new_n17329), .B(new_n23692), .C(new_n11987), .Y(new_n23693));
  O2A1O1Ixp33_ASAP7_75t_L   g23437(.A1(new_n11998), .A2(new_n12993), .B(new_n23690), .C(\a[62] ), .Y(new_n23694));
  OAI21xp33_ASAP7_75t_L     g23438(.A1(new_n23694), .A2(new_n23693), .B(new_n23688), .Y(new_n23695));
  OR3x1_ASAP7_75t_L         g23439(.A(new_n23693), .B(new_n23688), .C(new_n23694), .Y(new_n23696));
  AND2x2_ASAP7_75t_L        g23440(.A(new_n23695), .B(new_n23696), .Y(new_n23697));
  OAI21xp33_ASAP7_75t_L     g23441(.A1(new_n23661), .A2(new_n23664), .B(new_n23697), .Y(new_n23698));
  A2O1A1O1Ixp25_ASAP7_75t_L g23442(.A1(new_n23663), .A2(new_n23655), .B(new_n23611), .C(new_n23665), .D(new_n23697), .Y(new_n23699));
  AOI21xp33_ASAP7_75t_L     g23443(.A1(new_n23698), .A2(new_n23697), .B(new_n23699), .Y(new_n23700));
  A2O1A1O1Ixp25_ASAP7_75t_L g23444(.A1(new_n23672), .A2(new_n23644), .B(new_n23674), .C(new_n23670), .D(new_n23700), .Y(new_n23701));
  A2O1A1Ixp33_ASAP7_75t_L   g23445(.A1(new_n23672), .A2(new_n23644), .B(new_n23674), .C(new_n23670), .Y(new_n23702));
  AOI21xp33_ASAP7_75t_L     g23446(.A1(new_n23697), .A2(new_n23678), .B(new_n23702), .Y(new_n23703));
  O2A1O1Ixp33_ASAP7_75t_L   g23447(.A1(new_n23697), .A2(new_n23678), .B(new_n23703), .C(new_n23701), .Y(\f[124] ));
  O2A1O1Ixp33_ASAP7_75t_L   g23448(.A1(new_n23694), .A2(new_n23693), .B(new_n23688), .C(new_n23684), .Y(new_n23705));
  A2O1A1O1Ixp25_ASAP7_75t_L g23449(.A1(new_n13028), .A2(\b[60] ), .B(new_n23649), .C(new_n23652), .D(new_n23682), .Y(new_n23706));
  NAND2xp33_ASAP7_75t_L     g23450(.A(\b[61] ), .B(new_n13029), .Y(new_n23707));
  O2A1O1Ixp33_ASAP7_75t_L   g23451(.A1(new_n12672), .A2(new_n12603), .B(new_n23707), .C(new_n23681), .Y(new_n23708));
  A2O1A1Ixp33_ASAP7_75t_L   g23452(.A1(new_n12685), .A2(new_n12686), .B(new_n12603), .C(new_n23707), .Y(new_n23709));
  O2A1O1Ixp33_ASAP7_75t_L   g23453(.A1(new_n12258), .A2(new_n12672), .B(new_n23685), .C(new_n23709), .Y(new_n23710));
  NOR2xp33_ASAP7_75t_L      g23454(.A(new_n23710), .B(new_n23708), .Y(new_n23711));
  NOR2xp33_ASAP7_75t_L      g23455(.A(new_n12956), .B(new_n12320), .Y(new_n23712));
  INVx1_ASAP7_75t_L         g23456(.A(new_n23712), .Y(new_n23713));
  A2O1A1Ixp33_ASAP7_75t_L   g23457(.A1(new_n14444), .A2(new_n12603), .B(new_n12956), .C(new_n23713), .Y(new_n23714));
  O2A1O1Ixp33_ASAP7_75t_L   g23458(.A1(new_n11997), .A2(new_n23712), .B(new_n23714), .C(new_n11987), .Y(new_n23715));
  INVx1_ASAP7_75t_L         g23459(.A(new_n23715), .Y(new_n23716));
  O2A1O1Ixp33_ASAP7_75t_L   g23460(.A1(new_n11998), .A2(new_n13573), .B(new_n23713), .C(\a[62] ), .Y(new_n23717));
  INVx1_ASAP7_75t_L         g23461(.A(new_n23717), .Y(new_n23718));
  NAND2xp33_ASAP7_75t_L     g23462(.A(new_n23718), .B(new_n23716), .Y(new_n23719));
  NAND2xp33_ASAP7_75t_L     g23463(.A(new_n23711), .B(new_n23719), .Y(new_n23720));
  OR3x1_ASAP7_75t_L         g23464(.A(new_n23715), .B(new_n23711), .C(new_n23717), .Y(new_n23721));
  AND2x2_ASAP7_75t_L        g23465(.A(new_n23721), .B(new_n23720), .Y(new_n23722));
  INVx1_ASAP7_75t_L         g23466(.A(new_n23722), .Y(new_n23723));
  O2A1O1Ixp33_ASAP7_75t_L   g23467(.A1(new_n23681), .A2(new_n23706), .B(new_n23695), .C(new_n23723), .Y(new_n23724));
  A2O1A1Ixp33_ASAP7_75t_L   g23468(.A1(new_n23637), .A2(new_n23636), .B(new_n23632), .C(new_n23673), .Y(new_n23725));
  O2A1O1Ixp33_ASAP7_75t_L   g23469(.A1(new_n23681), .A2(new_n23706), .B(new_n23695), .C(new_n23722), .Y(new_n23726));
  NOR2xp33_ASAP7_75t_L      g23470(.A(new_n23723), .B(new_n23724), .Y(new_n23727));
  NOR2xp33_ASAP7_75t_L      g23471(.A(new_n23726), .B(new_n23727), .Y(new_n23728));
  A2O1A1O1Ixp25_ASAP7_75t_L g23472(.A1(new_n23670), .A2(new_n23725), .B(new_n23700), .C(new_n23698), .D(new_n23728), .Y(new_n23729));
  A2O1A1Ixp33_ASAP7_75t_L   g23473(.A1(new_n23725), .A2(new_n23670), .B(new_n23700), .C(new_n23698), .Y(new_n23730));
  NOR2xp33_ASAP7_75t_L      g23474(.A(new_n23727), .B(new_n23730), .Y(new_n23731));
  O2A1O1Ixp33_ASAP7_75t_L   g23475(.A1(new_n23724), .A2(new_n23705), .B(new_n23731), .C(new_n23729), .Y(\f[125] ));
  O2A1O1Ixp33_ASAP7_75t_L   g23476(.A1(new_n23726), .A2(new_n23722), .B(new_n23730), .C(new_n23724), .Y(new_n23733));
  O2A1O1Ixp33_ASAP7_75t_L   g23477(.A1(new_n23717), .A2(new_n23715), .B(new_n23711), .C(new_n23708), .Y(new_n23734));
  NOR2xp33_ASAP7_75t_L      g23478(.A(new_n12603), .B(new_n13030), .Y(new_n23735));
  A2O1A1Ixp33_ASAP7_75t_L   g23479(.A1(\a[63] ), .A2(\b[63] ), .B(new_n23735), .C(new_n11987), .Y(new_n23736));
  O2A1O1Ixp33_ASAP7_75t_L   g23480(.A1(new_n12669), .A2(new_n12671), .B(\b[63] ), .C(new_n23735), .Y(new_n23737));
  NAND2xp33_ASAP7_75t_L     g23481(.A(\a[62] ), .B(new_n23737), .Y(new_n23738));
  NAND2xp33_ASAP7_75t_L     g23482(.A(new_n23736), .B(new_n23738), .Y(new_n23739));
  INVx1_ASAP7_75t_L         g23483(.A(new_n23739), .Y(new_n23740));
  A2O1A1Ixp33_ASAP7_75t_L   g23484(.A1(new_n13028), .A2(\b[61] ), .B(new_n23679), .C(new_n23740), .Y(new_n23741));
  NAND2xp33_ASAP7_75t_L     g23485(.A(new_n23680), .B(new_n23739), .Y(new_n23742));
  AND2x2_ASAP7_75t_L        g23486(.A(new_n23742), .B(new_n23741), .Y(new_n23743));
  XNOR2x2_ASAP7_75t_L       g23487(.A(new_n23743), .B(new_n23734), .Y(new_n23744));
  XNOR2x2_ASAP7_75t_L       g23488(.A(new_n23744), .B(new_n23733), .Y(\f[126] ));
  NAND2xp33_ASAP7_75t_L     g23489(.A(\b[63] ), .B(new_n13029), .Y(new_n23746));
  O2A1O1Ixp33_ASAP7_75t_L   g23490(.A1(new_n23680), .A2(new_n23739), .B(new_n23736), .C(new_n23746), .Y(new_n23747));
  AND3x1_ASAP7_75t_L        g23491(.A(new_n23741), .B(new_n23746), .C(new_n23736), .Y(new_n23748));
  NOR2xp33_ASAP7_75t_L      g23492(.A(new_n23747), .B(new_n23748), .Y(new_n23749));
  INVx1_ASAP7_75t_L         g23493(.A(new_n23728), .Y(new_n23750));
  A2O1A1Ixp33_ASAP7_75t_L   g23494(.A1(new_n23719), .A2(new_n23711), .B(new_n23708), .C(new_n23743), .Y(new_n23751));
  INVx1_ASAP7_75t_L         g23495(.A(new_n23751), .Y(new_n23752));
  A2O1A1O1Ixp25_ASAP7_75t_L g23496(.A1(new_n23750), .A2(new_n23730), .B(new_n23724), .C(new_n23744), .D(new_n23752), .Y(new_n23753));
  XOR2x2_ASAP7_75t_L        g23497(.A(new_n23749), .B(new_n23753), .Y(\f[127] ));
endmodule


