// Benchmark "top" written by ABC on Mon Dec 25 16:29:22 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n423, new_n424, new_n425,
    new_n426, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n451, new_n452, new_n453, new_n454, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1235, new_n1236, new_n1237, new_n1238, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1357, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1403, new_n1404, new_n1405, new_n1406, new_n1408,
    new_n1409, new_n1410, new_n1411, new_n1412, new_n1413, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1418, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1464, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1469, new_n1470, new_n1471, new_n1472, new_n1473, new_n1474,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1524, new_n1525, new_n1526, new_n1527, new_n1528,
    new_n1529, new_n1530, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1558;
  XOR2x2_ASAP7_75t_L        g0000(.A(\b[0] ), .B(\a[0] ), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g0001(.A(\b[0] ), .B(\a[0] ), .Y(new_n387));
  INVx1_ASAP7_75t_L         g0002(.A(\a[1] ), .Y(new_n388));
  INVx1_ASAP7_75t_L         g0003(.A(\b[1] ), .Y(new_n389));
  NAND2xp33_ASAP7_75t_L     g0004(.A(new_n389), .B(new_n388), .Y(new_n390));
  NAND2xp33_ASAP7_75t_L     g0005(.A(\b[1] ), .B(\a[1] ), .Y(new_n391));
  NAND2xp33_ASAP7_75t_L     g0006(.A(new_n391), .B(new_n390), .Y(new_n392));
  XOR2x2_ASAP7_75t_L        g0007(.A(new_n387), .B(new_n392), .Y(\f[1] ));
  NAND3xp33_ASAP7_75t_L     g0008(.A(new_n390), .B(\b[0] ), .C(\a[0] ), .Y(new_n394));
  NOR2xp33_ASAP7_75t_L      g0009(.A(\a[2] ), .B(\b[2] ), .Y(new_n395));
  INVx1_ASAP7_75t_L         g0010(.A(new_n395), .Y(new_n396));
  NAND2xp33_ASAP7_75t_L     g0011(.A(\b[2] ), .B(\a[2] ), .Y(new_n397));
  NAND2xp33_ASAP7_75t_L     g0012(.A(new_n397), .B(new_n396), .Y(new_n398));
  AND3x1_ASAP7_75t_L        g0013(.A(new_n394), .B(new_n398), .C(new_n391), .Y(new_n399));
  O2A1O1Ixp33_ASAP7_75t_L   g0014(.A1(new_n388), .A2(new_n389), .B(new_n394), .C(new_n398), .Y(new_n400));
  NOR2xp33_ASAP7_75t_L      g0015(.A(new_n400), .B(new_n399), .Y(\f[2] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0016(.A1(new_n394), .A2(new_n391), .B(new_n395), .C(new_n397), .Y(new_n402));
  INVx1_ASAP7_75t_L         g0017(.A(\a[3] ), .Y(new_n403));
  INVx1_ASAP7_75t_L         g0018(.A(\b[3] ), .Y(new_n404));
  NAND2xp33_ASAP7_75t_L     g0019(.A(new_n404), .B(new_n403), .Y(new_n405));
  NOR2xp33_ASAP7_75t_L      g0020(.A(new_n403), .B(new_n404), .Y(new_n406));
  INVx1_ASAP7_75t_L         g0021(.A(new_n406), .Y(new_n407));
  AOI21xp33_ASAP7_75t_L     g0022(.A1(new_n407), .A2(new_n405), .B(new_n402), .Y(new_n408));
  NAND2xp33_ASAP7_75t_L     g0023(.A(new_n405), .B(new_n407), .Y(new_n409));
  A2O1A1O1Ixp25_ASAP7_75t_L g0024(.A1(new_n394), .A2(new_n391), .B(new_n395), .C(new_n397), .D(new_n409), .Y(new_n410));
  NOR2xp33_ASAP7_75t_L      g0025(.A(new_n410), .B(new_n408), .Y(\f[3] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0026(.A1(new_n388), .A2(new_n389), .B(new_n394), .C(new_n395), .Y(new_n412));
  A2O1A1Ixp33_ASAP7_75t_L   g0027(.A1(\b[2] ), .A2(\a[2] ), .B(new_n412), .C(new_n405), .Y(new_n413));
  INVx1_ASAP7_75t_L         g0028(.A(\a[4] ), .Y(new_n414));
  INVx1_ASAP7_75t_L         g0029(.A(\b[4] ), .Y(new_n415));
  NAND2xp33_ASAP7_75t_L     g0030(.A(new_n415), .B(new_n414), .Y(new_n416));
  NOR2xp33_ASAP7_75t_L      g0031(.A(new_n414), .B(new_n415), .Y(new_n417));
  INVx1_ASAP7_75t_L         g0032(.A(new_n417), .Y(new_n418));
  NAND2xp33_ASAP7_75t_L     g0033(.A(new_n416), .B(new_n418), .Y(new_n419));
  AND3x1_ASAP7_75t_L        g0034(.A(new_n413), .B(new_n419), .C(new_n407), .Y(new_n420));
  O2A1O1Ixp33_ASAP7_75t_L   g0035(.A1(new_n403), .A2(new_n404), .B(new_n413), .C(new_n419), .Y(new_n421));
  NOR2xp33_ASAP7_75t_L      g0036(.A(new_n421), .B(new_n420), .Y(\f[4] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0037(.A1(new_n405), .A2(new_n402), .B(new_n406), .C(new_n416), .D(new_n417), .Y(new_n423));
  NOR2xp33_ASAP7_75t_L      g0038(.A(\a[5] ), .B(\b[5] ), .Y(new_n424));
  AND2x2_ASAP7_75t_L        g0039(.A(\a[5] ), .B(\b[5] ), .Y(new_n425));
  NOR2xp33_ASAP7_75t_L      g0040(.A(new_n424), .B(new_n425), .Y(new_n426));
  XNOR2x2_ASAP7_75t_L       g0041(.A(new_n426), .B(new_n423), .Y(\f[5] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0042(.A1(new_n402), .A2(new_n405), .B(new_n406), .C(new_n416), .Y(new_n428));
  NAND2xp33_ASAP7_75t_L     g0043(.A(\b[5] ), .B(\a[5] ), .Y(new_n429));
  A2O1A1Ixp33_ASAP7_75t_L   g0044(.A1(new_n428), .A2(new_n418), .B(new_n424), .C(new_n429), .Y(new_n430));
  INVx1_ASAP7_75t_L         g0045(.A(\a[6] ), .Y(new_n431));
  INVx1_ASAP7_75t_L         g0046(.A(\b[6] ), .Y(new_n432));
  NAND2xp33_ASAP7_75t_L     g0047(.A(new_n432), .B(new_n431), .Y(new_n433));
  NOR2xp33_ASAP7_75t_L      g0048(.A(new_n431), .B(new_n432), .Y(new_n434));
  INVx1_ASAP7_75t_L         g0049(.A(new_n434), .Y(new_n435));
  AOI21xp33_ASAP7_75t_L     g0050(.A1(new_n435), .A2(new_n433), .B(new_n430), .Y(new_n436));
  NAND2xp33_ASAP7_75t_L     g0051(.A(new_n433), .B(new_n435), .Y(new_n437));
  A2O1A1O1Ixp25_ASAP7_75t_L g0052(.A1(new_n418), .A2(new_n428), .B(new_n424), .C(new_n429), .D(new_n437), .Y(new_n438));
  NOR2xp33_ASAP7_75t_L      g0053(.A(new_n438), .B(new_n436), .Y(\f[6] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0054(.A1(new_n414), .A2(new_n415), .B(new_n428), .C(new_n424), .Y(new_n440));
  A2O1A1Ixp33_ASAP7_75t_L   g0055(.A1(\b[5] ), .A2(\a[5] ), .B(new_n440), .C(new_n433), .Y(new_n441));
  INVx1_ASAP7_75t_L         g0056(.A(\a[7] ), .Y(new_n442));
  INVx1_ASAP7_75t_L         g0057(.A(\b[7] ), .Y(new_n443));
  NAND2xp33_ASAP7_75t_L     g0058(.A(new_n443), .B(new_n442), .Y(new_n444));
  NOR2xp33_ASAP7_75t_L      g0059(.A(new_n442), .B(new_n443), .Y(new_n445));
  INVx1_ASAP7_75t_L         g0060(.A(new_n445), .Y(new_n446));
  NAND2xp33_ASAP7_75t_L     g0061(.A(new_n444), .B(new_n446), .Y(new_n447));
  AND3x1_ASAP7_75t_L        g0062(.A(new_n441), .B(new_n447), .C(new_n435), .Y(new_n448));
  O2A1O1Ixp33_ASAP7_75t_L   g0063(.A1(new_n431), .A2(new_n432), .B(new_n441), .C(new_n447), .Y(new_n449));
  NOR2xp33_ASAP7_75t_L      g0064(.A(new_n449), .B(new_n448), .Y(\f[7] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0065(.A1(new_n433), .A2(new_n430), .B(new_n434), .C(new_n444), .D(new_n445), .Y(new_n451));
  NOR2xp33_ASAP7_75t_L      g0066(.A(\a[8] ), .B(\b[8] ), .Y(new_n452));
  AND2x2_ASAP7_75t_L        g0067(.A(\a[8] ), .B(\b[8] ), .Y(new_n453));
  NOR2xp33_ASAP7_75t_L      g0068(.A(new_n452), .B(new_n453), .Y(new_n454));
  XNOR2x2_ASAP7_75t_L       g0069(.A(new_n454), .B(new_n451), .Y(\f[8] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0070(.A1(new_n430), .A2(new_n433), .B(new_n434), .C(new_n444), .Y(new_n456));
  NAND2xp33_ASAP7_75t_L     g0071(.A(\b[8] ), .B(\a[8] ), .Y(new_n457));
  A2O1A1Ixp33_ASAP7_75t_L   g0072(.A1(new_n456), .A2(new_n446), .B(new_n452), .C(new_n457), .Y(new_n458));
  INVx1_ASAP7_75t_L         g0073(.A(\a[9] ), .Y(new_n459));
  INVx1_ASAP7_75t_L         g0074(.A(\b[9] ), .Y(new_n460));
  NAND2xp33_ASAP7_75t_L     g0075(.A(new_n460), .B(new_n459), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g0076(.A(new_n459), .B(new_n460), .Y(new_n462));
  INVx1_ASAP7_75t_L         g0077(.A(new_n462), .Y(new_n463));
  AOI21xp33_ASAP7_75t_L     g0078(.A1(new_n463), .A2(new_n461), .B(new_n458), .Y(new_n464));
  NAND2xp33_ASAP7_75t_L     g0079(.A(new_n461), .B(new_n463), .Y(new_n465));
  A2O1A1O1Ixp25_ASAP7_75t_L g0080(.A1(new_n446), .A2(new_n456), .B(new_n452), .C(new_n457), .D(new_n465), .Y(new_n466));
  NOR2xp33_ASAP7_75t_L      g0081(.A(new_n466), .B(new_n464), .Y(\f[9] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0082(.A1(new_n442), .A2(new_n443), .B(new_n456), .C(new_n452), .Y(new_n468));
  A2O1A1Ixp33_ASAP7_75t_L   g0083(.A1(\b[8] ), .A2(\a[8] ), .B(new_n468), .C(new_n461), .Y(new_n469));
  INVx1_ASAP7_75t_L         g0084(.A(\a[10] ), .Y(new_n470));
  INVx1_ASAP7_75t_L         g0085(.A(\b[10] ), .Y(new_n471));
  NAND2xp33_ASAP7_75t_L     g0086(.A(new_n471), .B(new_n470), .Y(new_n472));
  NOR2xp33_ASAP7_75t_L      g0087(.A(new_n470), .B(new_n471), .Y(new_n473));
  INVx1_ASAP7_75t_L         g0088(.A(new_n473), .Y(new_n474));
  NAND2xp33_ASAP7_75t_L     g0089(.A(new_n472), .B(new_n474), .Y(new_n475));
  AND3x1_ASAP7_75t_L        g0090(.A(new_n469), .B(new_n475), .C(new_n463), .Y(new_n476));
  O2A1O1Ixp33_ASAP7_75t_L   g0091(.A1(new_n459), .A2(new_n460), .B(new_n469), .C(new_n475), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g0092(.A(new_n477), .B(new_n476), .Y(\f[10] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0093(.A1(new_n461), .A2(new_n458), .B(new_n462), .C(new_n472), .D(new_n473), .Y(new_n479));
  NOR2xp33_ASAP7_75t_L      g0094(.A(\a[11] ), .B(\b[11] ), .Y(new_n480));
  NAND2xp33_ASAP7_75t_L     g0095(.A(\b[11] ), .B(\a[11] ), .Y(new_n481));
  INVx1_ASAP7_75t_L         g0096(.A(new_n481), .Y(new_n482));
  NOR2xp33_ASAP7_75t_L      g0097(.A(new_n480), .B(new_n482), .Y(new_n483));
  XNOR2x2_ASAP7_75t_L       g0098(.A(new_n483), .B(new_n479), .Y(\f[11] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0099(.A1(new_n458), .A2(new_n461), .B(new_n462), .C(new_n472), .Y(new_n485));
  A2O1A1Ixp33_ASAP7_75t_L   g0100(.A1(new_n485), .A2(new_n474), .B(new_n480), .C(new_n481), .Y(new_n486));
  INVx1_ASAP7_75t_L         g0101(.A(\a[12] ), .Y(new_n487));
  INVx1_ASAP7_75t_L         g0102(.A(\b[12] ), .Y(new_n488));
  NAND2xp33_ASAP7_75t_L     g0103(.A(new_n488), .B(new_n487), .Y(new_n489));
  NOR2xp33_ASAP7_75t_L      g0104(.A(new_n487), .B(new_n488), .Y(new_n490));
  INVx1_ASAP7_75t_L         g0105(.A(new_n490), .Y(new_n491));
  AOI21xp33_ASAP7_75t_L     g0106(.A1(new_n491), .A2(new_n489), .B(new_n486), .Y(new_n492));
  NAND2xp33_ASAP7_75t_L     g0107(.A(new_n489), .B(new_n491), .Y(new_n493));
  A2O1A1O1Ixp25_ASAP7_75t_L g0108(.A1(new_n474), .A2(new_n485), .B(new_n480), .C(new_n481), .D(new_n493), .Y(new_n494));
  NOR2xp33_ASAP7_75t_L      g0109(.A(new_n494), .B(new_n492), .Y(\f[12] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0110(.A1(new_n470), .A2(new_n471), .B(new_n485), .C(new_n480), .Y(new_n496));
  A2O1A1Ixp33_ASAP7_75t_L   g0111(.A1(\b[11] ), .A2(\a[11] ), .B(new_n496), .C(new_n489), .Y(new_n497));
  INVx1_ASAP7_75t_L         g0112(.A(\a[13] ), .Y(new_n498));
  INVx1_ASAP7_75t_L         g0113(.A(\b[13] ), .Y(new_n499));
  NAND2xp33_ASAP7_75t_L     g0114(.A(new_n499), .B(new_n498), .Y(new_n500));
  NOR2xp33_ASAP7_75t_L      g0115(.A(new_n498), .B(new_n499), .Y(new_n501));
  INVx1_ASAP7_75t_L         g0116(.A(new_n501), .Y(new_n502));
  NAND2xp33_ASAP7_75t_L     g0117(.A(new_n500), .B(new_n502), .Y(new_n503));
  AND3x1_ASAP7_75t_L        g0118(.A(new_n497), .B(new_n503), .C(new_n491), .Y(new_n504));
  O2A1O1Ixp33_ASAP7_75t_L   g0119(.A1(new_n487), .A2(new_n488), .B(new_n497), .C(new_n503), .Y(new_n505));
  NOR2xp33_ASAP7_75t_L      g0120(.A(new_n505), .B(new_n504), .Y(\f[13] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0121(.A1(new_n489), .A2(new_n486), .B(new_n490), .C(new_n500), .D(new_n501), .Y(new_n507));
  NOR2xp33_ASAP7_75t_L      g0122(.A(\a[14] ), .B(\b[14] ), .Y(new_n508));
  AND2x2_ASAP7_75t_L        g0123(.A(\a[14] ), .B(\b[14] ), .Y(new_n509));
  NOR2xp33_ASAP7_75t_L      g0124(.A(new_n508), .B(new_n509), .Y(new_n510));
  XNOR2x2_ASAP7_75t_L       g0125(.A(new_n510), .B(new_n507), .Y(\f[14] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0126(.A1(new_n486), .A2(new_n489), .B(new_n490), .C(new_n500), .Y(new_n512));
  NAND2xp33_ASAP7_75t_L     g0127(.A(\b[14] ), .B(\a[14] ), .Y(new_n513));
  A2O1A1Ixp33_ASAP7_75t_L   g0128(.A1(new_n512), .A2(new_n502), .B(new_n508), .C(new_n513), .Y(new_n514));
  INVx1_ASAP7_75t_L         g0129(.A(\a[15] ), .Y(new_n515));
  INVx1_ASAP7_75t_L         g0130(.A(\b[15] ), .Y(new_n516));
  NAND2xp33_ASAP7_75t_L     g0131(.A(new_n516), .B(new_n515), .Y(new_n517));
  NOR2xp33_ASAP7_75t_L      g0132(.A(new_n515), .B(new_n516), .Y(new_n518));
  INVx1_ASAP7_75t_L         g0133(.A(new_n518), .Y(new_n519));
  AOI21xp33_ASAP7_75t_L     g0134(.A1(new_n519), .A2(new_n517), .B(new_n514), .Y(new_n520));
  NAND2xp33_ASAP7_75t_L     g0135(.A(new_n517), .B(new_n519), .Y(new_n521));
  A2O1A1O1Ixp25_ASAP7_75t_L g0136(.A1(new_n502), .A2(new_n512), .B(new_n508), .C(new_n513), .D(new_n521), .Y(new_n522));
  NOR2xp33_ASAP7_75t_L      g0137(.A(new_n522), .B(new_n520), .Y(\f[15] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0138(.A1(new_n498), .A2(new_n499), .B(new_n512), .C(new_n508), .Y(new_n524));
  A2O1A1Ixp33_ASAP7_75t_L   g0139(.A1(\b[14] ), .A2(\a[14] ), .B(new_n524), .C(new_n517), .Y(new_n525));
  INVx1_ASAP7_75t_L         g0140(.A(\a[16] ), .Y(new_n526));
  INVx1_ASAP7_75t_L         g0141(.A(\b[16] ), .Y(new_n527));
  NAND2xp33_ASAP7_75t_L     g0142(.A(new_n527), .B(new_n526), .Y(new_n528));
  NOR2xp33_ASAP7_75t_L      g0143(.A(new_n526), .B(new_n527), .Y(new_n529));
  INVx1_ASAP7_75t_L         g0144(.A(new_n529), .Y(new_n530));
  NAND2xp33_ASAP7_75t_L     g0145(.A(new_n528), .B(new_n530), .Y(new_n531));
  AND3x1_ASAP7_75t_L        g0146(.A(new_n525), .B(new_n531), .C(new_n519), .Y(new_n532));
  O2A1O1Ixp33_ASAP7_75t_L   g0147(.A1(new_n515), .A2(new_n516), .B(new_n525), .C(new_n531), .Y(new_n533));
  NOR2xp33_ASAP7_75t_L      g0148(.A(new_n533), .B(new_n532), .Y(\f[16] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0149(.A1(new_n517), .A2(new_n514), .B(new_n518), .C(new_n528), .D(new_n529), .Y(new_n535));
  NOR2xp33_ASAP7_75t_L      g0150(.A(\a[17] ), .B(\b[17] ), .Y(new_n536));
  AND2x2_ASAP7_75t_L        g0151(.A(\a[17] ), .B(\b[17] ), .Y(new_n537));
  NOR2xp33_ASAP7_75t_L      g0152(.A(new_n536), .B(new_n537), .Y(new_n538));
  XNOR2x2_ASAP7_75t_L       g0153(.A(new_n538), .B(new_n535), .Y(\f[17] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0154(.A1(new_n514), .A2(new_n517), .B(new_n518), .C(new_n528), .Y(new_n540));
  NAND2xp33_ASAP7_75t_L     g0155(.A(\b[17] ), .B(\a[17] ), .Y(new_n541));
  A2O1A1Ixp33_ASAP7_75t_L   g0156(.A1(new_n540), .A2(new_n530), .B(new_n536), .C(new_n541), .Y(new_n542));
  INVx1_ASAP7_75t_L         g0157(.A(\a[18] ), .Y(new_n543));
  INVx1_ASAP7_75t_L         g0158(.A(\b[18] ), .Y(new_n544));
  NAND2xp33_ASAP7_75t_L     g0159(.A(new_n544), .B(new_n543), .Y(new_n545));
  NOR2xp33_ASAP7_75t_L      g0160(.A(new_n543), .B(new_n544), .Y(new_n546));
  INVx1_ASAP7_75t_L         g0161(.A(new_n546), .Y(new_n547));
  AOI21xp33_ASAP7_75t_L     g0162(.A1(new_n547), .A2(new_n545), .B(new_n542), .Y(new_n548));
  NAND2xp33_ASAP7_75t_L     g0163(.A(new_n545), .B(new_n547), .Y(new_n549));
  A2O1A1O1Ixp25_ASAP7_75t_L g0164(.A1(new_n530), .A2(new_n540), .B(new_n536), .C(new_n541), .D(new_n549), .Y(new_n550));
  NOR2xp33_ASAP7_75t_L      g0165(.A(new_n550), .B(new_n548), .Y(\f[18] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0166(.A1(new_n526), .A2(new_n527), .B(new_n540), .C(new_n536), .Y(new_n552));
  A2O1A1Ixp33_ASAP7_75t_L   g0167(.A1(\b[17] ), .A2(\a[17] ), .B(new_n552), .C(new_n545), .Y(new_n553));
  INVx1_ASAP7_75t_L         g0168(.A(\a[19] ), .Y(new_n554));
  INVx1_ASAP7_75t_L         g0169(.A(\b[19] ), .Y(new_n555));
  NAND2xp33_ASAP7_75t_L     g0170(.A(new_n555), .B(new_n554), .Y(new_n556));
  NOR2xp33_ASAP7_75t_L      g0171(.A(new_n554), .B(new_n555), .Y(new_n557));
  INVx1_ASAP7_75t_L         g0172(.A(new_n557), .Y(new_n558));
  NAND2xp33_ASAP7_75t_L     g0173(.A(new_n556), .B(new_n558), .Y(new_n559));
  AND3x1_ASAP7_75t_L        g0174(.A(new_n553), .B(new_n559), .C(new_n547), .Y(new_n560));
  O2A1O1Ixp33_ASAP7_75t_L   g0175(.A1(new_n543), .A2(new_n544), .B(new_n553), .C(new_n559), .Y(new_n561));
  NOR2xp33_ASAP7_75t_L      g0176(.A(new_n561), .B(new_n560), .Y(\f[19] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0177(.A1(new_n545), .A2(new_n542), .B(new_n546), .C(new_n556), .D(new_n557), .Y(new_n563));
  NOR2xp33_ASAP7_75t_L      g0178(.A(\a[20] ), .B(\b[20] ), .Y(new_n564));
  AND2x2_ASAP7_75t_L        g0179(.A(\a[20] ), .B(\b[20] ), .Y(new_n565));
  NOR2xp33_ASAP7_75t_L      g0180(.A(new_n564), .B(new_n565), .Y(new_n566));
  XNOR2x2_ASAP7_75t_L       g0181(.A(new_n566), .B(new_n563), .Y(\f[20] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0182(.A1(new_n542), .A2(new_n545), .B(new_n546), .C(new_n556), .Y(new_n568));
  NAND2xp33_ASAP7_75t_L     g0183(.A(\b[20] ), .B(\a[20] ), .Y(new_n569));
  A2O1A1Ixp33_ASAP7_75t_L   g0184(.A1(new_n568), .A2(new_n558), .B(new_n564), .C(new_n569), .Y(new_n570));
  INVx1_ASAP7_75t_L         g0185(.A(\a[21] ), .Y(new_n571));
  INVx1_ASAP7_75t_L         g0186(.A(\b[21] ), .Y(new_n572));
  NAND2xp33_ASAP7_75t_L     g0187(.A(new_n572), .B(new_n571), .Y(new_n573));
  NOR2xp33_ASAP7_75t_L      g0188(.A(new_n571), .B(new_n572), .Y(new_n574));
  INVx1_ASAP7_75t_L         g0189(.A(new_n574), .Y(new_n575));
  AOI21xp33_ASAP7_75t_L     g0190(.A1(new_n575), .A2(new_n573), .B(new_n570), .Y(new_n576));
  NAND2xp33_ASAP7_75t_L     g0191(.A(new_n573), .B(new_n575), .Y(new_n577));
  A2O1A1O1Ixp25_ASAP7_75t_L g0192(.A1(new_n558), .A2(new_n568), .B(new_n564), .C(new_n569), .D(new_n577), .Y(new_n578));
  NOR2xp33_ASAP7_75t_L      g0193(.A(new_n578), .B(new_n576), .Y(\f[21] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0194(.A1(new_n554), .A2(new_n555), .B(new_n568), .C(new_n564), .Y(new_n580));
  A2O1A1Ixp33_ASAP7_75t_L   g0195(.A1(\b[20] ), .A2(\a[20] ), .B(new_n580), .C(new_n573), .Y(new_n581));
  INVx1_ASAP7_75t_L         g0196(.A(\a[22] ), .Y(new_n582));
  INVx1_ASAP7_75t_L         g0197(.A(\b[22] ), .Y(new_n583));
  NAND2xp33_ASAP7_75t_L     g0198(.A(new_n583), .B(new_n582), .Y(new_n584));
  NOR2xp33_ASAP7_75t_L      g0199(.A(new_n582), .B(new_n583), .Y(new_n585));
  INVx1_ASAP7_75t_L         g0200(.A(new_n585), .Y(new_n586));
  NAND2xp33_ASAP7_75t_L     g0201(.A(new_n584), .B(new_n586), .Y(new_n587));
  AND3x1_ASAP7_75t_L        g0202(.A(new_n581), .B(new_n587), .C(new_n575), .Y(new_n588));
  O2A1O1Ixp33_ASAP7_75t_L   g0203(.A1(new_n571), .A2(new_n572), .B(new_n581), .C(new_n587), .Y(new_n589));
  NOR2xp33_ASAP7_75t_L      g0204(.A(new_n589), .B(new_n588), .Y(\f[22] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0205(.A1(new_n573), .A2(new_n570), .B(new_n574), .C(new_n584), .D(new_n585), .Y(new_n591));
  NOR2xp33_ASAP7_75t_L      g0206(.A(\a[23] ), .B(\b[23] ), .Y(new_n592));
  AND2x2_ASAP7_75t_L        g0207(.A(\a[23] ), .B(\b[23] ), .Y(new_n593));
  NOR2xp33_ASAP7_75t_L      g0208(.A(new_n592), .B(new_n593), .Y(new_n594));
  XNOR2x2_ASAP7_75t_L       g0209(.A(new_n594), .B(new_n591), .Y(\f[23] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0210(.A1(new_n570), .A2(new_n573), .B(new_n574), .C(new_n584), .Y(new_n596));
  NAND2xp33_ASAP7_75t_L     g0211(.A(\b[23] ), .B(\a[23] ), .Y(new_n597));
  A2O1A1Ixp33_ASAP7_75t_L   g0212(.A1(new_n596), .A2(new_n586), .B(new_n592), .C(new_n597), .Y(new_n598));
  INVx1_ASAP7_75t_L         g0213(.A(\a[24] ), .Y(new_n599));
  INVx1_ASAP7_75t_L         g0214(.A(\b[24] ), .Y(new_n600));
  NAND2xp33_ASAP7_75t_L     g0215(.A(new_n600), .B(new_n599), .Y(new_n601));
  NOR2xp33_ASAP7_75t_L      g0216(.A(new_n599), .B(new_n600), .Y(new_n602));
  INVx1_ASAP7_75t_L         g0217(.A(new_n602), .Y(new_n603));
  AOI21xp33_ASAP7_75t_L     g0218(.A1(new_n603), .A2(new_n601), .B(new_n598), .Y(new_n604));
  NAND2xp33_ASAP7_75t_L     g0219(.A(new_n601), .B(new_n603), .Y(new_n605));
  A2O1A1O1Ixp25_ASAP7_75t_L g0220(.A1(new_n586), .A2(new_n596), .B(new_n592), .C(new_n597), .D(new_n605), .Y(new_n606));
  NOR2xp33_ASAP7_75t_L      g0221(.A(new_n606), .B(new_n604), .Y(\f[24] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0222(.A1(new_n582), .A2(new_n583), .B(new_n596), .C(new_n592), .Y(new_n608));
  A2O1A1Ixp33_ASAP7_75t_L   g0223(.A1(\b[23] ), .A2(\a[23] ), .B(new_n608), .C(new_n601), .Y(new_n609));
  INVx1_ASAP7_75t_L         g0224(.A(\a[25] ), .Y(new_n610));
  INVx1_ASAP7_75t_L         g0225(.A(\b[25] ), .Y(new_n611));
  NAND2xp33_ASAP7_75t_L     g0226(.A(new_n611), .B(new_n610), .Y(new_n612));
  NOR2xp33_ASAP7_75t_L      g0227(.A(new_n610), .B(new_n611), .Y(new_n613));
  INVx1_ASAP7_75t_L         g0228(.A(new_n613), .Y(new_n614));
  NAND2xp33_ASAP7_75t_L     g0229(.A(new_n612), .B(new_n614), .Y(new_n615));
  AND3x1_ASAP7_75t_L        g0230(.A(new_n609), .B(new_n615), .C(new_n603), .Y(new_n616));
  O2A1O1Ixp33_ASAP7_75t_L   g0231(.A1(new_n599), .A2(new_n600), .B(new_n609), .C(new_n615), .Y(new_n617));
  NOR2xp33_ASAP7_75t_L      g0232(.A(new_n617), .B(new_n616), .Y(\f[25] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0233(.A1(new_n601), .A2(new_n598), .B(new_n602), .C(new_n612), .D(new_n613), .Y(new_n619));
  NOR2xp33_ASAP7_75t_L      g0234(.A(\a[26] ), .B(\b[26] ), .Y(new_n620));
  AND2x2_ASAP7_75t_L        g0235(.A(\a[26] ), .B(\b[26] ), .Y(new_n621));
  NOR2xp33_ASAP7_75t_L      g0236(.A(new_n620), .B(new_n621), .Y(new_n622));
  XNOR2x2_ASAP7_75t_L       g0237(.A(new_n622), .B(new_n619), .Y(\f[26] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0238(.A1(new_n598), .A2(new_n601), .B(new_n602), .C(new_n612), .Y(new_n624));
  NAND2xp33_ASAP7_75t_L     g0239(.A(\b[26] ), .B(\a[26] ), .Y(new_n625));
  A2O1A1Ixp33_ASAP7_75t_L   g0240(.A1(new_n624), .A2(new_n614), .B(new_n620), .C(new_n625), .Y(new_n626));
  INVx1_ASAP7_75t_L         g0241(.A(\a[27] ), .Y(new_n627));
  INVx1_ASAP7_75t_L         g0242(.A(\b[27] ), .Y(new_n628));
  NAND2xp33_ASAP7_75t_L     g0243(.A(new_n628), .B(new_n627), .Y(new_n629));
  NOR2xp33_ASAP7_75t_L      g0244(.A(new_n627), .B(new_n628), .Y(new_n630));
  INVx1_ASAP7_75t_L         g0245(.A(new_n630), .Y(new_n631));
  AOI21xp33_ASAP7_75t_L     g0246(.A1(new_n631), .A2(new_n629), .B(new_n626), .Y(new_n632));
  NAND2xp33_ASAP7_75t_L     g0247(.A(new_n629), .B(new_n631), .Y(new_n633));
  A2O1A1O1Ixp25_ASAP7_75t_L g0248(.A1(new_n614), .A2(new_n624), .B(new_n620), .C(new_n625), .D(new_n633), .Y(new_n634));
  NOR2xp33_ASAP7_75t_L      g0249(.A(new_n634), .B(new_n632), .Y(\f[27] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0250(.A1(new_n610), .A2(new_n611), .B(new_n624), .C(new_n620), .Y(new_n636));
  A2O1A1Ixp33_ASAP7_75t_L   g0251(.A1(\b[26] ), .A2(\a[26] ), .B(new_n636), .C(new_n629), .Y(new_n637));
  INVx1_ASAP7_75t_L         g0252(.A(\a[28] ), .Y(new_n638));
  INVx1_ASAP7_75t_L         g0253(.A(\b[28] ), .Y(new_n639));
  NAND2xp33_ASAP7_75t_L     g0254(.A(new_n639), .B(new_n638), .Y(new_n640));
  NOR2xp33_ASAP7_75t_L      g0255(.A(new_n638), .B(new_n639), .Y(new_n641));
  INVx1_ASAP7_75t_L         g0256(.A(new_n641), .Y(new_n642));
  NAND2xp33_ASAP7_75t_L     g0257(.A(new_n640), .B(new_n642), .Y(new_n643));
  AND3x1_ASAP7_75t_L        g0258(.A(new_n637), .B(new_n643), .C(new_n631), .Y(new_n644));
  O2A1O1Ixp33_ASAP7_75t_L   g0259(.A1(new_n627), .A2(new_n628), .B(new_n637), .C(new_n643), .Y(new_n645));
  NOR2xp33_ASAP7_75t_L      g0260(.A(new_n645), .B(new_n644), .Y(\f[28] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0261(.A1(new_n629), .A2(new_n626), .B(new_n630), .C(new_n640), .D(new_n641), .Y(new_n647));
  NOR2xp33_ASAP7_75t_L      g0262(.A(\a[29] ), .B(\b[29] ), .Y(new_n648));
  AND2x2_ASAP7_75t_L        g0263(.A(\a[29] ), .B(\b[29] ), .Y(new_n649));
  NOR2xp33_ASAP7_75t_L      g0264(.A(new_n648), .B(new_n649), .Y(new_n650));
  XNOR2x2_ASAP7_75t_L       g0265(.A(new_n650), .B(new_n647), .Y(\f[29] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0266(.A1(new_n626), .A2(new_n629), .B(new_n630), .C(new_n640), .Y(new_n652));
  NAND2xp33_ASAP7_75t_L     g0267(.A(\b[29] ), .B(\a[29] ), .Y(new_n653));
  A2O1A1Ixp33_ASAP7_75t_L   g0268(.A1(new_n652), .A2(new_n642), .B(new_n648), .C(new_n653), .Y(new_n654));
  INVx1_ASAP7_75t_L         g0269(.A(\a[30] ), .Y(new_n655));
  INVx1_ASAP7_75t_L         g0270(.A(\b[30] ), .Y(new_n656));
  NAND2xp33_ASAP7_75t_L     g0271(.A(new_n656), .B(new_n655), .Y(new_n657));
  NOR2xp33_ASAP7_75t_L      g0272(.A(new_n655), .B(new_n656), .Y(new_n658));
  INVx1_ASAP7_75t_L         g0273(.A(new_n658), .Y(new_n659));
  AOI21xp33_ASAP7_75t_L     g0274(.A1(new_n659), .A2(new_n657), .B(new_n654), .Y(new_n660));
  NAND2xp33_ASAP7_75t_L     g0275(.A(new_n657), .B(new_n659), .Y(new_n661));
  A2O1A1O1Ixp25_ASAP7_75t_L g0276(.A1(new_n642), .A2(new_n652), .B(new_n648), .C(new_n653), .D(new_n661), .Y(new_n662));
  NOR2xp33_ASAP7_75t_L      g0277(.A(new_n662), .B(new_n660), .Y(\f[30] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0278(.A1(new_n638), .A2(new_n639), .B(new_n652), .C(new_n648), .Y(new_n664));
  A2O1A1Ixp33_ASAP7_75t_L   g0279(.A1(\b[29] ), .A2(\a[29] ), .B(new_n664), .C(new_n657), .Y(new_n665));
  INVx1_ASAP7_75t_L         g0280(.A(\a[31] ), .Y(new_n666));
  INVx1_ASAP7_75t_L         g0281(.A(\b[31] ), .Y(new_n667));
  NAND2xp33_ASAP7_75t_L     g0282(.A(new_n667), .B(new_n666), .Y(new_n668));
  NOR2xp33_ASAP7_75t_L      g0283(.A(new_n666), .B(new_n667), .Y(new_n669));
  INVx1_ASAP7_75t_L         g0284(.A(new_n669), .Y(new_n670));
  NAND2xp33_ASAP7_75t_L     g0285(.A(new_n668), .B(new_n670), .Y(new_n671));
  AND3x1_ASAP7_75t_L        g0286(.A(new_n665), .B(new_n671), .C(new_n659), .Y(new_n672));
  O2A1O1Ixp33_ASAP7_75t_L   g0287(.A1(new_n655), .A2(new_n656), .B(new_n665), .C(new_n671), .Y(new_n673));
  NOR2xp33_ASAP7_75t_L      g0288(.A(new_n673), .B(new_n672), .Y(\f[31] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0289(.A1(new_n657), .A2(new_n654), .B(new_n658), .C(new_n668), .D(new_n669), .Y(new_n675));
  NOR2xp33_ASAP7_75t_L      g0290(.A(\a[32] ), .B(\b[32] ), .Y(new_n676));
  AND2x2_ASAP7_75t_L        g0291(.A(\a[32] ), .B(\b[32] ), .Y(new_n677));
  NOR2xp33_ASAP7_75t_L      g0292(.A(new_n676), .B(new_n677), .Y(new_n678));
  XNOR2x2_ASAP7_75t_L       g0293(.A(new_n678), .B(new_n675), .Y(\f[32] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0294(.A1(new_n654), .A2(new_n657), .B(new_n658), .C(new_n668), .Y(new_n680));
  NAND2xp33_ASAP7_75t_L     g0295(.A(\b[32] ), .B(\a[32] ), .Y(new_n681));
  A2O1A1Ixp33_ASAP7_75t_L   g0296(.A1(new_n680), .A2(new_n670), .B(new_n676), .C(new_n681), .Y(new_n682));
  INVx1_ASAP7_75t_L         g0297(.A(\a[33] ), .Y(new_n683));
  INVx1_ASAP7_75t_L         g0298(.A(\b[33] ), .Y(new_n684));
  NAND2xp33_ASAP7_75t_L     g0299(.A(new_n684), .B(new_n683), .Y(new_n685));
  NOR2xp33_ASAP7_75t_L      g0300(.A(new_n683), .B(new_n684), .Y(new_n686));
  INVx1_ASAP7_75t_L         g0301(.A(new_n686), .Y(new_n687));
  AOI21xp33_ASAP7_75t_L     g0302(.A1(new_n687), .A2(new_n685), .B(new_n682), .Y(new_n688));
  NAND2xp33_ASAP7_75t_L     g0303(.A(new_n685), .B(new_n687), .Y(new_n689));
  A2O1A1O1Ixp25_ASAP7_75t_L g0304(.A1(new_n670), .A2(new_n680), .B(new_n676), .C(new_n681), .D(new_n689), .Y(new_n690));
  NOR2xp33_ASAP7_75t_L      g0305(.A(new_n690), .B(new_n688), .Y(\f[33] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0306(.A1(new_n666), .A2(new_n667), .B(new_n680), .C(new_n676), .Y(new_n692));
  A2O1A1Ixp33_ASAP7_75t_L   g0307(.A1(\b[32] ), .A2(\a[32] ), .B(new_n692), .C(new_n685), .Y(new_n693));
  INVx1_ASAP7_75t_L         g0308(.A(\a[34] ), .Y(new_n694));
  INVx1_ASAP7_75t_L         g0309(.A(\b[34] ), .Y(new_n695));
  NAND2xp33_ASAP7_75t_L     g0310(.A(new_n695), .B(new_n694), .Y(new_n696));
  NOR2xp33_ASAP7_75t_L      g0311(.A(new_n694), .B(new_n695), .Y(new_n697));
  INVx1_ASAP7_75t_L         g0312(.A(new_n697), .Y(new_n698));
  NAND2xp33_ASAP7_75t_L     g0313(.A(new_n696), .B(new_n698), .Y(new_n699));
  AND3x1_ASAP7_75t_L        g0314(.A(new_n693), .B(new_n699), .C(new_n687), .Y(new_n700));
  O2A1O1Ixp33_ASAP7_75t_L   g0315(.A1(new_n683), .A2(new_n684), .B(new_n693), .C(new_n699), .Y(new_n701));
  NOR2xp33_ASAP7_75t_L      g0316(.A(new_n701), .B(new_n700), .Y(\f[34] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0317(.A1(new_n685), .A2(new_n682), .B(new_n686), .C(new_n696), .D(new_n697), .Y(new_n703));
  NOR2xp33_ASAP7_75t_L      g0318(.A(\a[35] ), .B(\b[35] ), .Y(new_n704));
  AND2x2_ASAP7_75t_L        g0319(.A(\a[35] ), .B(\b[35] ), .Y(new_n705));
  NOR2xp33_ASAP7_75t_L      g0320(.A(new_n704), .B(new_n705), .Y(new_n706));
  XNOR2x2_ASAP7_75t_L       g0321(.A(new_n706), .B(new_n703), .Y(\f[35] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0322(.A1(new_n682), .A2(new_n685), .B(new_n686), .C(new_n696), .Y(new_n708));
  NAND2xp33_ASAP7_75t_L     g0323(.A(\b[35] ), .B(\a[35] ), .Y(new_n709));
  A2O1A1Ixp33_ASAP7_75t_L   g0324(.A1(new_n708), .A2(new_n698), .B(new_n704), .C(new_n709), .Y(new_n710));
  INVx1_ASAP7_75t_L         g0325(.A(\a[36] ), .Y(new_n711));
  INVx1_ASAP7_75t_L         g0326(.A(\b[36] ), .Y(new_n712));
  NAND2xp33_ASAP7_75t_L     g0327(.A(new_n712), .B(new_n711), .Y(new_n713));
  NOR2xp33_ASAP7_75t_L      g0328(.A(new_n711), .B(new_n712), .Y(new_n714));
  INVx1_ASAP7_75t_L         g0329(.A(new_n714), .Y(new_n715));
  AOI21xp33_ASAP7_75t_L     g0330(.A1(new_n715), .A2(new_n713), .B(new_n710), .Y(new_n716));
  NAND2xp33_ASAP7_75t_L     g0331(.A(new_n713), .B(new_n715), .Y(new_n717));
  A2O1A1O1Ixp25_ASAP7_75t_L g0332(.A1(new_n698), .A2(new_n708), .B(new_n704), .C(new_n709), .D(new_n717), .Y(new_n718));
  NOR2xp33_ASAP7_75t_L      g0333(.A(new_n718), .B(new_n716), .Y(\f[36] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0334(.A1(new_n694), .A2(new_n695), .B(new_n708), .C(new_n704), .Y(new_n720));
  A2O1A1Ixp33_ASAP7_75t_L   g0335(.A1(\b[35] ), .A2(\a[35] ), .B(new_n720), .C(new_n713), .Y(new_n721));
  INVx1_ASAP7_75t_L         g0336(.A(\a[37] ), .Y(new_n722));
  INVx1_ASAP7_75t_L         g0337(.A(\b[37] ), .Y(new_n723));
  NAND2xp33_ASAP7_75t_L     g0338(.A(new_n723), .B(new_n722), .Y(new_n724));
  NOR2xp33_ASAP7_75t_L      g0339(.A(new_n722), .B(new_n723), .Y(new_n725));
  INVx1_ASAP7_75t_L         g0340(.A(new_n725), .Y(new_n726));
  NAND2xp33_ASAP7_75t_L     g0341(.A(new_n724), .B(new_n726), .Y(new_n727));
  AND3x1_ASAP7_75t_L        g0342(.A(new_n721), .B(new_n727), .C(new_n715), .Y(new_n728));
  O2A1O1Ixp33_ASAP7_75t_L   g0343(.A1(new_n711), .A2(new_n712), .B(new_n721), .C(new_n727), .Y(new_n729));
  NOR2xp33_ASAP7_75t_L      g0344(.A(new_n729), .B(new_n728), .Y(\f[37] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0345(.A1(new_n713), .A2(new_n710), .B(new_n714), .C(new_n724), .D(new_n725), .Y(new_n731));
  NOR2xp33_ASAP7_75t_L      g0346(.A(\a[38] ), .B(\b[38] ), .Y(new_n732));
  AND2x2_ASAP7_75t_L        g0347(.A(\a[38] ), .B(\b[38] ), .Y(new_n733));
  NOR2xp33_ASAP7_75t_L      g0348(.A(new_n732), .B(new_n733), .Y(new_n734));
  XNOR2x2_ASAP7_75t_L       g0349(.A(new_n734), .B(new_n731), .Y(\f[38] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0350(.A1(new_n710), .A2(new_n713), .B(new_n714), .C(new_n724), .Y(new_n736));
  NAND2xp33_ASAP7_75t_L     g0351(.A(\b[38] ), .B(\a[38] ), .Y(new_n737));
  A2O1A1Ixp33_ASAP7_75t_L   g0352(.A1(new_n736), .A2(new_n726), .B(new_n732), .C(new_n737), .Y(new_n738));
  INVx1_ASAP7_75t_L         g0353(.A(\a[39] ), .Y(new_n739));
  INVx1_ASAP7_75t_L         g0354(.A(\b[39] ), .Y(new_n740));
  NAND2xp33_ASAP7_75t_L     g0355(.A(new_n740), .B(new_n739), .Y(new_n741));
  NOR2xp33_ASAP7_75t_L      g0356(.A(new_n739), .B(new_n740), .Y(new_n742));
  INVx1_ASAP7_75t_L         g0357(.A(new_n742), .Y(new_n743));
  AOI21xp33_ASAP7_75t_L     g0358(.A1(new_n743), .A2(new_n741), .B(new_n738), .Y(new_n744));
  NAND2xp33_ASAP7_75t_L     g0359(.A(new_n741), .B(new_n743), .Y(new_n745));
  A2O1A1O1Ixp25_ASAP7_75t_L g0360(.A1(new_n726), .A2(new_n736), .B(new_n732), .C(new_n737), .D(new_n745), .Y(new_n746));
  NOR2xp33_ASAP7_75t_L      g0361(.A(new_n746), .B(new_n744), .Y(\f[39] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0362(.A1(new_n722), .A2(new_n723), .B(new_n736), .C(new_n732), .Y(new_n748));
  A2O1A1Ixp33_ASAP7_75t_L   g0363(.A1(\b[38] ), .A2(\a[38] ), .B(new_n748), .C(new_n741), .Y(new_n749));
  INVx1_ASAP7_75t_L         g0364(.A(\a[40] ), .Y(new_n750));
  INVx1_ASAP7_75t_L         g0365(.A(\b[40] ), .Y(new_n751));
  NAND2xp33_ASAP7_75t_L     g0366(.A(new_n751), .B(new_n750), .Y(new_n752));
  NOR2xp33_ASAP7_75t_L      g0367(.A(new_n750), .B(new_n751), .Y(new_n753));
  INVx1_ASAP7_75t_L         g0368(.A(new_n753), .Y(new_n754));
  NAND2xp33_ASAP7_75t_L     g0369(.A(new_n752), .B(new_n754), .Y(new_n755));
  AND3x1_ASAP7_75t_L        g0370(.A(new_n749), .B(new_n755), .C(new_n743), .Y(new_n756));
  O2A1O1Ixp33_ASAP7_75t_L   g0371(.A1(new_n739), .A2(new_n740), .B(new_n749), .C(new_n755), .Y(new_n757));
  NOR2xp33_ASAP7_75t_L      g0372(.A(new_n757), .B(new_n756), .Y(\f[40] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0373(.A1(new_n741), .A2(new_n738), .B(new_n742), .C(new_n752), .D(new_n753), .Y(new_n759));
  NOR2xp33_ASAP7_75t_L      g0374(.A(\a[41] ), .B(\b[41] ), .Y(new_n760));
  AND2x2_ASAP7_75t_L        g0375(.A(\a[41] ), .B(\b[41] ), .Y(new_n761));
  NOR2xp33_ASAP7_75t_L      g0376(.A(new_n760), .B(new_n761), .Y(new_n762));
  XNOR2x2_ASAP7_75t_L       g0377(.A(new_n762), .B(new_n759), .Y(\f[41] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0378(.A1(new_n738), .A2(new_n741), .B(new_n742), .C(new_n752), .Y(new_n764));
  NAND2xp33_ASAP7_75t_L     g0379(.A(\b[41] ), .B(\a[41] ), .Y(new_n765));
  A2O1A1Ixp33_ASAP7_75t_L   g0380(.A1(new_n764), .A2(new_n754), .B(new_n760), .C(new_n765), .Y(new_n766));
  INVx1_ASAP7_75t_L         g0381(.A(\a[42] ), .Y(new_n767));
  INVx1_ASAP7_75t_L         g0382(.A(\b[42] ), .Y(new_n768));
  NAND2xp33_ASAP7_75t_L     g0383(.A(new_n768), .B(new_n767), .Y(new_n769));
  NOR2xp33_ASAP7_75t_L      g0384(.A(new_n767), .B(new_n768), .Y(new_n770));
  INVx1_ASAP7_75t_L         g0385(.A(new_n770), .Y(new_n771));
  AOI21xp33_ASAP7_75t_L     g0386(.A1(new_n771), .A2(new_n769), .B(new_n766), .Y(new_n772));
  NAND2xp33_ASAP7_75t_L     g0387(.A(new_n769), .B(new_n771), .Y(new_n773));
  A2O1A1O1Ixp25_ASAP7_75t_L g0388(.A1(new_n754), .A2(new_n764), .B(new_n760), .C(new_n765), .D(new_n773), .Y(new_n774));
  NOR2xp33_ASAP7_75t_L      g0389(.A(new_n774), .B(new_n772), .Y(\f[42] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0390(.A1(new_n750), .A2(new_n751), .B(new_n764), .C(new_n760), .Y(new_n776));
  A2O1A1Ixp33_ASAP7_75t_L   g0391(.A1(\b[41] ), .A2(\a[41] ), .B(new_n776), .C(new_n769), .Y(new_n777));
  INVx1_ASAP7_75t_L         g0392(.A(\a[43] ), .Y(new_n778));
  INVx1_ASAP7_75t_L         g0393(.A(\b[43] ), .Y(new_n779));
  NAND2xp33_ASAP7_75t_L     g0394(.A(new_n779), .B(new_n778), .Y(new_n780));
  NOR2xp33_ASAP7_75t_L      g0395(.A(new_n778), .B(new_n779), .Y(new_n781));
  INVx1_ASAP7_75t_L         g0396(.A(new_n781), .Y(new_n782));
  NAND2xp33_ASAP7_75t_L     g0397(.A(new_n780), .B(new_n782), .Y(new_n783));
  AND3x1_ASAP7_75t_L        g0398(.A(new_n777), .B(new_n783), .C(new_n771), .Y(new_n784));
  O2A1O1Ixp33_ASAP7_75t_L   g0399(.A1(new_n767), .A2(new_n768), .B(new_n777), .C(new_n783), .Y(new_n785));
  NOR2xp33_ASAP7_75t_L      g0400(.A(new_n785), .B(new_n784), .Y(\f[43] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0401(.A1(new_n769), .A2(new_n766), .B(new_n770), .C(new_n780), .D(new_n781), .Y(new_n787));
  NOR2xp33_ASAP7_75t_L      g0402(.A(\a[44] ), .B(\b[44] ), .Y(new_n788));
  AND2x2_ASAP7_75t_L        g0403(.A(\a[44] ), .B(\b[44] ), .Y(new_n789));
  NOR2xp33_ASAP7_75t_L      g0404(.A(new_n788), .B(new_n789), .Y(new_n790));
  XNOR2x2_ASAP7_75t_L       g0405(.A(new_n790), .B(new_n787), .Y(\f[44] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0406(.A1(new_n766), .A2(new_n769), .B(new_n770), .C(new_n780), .Y(new_n792));
  NAND2xp33_ASAP7_75t_L     g0407(.A(\b[44] ), .B(\a[44] ), .Y(new_n793));
  A2O1A1Ixp33_ASAP7_75t_L   g0408(.A1(new_n792), .A2(new_n782), .B(new_n788), .C(new_n793), .Y(new_n794));
  INVx1_ASAP7_75t_L         g0409(.A(\a[45] ), .Y(new_n795));
  INVx1_ASAP7_75t_L         g0410(.A(\b[45] ), .Y(new_n796));
  NAND2xp33_ASAP7_75t_L     g0411(.A(new_n796), .B(new_n795), .Y(new_n797));
  NOR2xp33_ASAP7_75t_L      g0412(.A(new_n795), .B(new_n796), .Y(new_n798));
  INVx1_ASAP7_75t_L         g0413(.A(new_n798), .Y(new_n799));
  AOI21xp33_ASAP7_75t_L     g0414(.A1(new_n799), .A2(new_n797), .B(new_n794), .Y(new_n800));
  NAND2xp33_ASAP7_75t_L     g0415(.A(new_n797), .B(new_n799), .Y(new_n801));
  A2O1A1O1Ixp25_ASAP7_75t_L g0416(.A1(new_n782), .A2(new_n792), .B(new_n788), .C(new_n793), .D(new_n801), .Y(new_n802));
  NOR2xp33_ASAP7_75t_L      g0417(.A(new_n802), .B(new_n800), .Y(\f[45] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0418(.A1(new_n778), .A2(new_n779), .B(new_n792), .C(new_n788), .Y(new_n804));
  A2O1A1Ixp33_ASAP7_75t_L   g0419(.A1(\b[44] ), .A2(\a[44] ), .B(new_n804), .C(new_n797), .Y(new_n805));
  INVx1_ASAP7_75t_L         g0420(.A(\a[46] ), .Y(new_n806));
  INVx1_ASAP7_75t_L         g0421(.A(\b[46] ), .Y(new_n807));
  NAND2xp33_ASAP7_75t_L     g0422(.A(new_n807), .B(new_n806), .Y(new_n808));
  NOR2xp33_ASAP7_75t_L      g0423(.A(new_n806), .B(new_n807), .Y(new_n809));
  INVx1_ASAP7_75t_L         g0424(.A(new_n809), .Y(new_n810));
  NAND2xp33_ASAP7_75t_L     g0425(.A(new_n808), .B(new_n810), .Y(new_n811));
  AND3x1_ASAP7_75t_L        g0426(.A(new_n805), .B(new_n811), .C(new_n799), .Y(new_n812));
  O2A1O1Ixp33_ASAP7_75t_L   g0427(.A1(new_n795), .A2(new_n796), .B(new_n805), .C(new_n811), .Y(new_n813));
  NOR2xp33_ASAP7_75t_L      g0428(.A(new_n813), .B(new_n812), .Y(\f[46] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0429(.A1(new_n797), .A2(new_n794), .B(new_n798), .C(new_n808), .D(new_n809), .Y(new_n815));
  NOR2xp33_ASAP7_75t_L      g0430(.A(\a[47] ), .B(\b[47] ), .Y(new_n816));
  AND2x2_ASAP7_75t_L        g0431(.A(\a[47] ), .B(\b[47] ), .Y(new_n817));
  NOR2xp33_ASAP7_75t_L      g0432(.A(new_n816), .B(new_n817), .Y(new_n818));
  XNOR2x2_ASAP7_75t_L       g0433(.A(new_n818), .B(new_n815), .Y(\f[47] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0434(.A1(new_n794), .A2(new_n797), .B(new_n798), .C(new_n808), .Y(new_n820));
  NAND2xp33_ASAP7_75t_L     g0435(.A(\b[47] ), .B(\a[47] ), .Y(new_n821));
  A2O1A1Ixp33_ASAP7_75t_L   g0436(.A1(new_n820), .A2(new_n810), .B(new_n816), .C(new_n821), .Y(new_n822));
  INVx1_ASAP7_75t_L         g0437(.A(\a[48] ), .Y(new_n823));
  INVx1_ASAP7_75t_L         g0438(.A(\b[48] ), .Y(new_n824));
  NAND2xp33_ASAP7_75t_L     g0439(.A(new_n824), .B(new_n823), .Y(new_n825));
  NOR2xp33_ASAP7_75t_L      g0440(.A(new_n823), .B(new_n824), .Y(new_n826));
  INVx1_ASAP7_75t_L         g0441(.A(new_n826), .Y(new_n827));
  AOI21xp33_ASAP7_75t_L     g0442(.A1(new_n827), .A2(new_n825), .B(new_n822), .Y(new_n828));
  NAND2xp33_ASAP7_75t_L     g0443(.A(new_n825), .B(new_n827), .Y(new_n829));
  A2O1A1O1Ixp25_ASAP7_75t_L g0444(.A1(new_n810), .A2(new_n820), .B(new_n816), .C(new_n821), .D(new_n829), .Y(new_n830));
  NOR2xp33_ASAP7_75t_L      g0445(.A(new_n830), .B(new_n828), .Y(\f[48] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0446(.A1(new_n806), .A2(new_n807), .B(new_n820), .C(new_n816), .Y(new_n832));
  A2O1A1Ixp33_ASAP7_75t_L   g0447(.A1(\b[47] ), .A2(\a[47] ), .B(new_n832), .C(new_n825), .Y(new_n833));
  INVx1_ASAP7_75t_L         g0448(.A(\a[49] ), .Y(new_n834));
  INVx1_ASAP7_75t_L         g0449(.A(\b[49] ), .Y(new_n835));
  NAND2xp33_ASAP7_75t_L     g0450(.A(new_n835), .B(new_n834), .Y(new_n836));
  NOR2xp33_ASAP7_75t_L      g0451(.A(new_n834), .B(new_n835), .Y(new_n837));
  INVx1_ASAP7_75t_L         g0452(.A(new_n837), .Y(new_n838));
  NAND2xp33_ASAP7_75t_L     g0453(.A(new_n836), .B(new_n838), .Y(new_n839));
  AND3x1_ASAP7_75t_L        g0454(.A(new_n833), .B(new_n839), .C(new_n827), .Y(new_n840));
  O2A1O1Ixp33_ASAP7_75t_L   g0455(.A1(new_n823), .A2(new_n824), .B(new_n833), .C(new_n839), .Y(new_n841));
  NOR2xp33_ASAP7_75t_L      g0456(.A(new_n841), .B(new_n840), .Y(\f[49] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0457(.A1(new_n825), .A2(new_n822), .B(new_n826), .C(new_n836), .D(new_n837), .Y(new_n843));
  NOR2xp33_ASAP7_75t_L      g0458(.A(\a[50] ), .B(\b[50] ), .Y(new_n844));
  AND2x2_ASAP7_75t_L        g0459(.A(\a[50] ), .B(\b[50] ), .Y(new_n845));
  NOR2xp33_ASAP7_75t_L      g0460(.A(new_n844), .B(new_n845), .Y(new_n846));
  XNOR2x2_ASAP7_75t_L       g0461(.A(new_n846), .B(new_n843), .Y(\f[50] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0462(.A1(new_n822), .A2(new_n825), .B(new_n826), .C(new_n836), .Y(new_n848));
  NAND2xp33_ASAP7_75t_L     g0463(.A(\b[50] ), .B(\a[50] ), .Y(new_n849));
  A2O1A1Ixp33_ASAP7_75t_L   g0464(.A1(new_n848), .A2(new_n838), .B(new_n844), .C(new_n849), .Y(new_n850));
  INVx1_ASAP7_75t_L         g0465(.A(\a[51] ), .Y(new_n851));
  INVx1_ASAP7_75t_L         g0466(.A(\b[51] ), .Y(new_n852));
  NAND2xp33_ASAP7_75t_L     g0467(.A(new_n852), .B(new_n851), .Y(new_n853));
  NOR2xp33_ASAP7_75t_L      g0468(.A(new_n851), .B(new_n852), .Y(new_n854));
  INVx1_ASAP7_75t_L         g0469(.A(new_n854), .Y(new_n855));
  AOI21xp33_ASAP7_75t_L     g0470(.A1(new_n855), .A2(new_n853), .B(new_n850), .Y(new_n856));
  NAND2xp33_ASAP7_75t_L     g0471(.A(new_n853), .B(new_n855), .Y(new_n857));
  A2O1A1O1Ixp25_ASAP7_75t_L g0472(.A1(new_n838), .A2(new_n848), .B(new_n844), .C(new_n849), .D(new_n857), .Y(new_n858));
  NOR2xp33_ASAP7_75t_L      g0473(.A(new_n858), .B(new_n856), .Y(\f[51] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0474(.A1(new_n834), .A2(new_n835), .B(new_n848), .C(new_n844), .Y(new_n860));
  A2O1A1Ixp33_ASAP7_75t_L   g0475(.A1(\b[50] ), .A2(\a[50] ), .B(new_n860), .C(new_n853), .Y(new_n861));
  INVx1_ASAP7_75t_L         g0476(.A(\a[52] ), .Y(new_n862));
  INVx1_ASAP7_75t_L         g0477(.A(\b[52] ), .Y(new_n863));
  NAND2xp33_ASAP7_75t_L     g0478(.A(new_n863), .B(new_n862), .Y(new_n864));
  NOR2xp33_ASAP7_75t_L      g0479(.A(new_n862), .B(new_n863), .Y(new_n865));
  INVx1_ASAP7_75t_L         g0480(.A(new_n865), .Y(new_n866));
  NAND2xp33_ASAP7_75t_L     g0481(.A(new_n864), .B(new_n866), .Y(new_n867));
  AND3x1_ASAP7_75t_L        g0482(.A(new_n861), .B(new_n867), .C(new_n855), .Y(new_n868));
  O2A1O1Ixp33_ASAP7_75t_L   g0483(.A1(new_n851), .A2(new_n852), .B(new_n861), .C(new_n867), .Y(new_n869));
  NOR2xp33_ASAP7_75t_L      g0484(.A(new_n869), .B(new_n868), .Y(\f[52] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0485(.A1(new_n853), .A2(new_n850), .B(new_n854), .C(new_n864), .D(new_n865), .Y(new_n871));
  NOR2xp33_ASAP7_75t_L      g0486(.A(\a[53] ), .B(\b[53] ), .Y(new_n872));
  AND2x2_ASAP7_75t_L        g0487(.A(\a[53] ), .B(\b[53] ), .Y(new_n873));
  NOR2xp33_ASAP7_75t_L      g0488(.A(new_n872), .B(new_n873), .Y(new_n874));
  XNOR2x2_ASAP7_75t_L       g0489(.A(new_n874), .B(new_n871), .Y(\f[53] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0490(.A1(new_n850), .A2(new_n853), .B(new_n854), .C(new_n864), .Y(new_n876));
  NAND2xp33_ASAP7_75t_L     g0491(.A(\b[53] ), .B(\a[53] ), .Y(new_n877));
  A2O1A1Ixp33_ASAP7_75t_L   g0492(.A1(new_n876), .A2(new_n866), .B(new_n872), .C(new_n877), .Y(new_n878));
  INVx1_ASAP7_75t_L         g0493(.A(\a[54] ), .Y(new_n879));
  INVx1_ASAP7_75t_L         g0494(.A(\b[54] ), .Y(new_n880));
  NAND2xp33_ASAP7_75t_L     g0495(.A(new_n880), .B(new_n879), .Y(new_n881));
  NOR2xp33_ASAP7_75t_L      g0496(.A(new_n879), .B(new_n880), .Y(new_n882));
  INVx1_ASAP7_75t_L         g0497(.A(new_n882), .Y(new_n883));
  AOI21xp33_ASAP7_75t_L     g0498(.A1(new_n883), .A2(new_n881), .B(new_n878), .Y(new_n884));
  NAND2xp33_ASAP7_75t_L     g0499(.A(new_n881), .B(new_n883), .Y(new_n885));
  A2O1A1O1Ixp25_ASAP7_75t_L g0500(.A1(new_n866), .A2(new_n876), .B(new_n872), .C(new_n877), .D(new_n885), .Y(new_n886));
  NOR2xp33_ASAP7_75t_L      g0501(.A(new_n886), .B(new_n884), .Y(\f[54] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0502(.A1(new_n862), .A2(new_n863), .B(new_n876), .C(new_n872), .Y(new_n888));
  A2O1A1Ixp33_ASAP7_75t_L   g0503(.A1(\b[53] ), .A2(\a[53] ), .B(new_n888), .C(new_n881), .Y(new_n889));
  INVx1_ASAP7_75t_L         g0504(.A(\a[55] ), .Y(new_n890));
  INVx1_ASAP7_75t_L         g0505(.A(\b[55] ), .Y(new_n891));
  NAND2xp33_ASAP7_75t_L     g0506(.A(new_n891), .B(new_n890), .Y(new_n892));
  NOR2xp33_ASAP7_75t_L      g0507(.A(new_n890), .B(new_n891), .Y(new_n893));
  INVx1_ASAP7_75t_L         g0508(.A(new_n893), .Y(new_n894));
  NAND2xp33_ASAP7_75t_L     g0509(.A(new_n892), .B(new_n894), .Y(new_n895));
  AND3x1_ASAP7_75t_L        g0510(.A(new_n889), .B(new_n895), .C(new_n883), .Y(new_n896));
  O2A1O1Ixp33_ASAP7_75t_L   g0511(.A1(new_n879), .A2(new_n880), .B(new_n889), .C(new_n895), .Y(new_n897));
  NOR2xp33_ASAP7_75t_L      g0512(.A(new_n897), .B(new_n896), .Y(\f[55] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0513(.A1(new_n881), .A2(new_n878), .B(new_n882), .C(new_n892), .D(new_n893), .Y(new_n899));
  NOR2xp33_ASAP7_75t_L      g0514(.A(\a[56] ), .B(\b[56] ), .Y(new_n900));
  AND2x2_ASAP7_75t_L        g0515(.A(\a[56] ), .B(\b[56] ), .Y(new_n901));
  NOR2xp33_ASAP7_75t_L      g0516(.A(new_n900), .B(new_n901), .Y(new_n902));
  XNOR2x2_ASAP7_75t_L       g0517(.A(new_n902), .B(new_n899), .Y(\f[56] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0518(.A1(new_n878), .A2(new_n881), .B(new_n882), .C(new_n892), .Y(new_n904));
  NAND2xp33_ASAP7_75t_L     g0519(.A(\b[56] ), .B(\a[56] ), .Y(new_n905));
  A2O1A1Ixp33_ASAP7_75t_L   g0520(.A1(new_n904), .A2(new_n894), .B(new_n900), .C(new_n905), .Y(new_n906));
  INVx1_ASAP7_75t_L         g0521(.A(\a[57] ), .Y(new_n907));
  INVx1_ASAP7_75t_L         g0522(.A(\b[57] ), .Y(new_n908));
  NAND2xp33_ASAP7_75t_L     g0523(.A(new_n908), .B(new_n907), .Y(new_n909));
  NOR2xp33_ASAP7_75t_L      g0524(.A(new_n907), .B(new_n908), .Y(new_n910));
  INVx1_ASAP7_75t_L         g0525(.A(new_n910), .Y(new_n911));
  AOI21xp33_ASAP7_75t_L     g0526(.A1(new_n911), .A2(new_n909), .B(new_n906), .Y(new_n912));
  NAND2xp33_ASAP7_75t_L     g0527(.A(new_n909), .B(new_n911), .Y(new_n913));
  A2O1A1O1Ixp25_ASAP7_75t_L g0528(.A1(new_n894), .A2(new_n904), .B(new_n900), .C(new_n905), .D(new_n913), .Y(new_n914));
  NOR2xp33_ASAP7_75t_L      g0529(.A(new_n914), .B(new_n912), .Y(\f[57] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0530(.A1(new_n890), .A2(new_n891), .B(new_n904), .C(new_n900), .Y(new_n916));
  A2O1A1Ixp33_ASAP7_75t_L   g0531(.A1(\b[56] ), .A2(\a[56] ), .B(new_n916), .C(new_n909), .Y(new_n917));
  INVx1_ASAP7_75t_L         g0532(.A(\a[58] ), .Y(new_n918));
  INVx1_ASAP7_75t_L         g0533(.A(\b[58] ), .Y(new_n919));
  NAND2xp33_ASAP7_75t_L     g0534(.A(new_n919), .B(new_n918), .Y(new_n920));
  NOR2xp33_ASAP7_75t_L      g0535(.A(new_n918), .B(new_n919), .Y(new_n921));
  INVx1_ASAP7_75t_L         g0536(.A(new_n921), .Y(new_n922));
  NAND2xp33_ASAP7_75t_L     g0537(.A(new_n920), .B(new_n922), .Y(new_n923));
  AND3x1_ASAP7_75t_L        g0538(.A(new_n917), .B(new_n923), .C(new_n911), .Y(new_n924));
  O2A1O1Ixp33_ASAP7_75t_L   g0539(.A1(new_n907), .A2(new_n908), .B(new_n917), .C(new_n923), .Y(new_n925));
  NOR2xp33_ASAP7_75t_L      g0540(.A(new_n925), .B(new_n924), .Y(\f[58] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0541(.A1(new_n909), .A2(new_n906), .B(new_n910), .C(new_n920), .D(new_n921), .Y(new_n927));
  NOR2xp33_ASAP7_75t_L      g0542(.A(\a[59] ), .B(\b[59] ), .Y(new_n928));
  AND2x2_ASAP7_75t_L        g0543(.A(\a[59] ), .B(\b[59] ), .Y(new_n929));
  NOR2xp33_ASAP7_75t_L      g0544(.A(new_n928), .B(new_n929), .Y(new_n930));
  XNOR2x2_ASAP7_75t_L       g0545(.A(new_n930), .B(new_n927), .Y(\f[59] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0546(.A1(new_n906), .A2(new_n909), .B(new_n910), .C(new_n920), .Y(new_n932));
  NAND2xp33_ASAP7_75t_L     g0547(.A(\b[59] ), .B(\a[59] ), .Y(new_n933));
  A2O1A1Ixp33_ASAP7_75t_L   g0548(.A1(new_n932), .A2(new_n922), .B(new_n928), .C(new_n933), .Y(new_n934));
  INVx1_ASAP7_75t_L         g0549(.A(\a[60] ), .Y(new_n935));
  INVx1_ASAP7_75t_L         g0550(.A(\b[60] ), .Y(new_n936));
  NAND2xp33_ASAP7_75t_L     g0551(.A(new_n936), .B(new_n935), .Y(new_n937));
  NOR2xp33_ASAP7_75t_L      g0552(.A(new_n935), .B(new_n936), .Y(new_n938));
  INVx1_ASAP7_75t_L         g0553(.A(new_n938), .Y(new_n939));
  AOI21xp33_ASAP7_75t_L     g0554(.A1(new_n939), .A2(new_n937), .B(new_n934), .Y(new_n940));
  NAND2xp33_ASAP7_75t_L     g0555(.A(new_n937), .B(new_n939), .Y(new_n941));
  A2O1A1O1Ixp25_ASAP7_75t_L g0556(.A1(new_n922), .A2(new_n932), .B(new_n928), .C(new_n933), .D(new_n941), .Y(new_n942));
  NOR2xp33_ASAP7_75t_L      g0557(.A(new_n942), .B(new_n940), .Y(\f[60] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0558(.A1(new_n918), .A2(new_n919), .B(new_n932), .C(new_n928), .Y(new_n944));
  A2O1A1Ixp33_ASAP7_75t_L   g0559(.A1(\b[59] ), .A2(\a[59] ), .B(new_n944), .C(new_n937), .Y(new_n945));
  INVx1_ASAP7_75t_L         g0560(.A(\a[61] ), .Y(new_n946));
  INVx1_ASAP7_75t_L         g0561(.A(\b[61] ), .Y(new_n947));
  NAND2xp33_ASAP7_75t_L     g0562(.A(new_n947), .B(new_n946), .Y(new_n948));
  NOR2xp33_ASAP7_75t_L      g0563(.A(new_n946), .B(new_n947), .Y(new_n949));
  INVx1_ASAP7_75t_L         g0564(.A(new_n949), .Y(new_n950));
  NAND2xp33_ASAP7_75t_L     g0565(.A(new_n948), .B(new_n950), .Y(new_n951));
  AND3x1_ASAP7_75t_L        g0566(.A(new_n945), .B(new_n951), .C(new_n939), .Y(new_n952));
  O2A1O1Ixp33_ASAP7_75t_L   g0567(.A1(new_n935), .A2(new_n936), .B(new_n945), .C(new_n951), .Y(new_n953));
  NOR2xp33_ASAP7_75t_L      g0568(.A(new_n953), .B(new_n952), .Y(\f[61] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0569(.A1(new_n937), .A2(new_n934), .B(new_n938), .C(new_n948), .D(new_n949), .Y(new_n955));
  NOR2xp33_ASAP7_75t_L      g0570(.A(\a[62] ), .B(\b[62] ), .Y(new_n956));
  AND2x2_ASAP7_75t_L        g0571(.A(\a[62] ), .B(\b[62] ), .Y(new_n957));
  NOR2xp33_ASAP7_75t_L      g0572(.A(new_n956), .B(new_n957), .Y(new_n958));
  XNOR2x2_ASAP7_75t_L       g0573(.A(new_n958), .B(new_n955), .Y(\f[62] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0574(.A1(new_n934), .A2(new_n937), .B(new_n938), .C(new_n948), .Y(new_n960));
  NAND2xp33_ASAP7_75t_L     g0575(.A(\b[62] ), .B(\a[62] ), .Y(new_n961));
  A2O1A1Ixp33_ASAP7_75t_L   g0576(.A1(new_n960), .A2(new_n950), .B(new_n956), .C(new_n961), .Y(new_n962));
  INVx1_ASAP7_75t_L         g0577(.A(\a[63] ), .Y(new_n963));
  INVx1_ASAP7_75t_L         g0578(.A(\b[63] ), .Y(new_n964));
  NAND2xp33_ASAP7_75t_L     g0579(.A(new_n964), .B(new_n963), .Y(new_n965));
  NOR2xp33_ASAP7_75t_L      g0580(.A(new_n963), .B(new_n964), .Y(new_n966));
  INVx1_ASAP7_75t_L         g0581(.A(new_n966), .Y(new_n967));
  AOI21xp33_ASAP7_75t_L     g0582(.A1(new_n967), .A2(new_n965), .B(new_n962), .Y(new_n968));
  NAND2xp33_ASAP7_75t_L     g0583(.A(new_n965), .B(new_n967), .Y(new_n969));
  A2O1A1O1Ixp25_ASAP7_75t_L g0584(.A1(new_n950), .A2(new_n960), .B(new_n956), .C(new_n961), .D(new_n969), .Y(new_n970));
  NOR2xp33_ASAP7_75t_L      g0585(.A(new_n970), .B(new_n968), .Y(\f[63] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0586(.A1(new_n946), .A2(new_n947), .B(new_n960), .C(new_n956), .Y(new_n972));
  A2O1A1Ixp33_ASAP7_75t_L   g0587(.A1(\b[62] ), .A2(\a[62] ), .B(new_n972), .C(new_n965), .Y(new_n973));
  INVx1_ASAP7_75t_L         g0588(.A(\a[64] ), .Y(new_n974));
  INVx1_ASAP7_75t_L         g0589(.A(\b[64] ), .Y(new_n975));
  NAND2xp33_ASAP7_75t_L     g0590(.A(new_n975), .B(new_n974), .Y(new_n976));
  NOR2xp33_ASAP7_75t_L      g0591(.A(new_n974), .B(new_n975), .Y(new_n977));
  INVx1_ASAP7_75t_L         g0592(.A(new_n977), .Y(new_n978));
  NAND2xp33_ASAP7_75t_L     g0593(.A(new_n976), .B(new_n978), .Y(new_n979));
  AND3x1_ASAP7_75t_L        g0594(.A(new_n973), .B(new_n979), .C(new_n967), .Y(new_n980));
  O2A1O1Ixp33_ASAP7_75t_L   g0595(.A1(new_n963), .A2(new_n964), .B(new_n973), .C(new_n979), .Y(new_n981));
  NOR2xp33_ASAP7_75t_L      g0596(.A(new_n981), .B(new_n980), .Y(\f[64] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0597(.A1(new_n965), .A2(new_n962), .B(new_n966), .C(new_n976), .D(new_n977), .Y(new_n983));
  NOR2xp33_ASAP7_75t_L      g0598(.A(\a[65] ), .B(\b[65] ), .Y(new_n984));
  AND2x2_ASAP7_75t_L        g0599(.A(\a[65] ), .B(\b[65] ), .Y(new_n985));
  NOR2xp33_ASAP7_75t_L      g0600(.A(new_n984), .B(new_n985), .Y(new_n986));
  XNOR2x2_ASAP7_75t_L       g0601(.A(new_n986), .B(new_n983), .Y(\f[65] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0602(.A1(new_n962), .A2(new_n965), .B(new_n966), .C(new_n976), .Y(new_n988));
  NAND2xp33_ASAP7_75t_L     g0603(.A(\b[65] ), .B(\a[65] ), .Y(new_n989));
  A2O1A1Ixp33_ASAP7_75t_L   g0604(.A1(new_n988), .A2(new_n978), .B(new_n984), .C(new_n989), .Y(new_n990));
  INVx1_ASAP7_75t_L         g0605(.A(\a[66] ), .Y(new_n991));
  INVx1_ASAP7_75t_L         g0606(.A(\b[66] ), .Y(new_n992));
  NAND2xp33_ASAP7_75t_L     g0607(.A(new_n992), .B(new_n991), .Y(new_n993));
  NOR2xp33_ASAP7_75t_L      g0608(.A(new_n991), .B(new_n992), .Y(new_n994));
  INVx1_ASAP7_75t_L         g0609(.A(new_n994), .Y(new_n995));
  AOI21xp33_ASAP7_75t_L     g0610(.A1(new_n995), .A2(new_n993), .B(new_n990), .Y(new_n996));
  NAND2xp33_ASAP7_75t_L     g0611(.A(new_n993), .B(new_n995), .Y(new_n997));
  A2O1A1O1Ixp25_ASAP7_75t_L g0612(.A1(new_n978), .A2(new_n988), .B(new_n984), .C(new_n989), .D(new_n997), .Y(new_n998));
  NOR2xp33_ASAP7_75t_L      g0613(.A(new_n998), .B(new_n996), .Y(\f[66] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0614(.A1(new_n974), .A2(new_n975), .B(new_n988), .C(new_n984), .Y(new_n1000));
  A2O1A1Ixp33_ASAP7_75t_L   g0615(.A1(\b[65] ), .A2(\a[65] ), .B(new_n1000), .C(new_n993), .Y(new_n1001));
  INVx1_ASAP7_75t_L         g0616(.A(\a[67] ), .Y(new_n1002));
  INVx1_ASAP7_75t_L         g0617(.A(\b[67] ), .Y(new_n1003));
  NAND2xp33_ASAP7_75t_L     g0618(.A(new_n1003), .B(new_n1002), .Y(new_n1004));
  NOR2xp33_ASAP7_75t_L      g0619(.A(new_n1002), .B(new_n1003), .Y(new_n1005));
  INVx1_ASAP7_75t_L         g0620(.A(new_n1005), .Y(new_n1006));
  NAND2xp33_ASAP7_75t_L     g0621(.A(new_n1004), .B(new_n1006), .Y(new_n1007));
  AND3x1_ASAP7_75t_L        g0622(.A(new_n1001), .B(new_n1007), .C(new_n995), .Y(new_n1008));
  O2A1O1Ixp33_ASAP7_75t_L   g0623(.A1(new_n991), .A2(new_n992), .B(new_n1001), .C(new_n1007), .Y(new_n1009));
  NOR2xp33_ASAP7_75t_L      g0624(.A(new_n1009), .B(new_n1008), .Y(\f[67] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0625(.A1(new_n993), .A2(new_n990), .B(new_n994), .C(new_n1004), .D(new_n1005), .Y(new_n1011));
  NOR2xp33_ASAP7_75t_L      g0626(.A(\a[68] ), .B(\b[68] ), .Y(new_n1012));
  AND2x2_ASAP7_75t_L        g0627(.A(\a[68] ), .B(\b[68] ), .Y(new_n1013));
  NOR2xp33_ASAP7_75t_L      g0628(.A(new_n1012), .B(new_n1013), .Y(new_n1014));
  XNOR2x2_ASAP7_75t_L       g0629(.A(new_n1014), .B(new_n1011), .Y(\f[68] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0630(.A1(new_n990), .A2(new_n993), .B(new_n994), .C(new_n1004), .Y(new_n1016));
  NAND2xp33_ASAP7_75t_L     g0631(.A(\b[68] ), .B(\a[68] ), .Y(new_n1017));
  A2O1A1Ixp33_ASAP7_75t_L   g0632(.A1(new_n1016), .A2(new_n1006), .B(new_n1012), .C(new_n1017), .Y(new_n1018));
  INVx1_ASAP7_75t_L         g0633(.A(\a[69] ), .Y(new_n1019));
  INVx1_ASAP7_75t_L         g0634(.A(\b[69] ), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g0635(.A(new_n1020), .B(new_n1019), .Y(new_n1021));
  NOR2xp33_ASAP7_75t_L      g0636(.A(new_n1019), .B(new_n1020), .Y(new_n1022));
  INVx1_ASAP7_75t_L         g0637(.A(new_n1022), .Y(new_n1023));
  AOI21xp33_ASAP7_75t_L     g0638(.A1(new_n1023), .A2(new_n1021), .B(new_n1018), .Y(new_n1024));
  NAND2xp33_ASAP7_75t_L     g0639(.A(new_n1021), .B(new_n1023), .Y(new_n1025));
  A2O1A1O1Ixp25_ASAP7_75t_L g0640(.A1(new_n1006), .A2(new_n1016), .B(new_n1012), .C(new_n1017), .D(new_n1025), .Y(new_n1026));
  NOR2xp33_ASAP7_75t_L      g0641(.A(new_n1026), .B(new_n1024), .Y(\f[69] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0642(.A1(new_n1002), .A2(new_n1003), .B(new_n1016), .C(new_n1012), .Y(new_n1028));
  A2O1A1Ixp33_ASAP7_75t_L   g0643(.A1(\b[68] ), .A2(\a[68] ), .B(new_n1028), .C(new_n1021), .Y(new_n1029));
  INVx1_ASAP7_75t_L         g0644(.A(\a[70] ), .Y(new_n1030));
  INVx1_ASAP7_75t_L         g0645(.A(\b[70] ), .Y(new_n1031));
  NAND2xp33_ASAP7_75t_L     g0646(.A(new_n1031), .B(new_n1030), .Y(new_n1032));
  NOR2xp33_ASAP7_75t_L      g0647(.A(new_n1030), .B(new_n1031), .Y(new_n1033));
  INVx1_ASAP7_75t_L         g0648(.A(new_n1033), .Y(new_n1034));
  NAND2xp33_ASAP7_75t_L     g0649(.A(new_n1032), .B(new_n1034), .Y(new_n1035));
  AND3x1_ASAP7_75t_L        g0650(.A(new_n1029), .B(new_n1035), .C(new_n1023), .Y(new_n1036));
  O2A1O1Ixp33_ASAP7_75t_L   g0651(.A1(new_n1019), .A2(new_n1020), .B(new_n1029), .C(new_n1035), .Y(new_n1037));
  NOR2xp33_ASAP7_75t_L      g0652(.A(new_n1037), .B(new_n1036), .Y(\f[70] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0653(.A1(new_n1021), .A2(new_n1018), .B(new_n1022), .C(new_n1032), .D(new_n1033), .Y(new_n1039));
  NOR2xp33_ASAP7_75t_L      g0654(.A(\a[71] ), .B(\b[71] ), .Y(new_n1040));
  AND2x2_ASAP7_75t_L        g0655(.A(\a[71] ), .B(\b[71] ), .Y(new_n1041));
  NOR2xp33_ASAP7_75t_L      g0656(.A(new_n1040), .B(new_n1041), .Y(new_n1042));
  XNOR2x2_ASAP7_75t_L       g0657(.A(new_n1042), .B(new_n1039), .Y(\f[71] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0658(.A1(new_n1018), .A2(new_n1021), .B(new_n1022), .C(new_n1032), .Y(new_n1044));
  NAND2xp33_ASAP7_75t_L     g0659(.A(\b[71] ), .B(\a[71] ), .Y(new_n1045));
  A2O1A1Ixp33_ASAP7_75t_L   g0660(.A1(new_n1044), .A2(new_n1034), .B(new_n1040), .C(new_n1045), .Y(new_n1046));
  INVx1_ASAP7_75t_L         g0661(.A(\a[72] ), .Y(new_n1047));
  INVx1_ASAP7_75t_L         g0662(.A(\b[72] ), .Y(new_n1048));
  NAND2xp33_ASAP7_75t_L     g0663(.A(new_n1048), .B(new_n1047), .Y(new_n1049));
  NOR2xp33_ASAP7_75t_L      g0664(.A(new_n1047), .B(new_n1048), .Y(new_n1050));
  INVx1_ASAP7_75t_L         g0665(.A(new_n1050), .Y(new_n1051));
  AOI21xp33_ASAP7_75t_L     g0666(.A1(new_n1051), .A2(new_n1049), .B(new_n1046), .Y(new_n1052));
  NAND2xp33_ASAP7_75t_L     g0667(.A(new_n1049), .B(new_n1051), .Y(new_n1053));
  A2O1A1O1Ixp25_ASAP7_75t_L g0668(.A1(new_n1034), .A2(new_n1044), .B(new_n1040), .C(new_n1045), .D(new_n1053), .Y(new_n1054));
  NOR2xp33_ASAP7_75t_L      g0669(.A(new_n1054), .B(new_n1052), .Y(\f[72] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0670(.A1(new_n1030), .A2(new_n1031), .B(new_n1044), .C(new_n1040), .Y(new_n1056));
  A2O1A1Ixp33_ASAP7_75t_L   g0671(.A1(\b[71] ), .A2(\a[71] ), .B(new_n1056), .C(new_n1049), .Y(new_n1057));
  INVx1_ASAP7_75t_L         g0672(.A(\a[73] ), .Y(new_n1058));
  INVx1_ASAP7_75t_L         g0673(.A(\b[73] ), .Y(new_n1059));
  NAND2xp33_ASAP7_75t_L     g0674(.A(new_n1059), .B(new_n1058), .Y(new_n1060));
  NOR2xp33_ASAP7_75t_L      g0675(.A(new_n1058), .B(new_n1059), .Y(new_n1061));
  INVx1_ASAP7_75t_L         g0676(.A(new_n1061), .Y(new_n1062));
  NAND2xp33_ASAP7_75t_L     g0677(.A(new_n1060), .B(new_n1062), .Y(new_n1063));
  AND3x1_ASAP7_75t_L        g0678(.A(new_n1057), .B(new_n1063), .C(new_n1051), .Y(new_n1064));
  O2A1O1Ixp33_ASAP7_75t_L   g0679(.A1(new_n1047), .A2(new_n1048), .B(new_n1057), .C(new_n1063), .Y(new_n1065));
  NOR2xp33_ASAP7_75t_L      g0680(.A(new_n1065), .B(new_n1064), .Y(\f[73] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0681(.A1(new_n1049), .A2(new_n1046), .B(new_n1050), .C(new_n1060), .D(new_n1061), .Y(new_n1067));
  NOR2xp33_ASAP7_75t_L      g0682(.A(\a[74] ), .B(\b[74] ), .Y(new_n1068));
  AND2x2_ASAP7_75t_L        g0683(.A(\a[74] ), .B(\b[74] ), .Y(new_n1069));
  NOR2xp33_ASAP7_75t_L      g0684(.A(new_n1068), .B(new_n1069), .Y(new_n1070));
  XNOR2x2_ASAP7_75t_L       g0685(.A(new_n1070), .B(new_n1067), .Y(\f[74] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0686(.A1(new_n1046), .A2(new_n1049), .B(new_n1050), .C(new_n1060), .Y(new_n1072));
  NAND2xp33_ASAP7_75t_L     g0687(.A(\b[74] ), .B(\a[74] ), .Y(new_n1073));
  A2O1A1Ixp33_ASAP7_75t_L   g0688(.A1(new_n1072), .A2(new_n1062), .B(new_n1068), .C(new_n1073), .Y(new_n1074));
  INVx1_ASAP7_75t_L         g0689(.A(\a[75] ), .Y(new_n1075));
  INVx1_ASAP7_75t_L         g0690(.A(\b[75] ), .Y(new_n1076));
  NAND2xp33_ASAP7_75t_L     g0691(.A(new_n1076), .B(new_n1075), .Y(new_n1077));
  NOR2xp33_ASAP7_75t_L      g0692(.A(new_n1075), .B(new_n1076), .Y(new_n1078));
  INVx1_ASAP7_75t_L         g0693(.A(new_n1078), .Y(new_n1079));
  AOI21xp33_ASAP7_75t_L     g0694(.A1(new_n1079), .A2(new_n1077), .B(new_n1074), .Y(new_n1080));
  NAND2xp33_ASAP7_75t_L     g0695(.A(new_n1077), .B(new_n1079), .Y(new_n1081));
  A2O1A1O1Ixp25_ASAP7_75t_L g0696(.A1(new_n1062), .A2(new_n1072), .B(new_n1068), .C(new_n1073), .D(new_n1081), .Y(new_n1082));
  NOR2xp33_ASAP7_75t_L      g0697(.A(new_n1082), .B(new_n1080), .Y(\f[75] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0698(.A1(new_n1058), .A2(new_n1059), .B(new_n1072), .C(new_n1068), .Y(new_n1084));
  A2O1A1Ixp33_ASAP7_75t_L   g0699(.A1(\b[74] ), .A2(\a[74] ), .B(new_n1084), .C(new_n1077), .Y(new_n1085));
  INVx1_ASAP7_75t_L         g0700(.A(\a[76] ), .Y(new_n1086));
  INVx1_ASAP7_75t_L         g0701(.A(\b[76] ), .Y(new_n1087));
  NAND2xp33_ASAP7_75t_L     g0702(.A(new_n1087), .B(new_n1086), .Y(new_n1088));
  NOR2xp33_ASAP7_75t_L      g0703(.A(new_n1086), .B(new_n1087), .Y(new_n1089));
  INVx1_ASAP7_75t_L         g0704(.A(new_n1089), .Y(new_n1090));
  NAND2xp33_ASAP7_75t_L     g0705(.A(new_n1088), .B(new_n1090), .Y(new_n1091));
  AND3x1_ASAP7_75t_L        g0706(.A(new_n1085), .B(new_n1091), .C(new_n1079), .Y(new_n1092));
  O2A1O1Ixp33_ASAP7_75t_L   g0707(.A1(new_n1075), .A2(new_n1076), .B(new_n1085), .C(new_n1091), .Y(new_n1093));
  NOR2xp33_ASAP7_75t_L      g0708(.A(new_n1093), .B(new_n1092), .Y(\f[76] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0709(.A1(new_n1077), .A2(new_n1074), .B(new_n1078), .C(new_n1088), .D(new_n1089), .Y(new_n1095));
  NOR2xp33_ASAP7_75t_L      g0710(.A(\a[77] ), .B(\b[77] ), .Y(new_n1096));
  AND2x2_ASAP7_75t_L        g0711(.A(\a[77] ), .B(\b[77] ), .Y(new_n1097));
  NOR2xp33_ASAP7_75t_L      g0712(.A(new_n1096), .B(new_n1097), .Y(new_n1098));
  XNOR2x2_ASAP7_75t_L       g0713(.A(new_n1098), .B(new_n1095), .Y(\f[77] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0714(.A1(new_n1074), .A2(new_n1077), .B(new_n1078), .C(new_n1088), .Y(new_n1100));
  NAND2xp33_ASAP7_75t_L     g0715(.A(\b[77] ), .B(\a[77] ), .Y(new_n1101));
  A2O1A1Ixp33_ASAP7_75t_L   g0716(.A1(new_n1100), .A2(new_n1090), .B(new_n1096), .C(new_n1101), .Y(new_n1102));
  INVx1_ASAP7_75t_L         g0717(.A(\a[78] ), .Y(new_n1103));
  INVx1_ASAP7_75t_L         g0718(.A(\b[78] ), .Y(new_n1104));
  NAND2xp33_ASAP7_75t_L     g0719(.A(new_n1104), .B(new_n1103), .Y(new_n1105));
  NOR2xp33_ASAP7_75t_L      g0720(.A(new_n1103), .B(new_n1104), .Y(new_n1106));
  INVx1_ASAP7_75t_L         g0721(.A(new_n1106), .Y(new_n1107));
  AOI21xp33_ASAP7_75t_L     g0722(.A1(new_n1107), .A2(new_n1105), .B(new_n1102), .Y(new_n1108));
  NAND2xp33_ASAP7_75t_L     g0723(.A(new_n1105), .B(new_n1107), .Y(new_n1109));
  A2O1A1O1Ixp25_ASAP7_75t_L g0724(.A1(new_n1090), .A2(new_n1100), .B(new_n1096), .C(new_n1101), .D(new_n1109), .Y(new_n1110));
  NOR2xp33_ASAP7_75t_L      g0725(.A(new_n1110), .B(new_n1108), .Y(\f[78] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0726(.A1(new_n1086), .A2(new_n1087), .B(new_n1100), .C(new_n1096), .Y(new_n1112));
  A2O1A1Ixp33_ASAP7_75t_L   g0727(.A1(\b[77] ), .A2(\a[77] ), .B(new_n1112), .C(new_n1105), .Y(new_n1113));
  INVx1_ASAP7_75t_L         g0728(.A(\a[79] ), .Y(new_n1114));
  INVx1_ASAP7_75t_L         g0729(.A(\b[79] ), .Y(new_n1115));
  NAND2xp33_ASAP7_75t_L     g0730(.A(new_n1115), .B(new_n1114), .Y(new_n1116));
  NOR2xp33_ASAP7_75t_L      g0731(.A(new_n1114), .B(new_n1115), .Y(new_n1117));
  INVx1_ASAP7_75t_L         g0732(.A(new_n1117), .Y(new_n1118));
  NAND2xp33_ASAP7_75t_L     g0733(.A(new_n1116), .B(new_n1118), .Y(new_n1119));
  AND3x1_ASAP7_75t_L        g0734(.A(new_n1113), .B(new_n1119), .C(new_n1107), .Y(new_n1120));
  O2A1O1Ixp33_ASAP7_75t_L   g0735(.A1(new_n1103), .A2(new_n1104), .B(new_n1113), .C(new_n1119), .Y(new_n1121));
  NOR2xp33_ASAP7_75t_L      g0736(.A(new_n1121), .B(new_n1120), .Y(\f[79] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0737(.A1(new_n1105), .A2(new_n1102), .B(new_n1106), .C(new_n1116), .D(new_n1117), .Y(new_n1123));
  NOR2xp33_ASAP7_75t_L      g0738(.A(\a[80] ), .B(\b[80] ), .Y(new_n1124));
  AND2x2_ASAP7_75t_L        g0739(.A(\a[80] ), .B(\b[80] ), .Y(new_n1125));
  NOR2xp33_ASAP7_75t_L      g0740(.A(new_n1124), .B(new_n1125), .Y(new_n1126));
  XNOR2x2_ASAP7_75t_L       g0741(.A(new_n1126), .B(new_n1123), .Y(\f[80] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0742(.A1(new_n1102), .A2(new_n1105), .B(new_n1106), .C(new_n1116), .Y(new_n1128));
  NAND2xp33_ASAP7_75t_L     g0743(.A(\b[80] ), .B(\a[80] ), .Y(new_n1129));
  A2O1A1Ixp33_ASAP7_75t_L   g0744(.A1(new_n1128), .A2(new_n1118), .B(new_n1124), .C(new_n1129), .Y(new_n1130));
  INVx1_ASAP7_75t_L         g0745(.A(\a[81] ), .Y(new_n1131));
  INVx1_ASAP7_75t_L         g0746(.A(\b[81] ), .Y(new_n1132));
  NAND2xp33_ASAP7_75t_L     g0747(.A(new_n1132), .B(new_n1131), .Y(new_n1133));
  NOR2xp33_ASAP7_75t_L      g0748(.A(new_n1131), .B(new_n1132), .Y(new_n1134));
  INVx1_ASAP7_75t_L         g0749(.A(new_n1134), .Y(new_n1135));
  AOI21xp33_ASAP7_75t_L     g0750(.A1(new_n1135), .A2(new_n1133), .B(new_n1130), .Y(new_n1136));
  NAND2xp33_ASAP7_75t_L     g0751(.A(new_n1133), .B(new_n1135), .Y(new_n1137));
  A2O1A1O1Ixp25_ASAP7_75t_L g0752(.A1(new_n1118), .A2(new_n1128), .B(new_n1124), .C(new_n1129), .D(new_n1137), .Y(new_n1138));
  NOR2xp33_ASAP7_75t_L      g0753(.A(new_n1138), .B(new_n1136), .Y(\f[81] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0754(.A1(new_n1114), .A2(new_n1115), .B(new_n1128), .C(new_n1124), .Y(new_n1140));
  A2O1A1Ixp33_ASAP7_75t_L   g0755(.A1(\b[80] ), .A2(\a[80] ), .B(new_n1140), .C(new_n1133), .Y(new_n1141));
  INVx1_ASAP7_75t_L         g0756(.A(\a[82] ), .Y(new_n1142));
  INVx1_ASAP7_75t_L         g0757(.A(\b[82] ), .Y(new_n1143));
  NAND2xp33_ASAP7_75t_L     g0758(.A(new_n1143), .B(new_n1142), .Y(new_n1144));
  NOR2xp33_ASAP7_75t_L      g0759(.A(new_n1142), .B(new_n1143), .Y(new_n1145));
  INVx1_ASAP7_75t_L         g0760(.A(new_n1145), .Y(new_n1146));
  NAND2xp33_ASAP7_75t_L     g0761(.A(new_n1144), .B(new_n1146), .Y(new_n1147));
  AND3x1_ASAP7_75t_L        g0762(.A(new_n1141), .B(new_n1147), .C(new_n1135), .Y(new_n1148));
  O2A1O1Ixp33_ASAP7_75t_L   g0763(.A1(new_n1131), .A2(new_n1132), .B(new_n1141), .C(new_n1147), .Y(new_n1149));
  NOR2xp33_ASAP7_75t_L      g0764(.A(new_n1149), .B(new_n1148), .Y(\f[82] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0765(.A1(new_n1133), .A2(new_n1130), .B(new_n1134), .C(new_n1144), .D(new_n1145), .Y(new_n1151));
  NOR2xp33_ASAP7_75t_L      g0766(.A(\a[83] ), .B(\b[83] ), .Y(new_n1152));
  AND2x2_ASAP7_75t_L        g0767(.A(\a[83] ), .B(\b[83] ), .Y(new_n1153));
  NOR2xp33_ASAP7_75t_L      g0768(.A(new_n1152), .B(new_n1153), .Y(new_n1154));
  XNOR2x2_ASAP7_75t_L       g0769(.A(new_n1154), .B(new_n1151), .Y(\f[83] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0770(.A1(new_n1130), .A2(new_n1133), .B(new_n1134), .C(new_n1144), .Y(new_n1156));
  NAND2xp33_ASAP7_75t_L     g0771(.A(\b[83] ), .B(\a[83] ), .Y(new_n1157));
  A2O1A1Ixp33_ASAP7_75t_L   g0772(.A1(new_n1156), .A2(new_n1146), .B(new_n1152), .C(new_n1157), .Y(new_n1158));
  INVx1_ASAP7_75t_L         g0773(.A(\a[84] ), .Y(new_n1159));
  INVx1_ASAP7_75t_L         g0774(.A(\b[84] ), .Y(new_n1160));
  NAND2xp33_ASAP7_75t_L     g0775(.A(new_n1160), .B(new_n1159), .Y(new_n1161));
  NOR2xp33_ASAP7_75t_L      g0776(.A(new_n1159), .B(new_n1160), .Y(new_n1162));
  INVx1_ASAP7_75t_L         g0777(.A(new_n1162), .Y(new_n1163));
  AOI21xp33_ASAP7_75t_L     g0778(.A1(new_n1163), .A2(new_n1161), .B(new_n1158), .Y(new_n1164));
  NAND2xp33_ASAP7_75t_L     g0779(.A(new_n1161), .B(new_n1163), .Y(new_n1165));
  A2O1A1O1Ixp25_ASAP7_75t_L g0780(.A1(new_n1146), .A2(new_n1156), .B(new_n1152), .C(new_n1157), .D(new_n1165), .Y(new_n1166));
  NOR2xp33_ASAP7_75t_L      g0781(.A(new_n1166), .B(new_n1164), .Y(\f[84] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0782(.A1(new_n1142), .A2(new_n1143), .B(new_n1156), .C(new_n1152), .Y(new_n1168));
  A2O1A1Ixp33_ASAP7_75t_L   g0783(.A1(\b[83] ), .A2(\a[83] ), .B(new_n1168), .C(new_n1161), .Y(new_n1169));
  INVx1_ASAP7_75t_L         g0784(.A(\a[85] ), .Y(new_n1170));
  INVx1_ASAP7_75t_L         g0785(.A(\b[85] ), .Y(new_n1171));
  NAND2xp33_ASAP7_75t_L     g0786(.A(new_n1171), .B(new_n1170), .Y(new_n1172));
  NOR2xp33_ASAP7_75t_L      g0787(.A(new_n1170), .B(new_n1171), .Y(new_n1173));
  INVx1_ASAP7_75t_L         g0788(.A(new_n1173), .Y(new_n1174));
  NAND2xp33_ASAP7_75t_L     g0789(.A(new_n1172), .B(new_n1174), .Y(new_n1175));
  AND3x1_ASAP7_75t_L        g0790(.A(new_n1169), .B(new_n1175), .C(new_n1163), .Y(new_n1176));
  O2A1O1Ixp33_ASAP7_75t_L   g0791(.A1(new_n1159), .A2(new_n1160), .B(new_n1169), .C(new_n1175), .Y(new_n1177));
  NOR2xp33_ASAP7_75t_L      g0792(.A(new_n1177), .B(new_n1176), .Y(\f[85] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0793(.A1(new_n1161), .A2(new_n1158), .B(new_n1162), .C(new_n1172), .D(new_n1173), .Y(new_n1179));
  NOR2xp33_ASAP7_75t_L      g0794(.A(\a[86] ), .B(\b[86] ), .Y(new_n1180));
  AND2x2_ASAP7_75t_L        g0795(.A(\a[86] ), .B(\b[86] ), .Y(new_n1181));
  NOR2xp33_ASAP7_75t_L      g0796(.A(new_n1180), .B(new_n1181), .Y(new_n1182));
  XNOR2x2_ASAP7_75t_L       g0797(.A(new_n1182), .B(new_n1179), .Y(\f[86] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0798(.A1(new_n1158), .A2(new_n1161), .B(new_n1162), .C(new_n1172), .Y(new_n1184));
  NAND2xp33_ASAP7_75t_L     g0799(.A(\b[86] ), .B(\a[86] ), .Y(new_n1185));
  A2O1A1Ixp33_ASAP7_75t_L   g0800(.A1(new_n1184), .A2(new_n1174), .B(new_n1180), .C(new_n1185), .Y(new_n1186));
  INVx1_ASAP7_75t_L         g0801(.A(\a[87] ), .Y(new_n1187));
  INVx1_ASAP7_75t_L         g0802(.A(\b[87] ), .Y(new_n1188));
  NAND2xp33_ASAP7_75t_L     g0803(.A(new_n1188), .B(new_n1187), .Y(new_n1189));
  NOR2xp33_ASAP7_75t_L      g0804(.A(new_n1187), .B(new_n1188), .Y(new_n1190));
  INVx1_ASAP7_75t_L         g0805(.A(new_n1190), .Y(new_n1191));
  AOI21xp33_ASAP7_75t_L     g0806(.A1(new_n1191), .A2(new_n1189), .B(new_n1186), .Y(new_n1192));
  NAND2xp33_ASAP7_75t_L     g0807(.A(new_n1189), .B(new_n1191), .Y(new_n1193));
  A2O1A1O1Ixp25_ASAP7_75t_L g0808(.A1(new_n1174), .A2(new_n1184), .B(new_n1180), .C(new_n1185), .D(new_n1193), .Y(new_n1194));
  NOR2xp33_ASAP7_75t_L      g0809(.A(new_n1194), .B(new_n1192), .Y(\f[87] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0810(.A1(new_n1170), .A2(new_n1171), .B(new_n1184), .C(new_n1180), .Y(new_n1196));
  A2O1A1Ixp33_ASAP7_75t_L   g0811(.A1(\b[86] ), .A2(\a[86] ), .B(new_n1196), .C(new_n1189), .Y(new_n1197));
  INVx1_ASAP7_75t_L         g0812(.A(\a[88] ), .Y(new_n1198));
  INVx1_ASAP7_75t_L         g0813(.A(\b[88] ), .Y(new_n1199));
  NAND2xp33_ASAP7_75t_L     g0814(.A(new_n1199), .B(new_n1198), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g0815(.A(new_n1198), .B(new_n1199), .Y(new_n1201));
  INVx1_ASAP7_75t_L         g0816(.A(new_n1201), .Y(new_n1202));
  NAND2xp33_ASAP7_75t_L     g0817(.A(new_n1200), .B(new_n1202), .Y(new_n1203));
  AND3x1_ASAP7_75t_L        g0818(.A(new_n1197), .B(new_n1203), .C(new_n1191), .Y(new_n1204));
  O2A1O1Ixp33_ASAP7_75t_L   g0819(.A1(new_n1187), .A2(new_n1188), .B(new_n1197), .C(new_n1203), .Y(new_n1205));
  NOR2xp33_ASAP7_75t_L      g0820(.A(new_n1205), .B(new_n1204), .Y(\f[88] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0821(.A1(new_n1189), .A2(new_n1186), .B(new_n1190), .C(new_n1200), .D(new_n1201), .Y(new_n1207));
  NOR2xp33_ASAP7_75t_L      g0822(.A(\a[89] ), .B(\b[89] ), .Y(new_n1208));
  AND2x2_ASAP7_75t_L        g0823(.A(\a[89] ), .B(\b[89] ), .Y(new_n1209));
  NOR2xp33_ASAP7_75t_L      g0824(.A(new_n1208), .B(new_n1209), .Y(new_n1210));
  XNOR2x2_ASAP7_75t_L       g0825(.A(new_n1210), .B(new_n1207), .Y(\f[89] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0826(.A1(new_n1186), .A2(new_n1189), .B(new_n1190), .C(new_n1200), .Y(new_n1212));
  NAND2xp33_ASAP7_75t_L     g0827(.A(\b[89] ), .B(\a[89] ), .Y(new_n1213));
  A2O1A1Ixp33_ASAP7_75t_L   g0828(.A1(new_n1212), .A2(new_n1202), .B(new_n1208), .C(new_n1213), .Y(new_n1214));
  INVx1_ASAP7_75t_L         g0829(.A(\a[90] ), .Y(new_n1215));
  INVx1_ASAP7_75t_L         g0830(.A(\b[90] ), .Y(new_n1216));
  NAND2xp33_ASAP7_75t_L     g0831(.A(new_n1216), .B(new_n1215), .Y(new_n1217));
  NOR2xp33_ASAP7_75t_L      g0832(.A(new_n1215), .B(new_n1216), .Y(new_n1218));
  INVx1_ASAP7_75t_L         g0833(.A(new_n1218), .Y(new_n1219));
  AOI21xp33_ASAP7_75t_L     g0834(.A1(new_n1219), .A2(new_n1217), .B(new_n1214), .Y(new_n1220));
  NAND2xp33_ASAP7_75t_L     g0835(.A(new_n1217), .B(new_n1219), .Y(new_n1221));
  A2O1A1O1Ixp25_ASAP7_75t_L g0836(.A1(new_n1202), .A2(new_n1212), .B(new_n1208), .C(new_n1213), .D(new_n1221), .Y(new_n1222));
  NOR2xp33_ASAP7_75t_L      g0837(.A(new_n1222), .B(new_n1220), .Y(\f[90] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0838(.A1(new_n1198), .A2(new_n1199), .B(new_n1212), .C(new_n1208), .Y(new_n1224));
  A2O1A1Ixp33_ASAP7_75t_L   g0839(.A1(\b[89] ), .A2(\a[89] ), .B(new_n1224), .C(new_n1217), .Y(new_n1225));
  INVx1_ASAP7_75t_L         g0840(.A(\a[91] ), .Y(new_n1226));
  INVx1_ASAP7_75t_L         g0841(.A(\b[91] ), .Y(new_n1227));
  NAND2xp33_ASAP7_75t_L     g0842(.A(new_n1227), .B(new_n1226), .Y(new_n1228));
  NOR2xp33_ASAP7_75t_L      g0843(.A(new_n1226), .B(new_n1227), .Y(new_n1229));
  INVx1_ASAP7_75t_L         g0844(.A(new_n1229), .Y(new_n1230));
  NAND2xp33_ASAP7_75t_L     g0845(.A(new_n1228), .B(new_n1230), .Y(new_n1231));
  AND3x1_ASAP7_75t_L        g0846(.A(new_n1225), .B(new_n1231), .C(new_n1219), .Y(new_n1232));
  O2A1O1Ixp33_ASAP7_75t_L   g0847(.A1(new_n1215), .A2(new_n1216), .B(new_n1225), .C(new_n1231), .Y(new_n1233));
  NOR2xp33_ASAP7_75t_L      g0848(.A(new_n1233), .B(new_n1232), .Y(\f[91] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0849(.A1(new_n1217), .A2(new_n1214), .B(new_n1218), .C(new_n1228), .D(new_n1229), .Y(new_n1235));
  NOR2xp33_ASAP7_75t_L      g0850(.A(\a[92] ), .B(\b[92] ), .Y(new_n1236));
  AND2x2_ASAP7_75t_L        g0851(.A(\a[92] ), .B(\b[92] ), .Y(new_n1237));
  NOR2xp33_ASAP7_75t_L      g0852(.A(new_n1236), .B(new_n1237), .Y(new_n1238));
  XNOR2x2_ASAP7_75t_L       g0853(.A(new_n1238), .B(new_n1235), .Y(\f[92] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0854(.A1(new_n1214), .A2(new_n1217), .B(new_n1218), .C(new_n1228), .Y(new_n1240));
  NAND2xp33_ASAP7_75t_L     g0855(.A(\b[92] ), .B(\a[92] ), .Y(new_n1241));
  A2O1A1Ixp33_ASAP7_75t_L   g0856(.A1(new_n1240), .A2(new_n1230), .B(new_n1236), .C(new_n1241), .Y(new_n1242));
  INVx1_ASAP7_75t_L         g0857(.A(\a[93] ), .Y(new_n1243));
  INVx1_ASAP7_75t_L         g0858(.A(\b[93] ), .Y(new_n1244));
  NAND2xp33_ASAP7_75t_L     g0859(.A(new_n1244), .B(new_n1243), .Y(new_n1245));
  NOR2xp33_ASAP7_75t_L      g0860(.A(new_n1243), .B(new_n1244), .Y(new_n1246));
  INVx1_ASAP7_75t_L         g0861(.A(new_n1246), .Y(new_n1247));
  AOI21xp33_ASAP7_75t_L     g0862(.A1(new_n1247), .A2(new_n1245), .B(new_n1242), .Y(new_n1248));
  NAND2xp33_ASAP7_75t_L     g0863(.A(new_n1245), .B(new_n1247), .Y(new_n1249));
  A2O1A1O1Ixp25_ASAP7_75t_L g0864(.A1(new_n1230), .A2(new_n1240), .B(new_n1236), .C(new_n1241), .D(new_n1249), .Y(new_n1250));
  NOR2xp33_ASAP7_75t_L      g0865(.A(new_n1250), .B(new_n1248), .Y(\f[93] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0866(.A1(new_n1226), .A2(new_n1227), .B(new_n1240), .C(new_n1236), .Y(new_n1252));
  A2O1A1Ixp33_ASAP7_75t_L   g0867(.A1(\b[92] ), .A2(\a[92] ), .B(new_n1252), .C(new_n1245), .Y(new_n1253));
  INVx1_ASAP7_75t_L         g0868(.A(\a[94] ), .Y(new_n1254));
  INVx1_ASAP7_75t_L         g0869(.A(\b[94] ), .Y(new_n1255));
  NAND2xp33_ASAP7_75t_L     g0870(.A(new_n1255), .B(new_n1254), .Y(new_n1256));
  NOR2xp33_ASAP7_75t_L      g0871(.A(new_n1254), .B(new_n1255), .Y(new_n1257));
  INVx1_ASAP7_75t_L         g0872(.A(new_n1257), .Y(new_n1258));
  NAND2xp33_ASAP7_75t_L     g0873(.A(new_n1256), .B(new_n1258), .Y(new_n1259));
  AND3x1_ASAP7_75t_L        g0874(.A(new_n1253), .B(new_n1259), .C(new_n1247), .Y(new_n1260));
  O2A1O1Ixp33_ASAP7_75t_L   g0875(.A1(new_n1243), .A2(new_n1244), .B(new_n1253), .C(new_n1259), .Y(new_n1261));
  NOR2xp33_ASAP7_75t_L      g0876(.A(new_n1261), .B(new_n1260), .Y(\f[94] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0877(.A1(new_n1245), .A2(new_n1242), .B(new_n1246), .C(new_n1256), .D(new_n1257), .Y(new_n1263));
  NOR2xp33_ASAP7_75t_L      g0878(.A(\a[95] ), .B(\b[95] ), .Y(new_n1264));
  AND2x2_ASAP7_75t_L        g0879(.A(\a[95] ), .B(\b[95] ), .Y(new_n1265));
  NOR2xp33_ASAP7_75t_L      g0880(.A(new_n1264), .B(new_n1265), .Y(new_n1266));
  XNOR2x2_ASAP7_75t_L       g0881(.A(new_n1266), .B(new_n1263), .Y(\f[95] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0882(.A1(new_n1242), .A2(new_n1245), .B(new_n1246), .C(new_n1256), .Y(new_n1268));
  NAND2xp33_ASAP7_75t_L     g0883(.A(\b[95] ), .B(\a[95] ), .Y(new_n1269));
  A2O1A1Ixp33_ASAP7_75t_L   g0884(.A1(new_n1268), .A2(new_n1258), .B(new_n1264), .C(new_n1269), .Y(new_n1270));
  INVx1_ASAP7_75t_L         g0885(.A(\a[96] ), .Y(new_n1271));
  INVx1_ASAP7_75t_L         g0886(.A(\b[96] ), .Y(new_n1272));
  NAND2xp33_ASAP7_75t_L     g0887(.A(new_n1272), .B(new_n1271), .Y(new_n1273));
  NOR2xp33_ASAP7_75t_L      g0888(.A(new_n1271), .B(new_n1272), .Y(new_n1274));
  INVx1_ASAP7_75t_L         g0889(.A(new_n1274), .Y(new_n1275));
  AOI21xp33_ASAP7_75t_L     g0890(.A1(new_n1275), .A2(new_n1273), .B(new_n1270), .Y(new_n1276));
  NAND2xp33_ASAP7_75t_L     g0891(.A(new_n1273), .B(new_n1275), .Y(new_n1277));
  A2O1A1O1Ixp25_ASAP7_75t_L g0892(.A1(new_n1258), .A2(new_n1268), .B(new_n1264), .C(new_n1269), .D(new_n1277), .Y(new_n1278));
  NOR2xp33_ASAP7_75t_L      g0893(.A(new_n1278), .B(new_n1276), .Y(\f[96] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0894(.A1(new_n1254), .A2(new_n1255), .B(new_n1268), .C(new_n1264), .Y(new_n1280));
  A2O1A1Ixp33_ASAP7_75t_L   g0895(.A1(\b[95] ), .A2(\a[95] ), .B(new_n1280), .C(new_n1273), .Y(new_n1281));
  INVx1_ASAP7_75t_L         g0896(.A(\a[97] ), .Y(new_n1282));
  INVx1_ASAP7_75t_L         g0897(.A(\b[97] ), .Y(new_n1283));
  NAND2xp33_ASAP7_75t_L     g0898(.A(new_n1283), .B(new_n1282), .Y(new_n1284));
  NOR2xp33_ASAP7_75t_L      g0899(.A(new_n1282), .B(new_n1283), .Y(new_n1285));
  INVx1_ASAP7_75t_L         g0900(.A(new_n1285), .Y(new_n1286));
  NAND2xp33_ASAP7_75t_L     g0901(.A(new_n1284), .B(new_n1286), .Y(new_n1287));
  AND3x1_ASAP7_75t_L        g0902(.A(new_n1281), .B(new_n1287), .C(new_n1275), .Y(new_n1288));
  O2A1O1Ixp33_ASAP7_75t_L   g0903(.A1(new_n1271), .A2(new_n1272), .B(new_n1281), .C(new_n1287), .Y(new_n1289));
  NOR2xp33_ASAP7_75t_L      g0904(.A(new_n1289), .B(new_n1288), .Y(\f[97] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0905(.A1(new_n1273), .A2(new_n1270), .B(new_n1274), .C(new_n1284), .D(new_n1285), .Y(new_n1291));
  NOR2xp33_ASAP7_75t_L      g0906(.A(\a[98] ), .B(\b[98] ), .Y(new_n1292));
  AND2x2_ASAP7_75t_L        g0907(.A(\a[98] ), .B(\b[98] ), .Y(new_n1293));
  NOR2xp33_ASAP7_75t_L      g0908(.A(new_n1292), .B(new_n1293), .Y(new_n1294));
  XNOR2x2_ASAP7_75t_L       g0909(.A(new_n1294), .B(new_n1291), .Y(\f[98] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0910(.A1(new_n1270), .A2(new_n1273), .B(new_n1274), .C(new_n1284), .Y(new_n1296));
  NAND2xp33_ASAP7_75t_L     g0911(.A(\b[98] ), .B(\a[98] ), .Y(new_n1297));
  A2O1A1Ixp33_ASAP7_75t_L   g0912(.A1(new_n1296), .A2(new_n1286), .B(new_n1292), .C(new_n1297), .Y(new_n1298));
  INVx1_ASAP7_75t_L         g0913(.A(\a[99] ), .Y(new_n1299));
  INVx1_ASAP7_75t_L         g0914(.A(\b[99] ), .Y(new_n1300));
  NAND2xp33_ASAP7_75t_L     g0915(.A(new_n1300), .B(new_n1299), .Y(new_n1301));
  NOR2xp33_ASAP7_75t_L      g0916(.A(new_n1299), .B(new_n1300), .Y(new_n1302));
  INVx1_ASAP7_75t_L         g0917(.A(new_n1302), .Y(new_n1303));
  AOI21xp33_ASAP7_75t_L     g0918(.A1(new_n1303), .A2(new_n1301), .B(new_n1298), .Y(new_n1304));
  NAND2xp33_ASAP7_75t_L     g0919(.A(new_n1301), .B(new_n1303), .Y(new_n1305));
  A2O1A1O1Ixp25_ASAP7_75t_L g0920(.A1(new_n1286), .A2(new_n1296), .B(new_n1292), .C(new_n1297), .D(new_n1305), .Y(new_n1306));
  NOR2xp33_ASAP7_75t_L      g0921(.A(new_n1306), .B(new_n1304), .Y(\f[99] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0922(.A1(new_n1282), .A2(new_n1283), .B(new_n1296), .C(new_n1292), .Y(new_n1308));
  A2O1A1Ixp33_ASAP7_75t_L   g0923(.A1(\b[98] ), .A2(\a[98] ), .B(new_n1308), .C(new_n1301), .Y(new_n1309));
  INVx1_ASAP7_75t_L         g0924(.A(\a[100] ), .Y(new_n1310));
  INVx1_ASAP7_75t_L         g0925(.A(\b[100] ), .Y(new_n1311));
  NAND2xp33_ASAP7_75t_L     g0926(.A(new_n1311), .B(new_n1310), .Y(new_n1312));
  NOR2xp33_ASAP7_75t_L      g0927(.A(new_n1310), .B(new_n1311), .Y(new_n1313));
  INVx1_ASAP7_75t_L         g0928(.A(new_n1313), .Y(new_n1314));
  NAND2xp33_ASAP7_75t_L     g0929(.A(new_n1312), .B(new_n1314), .Y(new_n1315));
  AND3x1_ASAP7_75t_L        g0930(.A(new_n1309), .B(new_n1315), .C(new_n1303), .Y(new_n1316));
  O2A1O1Ixp33_ASAP7_75t_L   g0931(.A1(new_n1299), .A2(new_n1300), .B(new_n1309), .C(new_n1315), .Y(new_n1317));
  NOR2xp33_ASAP7_75t_L      g0932(.A(new_n1317), .B(new_n1316), .Y(\f[100] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0933(.A1(new_n1301), .A2(new_n1298), .B(new_n1302), .C(new_n1312), .D(new_n1313), .Y(new_n1319));
  NOR2xp33_ASAP7_75t_L      g0934(.A(\a[101] ), .B(\b[101] ), .Y(new_n1320));
  AND2x2_ASAP7_75t_L        g0935(.A(\a[101] ), .B(\b[101] ), .Y(new_n1321));
  NOR2xp33_ASAP7_75t_L      g0936(.A(new_n1320), .B(new_n1321), .Y(new_n1322));
  XNOR2x2_ASAP7_75t_L       g0937(.A(new_n1322), .B(new_n1319), .Y(\f[101] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0938(.A1(new_n1298), .A2(new_n1301), .B(new_n1302), .C(new_n1312), .Y(new_n1324));
  NAND2xp33_ASAP7_75t_L     g0939(.A(\b[101] ), .B(\a[101] ), .Y(new_n1325));
  A2O1A1Ixp33_ASAP7_75t_L   g0940(.A1(new_n1324), .A2(new_n1314), .B(new_n1320), .C(new_n1325), .Y(new_n1326));
  INVx1_ASAP7_75t_L         g0941(.A(\a[102] ), .Y(new_n1327));
  INVx1_ASAP7_75t_L         g0942(.A(\b[102] ), .Y(new_n1328));
  NAND2xp33_ASAP7_75t_L     g0943(.A(new_n1328), .B(new_n1327), .Y(new_n1329));
  NOR2xp33_ASAP7_75t_L      g0944(.A(new_n1327), .B(new_n1328), .Y(new_n1330));
  INVx1_ASAP7_75t_L         g0945(.A(new_n1330), .Y(new_n1331));
  AOI21xp33_ASAP7_75t_L     g0946(.A1(new_n1331), .A2(new_n1329), .B(new_n1326), .Y(new_n1332));
  NAND2xp33_ASAP7_75t_L     g0947(.A(new_n1329), .B(new_n1331), .Y(new_n1333));
  A2O1A1O1Ixp25_ASAP7_75t_L g0948(.A1(new_n1314), .A2(new_n1324), .B(new_n1320), .C(new_n1325), .D(new_n1333), .Y(new_n1334));
  NOR2xp33_ASAP7_75t_L      g0949(.A(new_n1334), .B(new_n1332), .Y(\f[102] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0950(.A1(new_n1310), .A2(new_n1311), .B(new_n1324), .C(new_n1320), .Y(new_n1336));
  A2O1A1Ixp33_ASAP7_75t_L   g0951(.A1(\b[101] ), .A2(\a[101] ), .B(new_n1336), .C(new_n1329), .Y(new_n1337));
  INVx1_ASAP7_75t_L         g0952(.A(\a[103] ), .Y(new_n1338));
  INVx1_ASAP7_75t_L         g0953(.A(\b[103] ), .Y(new_n1339));
  NAND2xp33_ASAP7_75t_L     g0954(.A(new_n1339), .B(new_n1338), .Y(new_n1340));
  NOR2xp33_ASAP7_75t_L      g0955(.A(new_n1338), .B(new_n1339), .Y(new_n1341));
  INVx1_ASAP7_75t_L         g0956(.A(new_n1341), .Y(new_n1342));
  NAND2xp33_ASAP7_75t_L     g0957(.A(new_n1340), .B(new_n1342), .Y(new_n1343));
  AND3x1_ASAP7_75t_L        g0958(.A(new_n1337), .B(new_n1343), .C(new_n1331), .Y(new_n1344));
  O2A1O1Ixp33_ASAP7_75t_L   g0959(.A1(new_n1327), .A2(new_n1328), .B(new_n1337), .C(new_n1343), .Y(new_n1345));
  NOR2xp33_ASAP7_75t_L      g0960(.A(new_n1345), .B(new_n1344), .Y(\f[103] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0961(.A1(new_n1329), .A2(new_n1326), .B(new_n1330), .C(new_n1340), .D(new_n1341), .Y(new_n1347));
  NOR2xp33_ASAP7_75t_L      g0962(.A(\a[104] ), .B(\b[104] ), .Y(new_n1348));
  AND2x2_ASAP7_75t_L        g0963(.A(\a[104] ), .B(\b[104] ), .Y(new_n1349));
  NOR2xp33_ASAP7_75t_L      g0964(.A(new_n1348), .B(new_n1349), .Y(new_n1350));
  XNOR2x2_ASAP7_75t_L       g0965(.A(new_n1350), .B(new_n1347), .Y(\f[104] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0966(.A1(new_n1326), .A2(new_n1329), .B(new_n1330), .C(new_n1340), .Y(new_n1352));
  NAND2xp33_ASAP7_75t_L     g0967(.A(\b[104] ), .B(\a[104] ), .Y(new_n1353));
  A2O1A1Ixp33_ASAP7_75t_L   g0968(.A1(new_n1352), .A2(new_n1342), .B(new_n1348), .C(new_n1353), .Y(new_n1354));
  INVx1_ASAP7_75t_L         g0969(.A(\a[105] ), .Y(new_n1355));
  INVx1_ASAP7_75t_L         g0970(.A(\b[105] ), .Y(new_n1356));
  NAND2xp33_ASAP7_75t_L     g0971(.A(new_n1356), .B(new_n1355), .Y(new_n1357));
  NOR2xp33_ASAP7_75t_L      g0972(.A(new_n1355), .B(new_n1356), .Y(new_n1358));
  INVx1_ASAP7_75t_L         g0973(.A(new_n1358), .Y(new_n1359));
  AOI21xp33_ASAP7_75t_L     g0974(.A1(new_n1359), .A2(new_n1357), .B(new_n1354), .Y(new_n1360));
  NAND2xp33_ASAP7_75t_L     g0975(.A(new_n1357), .B(new_n1359), .Y(new_n1361));
  A2O1A1O1Ixp25_ASAP7_75t_L g0976(.A1(new_n1342), .A2(new_n1352), .B(new_n1348), .C(new_n1353), .D(new_n1361), .Y(new_n1362));
  NOR2xp33_ASAP7_75t_L      g0977(.A(new_n1362), .B(new_n1360), .Y(\f[105] ));
  O2A1O1Ixp33_ASAP7_75t_L   g0978(.A1(new_n1338), .A2(new_n1339), .B(new_n1352), .C(new_n1348), .Y(new_n1364));
  A2O1A1Ixp33_ASAP7_75t_L   g0979(.A1(\b[104] ), .A2(\a[104] ), .B(new_n1364), .C(new_n1357), .Y(new_n1365));
  INVx1_ASAP7_75t_L         g0980(.A(\a[106] ), .Y(new_n1366));
  INVx1_ASAP7_75t_L         g0981(.A(\b[106] ), .Y(new_n1367));
  NAND2xp33_ASAP7_75t_L     g0982(.A(new_n1367), .B(new_n1366), .Y(new_n1368));
  NOR2xp33_ASAP7_75t_L      g0983(.A(new_n1366), .B(new_n1367), .Y(new_n1369));
  INVx1_ASAP7_75t_L         g0984(.A(new_n1369), .Y(new_n1370));
  NAND2xp33_ASAP7_75t_L     g0985(.A(new_n1368), .B(new_n1370), .Y(new_n1371));
  AND3x1_ASAP7_75t_L        g0986(.A(new_n1365), .B(new_n1371), .C(new_n1359), .Y(new_n1372));
  O2A1O1Ixp33_ASAP7_75t_L   g0987(.A1(new_n1355), .A2(new_n1356), .B(new_n1365), .C(new_n1371), .Y(new_n1373));
  NOR2xp33_ASAP7_75t_L      g0988(.A(new_n1373), .B(new_n1372), .Y(\f[106] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g0989(.A1(new_n1357), .A2(new_n1354), .B(new_n1358), .C(new_n1368), .D(new_n1369), .Y(new_n1375));
  NOR2xp33_ASAP7_75t_L      g0990(.A(\a[107] ), .B(\b[107] ), .Y(new_n1376));
  AND2x2_ASAP7_75t_L        g0991(.A(\a[107] ), .B(\b[107] ), .Y(new_n1377));
  NOR2xp33_ASAP7_75t_L      g0992(.A(new_n1376), .B(new_n1377), .Y(new_n1378));
  XNOR2x2_ASAP7_75t_L       g0993(.A(new_n1378), .B(new_n1375), .Y(\f[107] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0994(.A1(new_n1354), .A2(new_n1357), .B(new_n1358), .C(new_n1368), .Y(new_n1380));
  NAND2xp33_ASAP7_75t_L     g0995(.A(\b[107] ), .B(\a[107] ), .Y(new_n1381));
  A2O1A1Ixp33_ASAP7_75t_L   g0996(.A1(new_n1380), .A2(new_n1370), .B(new_n1376), .C(new_n1381), .Y(new_n1382));
  INVx1_ASAP7_75t_L         g0997(.A(\a[108] ), .Y(new_n1383));
  INVx1_ASAP7_75t_L         g0998(.A(\b[108] ), .Y(new_n1384));
  NAND2xp33_ASAP7_75t_L     g0999(.A(new_n1384), .B(new_n1383), .Y(new_n1385));
  NOR2xp33_ASAP7_75t_L      g1000(.A(new_n1383), .B(new_n1384), .Y(new_n1386));
  INVx1_ASAP7_75t_L         g1001(.A(new_n1386), .Y(new_n1387));
  AOI21xp33_ASAP7_75t_L     g1002(.A1(new_n1387), .A2(new_n1385), .B(new_n1382), .Y(new_n1388));
  NAND2xp33_ASAP7_75t_L     g1003(.A(new_n1385), .B(new_n1387), .Y(new_n1389));
  A2O1A1O1Ixp25_ASAP7_75t_L g1004(.A1(new_n1370), .A2(new_n1380), .B(new_n1376), .C(new_n1381), .D(new_n1389), .Y(new_n1390));
  NOR2xp33_ASAP7_75t_L      g1005(.A(new_n1390), .B(new_n1388), .Y(\f[108] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1006(.A1(new_n1366), .A2(new_n1367), .B(new_n1380), .C(new_n1376), .Y(new_n1392));
  A2O1A1Ixp33_ASAP7_75t_L   g1007(.A1(\b[107] ), .A2(\a[107] ), .B(new_n1392), .C(new_n1385), .Y(new_n1393));
  INVx1_ASAP7_75t_L         g1008(.A(\a[109] ), .Y(new_n1394));
  INVx1_ASAP7_75t_L         g1009(.A(\b[109] ), .Y(new_n1395));
  NAND2xp33_ASAP7_75t_L     g1010(.A(new_n1395), .B(new_n1394), .Y(new_n1396));
  NOR2xp33_ASAP7_75t_L      g1011(.A(new_n1394), .B(new_n1395), .Y(new_n1397));
  INVx1_ASAP7_75t_L         g1012(.A(new_n1397), .Y(new_n1398));
  NAND2xp33_ASAP7_75t_L     g1013(.A(new_n1396), .B(new_n1398), .Y(new_n1399));
  AND3x1_ASAP7_75t_L        g1014(.A(new_n1393), .B(new_n1399), .C(new_n1387), .Y(new_n1400));
  O2A1O1Ixp33_ASAP7_75t_L   g1015(.A1(new_n1383), .A2(new_n1384), .B(new_n1393), .C(new_n1399), .Y(new_n1401));
  NOR2xp33_ASAP7_75t_L      g1016(.A(new_n1401), .B(new_n1400), .Y(\f[109] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1017(.A1(new_n1385), .A2(new_n1382), .B(new_n1386), .C(new_n1396), .D(new_n1397), .Y(new_n1403));
  NOR2xp33_ASAP7_75t_L      g1018(.A(\a[110] ), .B(\b[110] ), .Y(new_n1404));
  AND2x2_ASAP7_75t_L        g1019(.A(\a[110] ), .B(\b[110] ), .Y(new_n1405));
  NOR2xp33_ASAP7_75t_L      g1020(.A(new_n1404), .B(new_n1405), .Y(new_n1406));
  XNOR2x2_ASAP7_75t_L       g1021(.A(new_n1406), .B(new_n1403), .Y(\f[110] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1022(.A1(new_n1382), .A2(new_n1385), .B(new_n1386), .C(new_n1396), .Y(new_n1408));
  NAND2xp33_ASAP7_75t_L     g1023(.A(\b[110] ), .B(\a[110] ), .Y(new_n1409));
  A2O1A1Ixp33_ASAP7_75t_L   g1024(.A1(new_n1408), .A2(new_n1398), .B(new_n1404), .C(new_n1409), .Y(new_n1410));
  INVx1_ASAP7_75t_L         g1025(.A(\a[111] ), .Y(new_n1411));
  INVx1_ASAP7_75t_L         g1026(.A(\b[111] ), .Y(new_n1412));
  NAND2xp33_ASAP7_75t_L     g1027(.A(new_n1412), .B(new_n1411), .Y(new_n1413));
  NOR2xp33_ASAP7_75t_L      g1028(.A(new_n1411), .B(new_n1412), .Y(new_n1414));
  INVx1_ASAP7_75t_L         g1029(.A(new_n1414), .Y(new_n1415));
  AOI21xp33_ASAP7_75t_L     g1030(.A1(new_n1415), .A2(new_n1413), .B(new_n1410), .Y(new_n1416));
  NAND2xp33_ASAP7_75t_L     g1031(.A(new_n1413), .B(new_n1415), .Y(new_n1417));
  A2O1A1O1Ixp25_ASAP7_75t_L g1032(.A1(new_n1398), .A2(new_n1408), .B(new_n1404), .C(new_n1409), .D(new_n1417), .Y(new_n1418));
  NOR2xp33_ASAP7_75t_L      g1033(.A(new_n1418), .B(new_n1416), .Y(\f[111] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1034(.A1(new_n1394), .A2(new_n1395), .B(new_n1408), .C(new_n1404), .Y(new_n1420));
  A2O1A1Ixp33_ASAP7_75t_L   g1035(.A1(\b[110] ), .A2(\a[110] ), .B(new_n1420), .C(new_n1413), .Y(new_n1421));
  INVx1_ASAP7_75t_L         g1036(.A(\a[112] ), .Y(new_n1422));
  INVx1_ASAP7_75t_L         g1037(.A(\b[112] ), .Y(new_n1423));
  NAND2xp33_ASAP7_75t_L     g1038(.A(new_n1423), .B(new_n1422), .Y(new_n1424));
  NOR2xp33_ASAP7_75t_L      g1039(.A(new_n1422), .B(new_n1423), .Y(new_n1425));
  INVx1_ASAP7_75t_L         g1040(.A(new_n1425), .Y(new_n1426));
  NAND2xp33_ASAP7_75t_L     g1041(.A(new_n1424), .B(new_n1426), .Y(new_n1427));
  AND3x1_ASAP7_75t_L        g1042(.A(new_n1421), .B(new_n1427), .C(new_n1415), .Y(new_n1428));
  O2A1O1Ixp33_ASAP7_75t_L   g1043(.A1(new_n1411), .A2(new_n1412), .B(new_n1421), .C(new_n1427), .Y(new_n1429));
  NOR2xp33_ASAP7_75t_L      g1044(.A(new_n1429), .B(new_n1428), .Y(\f[112] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1045(.A1(new_n1413), .A2(new_n1410), .B(new_n1414), .C(new_n1424), .D(new_n1425), .Y(new_n1431));
  NOR2xp33_ASAP7_75t_L      g1046(.A(\a[113] ), .B(\b[113] ), .Y(new_n1432));
  AND2x2_ASAP7_75t_L        g1047(.A(\a[113] ), .B(\b[113] ), .Y(new_n1433));
  NOR2xp33_ASAP7_75t_L      g1048(.A(new_n1432), .B(new_n1433), .Y(new_n1434));
  XNOR2x2_ASAP7_75t_L       g1049(.A(new_n1434), .B(new_n1431), .Y(\f[113] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1050(.A1(new_n1410), .A2(new_n1413), .B(new_n1414), .C(new_n1424), .Y(new_n1436));
  NAND2xp33_ASAP7_75t_L     g1051(.A(\b[113] ), .B(\a[113] ), .Y(new_n1437));
  A2O1A1Ixp33_ASAP7_75t_L   g1052(.A1(new_n1436), .A2(new_n1426), .B(new_n1432), .C(new_n1437), .Y(new_n1438));
  INVx1_ASAP7_75t_L         g1053(.A(\a[114] ), .Y(new_n1439));
  INVx1_ASAP7_75t_L         g1054(.A(\b[114] ), .Y(new_n1440));
  NAND2xp33_ASAP7_75t_L     g1055(.A(new_n1440), .B(new_n1439), .Y(new_n1441));
  NOR2xp33_ASAP7_75t_L      g1056(.A(new_n1439), .B(new_n1440), .Y(new_n1442));
  INVx1_ASAP7_75t_L         g1057(.A(new_n1442), .Y(new_n1443));
  AOI21xp33_ASAP7_75t_L     g1058(.A1(new_n1443), .A2(new_n1441), .B(new_n1438), .Y(new_n1444));
  NAND2xp33_ASAP7_75t_L     g1059(.A(new_n1441), .B(new_n1443), .Y(new_n1445));
  A2O1A1O1Ixp25_ASAP7_75t_L g1060(.A1(new_n1426), .A2(new_n1436), .B(new_n1432), .C(new_n1437), .D(new_n1445), .Y(new_n1446));
  NOR2xp33_ASAP7_75t_L      g1061(.A(new_n1446), .B(new_n1444), .Y(\f[114] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1062(.A1(new_n1422), .A2(new_n1423), .B(new_n1436), .C(new_n1432), .Y(new_n1448));
  A2O1A1Ixp33_ASAP7_75t_L   g1063(.A1(\b[113] ), .A2(\a[113] ), .B(new_n1448), .C(new_n1441), .Y(new_n1449));
  INVx1_ASAP7_75t_L         g1064(.A(\a[115] ), .Y(new_n1450));
  INVx1_ASAP7_75t_L         g1065(.A(\b[115] ), .Y(new_n1451));
  NAND2xp33_ASAP7_75t_L     g1066(.A(new_n1451), .B(new_n1450), .Y(new_n1452));
  NOR2xp33_ASAP7_75t_L      g1067(.A(new_n1450), .B(new_n1451), .Y(new_n1453));
  INVx1_ASAP7_75t_L         g1068(.A(new_n1453), .Y(new_n1454));
  NAND2xp33_ASAP7_75t_L     g1069(.A(new_n1452), .B(new_n1454), .Y(new_n1455));
  AND3x1_ASAP7_75t_L        g1070(.A(new_n1449), .B(new_n1455), .C(new_n1443), .Y(new_n1456));
  O2A1O1Ixp33_ASAP7_75t_L   g1071(.A1(new_n1439), .A2(new_n1440), .B(new_n1449), .C(new_n1455), .Y(new_n1457));
  NOR2xp33_ASAP7_75t_L      g1072(.A(new_n1457), .B(new_n1456), .Y(\f[115] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1073(.A1(new_n1441), .A2(new_n1438), .B(new_n1442), .C(new_n1452), .D(new_n1453), .Y(new_n1459));
  NOR2xp33_ASAP7_75t_L      g1074(.A(\a[116] ), .B(\b[116] ), .Y(new_n1460));
  AND2x2_ASAP7_75t_L        g1075(.A(\a[116] ), .B(\b[116] ), .Y(new_n1461));
  NOR2xp33_ASAP7_75t_L      g1076(.A(new_n1460), .B(new_n1461), .Y(new_n1462));
  XNOR2x2_ASAP7_75t_L       g1077(.A(new_n1462), .B(new_n1459), .Y(\f[116] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1078(.A1(new_n1438), .A2(new_n1441), .B(new_n1442), .C(new_n1452), .Y(new_n1464));
  NAND2xp33_ASAP7_75t_L     g1079(.A(\b[116] ), .B(\a[116] ), .Y(new_n1465));
  A2O1A1Ixp33_ASAP7_75t_L   g1080(.A1(new_n1464), .A2(new_n1454), .B(new_n1460), .C(new_n1465), .Y(new_n1466));
  INVx1_ASAP7_75t_L         g1081(.A(\a[117] ), .Y(new_n1467));
  INVx1_ASAP7_75t_L         g1082(.A(\b[117] ), .Y(new_n1468));
  NAND2xp33_ASAP7_75t_L     g1083(.A(new_n1468), .B(new_n1467), .Y(new_n1469));
  NOR2xp33_ASAP7_75t_L      g1084(.A(new_n1467), .B(new_n1468), .Y(new_n1470));
  INVx1_ASAP7_75t_L         g1085(.A(new_n1470), .Y(new_n1471));
  AOI21xp33_ASAP7_75t_L     g1086(.A1(new_n1471), .A2(new_n1469), .B(new_n1466), .Y(new_n1472));
  NAND2xp33_ASAP7_75t_L     g1087(.A(new_n1469), .B(new_n1471), .Y(new_n1473));
  A2O1A1O1Ixp25_ASAP7_75t_L g1088(.A1(new_n1454), .A2(new_n1464), .B(new_n1460), .C(new_n1465), .D(new_n1473), .Y(new_n1474));
  NOR2xp33_ASAP7_75t_L      g1089(.A(new_n1474), .B(new_n1472), .Y(\f[117] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1090(.A1(new_n1450), .A2(new_n1451), .B(new_n1464), .C(new_n1460), .Y(new_n1476));
  A2O1A1Ixp33_ASAP7_75t_L   g1091(.A1(\b[116] ), .A2(\a[116] ), .B(new_n1476), .C(new_n1469), .Y(new_n1477));
  INVx1_ASAP7_75t_L         g1092(.A(\a[118] ), .Y(new_n1478));
  INVx1_ASAP7_75t_L         g1093(.A(\b[118] ), .Y(new_n1479));
  NAND2xp33_ASAP7_75t_L     g1094(.A(new_n1479), .B(new_n1478), .Y(new_n1480));
  NOR2xp33_ASAP7_75t_L      g1095(.A(new_n1478), .B(new_n1479), .Y(new_n1481));
  INVx1_ASAP7_75t_L         g1096(.A(new_n1481), .Y(new_n1482));
  NAND2xp33_ASAP7_75t_L     g1097(.A(new_n1480), .B(new_n1482), .Y(new_n1483));
  AND3x1_ASAP7_75t_L        g1098(.A(new_n1477), .B(new_n1483), .C(new_n1471), .Y(new_n1484));
  O2A1O1Ixp33_ASAP7_75t_L   g1099(.A1(new_n1467), .A2(new_n1468), .B(new_n1477), .C(new_n1483), .Y(new_n1485));
  NOR2xp33_ASAP7_75t_L      g1100(.A(new_n1485), .B(new_n1484), .Y(\f[118] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1101(.A1(new_n1469), .A2(new_n1466), .B(new_n1470), .C(new_n1480), .D(new_n1481), .Y(new_n1487));
  NOR2xp33_ASAP7_75t_L      g1102(.A(\a[119] ), .B(\b[119] ), .Y(new_n1488));
  AND2x2_ASAP7_75t_L        g1103(.A(\a[119] ), .B(\b[119] ), .Y(new_n1489));
  NOR2xp33_ASAP7_75t_L      g1104(.A(new_n1488), .B(new_n1489), .Y(new_n1490));
  XNOR2x2_ASAP7_75t_L       g1105(.A(new_n1490), .B(new_n1487), .Y(\f[119] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1106(.A1(new_n1466), .A2(new_n1469), .B(new_n1470), .C(new_n1480), .Y(new_n1492));
  NAND2xp33_ASAP7_75t_L     g1107(.A(\b[119] ), .B(\a[119] ), .Y(new_n1493));
  A2O1A1Ixp33_ASAP7_75t_L   g1108(.A1(new_n1492), .A2(new_n1482), .B(new_n1488), .C(new_n1493), .Y(new_n1494));
  INVx1_ASAP7_75t_L         g1109(.A(\a[120] ), .Y(new_n1495));
  INVx1_ASAP7_75t_L         g1110(.A(\b[120] ), .Y(new_n1496));
  NAND2xp33_ASAP7_75t_L     g1111(.A(new_n1496), .B(new_n1495), .Y(new_n1497));
  NOR2xp33_ASAP7_75t_L      g1112(.A(new_n1495), .B(new_n1496), .Y(new_n1498));
  INVx1_ASAP7_75t_L         g1113(.A(new_n1498), .Y(new_n1499));
  AOI21xp33_ASAP7_75t_L     g1114(.A1(new_n1499), .A2(new_n1497), .B(new_n1494), .Y(new_n1500));
  NAND2xp33_ASAP7_75t_L     g1115(.A(new_n1497), .B(new_n1499), .Y(new_n1501));
  A2O1A1O1Ixp25_ASAP7_75t_L g1116(.A1(new_n1482), .A2(new_n1492), .B(new_n1488), .C(new_n1493), .D(new_n1501), .Y(new_n1502));
  NOR2xp33_ASAP7_75t_L      g1117(.A(new_n1502), .B(new_n1500), .Y(\f[120] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1118(.A1(new_n1478), .A2(new_n1479), .B(new_n1492), .C(new_n1488), .Y(new_n1504));
  A2O1A1Ixp33_ASAP7_75t_L   g1119(.A1(\b[119] ), .A2(\a[119] ), .B(new_n1504), .C(new_n1497), .Y(new_n1505));
  INVx1_ASAP7_75t_L         g1120(.A(\a[121] ), .Y(new_n1506));
  INVx1_ASAP7_75t_L         g1121(.A(\b[121] ), .Y(new_n1507));
  NAND2xp33_ASAP7_75t_L     g1122(.A(new_n1507), .B(new_n1506), .Y(new_n1508));
  NOR2xp33_ASAP7_75t_L      g1123(.A(new_n1506), .B(new_n1507), .Y(new_n1509));
  INVx1_ASAP7_75t_L         g1124(.A(new_n1509), .Y(new_n1510));
  NAND2xp33_ASAP7_75t_L     g1125(.A(new_n1508), .B(new_n1510), .Y(new_n1511));
  AND3x1_ASAP7_75t_L        g1126(.A(new_n1505), .B(new_n1511), .C(new_n1499), .Y(new_n1512));
  O2A1O1Ixp33_ASAP7_75t_L   g1127(.A1(new_n1495), .A2(new_n1496), .B(new_n1505), .C(new_n1511), .Y(new_n1513));
  NOR2xp33_ASAP7_75t_L      g1128(.A(new_n1513), .B(new_n1512), .Y(\f[121] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1129(.A1(new_n1497), .A2(new_n1494), .B(new_n1498), .C(new_n1508), .D(new_n1509), .Y(new_n1515));
  NOR2xp33_ASAP7_75t_L      g1130(.A(\a[122] ), .B(\b[122] ), .Y(new_n1516));
  AND2x2_ASAP7_75t_L        g1131(.A(\a[122] ), .B(\b[122] ), .Y(new_n1517));
  NOR2xp33_ASAP7_75t_L      g1132(.A(new_n1516), .B(new_n1517), .Y(new_n1518));
  XNOR2x2_ASAP7_75t_L       g1133(.A(new_n1518), .B(new_n1515), .Y(\f[122] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1134(.A1(new_n1494), .A2(new_n1497), .B(new_n1498), .C(new_n1508), .Y(new_n1520));
  NAND2xp33_ASAP7_75t_L     g1135(.A(\b[122] ), .B(\a[122] ), .Y(new_n1521));
  A2O1A1Ixp33_ASAP7_75t_L   g1136(.A1(new_n1520), .A2(new_n1510), .B(new_n1516), .C(new_n1521), .Y(new_n1522));
  INVx1_ASAP7_75t_L         g1137(.A(\a[123] ), .Y(new_n1523));
  INVx1_ASAP7_75t_L         g1138(.A(\b[123] ), .Y(new_n1524));
  NAND2xp33_ASAP7_75t_L     g1139(.A(new_n1524), .B(new_n1523), .Y(new_n1525));
  NOR2xp33_ASAP7_75t_L      g1140(.A(new_n1523), .B(new_n1524), .Y(new_n1526));
  INVx1_ASAP7_75t_L         g1141(.A(new_n1526), .Y(new_n1527));
  AOI21xp33_ASAP7_75t_L     g1142(.A1(new_n1527), .A2(new_n1525), .B(new_n1522), .Y(new_n1528));
  NAND2xp33_ASAP7_75t_L     g1143(.A(new_n1525), .B(new_n1527), .Y(new_n1529));
  A2O1A1O1Ixp25_ASAP7_75t_L g1144(.A1(new_n1510), .A2(new_n1520), .B(new_n1516), .C(new_n1521), .D(new_n1529), .Y(new_n1530));
  NOR2xp33_ASAP7_75t_L      g1145(.A(new_n1530), .B(new_n1528), .Y(\f[123] ));
  O2A1O1Ixp33_ASAP7_75t_L   g1146(.A1(new_n1506), .A2(new_n1507), .B(new_n1520), .C(new_n1516), .Y(new_n1532));
  A2O1A1Ixp33_ASAP7_75t_L   g1147(.A1(\b[122] ), .A2(\a[122] ), .B(new_n1532), .C(new_n1525), .Y(new_n1533));
  INVx1_ASAP7_75t_L         g1148(.A(\a[124] ), .Y(new_n1534));
  INVx1_ASAP7_75t_L         g1149(.A(\b[124] ), .Y(new_n1535));
  NAND2xp33_ASAP7_75t_L     g1150(.A(new_n1535), .B(new_n1534), .Y(new_n1536));
  NOR2xp33_ASAP7_75t_L      g1151(.A(new_n1534), .B(new_n1535), .Y(new_n1537));
  INVx1_ASAP7_75t_L         g1152(.A(new_n1537), .Y(new_n1538));
  NAND2xp33_ASAP7_75t_L     g1153(.A(new_n1536), .B(new_n1538), .Y(new_n1539));
  AND3x1_ASAP7_75t_L        g1154(.A(new_n1533), .B(new_n1539), .C(new_n1527), .Y(new_n1540));
  O2A1O1Ixp33_ASAP7_75t_L   g1155(.A1(new_n1523), .A2(new_n1524), .B(new_n1533), .C(new_n1539), .Y(new_n1541));
  NOR2xp33_ASAP7_75t_L      g1156(.A(new_n1541), .B(new_n1540), .Y(\f[124] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g1157(.A1(new_n1525), .A2(new_n1522), .B(new_n1526), .C(new_n1536), .D(new_n1537), .Y(new_n1543));
  NOR2xp33_ASAP7_75t_L      g1158(.A(\a[125] ), .B(\b[125] ), .Y(new_n1544));
  AND2x2_ASAP7_75t_L        g1159(.A(\a[125] ), .B(\b[125] ), .Y(new_n1545));
  NOR2xp33_ASAP7_75t_L      g1160(.A(new_n1544), .B(new_n1545), .Y(new_n1546));
  XNOR2x2_ASAP7_75t_L       g1161(.A(new_n1546), .B(new_n1543), .Y(\f[125] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1162(.A1(new_n1522), .A2(new_n1525), .B(new_n1526), .C(new_n1536), .Y(new_n1548));
  NAND2xp33_ASAP7_75t_L     g1163(.A(\b[125] ), .B(\a[125] ), .Y(new_n1549));
  A2O1A1Ixp33_ASAP7_75t_L   g1164(.A1(new_n1548), .A2(new_n1538), .B(new_n1544), .C(new_n1549), .Y(new_n1550));
  XNOR2x2_ASAP7_75t_L       g1165(.A(\b[126] ), .B(\a[126] ), .Y(new_n1551));
  XNOR2x2_ASAP7_75t_L       g1166(.A(new_n1551), .B(new_n1550), .Y(\f[126] ));
  MAJIxp5_ASAP7_75t_L       g1167(.A(new_n1550), .B(\a[126] ), .C(\b[126] ), .Y(new_n1553));
  NOR2xp33_ASAP7_75t_L      g1168(.A(\a[127] ), .B(\b[127] ), .Y(new_n1554));
  AND2x2_ASAP7_75t_L        g1169(.A(\a[127] ), .B(\b[127] ), .Y(new_n1555));
  NOR2xp33_ASAP7_75t_L      g1170(.A(new_n1554), .B(new_n1555), .Y(new_n1556));
  XNOR2x2_ASAP7_75t_L       g1171(.A(new_n1556), .B(new_n1553), .Y(\f[127] ));
  NAND2xp33_ASAP7_75t_L     g1172(.A(\b[127] ), .B(\a[127] ), .Y(new_n1558));
  OAI21xp33_ASAP7_75t_L     g1173(.A1(new_n1554), .A2(new_n1553), .B(new_n1558), .Y(cOut));
endmodule


