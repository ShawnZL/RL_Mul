// Benchmark "top" written by ABC on Mon Dec 25 16:29:26 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386, new_n387, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1378,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1404;
  assign new_n386 = \a[0]  & ~\b[0] ;
  assign new_n387 = ~\a[0]  & \b[0] ;
  assign \f[0]  = new_n386 | new_n387;
  assign new_n389 = \a[0]  & \b[0] ;
  assign new_n390 = ~\a[1]  & ~\b[1] ;
  assign new_n391 = \a[1]  & \b[1] ;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = new_n389 & ~new_n392;
  assign new_n394 = ~new_n389 & new_n392;
  assign \f[1]  = new_n393 | new_n394;
  assign new_n396 = new_n389 & ~new_n390;
  assign new_n397 = ~new_n391 & ~new_n396;
  assign new_n398 = ~\a[2]  & ~\b[2] ;
  assign new_n399 = \a[2]  & \b[2] ;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = new_n397 & ~new_n400;
  assign new_n402 = ~new_n397 & new_n400;
  assign \f[2]  = ~new_n401 & ~new_n402;
  assign new_n404 = ~new_n397 & ~new_n398;
  assign new_n405 = ~new_n399 & ~new_n404;
  assign new_n406 = ~\a[3]  & ~\b[3] ;
  assign new_n407 = \a[3]  & \b[3] ;
  assign new_n408 = ~new_n406 & ~new_n407;
  assign new_n409 = new_n405 & ~new_n408;
  assign new_n410 = ~new_n405 & new_n408;
  assign \f[3]  = ~new_n409 & ~new_n410;
  assign new_n412 = ~new_n405 & ~new_n406;
  assign new_n413 = ~new_n407 & ~new_n412;
  assign new_n414 = ~\a[4]  & ~\b[4] ;
  assign new_n415 = \a[4]  & \b[4] ;
  assign new_n416 = ~new_n414 & ~new_n415;
  assign new_n417 = new_n413 & ~new_n416;
  assign new_n418 = ~new_n413 & new_n416;
  assign \f[4]  = ~new_n417 & ~new_n418;
  assign new_n420 = ~new_n413 & ~new_n414;
  assign new_n421 = ~new_n415 & ~new_n420;
  assign new_n422 = ~\a[5]  & ~\b[5] ;
  assign new_n423 = \a[5]  & \b[5] ;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = new_n421 & ~new_n424;
  assign new_n426 = ~new_n421 & new_n424;
  assign \f[5]  = ~new_n425 & ~new_n426;
  assign new_n428 = ~new_n421 & ~new_n422;
  assign new_n429 = ~new_n423 & ~new_n428;
  assign new_n430 = ~\a[6]  & ~\b[6] ;
  assign new_n431 = \a[6]  & \b[6] ;
  assign new_n432 = ~new_n430 & ~new_n431;
  assign new_n433 = new_n429 & ~new_n432;
  assign new_n434 = ~new_n429 & new_n432;
  assign \f[6]  = ~new_n433 & ~new_n434;
  assign new_n436 = ~new_n429 & ~new_n430;
  assign new_n437 = ~new_n431 & ~new_n436;
  assign new_n438 = ~\a[7]  & ~\b[7] ;
  assign new_n439 = \a[7]  & \b[7] ;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = new_n437 & ~new_n440;
  assign new_n442 = ~new_n437 & new_n440;
  assign \f[7]  = ~new_n441 & ~new_n442;
  assign new_n444 = ~new_n437 & ~new_n438;
  assign new_n445 = ~new_n439 & ~new_n444;
  assign new_n446 = ~\a[8]  & ~\b[8] ;
  assign new_n447 = \a[8]  & \b[8] ;
  assign new_n448 = ~new_n446 & ~new_n447;
  assign new_n449 = new_n445 & ~new_n448;
  assign new_n450 = ~new_n445 & new_n448;
  assign \f[8]  = ~new_n449 & ~new_n450;
  assign new_n452 = ~new_n445 & ~new_n446;
  assign new_n453 = ~new_n447 & ~new_n452;
  assign new_n454 = ~\a[9]  & ~\b[9] ;
  assign new_n455 = \a[9]  & \b[9] ;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457 = new_n453 & ~new_n456;
  assign new_n458 = ~new_n453 & new_n456;
  assign \f[9]  = ~new_n457 & ~new_n458;
  assign new_n460 = ~new_n453 & ~new_n454;
  assign new_n461 = ~new_n455 & ~new_n460;
  assign new_n462 = ~\a[10]  & ~\b[10] ;
  assign new_n463 = \a[10]  & \b[10] ;
  assign new_n464 = ~new_n462 & ~new_n463;
  assign new_n465 = new_n461 & ~new_n464;
  assign new_n466 = ~new_n461 & new_n464;
  assign \f[10]  = ~new_n465 & ~new_n466;
  assign new_n468 = ~new_n461 & ~new_n462;
  assign new_n469 = ~new_n463 & ~new_n468;
  assign new_n470 = ~\a[11]  & ~\b[11] ;
  assign new_n471 = \a[11]  & \b[11] ;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = new_n469 & ~new_n472;
  assign new_n474 = ~new_n469 & new_n472;
  assign \f[11]  = ~new_n473 & ~new_n474;
  assign new_n476 = ~new_n469 & ~new_n470;
  assign new_n477 = ~new_n471 & ~new_n476;
  assign new_n478 = ~\a[12]  & ~\b[12] ;
  assign new_n479 = \a[12]  & \b[12] ;
  assign new_n480 = ~new_n478 & ~new_n479;
  assign new_n481 = new_n477 & ~new_n480;
  assign new_n482 = ~new_n477 & new_n480;
  assign \f[12]  = ~new_n481 & ~new_n482;
  assign new_n484 = ~new_n477 & ~new_n478;
  assign new_n485 = ~new_n479 & ~new_n484;
  assign new_n486 = ~\a[13]  & ~\b[13] ;
  assign new_n487 = \a[13]  & \b[13] ;
  assign new_n488 = ~new_n486 & ~new_n487;
  assign new_n489 = new_n485 & ~new_n488;
  assign new_n490 = ~new_n485 & new_n488;
  assign \f[13]  = ~new_n489 & ~new_n490;
  assign new_n492 = ~new_n485 & ~new_n486;
  assign new_n493 = ~new_n487 & ~new_n492;
  assign new_n494 = ~\a[14]  & ~\b[14] ;
  assign new_n495 = \a[14]  & \b[14] ;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = new_n493 & ~new_n496;
  assign new_n498 = ~new_n493 & new_n496;
  assign \f[14]  = ~new_n497 & ~new_n498;
  assign new_n500 = ~new_n493 & ~new_n494;
  assign new_n501 = ~new_n495 & ~new_n500;
  assign new_n502 = ~\a[15]  & ~\b[15] ;
  assign new_n503 = \a[15]  & \b[15] ;
  assign new_n504 = ~new_n502 & ~new_n503;
  assign new_n505 = new_n501 & ~new_n504;
  assign new_n506 = ~new_n501 & new_n504;
  assign \f[15]  = ~new_n505 & ~new_n506;
  assign new_n508 = ~new_n501 & ~new_n502;
  assign new_n509 = ~new_n503 & ~new_n508;
  assign new_n510 = ~\a[16]  & ~\b[16] ;
  assign new_n511 = \a[16]  & \b[16] ;
  assign new_n512 = ~new_n510 & ~new_n511;
  assign new_n513 = new_n509 & ~new_n512;
  assign new_n514 = ~new_n509 & new_n512;
  assign \f[16]  = ~new_n513 & ~new_n514;
  assign new_n516 = ~new_n509 & ~new_n510;
  assign new_n517 = ~new_n511 & ~new_n516;
  assign new_n518 = ~\a[17]  & ~\b[17] ;
  assign new_n519 = \a[17]  & \b[17] ;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = new_n517 & ~new_n520;
  assign new_n522 = ~new_n517 & new_n520;
  assign \f[17]  = ~new_n521 & ~new_n522;
  assign new_n524 = ~new_n517 & ~new_n518;
  assign new_n525 = ~new_n519 & ~new_n524;
  assign new_n526 = ~\a[18]  & ~\b[18] ;
  assign new_n527 = \a[18]  & \b[18] ;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign new_n529 = new_n525 & ~new_n528;
  assign new_n530 = ~new_n525 & new_n528;
  assign \f[18]  = ~new_n529 & ~new_n530;
  assign new_n532 = ~new_n525 & ~new_n526;
  assign new_n533 = ~new_n527 & ~new_n532;
  assign new_n534 = ~\a[19]  & ~\b[19] ;
  assign new_n535 = \a[19]  & \b[19] ;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537 = new_n533 & ~new_n536;
  assign new_n538 = ~new_n533 & new_n536;
  assign \f[19]  = ~new_n537 & ~new_n538;
  assign new_n540 = ~new_n533 & ~new_n534;
  assign new_n541 = ~new_n535 & ~new_n540;
  assign new_n542 = ~\a[20]  & ~\b[20] ;
  assign new_n543 = \a[20]  & \b[20] ;
  assign new_n544 = ~new_n542 & ~new_n543;
  assign new_n545 = new_n541 & ~new_n544;
  assign new_n546 = ~new_n541 & new_n544;
  assign \f[20]  = ~new_n545 & ~new_n546;
  assign new_n548 = ~new_n541 & ~new_n542;
  assign new_n549 = ~new_n543 & ~new_n548;
  assign new_n550 = ~\a[21]  & ~\b[21] ;
  assign new_n551 = \a[21]  & \b[21] ;
  assign new_n552 = ~new_n550 & ~new_n551;
  assign new_n553 = new_n549 & ~new_n552;
  assign new_n554 = ~new_n549 & new_n552;
  assign \f[21]  = ~new_n553 & ~new_n554;
  assign new_n556 = ~new_n549 & ~new_n550;
  assign new_n557 = ~new_n551 & ~new_n556;
  assign new_n558 = ~\a[22]  & ~\b[22] ;
  assign new_n559 = \a[22]  & \b[22] ;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = new_n557 & ~new_n560;
  assign new_n562 = ~new_n557 & new_n560;
  assign \f[22]  = ~new_n561 & ~new_n562;
  assign new_n564 = ~new_n557 & ~new_n558;
  assign new_n565 = ~new_n559 & ~new_n564;
  assign new_n566 = ~\a[23]  & ~\b[23] ;
  assign new_n567 = \a[23]  & \b[23] ;
  assign new_n568 = ~new_n566 & ~new_n567;
  assign new_n569 = new_n565 & ~new_n568;
  assign new_n570 = ~new_n565 & new_n568;
  assign \f[23]  = ~new_n569 & ~new_n570;
  assign new_n572 = ~new_n565 & ~new_n566;
  assign new_n573 = ~new_n567 & ~new_n572;
  assign new_n574 = ~\a[24]  & ~\b[24] ;
  assign new_n575 = \a[24]  & \b[24] ;
  assign new_n576 = ~new_n574 & ~new_n575;
  assign new_n577 = new_n573 & ~new_n576;
  assign new_n578 = ~new_n573 & new_n576;
  assign \f[24]  = ~new_n577 & ~new_n578;
  assign new_n580 = ~new_n573 & ~new_n574;
  assign new_n581 = ~new_n575 & ~new_n580;
  assign new_n582 = ~\a[25]  & ~\b[25] ;
  assign new_n583 = \a[25]  & \b[25] ;
  assign new_n584 = ~new_n582 & ~new_n583;
  assign new_n585 = new_n581 & ~new_n584;
  assign new_n586 = ~new_n581 & new_n584;
  assign \f[25]  = ~new_n585 & ~new_n586;
  assign new_n588 = ~new_n581 & ~new_n582;
  assign new_n589 = ~new_n583 & ~new_n588;
  assign new_n590 = ~\a[26]  & ~\b[26] ;
  assign new_n591 = \a[26]  & \b[26] ;
  assign new_n592 = ~new_n590 & ~new_n591;
  assign new_n593 = new_n589 & ~new_n592;
  assign new_n594 = ~new_n589 & new_n592;
  assign \f[26]  = ~new_n593 & ~new_n594;
  assign new_n596 = ~new_n589 & ~new_n590;
  assign new_n597 = ~new_n591 & ~new_n596;
  assign new_n598 = ~\a[27]  & ~\b[27] ;
  assign new_n599 = \a[27]  & \b[27] ;
  assign new_n600 = ~new_n598 & ~new_n599;
  assign new_n601 = new_n597 & ~new_n600;
  assign new_n602 = ~new_n597 & new_n600;
  assign \f[27]  = ~new_n601 & ~new_n602;
  assign new_n604 = ~new_n597 & ~new_n598;
  assign new_n605 = ~new_n599 & ~new_n604;
  assign new_n606 = ~\a[28]  & ~\b[28] ;
  assign new_n607 = \a[28]  & \b[28] ;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = new_n605 & ~new_n608;
  assign new_n610 = ~new_n605 & new_n608;
  assign \f[28]  = ~new_n609 & ~new_n610;
  assign new_n612 = ~new_n605 & ~new_n606;
  assign new_n613 = ~new_n607 & ~new_n612;
  assign new_n614 = ~\a[29]  & ~\b[29] ;
  assign new_n615 = \a[29]  & \b[29] ;
  assign new_n616 = ~new_n614 & ~new_n615;
  assign new_n617 = new_n613 & ~new_n616;
  assign new_n618 = ~new_n613 & new_n616;
  assign \f[29]  = ~new_n617 & ~new_n618;
  assign new_n620 = ~new_n613 & ~new_n614;
  assign new_n621 = ~new_n615 & ~new_n620;
  assign new_n622 = ~\a[30]  & ~\b[30] ;
  assign new_n623 = \a[30]  & \b[30] ;
  assign new_n624 = ~new_n622 & ~new_n623;
  assign new_n625 = new_n621 & ~new_n624;
  assign new_n626 = ~new_n621 & new_n624;
  assign \f[30]  = ~new_n625 & ~new_n626;
  assign new_n628 = ~new_n621 & ~new_n622;
  assign new_n629 = ~new_n623 & ~new_n628;
  assign new_n630 = ~\a[31]  & ~\b[31] ;
  assign new_n631 = \a[31]  & \b[31] ;
  assign new_n632 = ~new_n630 & ~new_n631;
  assign new_n633 = new_n629 & ~new_n632;
  assign new_n634 = ~new_n629 & new_n632;
  assign \f[31]  = ~new_n633 & ~new_n634;
  assign new_n636 = ~new_n629 & ~new_n630;
  assign new_n637 = ~new_n631 & ~new_n636;
  assign new_n638 = ~\a[32]  & ~\b[32] ;
  assign new_n639 = \a[32]  & \b[32] ;
  assign new_n640 = ~new_n638 & ~new_n639;
  assign new_n641 = new_n637 & ~new_n640;
  assign new_n642 = ~new_n637 & new_n640;
  assign \f[32]  = ~new_n641 & ~new_n642;
  assign new_n644 = ~new_n637 & ~new_n638;
  assign new_n645 = ~new_n639 & ~new_n644;
  assign new_n646 = ~\a[33]  & ~\b[33] ;
  assign new_n647 = \a[33]  & \b[33] ;
  assign new_n648 = ~new_n646 & ~new_n647;
  assign new_n649 = new_n645 & ~new_n648;
  assign new_n650 = ~new_n645 & new_n648;
  assign \f[33]  = ~new_n649 & ~new_n650;
  assign new_n652 = ~new_n645 & ~new_n646;
  assign new_n653 = ~new_n647 & ~new_n652;
  assign new_n654 = ~\a[34]  & ~\b[34] ;
  assign new_n655 = \a[34]  & \b[34] ;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = new_n653 & ~new_n656;
  assign new_n658 = ~new_n653 & new_n656;
  assign \f[34]  = ~new_n657 & ~new_n658;
  assign new_n660 = ~new_n653 & ~new_n654;
  assign new_n661 = ~new_n655 & ~new_n660;
  assign new_n662 = ~\a[35]  & ~\b[35] ;
  assign new_n663 = \a[35]  & \b[35] ;
  assign new_n664 = ~new_n662 & ~new_n663;
  assign new_n665 = new_n661 & ~new_n664;
  assign new_n666 = ~new_n661 & new_n664;
  assign \f[35]  = ~new_n665 & ~new_n666;
  assign new_n668 = ~new_n661 & ~new_n662;
  assign new_n669 = ~new_n663 & ~new_n668;
  assign new_n670 = ~\a[36]  & ~\b[36] ;
  assign new_n671 = \a[36]  & \b[36] ;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = new_n669 & ~new_n672;
  assign new_n674 = ~new_n669 & new_n672;
  assign \f[36]  = ~new_n673 & ~new_n674;
  assign new_n676 = ~new_n669 & ~new_n670;
  assign new_n677 = ~new_n671 & ~new_n676;
  assign new_n678 = ~\a[37]  & ~\b[37] ;
  assign new_n679 = \a[37]  & \b[37] ;
  assign new_n680 = ~new_n678 & ~new_n679;
  assign new_n681 = new_n677 & ~new_n680;
  assign new_n682 = ~new_n677 & new_n680;
  assign \f[37]  = ~new_n681 & ~new_n682;
  assign new_n684 = ~new_n677 & ~new_n678;
  assign new_n685 = ~new_n679 & ~new_n684;
  assign new_n686 = ~\a[38]  & ~\b[38] ;
  assign new_n687 = \a[38]  & \b[38] ;
  assign new_n688 = ~new_n686 & ~new_n687;
  assign new_n689 = new_n685 & ~new_n688;
  assign new_n690 = ~new_n685 & new_n688;
  assign \f[38]  = ~new_n689 & ~new_n690;
  assign new_n692 = ~new_n685 & ~new_n686;
  assign new_n693 = ~new_n687 & ~new_n692;
  assign new_n694 = ~\a[39]  & ~\b[39] ;
  assign new_n695 = \a[39]  & \b[39] ;
  assign new_n696 = ~new_n694 & ~new_n695;
  assign new_n697 = new_n693 & ~new_n696;
  assign new_n698 = ~new_n693 & new_n696;
  assign \f[39]  = ~new_n697 & ~new_n698;
  assign new_n700 = ~new_n693 & ~new_n694;
  assign new_n701 = ~new_n695 & ~new_n700;
  assign new_n702 = ~\a[40]  & ~\b[40] ;
  assign new_n703 = \a[40]  & \b[40] ;
  assign new_n704 = ~new_n702 & ~new_n703;
  assign new_n705 = new_n701 & ~new_n704;
  assign new_n706 = ~new_n701 & new_n704;
  assign \f[40]  = ~new_n705 & ~new_n706;
  assign new_n708 = ~new_n701 & ~new_n702;
  assign new_n709 = ~new_n703 & ~new_n708;
  assign new_n710 = ~\a[41]  & ~\b[41] ;
  assign new_n711 = \a[41]  & \b[41] ;
  assign new_n712 = ~new_n710 & ~new_n711;
  assign new_n713 = new_n709 & ~new_n712;
  assign new_n714 = ~new_n709 & new_n712;
  assign \f[41]  = ~new_n713 & ~new_n714;
  assign new_n716 = ~new_n709 & ~new_n710;
  assign new_n717 = ~new_n711 & ~new_n716;
  assign new_n718 = ~\a[42]  & ~\b[42] ;
  assign new_n719 = \a[42]  & \b[42] ;
  assign new_n720 = ~new_n718 & ~new_n719;
  assign new_n721 = new_n717 & ~new_n720;
  assign new_n722 = ~new_n717 & new_n720;
  assign \f[42]  = ~new_n721 & ~new_n722;
  assign new_n724 = ~new_n717 & ~new_n718;
  assign new_n725 = ~new_n719 & ~new_n724;
  assign new_n726 = ~\a[43]  & ~\b[43] ;
  assign new_n727 = \a[43]  & \b[43] ;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = new_n725 & ~new_n728;
  assign new_n730 = ~new_n725 & new_n728;
  assign \f[43]  = ~new_n729 & ~new_n730;
  assign new_n732 = ~new_n725 & ~new_n726;
  assign new_n733 = ~new_n727 & ~new_n732;
  assign new_n734 = ~\a[44]  & ~\b[44] ;
  assign new_n735 = \a[44]  & \b[44] ;
  assign new_n736 = ~new_n734 & ~new_n735;
  assign new_n737 = new_n733 & ~new_n736;
  assign new_n738 = ~new_n733 & new_n736;
  assign \f[44]  = ~new_n737 & ~new_n738;
  assign new_n740 = ~new_n733 & ~new_n734;
  assign new_n741 = ~new_n735 & ~new_n740;
  assign new_n742 = ~\a[45]  & ~\b[45] ;
  assign new_n743 = \a[45]  & \b[45] ;
  assign new_n744 = ~new_n742 & ~new_n743;
  assign new_n745 = new_n741 & ~new_n744;
  assign new_n746 = ~new_n741 & new_n744;
  assign \f[45]  = ~new_n745 & ~new_n746;
  assign new_n748 = ~new_n741 & ~new_n742;
  assign new_n749 = ~new_n743 & ~new_n748;
  assign new_n750 = ~\a[46]  & ~\b[46] ;
  assign new_n751 = \a[46]  & \b[46] ;
  assign new_n752 = ~new_n750 & ~new_n751;
  assign new_n753 = new_n749 & ~new_n752;
  assign new_n754 = ~new_n749 & new_n752;
  assign \f[46]  = ~new_n753 & ~new_n754;
  assign new_n756 = ~new_n749 & ~new_n750;
  assign new_n757 = ~new_n751 & ~new_n756;
  assign new_n758 = ~\a[47]  & ~\b[47] ;
  assign new_n759 = \a[47]  & \b[47] ;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = new_n757 & ~new_n760;
  assign new_n762 = ~new_n757 & new_n760;
  assign \f[47]  = ~new_n761 & ~new_n762;
  assign new_n764 = ~new_n757 & ~new_n758;
  assign new_n765 = ~new_n759 & ~new_n764;
  assign new_n766 = ~\a[48]  & ~\b[48] ;
  assign new_n767 = \a[48]  & \b[48] ;
  assign new_n768 = ~new_n766 & ~new_n767;
  assign new_n769 = new_n765 & ~new_n768;
  assign new_n770 = ~new_n765 & new_n768;
  assign \f[48]  = ~new_n769 & ~new_n770;
  assign new_n772 = ~new_n765 & ~new_n766;
  assign new_n773 = ~new_n767 & ~new_n772;
  assign new_n774 = ~\a[49]  & ~\b[49] ;
  assign new_n775 = \a[49]  & \b[49] ;
  assign new_n776 = ~new_n774 & ~new_n775;
  assign new_n777 = new_n773 & ~new_n776;
  assign new_n778 = ~new_n773 & new_n776;
  assign \f[49]  = ~new_n777 & ~new_n778;
  assign new_n780 = ~new_n773 & ~new_n774;
  assign new_n781 = ~new_n775 & ~new_n780;
  assign new_n782 = ~\a[50]  & ~\b[50] ;
  assign new_n783 = \a[50]  & \b[50] ;
  assign new_n784 = ~new_n782 & ~new_n783;
  assign new_n785 = new_n781 & ~new_n784;
  assign new_n786 = ~new_n781 & new_n784;
  assign \f[50]  = ~new_n785 & ~new_n786;
  assign new_n788 = ~new_n781 & ~new_n782;
  assign new_n789 = ~new_n783 & ~new_n788;
  assign new_n790 = ~\a[51]  & ~\b[51] ;
  assign new_n791 = \a[51]  & \b[51] ;
  assign new_n792 = ~new_n790 & ~new_n791;
  assign new_n793 = new_n789 & ~new_n792;
  assign new_n794 = ~new_n789 & new_n792;
  assign \f[51]  = ~new_n793 & ~new_n794;
  assign new_n796 = ~new_n789 & ~new_n790;
  assign new_n797 = ~new_n791 & ~new_n796;
  assign new_n798 = ~\a[52]  & ~\b[52] ;
  assign new_n799 = \a[52]  & \b[52] ;
  assign new_n800 = ~new_n798 & ~new_n799;
  assign new_n801 = new_n797 & ~new_n800;
  assign new_n802 = ~new_n797 & new_n800;
  assign \f[52]  = ~new_n801 & ~new_n802;
  assign new_n804 = ~new_n797 & ~new_n798;
  assign new_n805 = ~new_n799 & ~new_n804;
  assign new_n806 = ~\a[53]  & ~\b[53] ;
  assign new_n807 = \a[53]  & \b[53] ;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = new_n805 & ~new_n808;
  assign new_n810 = ~new_n805 & new_n808;
  assign \f[53]  = ~new_n809 & ~new_n810;
  assign new_n812 = ~new_n805 & ~new_n806;
  assign new_n813 = ~new_n807 & ~new_n812;
  assign new_n814 = ~\a[54]  & ~\b[54] ;
  assign new_n815 = \a[54]  & \b[54] ;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817 = new_n813 & ~new_n816;
  assign new_n818 = ~new_n813 & new_n816;
  assign \f[54]  = ~new_n817 & ~new_n818;
  assign new_n820 = ~new_n813 & ~new_n814;
  assign new_n821 = ~new_n815 & ~new_n820;
  assign new_n822 = ~\a[55]  & ~\b[55] ;
  assign new_n823 = \a[55]  & \b[55] ;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = new_n821 & ~new_n824;
  assign new_n826 = ~new_n821 & new_n824;
  assign \f[55]  = ~new_n825 & ~new_n826;
  assign new_n828 = ~new_n821 & ~new_n822;
  assign new_n829 = ~new_n823 & ~new_n828;
  assign new_n830 = ~\a[56]  & ~\b[56] ;
  assign new_n831 = \a[56]  & \b[56] ;
  assign new_n832 = ~new_n830 & ~new_n831;
  assign new_n833 = new_n829 & ~new_n832;
  assign new_n834 = ~new_n829 & new_n832;
  assign \f[56]  = ~new_n833 & ~new_n834;
  assign new_n836 = ~new_n829 & ~new_n830;
  assign new_n837 = ~new_n831 & ~new_n836;
  assign new_n838 = ~\a[57]  & ~\b[57] ;
  assign new_n839 = \a[57]  & \b[57] ;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = new_n837 & ~new_n840;
  assign new_n842 = ~new_n837 & new_n840;
  assign \f[57]  = ~new_n841 & ~new_n842;
  assign new_n844 = ~new_n837 & ~new_n838;
  assign new_n845 = ~new_n839 & ~new_n844;
  assign new_n846 = ~\a[58]  & ~\b[58] ;
  assign new_n847 = \a[58]  & \b[58] ;
  assign new_n848 = ~new_n846 & ~new_n847;
  assign new_n849 = new_n845 & ~new_n848;
  assign new_n850 = ~new_n845 & new_n848;
  assign \f[58]  = ~new_n849 & ~new_n850;
  assign new_n852 = ~new_n845 & ~new_n846;
  assign new_n853 = ~new_n847 & ~new_n852;
  assign new_n854 = ~\a[59]  & ~\b[59] ;
  assign new_n855 = \a[59]  & \b[59] ;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = new_n853 & ~new_n856;
  assign new_n858 = ~new_n853 & new_n856;
  assign \f[59]  = ~new_n857 & ~new_n858;
  assign new_n860 = ~new_n853 & ~new_n854;
  assign new_n861 = ~new_n855 & ~new_n860;
  assign new_n862 = ~\a[60]  & ~\b[60] ;
  assign new_n863 = \a[60]  & \b[60] ;
  assign new_n864 = ~new_n862 & ~new_n863;
  assign new_n865 = new_n861 & ~new_n864;
  assign new_n866 = ~new_n861 & new_n864;
  assign \f[60]  = ~new_n865 & ~new_n866;
  assign new_n868 = ~new_n861 & ~new_n862;
  assign new_n869 = ~new_n863 & ~new_n868;
  assign new_n870 = ~\a[61]  & ~\b[61] ;
  assign new_n871 = \a[61]  & \b[61] ;
  assign new_n872 = ~new_n870 & ~new_n871;
  assign new_n873 = new_n869 & ~new_n872;
  assign new_n874 = ~new_n869 & new_n872;
  assign \f[61]  = ~new_n873 & ~new_n874;
  assign new_n876 = ~new_n869 & ~new_n870;
  assign new_n877 = ~new_n871 & ~new_n876;
  assign new_n878 = ~\a[62]  & ~\b[62] ;
  assign new_n879 = \a[62]  & \b[62] ;
  assign new_n880 = ~new_n878 & ~new_n879;
  assign new_n881 = new_n877 & ~new_n880;
  assign new_n882 = ~new_n877 & new_n880;
  assign \f[62]  = ~new_n881 & ~new_n882;
  assign new_n884 = ~new_n877 & ~new_n878;
  assign new_n885 = ~new_n879 & ~new_n884;
  assign new_n886 = ~\a[63]  & ~\b[63] ;
  assign new_n887 = \a[63]  & \b[63] ;
  assign new_n888 = ~new_n886 & ~new_n887;
  assign new_n889 = new_n885 & ~new_n888;
  assign new_n890 = ~new_n885 & new_n888;
  assign \f[63]  = ~new_n889 & ~new_n890;
  assign new_n892 = ~new_n885 & ~new_n886;
  assign new_n893 = ~new_n887 & ~new_n892;
  assign new_n894 = ~\a[64]  & ~\b[64] ;
  assign new_n895 = \a[64]  & \b[64] ;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = new_n893 & ~new_n896;
  assign new_n898 = ~new_n893 & new_n896;
  assign \f[64]  = ~new_n897 & ~new_n898;
  assign new_n900 = ~new_n893 & ~new_n894;
  assign new_n901 = ~new_n895 & ~new_n900;
  assign new_n902 = ~\a[65]  & ~\b[65] ;
  assign new_n903 = \a[65]  & \b[65] ;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = new_n901 & ~new_n904;
  assign new_n906 = ~new_n901 & new_n904;
  assign \f[65]  = ~new_n905 & ~new_n906;
  assign new_n908 = ~new_n901 & ~new_n902;
  assign new_n909 = ~new_n903 & ~new_n908;
  assign new_n910 = ~\a[66]  & ~\b[66] ;
  assign new_n911 = \a[66]  & \b[66] ;
  assign new_n912 = ~new_n910 & ~new_n911;
  assign new_n913 = new_n909 & ~new_n912;
  assign new_n914 = ~new_n909 & new_n912;
  assign \f[66]  = ~new_n913 & ~new_n914;
  assign new_n916 = ~new_n909 & ~new_n910;
  assign new_n917 = ~new_n911 & ~new_n916;
  assign new_n918 = ~\a[67]  & ~\b[67] ;
  assign new_n919 = \a[67]  & \b[67] ;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = new_n917 & ~new_n920;
  assign new_n922 = ~new_n917 & new_n920;
  assign \f[67]  = ~new_n921 & ~new_n922;
  assign new_n924 = ~new_n917 & ~new_n918;
  assign new_n925 = ~new_n919 & ~new_n924;
  assign new_n926 = ~\a[68]  & ~\b[68] ;
  assign new_n927 = \a[68]  & \b[68] ;
  assign new_n928 = ~new_n926 & ~new_n927;
  assign new_n929 = new_n925 & ~new_n928;
  assign new_n930 = ~new_n925 & new_n928;
  assign \f[68]  = ~new_n929 & ~new_n930;
  assign new_n932 = ~new_n925 & ~new_n926;
  assign new_n933 = ~new_n927 & ~new_n932;
  assign new_n934 = ~\a[69]  & ~\b[69] ;
  assign new_n935 = \a[69]  & \b[69] ;
  assign new_n936 = ~new_n934 & ~new_n935;
  assign new_n937 = new_n933 & ~new_n936;
  assign new_n938 = ~new_n933 & new_n936;
  assign \f[69]  = ~new_n937 & ~new_n938;
  assign new_n940 = ~new_n933 & ~new_n934;
  assign new_n941 = ~new_n935 & ~new_n940;
  assign new_n942 = ~\a[70]  & ~\b[70] ;
  assign new_n943 = \a[70]  & \b[70] ;
  assign new_n944 = ~new_n942 & ~new_n943;
  assign new_n945 = new_n941 & ~new_n944;
  assign new_n946 = ~new_n941 & new_n944;
  assign \f[70]  = ~new_n945 & ~new_n946;
  assign new_n948 = ~new_n941 & ~new_n942;
  assign new_n949 = ~new_n943 & ~new_n948;
  assign new_n950 = ~\a[71]  & ~\b[71] ;
  assign new_n951 = \a[71]  & \b[71] ;
  assign new_n952 = ~new_n950 & ~new_n951;
  assign new_n953 = new_n949 & ~new_n952;
  assign new_n954 = ~new_n949 & new_n952;
  assign \f[71]  = ~new_n953 & ~new_n954;
  assign new_n956 = ~new_n949 & ~new_n950;
  assign new_n957 = ~new_n951 & ~new_n956;
  assign new_n958 = ~\a[72]  & ~\b[72] ;
  assign new_n959 = \a[72]  & \b[72] ;
  assign new_n960 = ~new_n958 & ~new_n959;
  assign new_n961 = new_n957 & ~new_n960;
  assign new_n962 = ~new_n957 & new_n960;
  assign \f[72]  = ~new_n961 & ~new_n962;
  assign new_n964 = ~new_n957 & ~new_n958;
  assign new_n965 = ~new_n959 & ~new_n964;
  assign new_n966 = ~\a[73]  & ~\b[73] ;
  assign new_n967 = \a[73]  & \b[73] ;
  assign new_n968 = ~new_n966 & ~new_n967;
  assign new_n969 = new_n965 & ~new_n968;
  assign new_n970 = ~new_n965 & new_n968;
  assign \f[73]  = ~new_n969 & ~new_n970;
  assign new_n972 = ~new_n965 & ~new_n966;
  assign new_n973 = ~new_n967 & ~new_n972;
  assign new_n974 = ~\a[74]  & ~\b[74] ;
  assign new_n975 = \a[74]  & \b[74] ;
  assign new_n976 = ~new_n974 & ~new_n975;
  assign new_n977 = new_n973 & ~new_n976;
  assign new_n978 = ~new_n973 & new_n976;
  assign \f[74]  = ~new_n977 & ~new_n978;
  assign new_n980 = ~new_n973 & ~new_n974;
  assign new_n981 = ~new_n975 & ~new_n980;
  assign new_n982 = ~\a[75]  & ~\b[75] ;
  assign new_n983 = \a[75]  & \b[75] ;
  assign new_n984 = ~new_n982 & ~new_n983;
  assign new_n985 = new_n981 & ~new_n984;
  assign new_n986 = ~new_n981 & new_n984;
  assign \f[75]  = ~new_n985 & ~new_n986;
  assign new_n988 = ~new_n981 & ~new_n982;
  assign new_n989 = ~new_n983 & ~new_n988;
  assign new_n990 = ~\a[76]  & ~\b[76] ;
  assign new_n991 = \a[76]  & \b[76] ;
  assign new_n992 = ~new_n990 & ~new_n991;
  assign new_n993 = new_n989 & ~new_n992;
  assign new_n994 = ~new_n989 & new_n992;
  assign \f[76]  = ~new_n993 & ~new_n994;
  assign new_n996 = ~new_n989 & ~new_n990;
  assign new_n997 = ~new_n991 & ~new_n996;
  assign new_n998 = ~\a[77]  & ~\b[77] ;
  assign new_n999 = \a[77]  & \b[77] ;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = new_n997 & ~new_n1000;
  assign new_n1002 = ~new_n997 & new_n1000;
  assign \f[77]  = ~new_n1001 & ~new_n1002;
  assign new_n1004 = ~new_n997 & ~new_n998;
  assign new_n1005 = ~new_n999 & ~new_n1004;
  assign new_n1006 = ~\a[78]  & ~\b[78] ;
  assign new_n1007 = \a[78]  & \b[78] ;
  assign new_n1008 = ~new_n1006 & ~new_n1007;
  assign new_n1009 = new_n1005 & ~new_n1008;
  assign new_n1010 = ~new_n1005 & new_n1008;
  assign \f[78]  = ~new_n1009 & ~new_n1010;
  assign new_n1012 = ~new_n1005 & ~new_n1006;
  assign new_n1013 = ~new_n1007 & ~new_n1012;
  assign new_n1014 = ~\a[79]  & ~\b[79] ;
  assign new_n1015 = \a[79]  & \b[79] ;
  assign new_n1016 = ~new_n1014 & ~new_n1015;
  assign new_n1017 = new_n1013 & ~new_n1016;
  assign new_n1018 = ~new_n1013 & new_n1016;
  assign \f[79]  = ~new_n1017 & ~new_n1018;
  assign new_n1020 = ~new_n1013 & ~new_n1014;
  assign new_n1021 = ~new_n1015 & ~new_n1020;
  assign new_n1022 = ~\a[80]  & ~\b[80] ;
  assign new_n1023 = \a[80]  & \b[80] ;
  assign new_n1024 = ~new_n1022 & ~new_n1023;
  assign new_n1025 = new_n1021 & ~new_n1024;
  assign new_n1026 = ~new_n1021 & new_n1024;
  assign \f[80]  = ~new_n1025 & ~new_n1026;
  assign new_n1028 = ~new_n1021 & ~new_n1022;
  assign new_n1029 = ~new_n1023 & ~new_n1028;
  assign new_n1030 = ~\a[81]  & ~\b[81] ;
  assign new_n1031 = \a[81]  & \b[81] ;
  assign new_n1032 = ~new_n1030 & ~new_n1031;
  assign new_n1033 = new_n1029 & ~new_n1032;
  assign new_n1034 = ~new_n1029 & new_n1032;
  assign \f[81]  = ~new_n1033 & ~new_n1034;
  assign new_n1036 = ~new_n1029 & ~new_n1030;
  assign new_n1037 = ~new_n1031 & ~new_n1036;
  assign new_n1038 = ~\a[82]  & ~\b[82] ;
  assign new_n1039 = \a[82]  & \b[82] ;
  assign new_n1040 = ~new_n1038 & ~new_n1039;
  assign new_n1041 = new_n1037 & ~new_n1040;
  assign new_n1042 = ~new_n1037 & new_n1040;
  assign \f[82]  = ~new_n1041 & ~new_n1042;
  assign new_n1044 = ~new_n1037 & ~new_n1038;
  assign new_n1045 = ~new_n1039 & ~new_n1044;
  assign new_n1046 = ~\a[83]  & ~\b[83] ;
  assign new_n1047 = \a[83]  & \b[83] ;
  assign new_n1048 = ~new_n1046 & ~new_n1047;
  assign new_n1049 = new_n1045 & ~new_n1048;
  assign new_n1050 = ~new_n1045 & new_n1048;
  assign \f[83]  = ~new_n1049 & ~new_n1050;
  assign new_n1052 = ~new_n1045 & ~new_n1046;
  assign new_n1053 = ~new_n1047 & ~new_n1052;
  assign new_n1054 = ~\a[84]  & ~\b[84] ;
  assign new_n1055 = \a[84]  & \b[84] ;
  assign new_n1056 = ~new_n1054 & ~new_n1055;
  assign new_n1057 = new_n1053 & ~new_n1056;
  assign new_n1058 = ~new_n1053 & new_n1056;
  assign \f[84]  = ~new_n1057 & ~new_n1058;
  assign new_n1060 = ~new_n1053 & ~new_n1054;
  assign new_n1061 = ~new_n1055 & ~new_n1060;
  assign new_n1062 = ~\a[85]  & ~\b[85] ;
  assign new_n1063 = \a[85]  & \b[85] ;
  assign new_n1064 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = new_n1061 & ~new_n1064;
  assign new_n1066 = ~new_n1061 & new_n1064;
  assign \f[85]  = ~new_n1065 & ~new_n1066;
  assign new_n1068 = ~new_n1061 & ~new_n1062;
  assign new_n1069 = ~new_n1063 & ~new_n1068;
  assign new_n1070 = ~\a[86]  & ~\b[86] ;
  assign new_n1071 = \a[86]  & \b[86] ;
  assign new_n1072 = ~new_n1070 & ~new_n1071;
  assign new_n1073 = new_n1069 & ~new_n1072;
  assign new_n1074 = ~new_n1069 & new_n1072;
  assign \f[86]  = ~new_n1073 & ~new_n1074;
  assign new_n1076 = ~new_n1069 & ~new_n1070;
  assign new_n1077 = ~new_n1071 & ~new_n1076;
  assign new_n1078 = ~\a[87]  & ~\b[87] ;
  assign new_n1079 = \a[87]  & \b[87] ;
  assign new_n1080 = ~new_n1078 & ~new_n1079;
  assign new_n1081 = new_n1077 & ~new_n1080;
  assign new_n1082 = ~new_n1077 & new_n1080;
  assign \f[87]  = ~new_n1081 & ~new_n1082;
  assign new_n1084 = ~new_n1077 & ~new_n1078;
  assign new_n1085 = ~new_n1079 & ~new_n1084;
  assign new_n1086 = ~\a[88]  & ~\b[88] ;
  assign new_n1087 = \a[88]  & \b[88] ;
  assign new_n1088 = ~new_n1086 & ~new_n1087;
  assign new_n1089 = new_n1085 & ~new_n1088;
  assign new_n1090 = ~new_n1085 & new_n1088;
  assign \f[88]  = ~new_n1089 & ~new_n1090;
  assign new_n1092 = ~new_n1085 & ~new_n1086;
  assign new_n1093 = ~new_n1087 & ~new_n1092;
  assign new_n1094 = ~\a[89]  & ~\b[89] ;
  assign new_n1095 = \a[89]  & \b[89] ;
  assign new_n1096 = ~new_n1094 & ~new_n1095;
  assign new_n1097 = new_n1093 & ~new_n1096;
  assign new_n1098 = ~new_n1093 & new_n1096;
  assign \f[89]  = ~new_n1097 & ~new_n1098;
  assign new_n1100 = ~new_n1093 & ~new_n1094;
  assign new_n1101 = ~new_n1095 & ~new_n1100;
  assign new_n1102 = ~\a[90]  & ~\b[90] ;
  assign new_n1103 = \a[90]  & \b[90] ;
  assign new_n1104 = ~new_n1102 & ~new_n1103;
  assign new_n1105 = new_n1101 & ~new_n1104;
  assign new_n1106 = ~new_n1101 & new_n1104;
  assign \f[90]  = ~new_n1105 & ~new_n1106;
  assign new_n1108 = ~new_n1101 & ~new_n1102;
  assign new_n1109 = ~new_n1103 & ~new_n1108;
  assign new_n1110 = ~\a[91]  & ~\b[91] ;
  assign new_n1111 = \a[91]  & \b[91] ;
  assign new_n1112 = ~new_n1110 & ~new_n1111;
  assign new_n1113 = new_n1109 & ~new_n1112;
  assign new_n1114 = ~new_n1109 & new_n1112;
  assign \f[91]  = ~new_n1113 & ~new_n1114;
  assign new_n1116 = ~new_n1109 & ~new_n1110;
  assign new_n1117 = ~new_n1111 & ~new_n1116;
  assign new_n1118 = ~\a[92]  & ~\b[92] ;
  assign new_n1119 = \a[92]  & \b[92] ;
  assign new_n1120 = ~new_n1118 & ~new_n1119;
  assign new_n1121 = new_n1117 & ~new_n1120;
  assign new_n1122 = ~new_n1117 & new_n1120;
  assign \f[92]  = ~new_n1121 & ~new_n1122;
  assign new_n1124 = ~new_n1117 & ~new_n1118;
  assign new_n1125 = ~new_n1119 & ~new_n1124;
  assign new_n1126 = ~\a[93]  & ~\b[93] ;
  assign new_n1127 = \a[93]  & \b[93] ;
  assign new_n1128 = ~new_n1126 & ~new_n1127;
  assign new_n1129 = new_n1125 & ~new_n1128;
  assign new_n1130 = ~new_n1125 & new_n1128;
  assign \f[93]  = ~new_n1129 & ~new_n1130;
  assign new_n1132 = ~new_n1125 & ~new_n1126;
  assign new_n1133 = ~new_n1127 & ~new_n1132;
  assign new_n1134 = ~\a[94]  & ~\b[94] ;
  assign new_n1135 = \a[94]  & \b[94] ;
  assign new_n1136 = ~new_n1134 & ~new_n1135;
  assign new_n1137 = new_n1133 & ~new_n1136;
  assign new_n1138 = ~new_n1133 & new_n1136;
  assign \f[94]  = ~new_n1137 & ~new_n1138;
  assign new_n1140 = ~new_n1133 & ~new_n1134;
  assign new_n1141 = ~new_n1135 & ~new_n1140;
  assign new_n1142 = ~\a[95]  & ~\b[95] ;
  assign new_n1143 = \a[95]  & \b[95] ;
  assign new_n1144 = ~new_n1142 & ~new_n1143;
  assign new_n1145 = new_n1141 & ~new_n1144;
  assign new_n1146 = ~new_n1141 & new_n1144;
  assign \f[95]  = ~new_n1145 & ~new_n1146;
  assign new_n1148 = ~new_n1141 & ~new_n1142;
  assign new_n1149 = ~new_n1143 & ~new_n1148;
  assign new_n1150 = ~\a[96]  & ~\b[96] ;
  assign new_n1151 = \a[96]  & \b[96] ;
  assign new_n1152 = ~new_n1150 & ~new_n1151;
  assign new_n1153 = new_n1149 & ~new_n1152;
  assign new_n1154 = ~new_n1149 & new_n1152;
  assign \f[96]  = ~new_n1153 & ~new_n1154;
  assign new_n1156 = ~new_n1149 & ~new_n1150;
  assign new_n1157 = ~new_n1151 & ~new_n1156;
  assign new_n1158 = ~\a[97]  & ~\b[97] ;
  assign new_n1159 = \a[97]  & \b[97] ;
  assign new_n1160 = ~new_n1158 & ~new_n1159;
  assign new_n1161 = new_n1157 & ~new_n1160;
  assign new_n1162 = ~new_n1157 & new_n1160;
  assign \f[97]  = ~new_n1161 & ~new_n1162;
  assign new_n1164 = ~new_n1157 & ~new_n1158;
  assign new_n1165 = ~new_n1159 & ~new_n1164;
  assign new_n1166 = ~\a[98]  & ~\b[98] ;
  assign new_n1167 = \a[98]  & \b[98] ;
  assign new_n1168 = ~new_n1166 & ~new_n1167;
  assign new_n1169 = new_n1165 & ~new_n1168;
  assign new_n1170 = ~new_n1165 & new_n1168;
  assign \f[98]  = ~new_n1169 & ~new_n1170;
  assign new_n1172 = ~new_n1165 & ~new_n1166;
  assign new_n1173 = ~new_n1167 & ~new_n1172;
  assign new_n1174 = ~\a[99]  & ~\b[99] ;
  assign new_n1175 = \a[99]  & \b[99] ;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = new_n1173 & ~new_n1176;
  assign new_n1178 = ~new_n1173 & new_n1176;
  assign \f[99]  = ~new_n1177 & ~new_n1178;
  assign new_n1180 = ~new_n1173 & ~new_n1174;
  assign new_n1181 = ~new_n1175 & ~new_n1180;
  assign new_n1182 = ~\a[100]  & ~\b[100] ;
  assign new_n1183 = \a[100]  & \b[100] ;
  assign new_n1184 = ~new_n1182 & ~new_n1183;
  assign new_n1185 = new_n1181 & ~new_n1184;
  assign new_n1186 = ~new_n1181 & new_n1184;
  assign \f[100]  = ~new_n1185 & ~new_n1186;
  assign new_n1188 = ~new_n1181 & ~new_n1182;
  assign new_n1189 = ~new_n1183 & ~new_n1188;
  assign new_n1190 = ~\a[101]  & ~\b[101] ;
  assign new_n1191 = \a[101]  & \b[101] ;
  assign new_n1192 = ~new_n1190 & ~new_n1191;
  assign new_n1193 = new_n1189 & ~new_n1192;
  assign new_n1194 = ~new_n1189 & new_n1192;
  assign \f[101]  = ~new_n1193 & ~new_n1194;
  assign new_n1196 = ~new_n1189 & ~new_n1190;
  assign new_n1197 = ~new_n1191 & ~new_n1196;
  assign new_n1198 = ~\a[102]  & ~\b[102] ;
  assign new_n1199 = \a[102]  & \b[102] ;
  assign new_n1200 = ~new_n1198 & ~new_n1199;
  assign new_n1201 = new_n1197 & ~new_n1200;
  assign new_n1202 = ~new_n1197 & new_n1200;
  assign \f[102]  = ~new_n1201 & ~new_n1202;
  assign new_n1204 = ~new_n1197 & ~new_n1198;
  assign new_n1205 = ~new_n1199 & ~new_n1204;
  assign new_n1206 = ~\a[103]  & ~\b[103] ;
  assign new_n1207 = \a[103]  & \b[103] ;
  assign new_n1208 = ~new_n1206 & ~new_n1207;
  assign new_n1209 = new_n1205 & ~new_n1208;
  assign new_n1210 = ~new_n1205 & new_n1208;
  assign \f[103]  = ~new_n1209 & ~new_n1210;
  assign new_n1212 = ~new_n1205 & ~new_n1206;
  assign new_n1213 = ~new_n1207 & ~new_n1212;
  assign new_n1214 = ~\a[104]  & ~\b[104] ;
  assign new_n1215 = \a[104]  & \b[104] ;
  assign new_n1216 = ~new_n1214 & ~new_n1215;
  assign new_n1217 = new_n1213 & ~new_n1216;
  assign new_n1218 = ~new_n1213 & new_n1216;
  assign \f[104]  = ~new_n1217 & ~new_n1218;
  assign new_n1220 = ~new_n1213 & ~new_n1214;
  assign new_n1221 = ~new_n1215 & ~new_n1220;
  assign new_n1222 = ~\a[105]  & ~\b[105] ;
  assign new_n1223 = \a[105]  & \b[105] ;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = new_n1221 & ~new_n1224;
  assign new_n1226 = ~new_n1221 & new_n1224;
  assign \f[105]  = ~new_n1225 & ~new_n1226;
  assign new_n1228 = ~new_n1221 & ~new_n1222;
  assign new_n1229 = ~new_n1223 & ~new_n1228;
  assign new_n1230 = ~\a[106]  & ~\b[106] ;
  assign new_n1231 = \a[106]  & \b[106] ;
  assign new_n1232 = ~new_n1230 & ~new_n1231;
  assign new_n1233 = new_n1229 & ~new_n1232;
  assign new_n1234 = ~new_n1229 & new_n1232;
  assign \f[106]  = ~new_n1233 & ~new_n1234;
  assign new_n1236 = ~new_n1229 & ~new_n1230;
  assign new_n1237 = ~new_n1231 & ~new_n1236;
  assign new_n1238 = ~\a[107]  & ~\b[107] ;
  assign new_n1239 = \a[107]  & \b[107] ;
  assign new_n1240 = ~new_n1238 & ~new_n1239;
  assign new_n1241 = new_n1237 & ~new_n1240;
  assign new_n1242 = ~new_n1237 & new_n1240;
  assign \f[107]  = ~new_n1241 & ~new_n1242;
  assign new_n1244 = ~new_n1237 & ~new_n1238;
  assign new_n1245 = ~new_n1239 & ~new_n1244;
  assign new_n1246 = ~\a[108]  & ~\b[108] ;
  assign new_n1247 = \a[108]  & \b[108] ;
  assign new_n1248 = ~new_n1246 & ~new_n1247;
  assign new_n1249 = new_n1245 & ~new_n1248;
  assign new_n1250 = ~new_n1245 & new_n1248;
  assign \f[108]  = ~new_n1249 & ~new_n1250;
  assign new_n1252 = ~new_n1245 & ~new_n1246;
  assign new_n1253 = ~new_n1247 & ~new_n1252;
  assign new_n1254 = ~\a[109]  & ~\b[109] ;
  assign new_n1255 = \a[109]  & \b[109] ;
  assign new_n1256 = ~new_n1254 & ~new_n1255;
  assign new_n1257 = new_n1253 & ~new_n1256;
  assign new_n1258 = ~new_n1253 & new_n1256;
  assign \f[109]  = ~new_n1257 & ~new_n1258;
  assign new_n1260 = ~new_n1253 & ~new_n1254;
  assign new_n1261 = ~new_n1255 & ~new_n1260;
  assign new_n1262 = ~\a[110]  & ~\b[110] ;
  assign new_n1263 = \a[110]  & \b[110] ;
  assign new_n1264 = ~new_n1262 & ~new_n1263;
  assign new_n1265 = new_n1261 & ~new_n1264;
  assign new_n1266 = ~new_n1261 & new_n1264;
  assign \f[110]  = ~new_n1265 & ~new_n1266;
  assign new_n1268 = ~new_n1261 & ~new_n1262;
  assign new_n1269 = ~new_n1263 & ~new_n1268;
  assign new_n1270 = ~\a[111]  & ~\b[111] ;
  assign new_n1271 = \a[111]  & \b[111] ;
  assign new_n1272 = ~new_n1270 & ~new_n1271;
  assign new_n1273 = new_n1269 & ~new_n1272;
  assign new_n1274 = ~new_n1269 & new_n1272;
  assign \f[111]  = ~new_n1273 & ~new_n1274;
  assign new_n1276 = ~new_n1269 & ~new_n1270;
  assign new_n1277 = ~new_n1271 & ~new_n1276;
  assign new_n1278 = ~\a[112]  & ~\b[112] ;
  assign new_n1279 = \a[112]  & \b[112] ;
  assign new_n1280 = ~new_n1278 & ~new_n1279;
  assign new_n1281 = new_n1277 & ~new_n1280;
  assign new_n1282 = ~new_n1277 & new_n1280;
  assign \f[112]  = ~new_n1281 & ~new_n1282;
  assign new_n1284 = ~new_n1277 & ~new_n1278;
  assign new_n1285 = ~new_n1279 & ~new_n1284;
  assign new_n1286 = ~\a[113]  & ~\b[113] ;
  assign new_n1287 = \a[113]  & \b[113] ;
  assign new_n1288 = ~new_n1286 & ~new_n1287;
  assign new_n1289 = new_n1285 & ~new_n1288;
  assign new_n1290 = ~new_n1285 & new_n1288;
  assign \f[113]  = ~new_n1289 & ~new_n1290;
  assign new_n1292 = ~new_n1285 & ~new_n1286;
  assign new_n1293 = ~new_n1287 & ~new_n1292;
  assign new_n1294 = ~\a[114]  & ~\b[114] ;
  assign new_n1295 = \a[114]  & \b[114] ;
  assign new_n1296 = ~new_n1294 & ~new_n1295;
  assign new_n1297 = new_n1293 & ~new_n1296;
  assign new_n1298 = ~new_n1293 & new_n1296;
  assign \f[114]  = ~new_n1297 & ~new_n1298;
  assign new_n1300 = ~new_n1293 & ~new_n1294;
  assign new_n1301 = ~new_n1295 & ~new_n1300;
  assign new_n1302 = ~\a[115]  & ~\b[115] ;
  assign new_n1303 = \a[115]  & \b[115] ;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = new_n1301 & ~new_n1304;
  assign new_n1306 = ~new_n1301 & new_n1304;
  assign \f[115]  = ~new_n1305 & ~new_n1306;
  assign new_n1308 = ~new_n1301 & ~new_n1302;
  assign new_n1309 = ~new_n1303 & ~new_n1308;
  assign new_n1310 = ~\a[116]  & ~\b[116] ;
  assign new_n1311 = \a[116]  & \b[116] ;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = new_n1309 & ~new_n1312;
  assign new_n1314 = ~new_n1309 & new_n1312;
  assign \f[116]  = ~new_n1313 & ~new_n1314;
  assign new_n1316 = ~new_n1309 & ~new_n1310;
  assign new_n1317 = ~new_n1311 & ~new_n1316;
  assign new_n1318 = ~\a[117]  & ~\b[117] ;
  assign new_n1319 = \a[117]  & \b[117] ;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = new_n1317 & ~new_n1320;
  assign new_n1322 = ~new_n1317 & new_n1320;
  assign \f[117]  = ~new_n1321 & ~new_n1322;
  assign new_n1324 = ~new_n1317 & ~new_n1318;
  assign new_n1325 = ~new_n1319 & ~new_n1324;
  assign new_n1326 = ~\a[118]  & ~\b[118] ;
  assign new_n1327 = \a[118]  & \b[118] ;
  assign new_n1328 = ~new_n1326 & ~new_n1327;
  assign new_n1329 = new_n1325 & ~new_n1328;
  assign new_n1330 = ~new_n1325 & new_n1328;
  assign \f[118]  = ~new_n1329 & ~new_n1330;
  assign new_n1332 = ~new_n1325 & ~new_n1326;
  assign new_n1333 = ~new_n1327 & ~new_n1332;
  assign new_n1334 = ~\a[119]  & ~\b[119] ;
  assign new_n1335 = \a[119]  & \b[119] ;
  assign new_n1336 = ~new_n1334 & ~new_n1335;
  assign new_n1337 = new_n1333 & ~new_n1336;
  assign new_n1338 = ~new_n1333 & new_n1336;
  assign \f[119]  = ~new_n1337 & ~new_n1338;
  assign new_n1340 = ~new_n1333 & ~new_n1334;
  assign new_n1341 = ~new_n1335 & ~new_n1340;
  assign new_n1342 = ~\a[120]  & ~\b[120] ;
  assign new_n1343 = \a[120]  & \b[120] ;
  assign new_n1344 = ~new_n1342 & ~new_n1343;
  assign new_n1345 = new_n1341 & ~new_n1344;
  assign new_n1346 = ~new_n1341 & new_n1344;
  assign \f[120]  = ~new_n1345 & ~new_n1346;
  assign new_n1348 = ~new_n1341 & ~new_n1342;
  assign new_n1349 = ~new_n1343 & ~new_n1348;
  assign new_n1350 = ~\a[121]  & ~\b[121] ;
  assign new_n1351 = \a[121]  & \b[121] ;
  assign new_n1352 = ~new_n1350 & ~new_n1351;
  assign new_n1353 = new_n1349 & ~new_n1352;
  assign new_n1354 = ~new_n1349 & new_n1352;
  assign \f[121]  = ~new_n1353 & ~new_n1354;
  assign new_n1356 = ~new_n1349 & ~new_n1350;
  assign new_n1357 = ~new_n1351 & ~new_n1356;
  assign new_n1358 = ~\a[122]  & ~\b[122] ;
  assign new_n1359 = \a[122]  & \b[122] ;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = new_n1357 & ~new_n1360;
  assign new_n1362 = ~new_n1357 & new_n1360;
  assign \f[122]  = ~new_n1361 & ~new_n1362;
  assign new_n1364 = ~new_n1357 & ~new_n1358;
  assign new_n1365 = ~new_n1359 & ~new_n1364;
  assign new_n1366 = ~\a[123]  & ~\b[123] ;
  assign new_n1367 = \a[123]  & \b[123] ;
  assign new_n1368 = ~new_n1366 & ~new_n1367;
  assign new_n1369 = new_n1365 & ~new_n1368;
  assign new_n1370 = ~new_n1365 & new_n1368;
  assign \f[123]  = ~new_n1369 & ~new_n1370;
  assign new_n1372 = ~new_n1365 & ~new_n1366;
  assign new_n1373 = ~new_n1367 & ~new_n1372;
  assign new_n1374 = ~\a[124]  & ~\b[124] ;
  assign new_n1375 = \a[124]  & \b[124] ;
  assign new_n1376 = ~new_n1374 & ~new_n1375;
  assign new_n1377 = new_n1373 & ~new_n1376;
  assign new_n1378 = ~new_n1373 & new_n1376;
  assign \f[124]  = ~new_n1377 & ~new_n1378;
  assign new_n1380 = ~new_n1373 & ~new_n1374;
  assign new_n1381 = ~new_n1375 & ~new_n1380;
  assign new_n1382 = ~\a[125]  & ~\b[125] ;
  assign new_n1383 = \a[125]  & \b[125] ;
  assign new_n1384 = ~new_n1382 & ~new_n1383;
  assign new_n1385 = new_n1381 & ~new_n1384;
  assign new_n1386 = ~new_n1381 & new_n1384;
  assign \f[125]  = ~new_n1385 & ~new_n1386;
  assign new_n1388 = ~new_n1381 & ~new_n1382;
  assign new_n1389 = ~new_n1383 & ~new_n1388;
  assign new_n1390 = ~\a[126]  & ~\b[126] ;
  assign new_n1391 = \a[126]  & \b[126] ;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = new_n1389 & ~new_n1392;
  assign new_n1394 = ~new_n1389 & new_n1392;
  assign \f[126]  = ~new_n1393 & ~new_n1394;
  assign new_n1396 = ~new_n1389 & ~new_n1390;
  assign new_n1397 = ~new_n1391 & ~new_n1396;
  assign new_n1398 = ~\a[127]  & ~\b[127] ;
  assign new_n1399 = \a[127]  & \b[127] ;
  assign new_n1400 = ~new_n1398 & ~new_n1399;
  assign new_n1401 = new_n1397 & ~new_n1400;
  assign new_n1402 = ~new_n1397 & new_n1400;
  assign \f[127]  = ~new_n1401 & ~new_n1402;
  assign new_n1404 = ~new_n1397 & ~new_n1398;
  assign cOut = new_n1399 | new_n1404;
endmodule


