// Benchmark "top" written by ABC on Mon Dec 25 17:56:53 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1750,
    new_n1751, new_n1752, new_n1753, new_n1754, new_n1755, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1830, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1837, new_n1838, new_n1839, new_n1840,
    new_n1841, new_n1842, new_n1843, new_n1844, new_n1845, new_n1846,
    new_n1847, new_n1848, new_n1849, new_n1850, new_n1851, new_n1852,
    new_n1853, new_n1854, new_n1855, new_n1856, new_n1857, new_n1858,
    new_n1859, new_n1860, new_n1861, new_n1862, new_n1863, new_n1864,
    new_n1865, new_n1866, new_n1867, new_n1868, new_n1869, new_n1870,
    new_n1871, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979,
    new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978, new_n2979, new_n2980, new_n2981,
    new_n2982, new_n2983, new_n2984, new_n2985, new_n2986, new_n2987,
    new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993,
    new_n2994, new_n2995, new_n2996, new_n2997, new_n2998, new_n2999,
    new_n3000, new_n3001, new_n3002, new_n3003, new_n3004, new_n3005,
    new_n3006, new_n3007, new_n3008, new_n3009, new_n3010, new_n3011,
    new_n3012, new_n3013, new_n3014, new_n3015, new_n3016, new_n3017,
    new_n3018, new_n3019, new_n3020, new_n3021, new_n3022, new_n3023,
    new_n3024, new_n3025, new_n3026, new_n3027, new_n3028, new_n3029,
    new_n3030, new_n3031, new_n3032, new_n3033, new_n3034, new_n3035,
    new_n3036, new_n3037, new_n3038, new_n3039, new_n3040, new_n3041,
    new_n3042, new_n3043, new_n3044, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3228, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055,
    new_n4056, new_n4057, new_n4058, new_n4059, new_n4060, new_n4061,
    new_n4062, new_n4063, new_n4064, new_n4065, new_n4066, new_n4067,
    new_n4068, new_n4069, new_n4070, new_n4071, new_n4072, new_n4073,
    new_n4074, new_n4075, new_n4076, new_n4077, new_n4078, new_n4079,
    new_n4080, new_n4081, new_n4082, new_n4083, new_n4084, new_n4085,
    new_n4086, new_n4087, new_n4088, new_n4089, new_n4090, new_n4091,
    new_n4092, new_n4093, new_n4094, new_n4095, new_n4096, new_n4097,
    new_n4098, new_n4099, new_n4100, new_n4101, new_n4102, new_n4103,
    new_n4104, new_n4105, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119, new_n4120, new_n4121,
    new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187,
    new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211,
    new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4482, new_n4483,
    new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489,
    new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495,
    new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588, new_n4589, new_n4590, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659, new_n4660, new_n4661, new_n4662, new_n4663,
    new_n4664, new_n4665, new_n4666, new_n4667, new_n4668, new_n4669,
    new_n4670, new_n4671, new_n4672, new_n4673, new_n4674, new_n4675,
    new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687,
    new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693,
    new_n4694, new_n4695, new_n4696, new_n4697, new_n4698, new_n4699,
    new_n4700, new_n4701, new_n4702, new_n4703, new_n4704, new_n4705,
    new_n4706, new_n4707, new_n4708, new_n4709, new_n4710, new_n4711,
    new_n4712, new_n4713, new_n4714, new_n4715, new_n4716, new_n4717,
    new_n4718, new_n4719, new_n4720, new_n4721, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766,
    new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772,
    new_n4773, new_n4774, new_n4775, new_n4776, new_n4777, new_n4778,
    new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784,
    new_n4785, new_n4786, new_n4787, new_n4788, new_n4789, new_n4790,
    new_n4791, new_n4792, new_n4793, new_n4794, new_n4795, new_n4796,
    new_n4797, new_n4798, new_n4799, new_n4800, new_n4801, new_n4802,
    new_n4803, new_n4804, new_n4805, new_n4806, new_n4807, new_n4808,
    new_n4809, new_n4810, new_n4811, new_n4812, new_n4813, new_n4814,
    new_n4815, new_n4816, new_n4817, new_n4818, new_n4819, new_n4820,
    new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826,
    new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031,
    new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5443, new_n5444, new_n5445, new_n5446, new_n5447,
    new_n5448, new_n5449, new_n5450, new_n5451, new_n5452, new_n5453,
    new_n5454, new_n5455, new_n5456, new_n5457, new_n5458, new_n5459,
    new_n5460, new_n5461, new_n5462, new_n5463, new_n5464, new_n5465,
    new_n5466, new_n5467, new_n5468, new_n5469, new_n5470, new_n5471,
    new_n5472, new_n5473, new_n5474, new_n5475, new_n5476, new_n5477,
    new_n5478, new_n5479, new_n5480, new_n5481, new_n5482, new_n5483,
    new_n5484, new_n5485, new_n5486, new_n5487, new_n5488, new_n5489,
    new_n5490, new_n5491, new_n5492, new_n5493, new_n5494, new_n5495,
    new_n5496, new_n5497, new_n5498, new_n5499, new_n5500, new_n5501,
    new_n5502, new_n5503, new_n5504, new_n5505, new_n5506, new_n5507,
    new_n5508, new_n5509, new_n5510, new_n5511, new_n5512, new_n5513,
    new_n5514, new_n5515, new_n5516, new_n5517, new_n5518, new_n5519,
    new_n5520, new_n5521, new_n5522, new_n5523, new_n5524, new_n5525,
    new_n5526, new_n5527, new_n5528, new_n5529, new_n5530, new_n5531,
    new_n5532, new_n5533, new_n5534, new_n5535, new_n5536, new_n5537,
    new_n5538, new_n5539, new_n5540, new_n5541, new_n5542, new_n5543,
    new_n5544, new_n5545, new_n5546, new_n5547, new_n5548, new_n5549,
    new_n5550, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555,
    new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561,
    new_n5562, new_n5563, new_n5564, new_n5565, new_n5566, new_n5567,
    new_n5568, new_n5569, new_n5570, new_n5571, new_n5572, new_n5573,
    new_n5574, new_n5575, new_n5576, new_n5577, new_n5578, new_n5579,
    new_n5580, new_n5581, new_n5582, new_n5583, new_n5584, new_n5585,
    new_n5586, new_n5587, new_n5588, new_n5589, new_n5590, new_n5591,
    new_n5592, new_n5593, new_n5594, new_n5595, new_n5596, new_n5597,
    new_n5598, new_n5599, new_n5600, new_n5601, new_n5602, new_n5603,
    new_n5604, new_n5605, new_n5606, new_n5607, new_n5608, new_n5609,
    new_n5610, new_n5611, new_n5612, new_n5613, new_n5614, new_n5615,
    new_n5616, new_n5617, new_n5618, new_n5619, new_n5620, new_n5621,
    new_n5622, new_n5623, new_n5624, new_n5625, new_n5626, new_n5627,
    new_n5628, new_n5629, new_n5630, new_n5631, new_n5632, new_n5633,
    new_n5634, new_n5635, new_n5636, new_n5637, new_n5638, new_n5639,
    new_n5640, new_n5641, new_n5642, new_n5643, new_n5644, new_n5645,
    new_n5646, new_n5647, new_n5648, new_n5649, new_n5650, new_n5651,
    new_n5652, new_n5653, new_n5654, new_n5655, new_n5656, new_n5657,
    new_n5658, new_n5659, new_n5660, new_n5661, new_n5662, new_n5663,
    new_n5664, new_n5665, new_n5666, new_n5667, new_n5668, new_n5669,
    new_n5670, new_n5671, new_n5672, new_n5673, new_n5674, new_n5675,
    new_n5676, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5947,
    new_n5948, new_n5949, new_n5950, new_n5951, new_n5952, new_n5953,
    new_n5954, new_n5955, new_n5956, new_n5957, new_n5958, new_n5959,
    new_n5960, new_n5961, new_n5962, new_n5963, new_n5964, new_n5965,
    new_n5966, new_n5967, new_n5968, new_n5969, new_n5970, new_n5971,
    new_n5972, new_n5973, new_n5974, new_n5975, new_n5976, new_n5977,
    new_n5978, new_n5979, new_n5980, new_n5981, new_n5982, new_n5983,
    new_n5984, new_n5985, new_n5986, new_n5987, new_n5988, new_n5989,
    new_n5990, new_n5991, new_n5992, new_n5993, new_n5994, new_n5995,
    new_n5996, new_n5997, new_n5998, new_n5999, new_n6000, new_n6001,
    new_n6002, new_n6003, new_n6004, new_n6005, new_n6006, new_n6007,
    new_n6008, new_n6009, new_n6010, new_n6011, new_n6012, new_n6013,
    new_n6014, new_n6015, new_n6016, new_n6017, new_n6018, new_n6019,
    new_n6020, new_n6021, new_n6022, new_n6023, new_n6024, new_n6025,
    new_n6026, new_n6027, new_n6028, new_n6029, new_n6030, new_n6031,
    new_n6032, new_n6033, new_n6034, new_n6035, new_n6036, new_n6037,
    new_n6038, new_n6039, new_n6040, new_n6041, new_n6042, new_n6043,
    new_n6044, new_n6045, new_n6046, new_n6047, new_n6048, new_n6049,
    new_n6050, new_n6051, new_n6052, new_n6053, new_n6054, new_n6055,
    new_n6056, new_n6057, new_n6058, new_n6059, new_n6060, new_n6061,
    new_n6062, new_n6063, new_n6064, new_n6065, new_n6066, new_n6067,
    new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073,
    new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079,
    new_n6080, new_n6081, new_n6082, new_n6083, new_n6084, new_n6085,
    new_n6086, new_n6087, new_n6088, new_n6089, new_n6090, new_n6091,
    new_n6092, new_n6093, new_n6094, new_n6095, new_n6096, new_n6097,
    new_n6098, new_n6099, new_n6100, new_n6101, new_n6102, new_n6103,
    new_n6104, new_n6105, new_n6106, new_n6107, new_n6108, new_n6109,
    new_n6110, new_n6111, new_n6112, new_n6113, new_n6114, new_n6115,
    new_n6116, new_n6117, new_n6118, new_n6119, new_n6120, new_n6121,
    new_n6122, new_n6123, new_n6124, new_n6125, new_n6126, new_n6127,
    new_n6128, new_n6129, new_n6130, new_n6131, new_n6132, new_n6133,
    new_n6134, new_n6135, new_n6136, new_n6137, new_n6138, new_n6139,
    new_n6140, new_n6141, new_n6142, new_n6143, new_n6144, new_n6145,
    new_n6146, new_n6147, new_n6148, new_n6149, new_n6150, new_n6151,
    new_n6152, new_n6153, new_n6154, new_n6155, new_n6156, new_n6157,
    new_n6158, new_n6159, new_n6160, new_n6161, new_n6162, new_n6163,
    new_n6164, new_n6165, new_n6166, new_n6167, new_n6168, new_n6169,
    new_n6170, new_n6171, new_n6172, new_n6173, new_n6174, new_n6175,
    new_n6176, new_n6177, new_n6178, new_n6179, new_n6180, new_n6181,
    new_n6182, new_n6183, new_n6184, new_n6185, new_n6186, new_n6187,
    new_n6188, new_n6189, new_n6190, new_n6191, new_n6192, new_n6193,
    new_n6194, new_n6195, new_n6196, new_n6197, new_n6198, new_n6199,
    new_n6200, new_n6201, new_n6202, new_n6203, new_n6204, new_n6205,
    new_n6206, new_n6207, new_n6208, new_n6209, new_n6210, new_n6211,
    new_n6212, new_n6213, new_n6214, new_n6216, new_n6217, new_n6218,
    new_n6219, new_n6220, new_n6221, new_n6222, new_n6223, new_n6224,
    new_n6225, new_n6226, new_n6227, new_n6228, new_n6229, new_n6230,
    new_n6231, new_n6232, new_n6233, new_n6234, new_n6235, new_n6236,
    new_n6237, new_n6238, new_n6239, new_n6240, new_n6241, new_n6242,
    new_n6243, new_n6244, new_n6245, new_n6246, new_n6247, new_n6248,
    new_n6249, new_n6250, new_n6251, new_n6252, new_n6253, new_n6254,
    new_n6255, new_n6256, new_n6257, new_n6258, new_n6259, new_n6260,
    new_n6261, new_n6262, new_n6263, new_n6264, new_n6265, new_n6266,
    new_n6267, new_n6268, new_n6269, new_n6270, new_n6271, new_n6272,
    new_n6273, new_n6274, new_n6275, new_n6276, new_n6277, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284,
    new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290,
    new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296,
    new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302,
    new_n6303, new_n6304, new_n6305, new_n6306, new_n6307, new_n6308,
    new_n6309, new_n6310, new_n6311, new_n6312, new_n6313, new_n6314,
    new_n6315, new_n6316, new_n6317, new_n6318, new_n6319, new_n6320,
    new_n6321, new_n6322, new_n6323, new_n6324, new_n6325, new_n6326,
    new_n6327, new_n6328, new_n6329, new_n6330, new_n6331, new_n6332,
    new_n6333, new_n6334, new_n6335, new_n6336, new_n6337, new_n6338,
    new_n6339, new_n6340, new_n6341, new_n6342, new_n6343, new_n6344,
    new_n6345, new_n6346, new_n6347, new_n6348, new_n6349, new_n6350,
    new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356,
    new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362,
    new_n6363, new_n6364, new_n6365, new_n6366, new_n6367, new_n6368,
    new_n6369, new_n6370, new_n6371, new_n6372, new_n6373, new_n6374,
    new_n6375, new_n6376, new_n6377, new_n6378, new_n6379, new_n6380,
    new_n6381, new_n6382, new_n6383, new_n6384, new_n6385, new_n6386,
    new_n6387, new_n6388, new_n6389, new_n6390, new_n6391, new_n6392,
    new_n6393, new_n6394, new_n6395, new_n6396, new_n6397, new_n6398,
    new_n6399, new_n6400, new_n6401, new_n6402, new_n6403, new_n6404,
    new_n6405, new_n6406, new_n6407, new_n6408, new_n6409, new_n6410,
    new_n6411, new_n6412, new_n6413, new_n6414, new_n6415, new_n6416,
    new_n6417, new_n6418, new_n6419, new_n6420, new_n6421, new_n6422,
    new_n6423, new_n6424, new_n6425, new_n6426, new_n6427, new_n6428,
    new_n6429, new_n6430, new_n6431, new_n6432, new_n6433, new_n6434,
    new_n6435, new_n6436, new_n6437, new_n6438, new_n6439, new_n6440,
    new_n6441, new_n6442, new_n6443, new_n6444, new_n6445, new_n6446,
    new_n6447, new_n6448, new_n6449, new_n6450, new_n6451, new_n6452,
    new_n6453, new_n6454, new_n6455, new_n6456, new_n6457, new_n6458,
    new_n6459, new_n6460, new_n6461, new_n6462, new_n6463, new_n6464,
    new_n6465, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470,
    new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476,
    new_n6477, new_n6478, new_n6479, new_n6480, new_n6481, new_n6482,
    new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488,
    new_n6489, new_n6490, new_n6491, new_n6493, new_n6494, new_n6495,
    new_n6496, new_n6497, new_n6498, new_n6499, new_n6500, new_n6501,
    new_n6502, new_n6503, new_n6504, new_n6505, new_n6506, new_n6507,
    new_n6508, new_n6509, new_n6510, new_n6511, new_n6512, new_n6513,
    new_n6514, new_n6515, new_n6516, new_n6517, new_n6518, new_n6519,
    new_n6520, new_n6521, new_n6522, new_n6523, new_n6524, new_n6525,
    new_n6526, new_n6527, new_n6528, new_n6529, new_n6530, new_n6531,
    new_n6532, new_n6533, new_n6534, new_n6535, new_n6536, new_n6537,
    new_n6538, new_n6539, new_n6540, new_n6541, new_n6542, new_n6543,
    new_n6544, new_n6545, new_n6546, new_n6547, new_n6548, new_n6549,
    new_n6550, new_n6551, new_n6552, new_n6553, new_n6554, new_n6555,
    new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561,
    new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790,
    new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814,
    new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820,
    new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826,
    new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832,
    new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838,
    new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844,
    new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850,
    new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856,
    new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862,
    new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868,
    new_n6869, new_n6870, new_n6871, new_n6872, new_n6873, new_n6874,
    new_n6875, new_n6876, new_n6877, new_n6878, new_n6879, new_n6880,
    new_n6881, new_n6882, new_n6883, new_n6884, new_n6885, new_n6886,
    new_n6887, new_n6888, new_n6889, new_n6890, new_n6891, new_n6892,
    new_n6893, new_n6894, new_n6895, new_n6896, new_n6897, new_n6898,
    new_n6899, new_n6900, new_n6901, new_n6902, new_n6903, new_n6904,
    new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910,
    new_n6911, new_n6912, new_n6913, new_n6914, new_n6915, new_n6916,
    new_n6917, new_n6918, new_n6919, new_n6920, new_n6921, new_n6922,
    new_n6923, new_n6924, new_n6925, new_n6926, new_n6927, new_n6928,
    new_n6929, new_n6930, new_n6931, new_n6932, new_n6933, new_n6934,
    new_n6935, new_n6936, new_n6937, new_n6938, new_n6939, new_n6940,
    new_n6941, new_n6942, new_n6943, new_n6944, new_n6945, new_n6946,
    new_n6947, new_n6948, new_n6949, new_n6950, new_n6951, new_n6952,
    new_n6953, new_n6954, new_n6955, new_n6956, new_n6957, new_n6958,
    new_n6959, new_n6960, new_n6961, new_n6962, new_n6963, new_n6964,
    new_n6965, new_n6966, new_n6967, new_n6968, new_n6969, new_n6970,
    new_n6971, new_n6972, new_n6973, new_n6974, new_n6975, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983, new_n6984, new_n6985, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7618, new_n7619, new_n7620, new_n7621,
    new_n7622, new_n7623, new_n7624, new_n7625, new_n7626, new_n7627,
    new_n7628, new_n7629, new_n7630, new_n7631, new_n7632, new_n7633,
    new_n7634, new_n7635, new_n7636, new_n7637, new_n7638, new_n7639,
    new_n7640, new_n7641, new_n7642, new_n7643, new_n7644, new_n7645,
    new_n7646, new_n7647, new_n7648, new_n7649, new_n7650, new_n7651,
    new_n7652, new_n7653, new_n7654, new_n7655, new_n7656, new_n7657,
    new_n7658, new_n7659, new_n7660, new_n7661, new_n7662, new_n7663,
    new_n7664, new_n7665, new_n7666, new_n7667, new_n7668, new_n7669,
    new_n7670, new_n7671, new_n7672, new_n7673, new_n7674, new_n7675,
    new_n7676, new_n7677, new_n7678, new_n7679, new_n7680, new_n7681,
    new_n7682, new_n7683, new_n7684, new_n7685, new_n7686, new_n7687,
    new_n7688, new_n7689, new_n7690, new_n7691, new_n7692, new_n7693,
    new_n7694, new_n7695, new_n7696, new_n7697, new_n7698, new_n7699,
    new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705,
    new_n7706, new_n7707, new_n7708, new_n7709, new_n7710, new_n7711,
    new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729,
    new_n7730, new_n7731, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741,
    new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747,
    new_n7748, new_n7749, new_n7750, new_n7751, new_n7752, new_n7753,
    new_n7754, new_n7755, new_n7756, new_n7757, new_n7758, new_n7759,
    new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765,
    new_n7766, new_n7767, new_n7768, new_n7769, new_n7770, new_n7771,
    new_n7772, new_n7773, new_n7774, new_n7775, new_n7776, new_n7777,
    new_n7778, new_n7779, new_n7780, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794, new_n7795,
    new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801,
    new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807,
    new_n7808, new_n7809, new_n7810, new_n7811, new_n7812, new_n7813,
    new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819,
    new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825,
    new_n7826, new_n7827, new_n7828, new_n7829, new_n7830, new_n7831,
    new_n7832, new_n7833, new_n7834, new_n7835, new_n7836, new_n7837,
    new_n7838, new_n7839, new_n7840, new_n7841, new_n7842, new_n7843,
    new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849,
    new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867,
    new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873,
    new_n7874, new_n7875, new_n7876, new_n7877, new_n7878, new_n7879,
    new_n7880, new_n7881, new_n7882, new_n7883, new_n7884, new_n7885,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8246, new_n8247,
    new_n8248, new_n8249, new_n8250, new_n8251, new_n8252, new_n8253,
    new_n8254, new_n8255, new_n8256, new_n8257, new_n8258, new_n8259,
    new_n8260, new_n8261, new_n8262, new_n8263, new_n8264, new_n8265,
    new_n8266, new_n8267, new_n8268, new_n8269, new_n8270, new_n8271,
    new_n8272, new_n8273, new_n8274, new_n8275, new_n8276, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285, new_n8286, new_n8287, new_n8288, new_n8289,
    new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295,
    new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301,
    new_n8302, new_n8303, new_n8304, new_n8305, new_n8306, new_n8307,
    new_n8308, new_n8309, new_n8310, new_n8311, new_n8312, new_n8313,
    new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319,
    new_n8320, new_n8321, new_n8322, new_n8323, new_n8324, new_n8325,
    new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331,
    new_n8332, new_n8333, new_n8334, new_n8335, new_n8336, new_n8337,
    new_n8338, new_n8339, new_n8340, new_n8341, new_n8342, new_n8343,
    new_n8344, new_n8345, new_n8346, new_n8347, new_n8348, new_n8349,
    new_n8350, new_n8351, new_n8352, new_n8353, new_n8354, new_n8355,
    new_n8356, new_n8357, new_n8358, new_n8359, new_n8360, new_n8361,
    new_n8362, new_n8363, new_n8364, new_n8365, new_n8366, new_n8367,
    new_n8368, new_n8369, new_n8370, new_n8371, new_n8372, new_n8373,
    new_n8374, new_n8375, new_n8376, new_n8377, new_n8378, new_n8379,
    new_n8380, new_n8381, new_n8382, new_n8383, new_n8384, new_n8385,
    new_n8386, new_n8387, new_n8388, new_n8389, new_n8390, new_n8391,
    new_n8392, new_n8393, new_n8394, new_n8395, new_n8396, new_n8397,
    new_n8398, new_n8399, new_n8400, new_n8401, new_n8402, new_n8403,
    new_n8404, new_n8405, new_n8406, new_n8407, new_n8408, new_n8409,
    new_n8410, new_n8411, new_n8412, new_n8413, new_n8414, new_n8415,
    new_n8416, new_n8417, new_n8418, new_n8419, new_n8420, new_n8421,
    new_n8422, new_n8423, new_n8424, new_n8425, new_n8426, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432, new_n8433,
    new_n8434, new_n8435, new_n8436, new_n8437, new_n8438, new_n8439,
    new_n8440, new_n8441, new_n8442, new_n8443, new_n8444, new_n8445,
    new_n8446, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451,
    new_n8452, new_n8453, new_n8454, new_n8455, new_n8456, new_n8457,
    new_n8458, new_n8459, new_n8460, new_n8461, new_n8462, new_n8463,
    new_n8464, new_n8465, new_n8466, new_n8467, new_n8468, new_n8469,
    new_n8470, new_n8471, new_n8472, new_n8473, new_n8474, new_n8475,
    new_n8476, new_n8477, new_n8478, new_n8479, new_n8480, new_n8481,
    new_n8482, new_n8483, new_n8484, new_n8485, new_n8486, new_n8487,
    new_n8488, new_n8489, new_n8490, new_n8491, new_n8492, new_n8493,
    new_n8494, new_n8495, new_n8496, new_n8497, new_n8498, new_n8499,
    new_n8500, new_n8501, new_n8502, new_n8503, new_n8504, new_n8505,
    new_n8506, new_n8507, new_n8508, new_n8509, new_n8510, new_n8511,
    new_n8512, new_n8513, new_n8514, new_n8515, new_n8516, new_n8517,
    new_n8518, new_n8519, new_n8520, new_n8521, new_n8522, new_n8523,
    new_n8524, new_n8525, new_n8526, new_n8527, new_n8528, new_n8529,
    new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535,
    new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541,
    new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547,
    new_n8548, new_n8549, new_n8550, new_n8551, new_n8552, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8566,
    new_n8567, new_n8568, new_n8569, new_n8570, new_n8571, new_n8572,
    new_n8573, new_n8574, new_n8575, new_n8576, new_n8577, new_n8578,
    new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584,
    new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590,
    new_n8591, new_n8592, new_n8593, new_n8594, new_n8595, new_n8596,
    new_n8597, new_n8598, new_n8599, new_n8600, new_n8601, new_n8602,
    new_n8603, new_n8604, new_n8605, new_n8606, new_n8607, new_n8608,
    new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614,
    new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620,
    new_n8621, new_n8622, new_n8623, new_n8624, new_n8625, new_n8626,
    new_n8627, new_n8628, new_n8629, new_n8630, new_n8631, new_n8632,
    new_n8633, new_n8634, new_n8635, new_n8636, new_n8637, new_n8638,
    new_n8639, new_n8640, new_n8641, new_n8642, new_n8643, new_n8644,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716,
    new_n8717, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803, new_n8804, new_n8805, new_n8806,
    new_n8807, new_n8808, new_n8809, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821, new_n8822, new_n8823, new_n8824,
    new_n8825, new_n8826, new_n8827, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861, new_n8862, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939,
    new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945,
    new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951,
    new_n8952, new_n8953, new_n8954, new_n8955, new_n8956, new_n8957,
    new_n8958, new_n8959, new_n8960, new_n8961, new_n8962, new_n8963,
    new_n8964, new_n8965, new_n8966, new_n8967, new_n8968, new_n8969,
    new_n8970, new_n8971, new_n8972, new_n8973, new_n8974, new_n8975,
    new_n8976, new_n8977, new_n8978, new_n8979, new_n8980, new_n8981,
    new_n8982, new_n8983, new_n8984, new_n8985, new_n8986, new_n8987,
    new_n8988, new_n8989, new_n8990, new_n8991, new_n8992, new_n8993,
    new_n8994, new_n8995, new_n8996, new_n8997, new_n8998, new_n8999,
    new_n9000, new_n9001, new_n9002, new_n9003, new_n9004, new_n9005,
    new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011,
    new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017,
    new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023,
    new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077,
    new_n9078, new_n9079, new_n9080, new_n9081, new_n9082, new_n9083,
    new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089,
    new_n9090, new_n9091, new_n9092, new_n9093, new_n9094, new_n9095,
    new_n9096, new_n9097, new_n9098, new_n9099, new_n9100, new_n9101,
    new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107,
    new_n9108, new_n9109, new_n9110, new_n9111, new_n9112, new_n9113,
    new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119,
    new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125,
    new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131,
    new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137,
    new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143,
    new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149,
    new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155,
    new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161,
    new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167,
    new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173,
    new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179,
    new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185,
    new_n9186, new_n9187, new_n9188, new_n9189, new_n9190, new_n9191,
    new_n9192, new_n9193, new_n9194, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9532, new_n9533, new_n9534, new_n9535,
    new_n9536, new_n9537, new_n9538, new_n9539, new_n9540, new_n9541,
    new_n9542, new_n9543, new_n9544, new_n9545, new_n9546, new_n9547,
    new_n9548, new_n9549, new_n9550, new_n9551, new_n9552, new_n9553,
    new_n9554, new_n9555, new_n9556, new_n9557, new_n9558, new_n9559,
    new_n9560, new_n9561, new_n9562, new_n9563, new_n9564, new_n9565,
    new_n9566, new_n9567, new_n9568, new_n9569, new_n9570, new_n9571,
    new_n9572, new_n9573, new_n9574, new_n9575, new_n9576, new_n9577,
    new_n9578, new_n9579, new_n9580, new_n9581, new_n9582, new_n9583,
    new_n9584, new_n9585, new_n9586, new_n9587, new_n9588, new_n9589,
    new_n9590, new_n9591, new_n9592, new_n9593, new_n9594, new_n9595,
    new_n9596, new_n9597, new_n9598, new_n9599, new_n9600, new_n9601,
    new_n9602, new_n9603, new_n9604, new_n9605, new_n9606, new_n9607,
    new_n9608, new_n9609, new_n9610, new_n9611, new_n9612, new_n9613,
    new_n9614, new_n9615, new_n9616, new_n9617, new_n9618, new_n9619,
    new_n9620, new_n9621, new_n9622, new_n9623, new_n9624, new_n9625,
    new_n9626, new_n9627, new_n9628, new_n9629, new_n9630, new_n9631,
    new_n9632, new_n9633, new_n9634, new_n9635, new_n9636, new_n9637,
    new_n9638, new_n9639, new_n9640, new_n9641, new_n9642, new_n9643,
    new_n9644, new_n9645, new_n9646, new_n9647, new_n9648, new_n9649,
    new_n9650, new_n9651, new_n9652, new_n9653, new_n9654, new_n9655,
    new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661,
    new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667,
    new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673,
    new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679,
    new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685,
    new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691,
    new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697,
    new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763,
    new_n9764, new_n9765, new_n9766, new_n9767, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820, new_n9821, new_n9822, new_n9823,
    new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829,
    new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917, new_n9918, new_n9919, new_n9920,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934, new_n9935, new_n9936, new_n9937, new_n9938,
    new_n9939, new_n9940, new_n9941, new_n9942, new_n9943, new_n9944,
    new_n9945, new_n9946, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967, new_n9968,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9987, new_n9988, new_n9989, new_n9990, new_n9991, new_n9992,
    new_n9993, new_n9994, new_n9995, new_n9996, new_n9997, new_n9998,
    new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004,
    new_n10005, new_n10006, new_n10007, new_n10008, new_n10009, new_n10010,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017, new_n10018, new_n10019, new_n10020, new_n10021, new_n10022,
    new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053, new_n10054, new_n10055, new_n10056, new_n10057, new_n10058,
    new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064,
    new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070,
    new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076,
    new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10096, new_n10097, new_n10098, new_n10099, new_n10100,
    new_n10101, new_n10102, new_n10103, new_n10104, new_n10105, new_n10106,
    new_n10107, new_n10108, new_n10109, new_n10110, new_n10111, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130,
    new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136,
    new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148,
    new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10156, new_n10157, new_n10158, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165, new_n10166,
    new_n10167, new_n10168, new_n10169, new_n10170, new_n10171, new_n10172,
    new_n10173, new_n10174, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197,
    new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10321, new_n10322, new_n10323,
    new_n10324, new_n10325, new_n10326, new_n10327, new_n10328, new_n10329,
    new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335,
    new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443,
    new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449,
    new_n10450, new_n10451, new_n10452, new_n10453, new_n10454, new_n10455,
    new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461,
    new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467,
    new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473,
    new_n10474, new_n10475, new_n10476, new_n10477, new_n10478, new_n10479,
    new_n10480, new_n10481, new_n10482, new_n10483, new_n10484, new_n10485,
    new_n10486, new_n10487, new_n10488, new_n10489, new_n10490, new_n10491,
    new_n10492, new_n10493, new_n10494, new_n10495, new_n10496, new_n10497,
    new_n10498, new_n10499, new_n10500, new_n10501, new_n10502, new_n10503,
    new_n10504, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540,
    new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546,
    new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582,
    new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593, new_n10594,
    new_n10595, new_n10596, new_n10597, new_n10598, new_n10599, new_n10600,
    new_n10601, new_n10602, new_n10603, new_n10604, new_n10605, new_n10606,
    new_n10607, new_n10608, new_n10609, new_n10610, new_n10611, new_n10612,
    new_n10613, new_n10614, new_n10615, new_n10616, new_n10617, new_n10618,
    new_n10619, new_n10620, new_n10621, new_n10622, new_n10623, new_n10624,
    new_n10625, new_n10626, new_n10627, new_n10628, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678,
    new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10684,
    new_n10685, new_n10686, new_n10687, new_n10688, new_n10689, new_n10690,
    new_n10691, new_n10692, new_n10693, new_n10694, new_n10695, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10877,
    new_n10878, new_n10879, new_n10880, new_n10881, new_n10882, new_n10883,
    new_n10884, new_n10885, new_n10886, new_n10887, new_n10888, new_n10889,
    new_n10890, new_n10891, new_n10892, new_n10893, new_n10894, new_n10895,
    new_n10896, new_n10897, new_n10898, new_n10899, new_n10900, new_n10901,
    new_n10902, new_n10903, new_n10904, new_n10905, new_n10906, new_n10907,
    new_n10908, new_n10909, new_n10910, new_n10911, new_n10912, new_n10913,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928, new_n10929, new_n10930, new_n10931,
    new_n10932, new_n10933, new_n10934, new_n10935, new_n10936, new_n10937,
    new_n10938, new_n10939, new_n10940, new_n10941, new_n10942, new_n10943,
    new_n10944, new_n10945, new_n10946, new_n10947, new_n10948, new_n10949,
    new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955,
    new_n10956, new_n10957, new_n10958, new_n10959, new_n10960, new_n10961,
    new_n10962, new_n10963, new_n10964, new_n10965, new_n10966, new_n10967,
    new_n10968, new_n10969, new_n10970, new_n10971, new_n10972, new_n10973,
    new_n10974, new_n10975, new_n10976, new_n10977, new_n10978, new_n10979,
    new_n10980, new_n10981, new_n10982, new_n10983, new_n10984, new_n10985,
    new_n10986, new_n10987, new_n10988, new_n10989, new_n10990, new_n10991,
    new_n10992, new_n10993, new_n10994, new_n10995, new_n10996, new_n10997,
    new_n10998, new_n10999, new_n11000, new_n11001, new_n11002, new_n11003,
    new_n11004, new_n11005, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011, new_n11012, new_n11013, new_n11014, new_n11015,
    new_n11016, new_n11017, new_n11018, new_n11019, new_n11020, new_n11021,
    new_n11022, new_n11023, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057,
    new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063,
    new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099,
    new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135,
    new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141,
    new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11153,
    new_n11154, new_n11155, new_n11156, new_n11157, new_n11158, new_n11159,
    new_n11160, new_n11161, new_n11162, new_n11163, new_n11164, new_n11165,
    new_n11166, new_n11167, new_n11168, new_n11169, new_n11170, new_n11171,
    new_n11172, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177,
    new_n11178, new_n11179, new_n11180, new_n11181, new_n11182, new_n11183,
    new_n11184, new_n11185, new_n11186, new_n11187, new_n11188, new_n11189,
    new_n11190, new_n11191, new_n11192, new_n11193, new_n11194, new_n11195,
    new_n11196, new_n11197, new_n11198, new_n11199, new_n11200, new_n11201,
    new_n11202, new_n11203, new_n11204, new_n11205, new_n11206, new_n11207,
    new_n11208, new_n11209, new_n11210, new_n11211, new_n11212, new_n11213,
    new_n11214, new_n11215, new_n11216, new_n11217, new_n11218, new_n11220,
    new_n11221, new_n11222, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257, new_n11258, new_n11259, new_n11260, new_n11261, new_n11262,
    new_n11263, new_n11264, new_n11265, new_n11266, new_n11267, new_n11268,
    new_n11269, new_n11270, new_n11271, new_n11272, new_n11273, new_n11274,
    new_n11275, new_n11276, new_n11277, new_n11278, new_n11279, new_n11280,
    new_n11281, new_n11282, new_n11283, new_n11284, new_n11285, new_n11286,
    new_n11287, new_n11288, new_n11289, new_n11290, new_n11291, new_n11292,
    new_n11293, new_n11294, new_n11295, new_n11296, new_n11297, new_n11298,
    new_n11299, new_n11300, new_n11301, new_n11302, new_n11303, new_n11304,
    new_n11305, new_n11306, new_n11307, new_n11308, new_n11309, new_n11310,
    new_n11311, new_n11312, new_n11313, new_n11314, new_n11315, new_n11316,
    new_n11317, new_n11318, new_n11319, new_n11320, new_n11321, new_n11322,
    new_n11323, new_n11324, new_n11325, new_n11326, new_n11327, new_n11328,
    new_n11329, new_n11330, new_n11331, new_n11332, new_n11333, new_n11334,
    new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347, new_n11348, new_n11349, new_n11350, new_n11351, new_n11352,
    new_n11353, new_n11354, new_n11355, new_n11356, new_n11357, new_n11358,
    new_n11359, new_n11360, new_n11361, new_n11362, new_n11363, new_n11364,
    new_n11365, new_n11366, new_n11367, new_n11368, new_n11369, new_n11370,
    new_n11371, new_n11372, new_n11373, new_n11374, new_n11375, new_n11376,
    new_n11377, new_n11378, new_n11379, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386, new_n11387, new_n11388,
    new_n11389, new_n11390, new_n11391, new_n11392, new_n11393, new_n11394,
    new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478,
    new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490,
    new_n11491, new_n11492, new_n11493, new_n11494, new_n11495, new_n11496,
    new_n11497, new_n11498, new_n11499, new_n11500, new_n11501, new_n11502,
    new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508,
    new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514,
    new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520,
    new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526,
    new_n11527, new_n11528, new_n11529, new_n11530, new_n11531, new_n11532,
    new_n11533, new_n11534, new_n11535, new_n11536, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574,
    new_n11576, new_n11577, new_n11578, new_n11579, new_n11580, new_n11581,
    new_n11582, new_n11583, new_n11584, new_n11585, new_n11586, new_n11587,
    new_n11588, new_n11589, new_n11590, new_n11591, new_n11592, new_n11593,
    new_n11594, new_n11595, new_n11596, new_n11597, new_n11598, new_n11599,
    new_n11600, new_n11601, new_n11602, new_n11603, new_n11604, new_n11605,
    new_n11606, new_n11607, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11615, new_n11616, new_n11617,
    new_n11618, new_n11619, new_n11620, new_n11621, new_n11622, new_n11623,
    new_n11624, new_n11625, new_n11626, new_n11627, new_n11628, new_n11629,
    new_n11630, new_n11631, new_n11632, new_n11633, new_n11634, new_n11635,
    new_n11636, new_n11637, new_n11638, new_n11639, new_n11640, new_n11641,
    new_n11642, new_n11643, new_n11644, new_n11645, new_n11646, new_n11647,
    new_n11648, new_n11649, new_n11650, new_n11651, new_n11652, new_n11653,
    new_n11654, new_n11655, new_n11656, new_n11657, new_n11658, new_n11659,
    new_n11660, new_n11661, new_n11662, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710, new_n11711, new_n11712, new_n11713,
    new_n11714, new_n11715, new_n11716, new_n11717, new_n11718, new_n11719,
    new_n11720, new_n11721, new_n11722, new_n11723, new_n11724, new_n11725,
    new_n11726, new_n11727, new_n11728, new_n11729, new_n11730, new_n11731,
    new_n11732, new_n11733, new_n11734, new_n11735, new_n11736, new_n11737,
    new_n11738, new_n11739, new_n11740, new_n11741, new_n11742, new_n11743,
    new_n11744, new_n11745, new_n11746, new_n11747, new_n11748, new_n11749,
    new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755,
    new_n11756, new_n11757, new_n11758, new_n11759, new_n11760, new_n11761,
    new_n11762, new_n11763, new_n11764, new_n11765, new_n11766, new_n11767,
    new_n11768, new_n11769, new_n11770, new_n11771, new_n11772, new_n11773,
    new_n11774, new_n11775, new_n11776, new_n11777, new_n11778, new_n11779,
    new_n11780, new_n11781, new_n11782, new_n11783, new_n11784, new_n11785,
    new_n11786, new_n11787, new_n11788, new_n11789, new_n11790, new_n11791,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820, new_n11821,
    new_n11822, new_n11823, new_n11824, new_n11825, new_n11826, new_n11827,
    new_n11828, new_n11829, new_n11830, new_n11831, new_n11832, new_n11833,
    new_n11834, new_n11835, new_n11836, new_n11837, new_n11838, new_n11839,
    new_n11840, new_n11841, new_n11842, new_n11843, new_n11844, new_n11845,
    new_n11846, new_n11847, new_n11848, new_n11849, new_n11850, new_n11851,
    new_n11852, new_n11853, new_n11854, new_n11855, new_n11856, new_n11857,
    new_n11858, new_n11859, new_n11860, new_n11861, new_n11862, new_n11863,
    new_n11864, new_n11865, new_n11866, new_n11867, new_n11868, new_n11869,
    new_n11870, new_n11871, new_n11872, new_n11873, new_n11874, new_n11875,
    new_n11876, new_n11877, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892, new_n11893,
    new_n11894, new_n11895, new_n11896, new_n11897, new_n11898, new_n11899,
    new_n11900, new_n11901, new_n11902, new_n11903, new_n11904, new_n11905,
    new_n11906, new_n11907, new_n11908, new_n11909, new_n11910, new_n11911,
    new_n11912, new_n11913, new_n11914, new_n11915, new_n11916, new_n11917,
    new_n11918, new_n11919, new_n11920, new_n11921, new_n11922, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948,
    new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954,
    new_n11955, new_n11956, new_n11957, new_n11958, new_n11959, new_n11960,
    new_n11961, new_n11962, new_n11963, new_n11964, new_n11965, new_n11966,
    new_n11967, new_n11968, new_n11969, new_n11970, new_n11971, new_n11972,
    new_n11973, new_n11974, new_n11975, new_n11976, new_n11977, new_n11978,
    new_n11979, new_n11980, new_n11981, new_n11982, new_n11983, new_n11984,
    new_n11985, new_n11986, new_n11987, new_n11988, new_n11989, new_n11990,
    new_n11991, new_n11992, new_n11993, new_n11994, new_n11995, new_n11996,
    new_n11997, new_n11998, new_n11999, new_n12000, new_n12001, new_n12002,
    new_n12003, new_n12004, new_n12005, new_n12006, new_n12007, new_n12008,
    new_n12009, new_n12010, new_n12011, new_n12012, new_n12013, new_n12014,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019, new_n12020,
    new_n12021, new_n12022, new_n12023, new_n12024, new_n12025, new_n12026,
    new_n12027, new_n12028, new_n12029, new_n12030, new_n12031, new_n12032,
    new_n12033, new_n12034, new_n12035, new_n12036, new_n12037, new_n12038,
    new_n12039, new_n12040, new_n12041, new_n12042, new_n12043, new_n12044,
    new_n12045, new_n12046, new_n12047, new_n12048, new_n12049, new_n12050,
    new_n12051, new_n12052, new_n12053, new_n12054, new_n12055, new_n12056,
    new_n12057, new_n12058, new_n12059, new_n12060, new_n12061, new_n12062,
    new_n12063, new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069, new_n12070, new_n12071, new_n12072, new_n12073, new_n12074,
    new_n12075, new_n12076, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111, new_n12112, new_n12113, new_n12114, new_n12115, new_n12116,
    new_n12117, new_n12118, new_n12119, new_n12120, new_n12121, new_n12122,
    new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128,
    new_n12129, new_n12130, new_n12131, new_n12132, new_n12133, new_n12134,
    new_n12135, new_n12136, new_n12137, new_n12138, new_n12139, new_n12140,
    new_n12141, new_n12142, new_n12143, new_n12144, new_n12145, new_n12146,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151, new_n12152,
    new_n12153, new_n12154, new_n12155, new_n12156, new_n12157, new_n12158,
    new_n12159, new_n12160, new_n12161, new_n12162, new_n12163, new_n12164,
    new_n12165, new_n12166, new_n12167, new_n12168, new_n12169, new_n12170,
    new_n12171, new_n12172, new_n12173, new_n12174, new_n12175, new_n12176,
    new_n12177, new_n12178, new_n12179, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188,
    new_n12189, new_n12190, new_n12191, new_n12192, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209, new_n12210, new_n12211, new_n12212,
    new_n12213, new_n12214, new_n12215, new_n12216, new_n12217, new_n12218,
    new_n12219, new_n12220, new_n12221, new_n12222, new_n12223, new_n12224,
    new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230,
    new_n12231, new_n12232, new_n12233, new_n12234, new_n12235, new_n12236,
    new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242,
    new_n12243, new_n12244, new_n12245, new_n12246, new_n12247, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12300, new_n12301, new_n12302, new_n12303,
    new_n12304, new_n12305, new_n12306, new_n12307, new_n12308, new_n12309,
    new_n12310, new_n12311, new_n12312, new_n12313, new_n12314, new_n12315,
    new_n12316, new_n12317, new_n12318, new_n12319, new_n12320, new_n12321,
    new_n12322, new_n12323, new_n12324, new_n12325, new_n12326, new_n12327,
    new_n12328, new_n12329, new_n12330, new_n12331, new_n12332, new_n12333,
    new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357,
    new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369,
    new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375,
    new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381,
    new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391, new_n12392, new_n12393,
    new_n12394, new_n12395, new_n12396, new_n12397, new_n12398, new_n12399,
    new_n12400, new_n12401, new_n12402, new_n12403, new_n12404, new_n12405,
    new_n12406, new_n12407, new_n12408, new_n12409, new_n12410, new_n12411,
    new_n12412, new_n12413, new_n12414, new_n12415, new_n12416, new_n12417,
    new_n12418, new_n12419, new_n12420, new_n12421, new_n12422, new_n12423,
    new_n12424, new_n12425, new_n12426, new_n12427, new_n12428, new_n12429,
    new_n12430, new_n12431, new_n12432, new_n12433, new_n12434, new_n12435,
    new_n12436, new_n12437, new_n12438, new_n12439, new_n12440, new_n12441,
    new_n12442, new_n12443, new_n12444, new_n12445, new_n12446, new_n12447,
    new_n12448, new_n12449, new_n12450, new_n12451, new_n12452, new_n12453,
    new_n12454, new_n12455, new_n12456, new_n12457, new_n12458, new_n12459,
    new_n12460, new_n12461, new_n12462, new_n12463, new_n12464, new_n12465,
    new_n12466, new_n12467, new_n12468, new_n12469, new_n12470, new_n12471,
    new_n12472, new_n12473, new_n12474, new_n12475, new_n12476, new_n12477,
    new_n12478, new_n12479, new_n12480, new_n12481, new_n12482, new_n12483,
    new_n12484, new_n12485, new_n12486, new_n12487, new_n12488, new_n12489,
    new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507,
    new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513,
    new_n12514, new_n12515, new_n12516, new_n12517, new_n12518, new_n12519,
    new_n12520, new_n12521, new_n12522, new_n12523, new_n12524, new_n12525,
    new_n12526, new_n12527, new_n12528, new_n12529, new_n12530, new_n12531,
    new_n12532, new_n12533, new_n12534, new_n12535, new_n12536, new_n12537,
    new_n12538, new_n12539, new_n12540, new_n12541, new_n12542, new_n12543,
    new_n12544, new_n12545, new_n12546, new_n12547, new_n12548, new_n12549,
    new_n12550, new_n12551, new_n12552, new_n12553, new_n12554, new_n12555,
    new_n12556, new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562, new_n12563, new_n12564, new_n12565, new_n12566, new_n12567,
    new_n12568, new_n12569, new_n12570, new_n12571, new_n12572, new_n12573,
    new_n12574, new_n12575, new_n12576, new_n12577, new_n12578, new_n12579,
    new_n12580, new_n12581, new_n12582, new_n12583, new_n12584, new_n12585,
    new_n12586, new_n12587, new_n12588, new_n12589, new_n12590, new_n12591,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12627, new_n12628,
    new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634,
    new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640,
    new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646,
    new_n12647, new_n12648, new_n12649, new_n12650, new_n12651, new_n12652,
    new_n12653, new_n12654, new_n12655, new_n12656, new_n12657, new_n12658,
    new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665, new_n12666, new_n12667, new_n12668, new_n12669, new_n12670,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694,
    new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700,
    new_n12701, new_n12702, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707, new_n12708, new_n12709, new_n12710, new_n12711, new_n12712,
    new_n12713, new_n12714, new_n12715, new_n12716, new_n12717, new_n12718,
    new_n12719, new_n12720, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740, new_n12741, new_n12742,
    new_n12743, new_n12744, new_n12745, new_n12746, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12751, new_n12752, new_n12753, new_n12754,
    new_n12755, new_n12756, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807, new_n12808,
    new_n12809, new_n12810, new_n12811, new_n12812, new_n12813, new_n12814,
    new_n12815, new_n12816, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821, new_n12822, new_n12823, new_n12824, new_n12825, new_n12826,
    new_n12827, new_n12828, new_n12829, new_n12830, new_n12831, new_n12832,
    new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838,
    new_n12839, new_n12840, new_n12841, new_n12842, new_n12843, new_n12844,
    new_n12845, new_n12846, new_n12847, new_n12848, new_n12849, new_n12850,
    new_n12851, new_n12852, new_n12853, new_n12854, new_n12855, new_n12856,
    new_n12857, new_n12858, new_n12859, new_n12860, new_n12861, new_n12862,
    new_n12863, new_n12864, new_n12865, new_n12866, new_n12867, new_n12868,
    new_n12869, new_n12870, new_n12871, new_n12872, new_n12873, new_n12874,
    new_n12875, new_n12876, new_n12877, new_n12878, new_n12879, new_n12880,
    new_n12881, new_n12882, new_n12883, new_n12884, new_n12885, new_n12886,
    new_n12887, new_n12888, new_n12889, new_n12890, new_n12891, new_n12892,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900, new_n12901, new_n12902, new_n12903, new_n12904,
    new_n12905, new_n12906, new_n12907, new_n12908, new_n12909, new_n12910,
    new_n12911, new_n12912, new_n12913, new_n12914, new_n12915, new_n12916,
    new_n12917, new_n12918, new_n12919, new_n12920, new_n12921, new_n12922,
    new_n12923, new_n12924, new_n12925, new_n12926, new_n12927, new_n12928,
    new_n12929, new_n12930, new_n12931, new_n12932, new_n12933, new_n12934,
    new_n12935, new_n12936, new_n12937, new_n12938, new_n12939, new_n12940,
    new_n12941, new_n12942, new_n12943, new_n12944, new_n12945, new_n12946,
    new_n12947, new_n12948, new_n12949, new_n12950, new_n12951, new_n12953,
    new_n12954, new_n12955, new_n12956, new_n12957, new_n12958, new_n12959,
    new_n12960, new_n12961, new_n12962, new_n12963, new_n12964, new_n12965,
    new_n12966, new_n12967, new_n12968, new_n12969, new_n12970, new_n12971,
    new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978, new_n12979, new_n12980, new_n12981, new_n12982, new_n12983,
    new_n12984, new_n12985, new_n12986, new_n12987, new_n12988, new_n12989,
    new_n12990, new_n12991, new_n12992, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005, new_n13006, new_n13007,
    new_n13008, new_n13009, new_n13010, new_n13011, new_n13012, new_n13013,
    new_n13014, new_n13015, new_n13016, new_n13017, new_n13018, new_n13019,
    new_n13020, new_n13021, new_n13022, new_n13023, new_n13024, new_n13025,
    new_n13026, new_n13027, new_n13028, new_n13029, new_n13030, new_n13031,
    new_n13032, new_n13033, new_n13034, new_n13035, new_n13036, new_n13037,
    new_n13038, new_n13039, new_n13040, new_n13041, new_n13042, new_n13043,
    new_n13044, new_n13045, new_n13046, new_n13047, new_n13048, new_n13049,
    new_n13050, new_n13051, new_n13052, new_n13053, new_n13054, new_n13055,
    new_n13056, new_n13057, new_n13058, new_n13059, new_n13060, new_n13061,
    new_n13062, new_n13063, new_n13064, new_n13065, new_n13066, new_n13067,
    new_n13068, new_n13069, new_n13070, new_n13071, new_n13072, new_n13073,
    new_n13074, new_n13075, new_n13076, new_n13077, new_n13078, new_n13079,
    new_n13080, new_n13081, new_n13082, new_n13083, new_n13084, new_n13085,
    new_n13086, new_n13087, new_n13088, new_n13089, new_n13090, new_n13091,
    new_n13092, new_n13093, new_n13094, new_n13095, new_n13096, new_n13097,
    new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103,
    new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109,
    new_n13110, new_n13111, new_n13112, new_n13113, new_n13114, new_n13115,
    new_n13116, new_n13117, new_n13118, new_n13119, new_n13120, new_n13121,
    new_n13122, new_n13123, new_n13124, new_n13125, new_n13126, new_n13127,
    new_n13128, new_n13129, new_n13130, new_n13131, new_n13132, new_n13133,
    new_n13134, new_n13135, new_n13136, new_n13137, new_n13138, new_n13139,
    new_n13140, new_n13141, new_n13142, new_n13143, new_n13144, new_n13145,
    new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151,
    new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157,
    new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163,
    new_n13164, new_n13165, new_n13166, new_n13167, new_n13168, new_n13169,
    new_n13170, new_n13171, new_n13172, new_n13173, new_n13174, new_n13175,
    new_n13176, new_n13177, new_n13178, new_n13179, new_n13180, new_n13181,
    new_n13182, new_n13183, new_n13184, new_n13185, new_n13186, new_n13187,
    new_n13188, new_n13189, new_n13190, new_n13191, new_n13192, new_n13193,
    new_n13194, new_n13195, new_n13196, new_n13197, new_n13198, new_n13199,
    new_n13200, new_n13201, new_n13202, new_n13203, new_n13204, new_n13205,
    new_n13206, new_n13207, new_n13208, new_n13209, new_n13210, new_n13211,
    new_n13212, new_n13213, new_n13214, new_n13215, new_n13216, new_n13217,
    new_n13218, new_n13219, new_n13220, new_n13221, new_n13222, new_n13223,
    new_n13224, new_n13225, new_n13226, new_n13227, new_n13228, new_n13229,
    new_n13230, new_n13231, new_n13232, new_n13233, new_n13234, new_n13235,
    new_n13236, new_n13237, new_n13238, new_n13239, new_n13240, new_n13241,
    new_n13242, new_n13243, new_n13244, new_n13245, new_n13246, new_n13247,
    new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253,
    new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259,
    new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404,
    new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13504, new_n13505, new_n13506, new_n13507,
    new_n13508, new_n13509, new_n13510, new_n13511, new_n13512, new_n13513,
    new_n13514, new_n13515, new_n13516, new_n13517, new_n13518, new_n13519,
    new_n13520, new_n13521, new_n13522, new_n13523, new_n13524, new_n13525,
    new_n13526, new_n13527, new_n13528, new_n13529, new_n13530, new_n13531,
    new_n13532, new_n13533, new_n13534, new_n13535, new_n13536, new_n13537,
    new_n13538, new_n13539, new_n13540, new_n13541, new_n13542, new_n13543,
    new_n13544, new_n13545, new_n13546, new_n13547, new_n13548, new_n13549,
    new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13722, new_n13723, new_n13724,
    new_n13725, new_n13726, new_n13727, new_n13728, new_n13729, new_n13730,
    new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736,
    new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742,
    new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748,
    new_n13749, new_n13750, new_n13751, new_n13752, new_n13753, new_n13754,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764, new_n13765, new_n13766,
    new_n13767, new_n13768, new_n13769, new_n13770, new_n13771, new_n13772,
    new_n13773, new_n13774, new_n13775, new_n13776, new_n13777, new_n13778,
    new_n13779, new_n13780, new_n13781, new_n13782, new_n13783, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850,
    new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856,
    new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862,
    new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868,
    new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874,
    new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880,
    new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886,
    new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892,
    new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898,
    new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904,
    new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910,
    new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13919, new_n13920, new_n13921, new_n13922,
    new_n13923, new_n13924, new_n13925, new_n13926, new_n13927, new_n13928,
    new_n13929, new_n13930, new_n13931, new_n13932, new_n13933, new_n13934,
    new_n13935, new_n13936, new_n13937, new_n13938, new_n13939, new_n13940,
    new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946,
    new_n13947, new_n13948, new_n13950, new_n13951, new_n13952, new_n13953,
    new_n13954, new_n13955, new_n13956, new_n13957, new_n13958, new_n13959,
    new_n13960, new_n13961, new_n13962, new_n13963, new_n13964, new_n13965,
    new_n13966, new_n13967, new_n13968, new_n13969, new_n13970, new_n13971,
    new_n13972, new_n13973, new_n13974, new_n13975, new_n13976, new_n13977,
    new_n13978, new_n13979, new_n13980, new_n13981, new_n13982, new_n13983,
    new_n13984, new_n13985, new_n13986, new_n13987, new_n13988, new_n13989,
    new_n13990, new_n13991, new_n13992, new_n13993, new_n13994, new_n13995,
    new_n13996, new_n13997, new_n13998, new_n13999, new_n14000, new_n14001,
    new_n14002, new_n14003, new_n14004, new_n14005, new_n14006, new_n14007,
    new_n14008, new_n14009, new_n14010, new_n14011, new_n14012, new_n14013,
    new_n14014, new_n14015, new_n14016, new_n14017, new_n14018, new_n14019,
    new_n14020, new_n14021, new_n14022, new_n14023, new_n14024, new_n14025,
    new_n14026, new_n14027, new_n14028, new_n14029, new_n14030, new_n14031,
    new_n14032, new_n14033, new_n14034, new_n14035, new_n14036, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059, new_n14060, new_n14061,
    new_n14062, new_n14063, new_n14064, new_n14065, new_n14066, new_n14067,
    new_n14068, new_n14069, new_n14070, new_n14071, new_n14072, new_n14073,
    new_n14074, new_n14075, new_n14076, new_n14077, new_n14078, new_n14079,
    new_n14080, new_n14081, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090, new_n14091,
    new_n14092, new_n14093, new_n14094, new_n14095, new_n14096, new_n14097,
    new_n14098, new_n14099, new_n14100, new_n14101, new_n14102, new_n14103,
    new_n14104, new_n14105, new_n14106, new_n14107, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120, new_n14121,
    new_n14122, new_n14123, new_n14124, new_n14125, new_n14126, new_n14127,
    new_n14128, new_n14129, new_n14130, new_n14131, new_n14132, new_n14133,
    new_n14134, new_n14135, new_n14136, new_n14137, new_n14138, new_n14139,
    new_n14140, new_n14141, new_n14142, new_n14143, new_n14144, new_n14145,
    new_n14146, new_n14147, new_n14148, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169,
    new_n14170, new_n14171, new_n14172, new_n14173, new_n14174, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14190, new_n14191, new_n14192, new_n14193, new_n14194,
    new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200,
    new_n14201, new_n14202, new_n14203, new_n14204, new_n14205, new_n14206,
    new_n14207, new_n14208, new_n14209, new_n14210, new_n14211, new_n14212,
    new_n14213, new_n14214, new_n14215, new_n14216, new_n14217, new_n14218,
    new_n14219, new_n14220, new_n14221, new_n14222, new_n14223, new_n14224,
    new_n14225, new_n14226, new_n14227, new_n14228, new_n14229, new_n14230,
    new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236,
    new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242,
    new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267, new_n14268, new_n14269, new_n14270, new_n14271, new_n14272,
    new_n14273, new_n14274, new_n14275, new_n14276, new_n14277, new_n14278,
    new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284,
    new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290,
    new_n14291, new_n14292, new_n14293, new_n14294, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310, new_n14311, new_n14312, new_n14313, new_n14314,
    new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320,
    new_n14321, new_n14322, new_n14323, new_n14324, new_n14325, new_n14326,
    new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332,
    new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342, new_n14343, new_n14344,
    new_n14345, new_n14346, new_n14347, new_n14348, new_n14349, new_n14350,
    new_n14351, new_n14352, new_n14353, new_n14354, new_n14355, new_n14356,
    new_n14357, new_n14358, new_n14359, new_n14360, new_n14361, new_n14362,
    new_n14363, new_n14364, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375, new_n14376, new_n14377, new_n14378, new_n14379, new_n14380,
    new_n14381, new_n14382, new_n14383, new_n14384, new_n14385, new_n14386,
    new_n14387, new_n14388, new_n14389, new_n14390, new_n14391, new_n14392,
    new_n14393, new_n14394, new_n14395, new_n14396, new_n14397, new_n14398,
    new_n14399, new_n14401, new_n14402, new_n14403, new_n14404, new_n14405,
    new_n14406, new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412, new_n14413, new_n14414, new_n14415, new_n14416, new_n14417,
    new_n14418, new_n14419, new_n14420, new_n14421, new_n14422, new_n14423,
    new_n14424, new_n14425, new_n14426, new_n14427, new_n14428, new_n14429,
    new_n14430, new_n14431, new_n14432, new_n14433, new_n14434, new_n14435,
    new_n14436, new_n14437, new_n14438, new_n14439, new_n14440, new_n14441,
    new_n14442, new_n14443, new_n14444, new_n14445, new_n14446, new_n14447,
    new_n14448, new_n14449, new_n14450, new_n14451, new_n14452, new_n14453,
    new_n14454, new_n14455, new_n14456, new_n14457, new_n14458, new_n14459,
    new_n14460, new_n14461, new_n14462, new_n14463, new_n14464, new_n14465,
    new_n14466, new_n14467, new_n14468, new_n14469, new_n14470, new_n14471,
    new_n14472, new_n14473, new_n14474, new_n14475, new_n14476, new_n14477,
    new_n14478, new_n14479, new_n14480, new_n14481, new_n14482, new_n14483,
    new_n14484, new_n14485, new_n14486, new_n14487, new_n14488, new_n14489,
    new_n14490, new_n14491, new_n14492, new_n14493, new_n14494, new_n14495,
    new_n14496, new_n14497, new_n14498, new_n14499, new_n14500, new_n14501,
    new_n14502, new_n14503, new_n14504, new_n14505, new_n14506, new_n14507,
    new_n14508, new_n14509, new_n14510, new_n14511, new_n14512, new_n14513,
    new_n14514, new_n14515, new_n14516, new_n14517, new_n14518, new_n14519,
    new_n14520, new_n14521, new_n14522, new_n14523, new_n14524, new_n14525,
    new_n14526, new_n14527, new_n14528, new_n14529, new_n14530, new_n14531,
    new_n14532, new_n14533, new_n14534, new_n14535, new_n14536, new_n14537,
    new_n14538, new_n14539, new_n14540, new_n14541, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546, new_n14547, new_n14548, new_n14549,
    new_n14550, new_n14551, new_n14552, new_n14553, new_n14554, new_n14555,
    new_n14556, new_n14557, new_n14558, new_n14559, new_n14560, new_n14561,
    new_n14562, new_n14563, new_n14564, new_n14565, new_n14566, new_n14567,
    new_n14568, new_n14569, new_n14570, new_n14571, new_n14572, new_n14573,
    new_n14574, new_n14575, new_n14576, new_n14577, new_n14578, new_n14579,
    new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585,
    new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591,
    new_n14592, new_n14593, new_n14594, new_n14595, new_n14596, new_n14597,
    new_n14598, new_n14599, new_n14600, new_n14601, new_n14602, new_n14603,
    new_n14604, new_n14605, new_n14606, new_n14607, new_n14608, new_n14609,
    new_n14610, new_n14611, new_n14612, new_n14613, new_n14614, new_n14615,
    new_n14616, new_n14617, new_n14619, new_n14620, new_n14621, new_n14622,
    new_n14623, new_n14624, new_n14625, new_n14626, new_n14627, new_n14628,
    new_n14629, new_n14630, new_n14631, new_n14632, new_n14633, new_n14634,
    new_n14635, new_n14636, new_n14637, new_n14638, new_n14639, new_n14640,
    new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646,
    new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652,
    new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658,
    new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664,
    new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670,
    new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676,
    new_n14677, new_n14678, new_n14679, new_n14680, new_n14681, new_n14682,
    new_n14683, new_n14684, new_n14685, new_n14686, new_n14687, new_n14688,
    new_n14689, new_n14690, new_n14691, new_n14692, new_n14693, new_n14694,
    new_n14695, new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701, new_n14702, new_n14703, new_n14704, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734, new_n14735, new_n14736,
    new_n14737, new_n14738, new_n14739, new_n14740, new_n14741, new_n14742,
    new_n14743, new_n14744, new_n14745, new_n14746, new_n14747, new_n14748,
    new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14761, new_n14762, new_n14763, new_n14764, new_n14765, new_n14766,
    new_n14767, new_n14768, new_n14769, new_n14770, new_n14771, new_n14772,
    new_n14773, new_n14774, new_n14775, new_n14776, new_n14777, new_n14778,
    new_n14779, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784,
    new_n14785, new_n14786, new_n14787, new_n14788, new_n14789, new_n14790,
    new_n14791, new_n14792, new_n14793, new_n14794, new_n14795, new_n14796,
    new_n14797, new_n14798, new_n14799, new_n14800, new_n14801, new_n14802,
    new_n14803, new_n14804, new_n14805, new_n14806, new_n14807, new_n14808,
    new_n14809, new_n14810, new_n14811, new_n14812, new_n14813, new_n14814,
    new_n14815, new_n14816, new_n14817, new_n14818, new_n14819, new_n14820,
    new_n14821, new_n14822, new_n14823, new_n14824, new_n14825, new_n14826,
    new_n14827, new_n14828, new_n14829, new_n14830, new_n14831, new_n14832,
    new_n14833, new_n14834, new_n14835, new_n14836, new_n14838, new_n14839,
    new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845,
    new_n14846, new_n14847, new_n14848, new_n14849, new_n14850, new_n14851,
    new_n14852, new_n14853, new_n14854, new_n14855, new_n14856, new_n14857,
    new_n14858, new_n14859, new_n14860, new_n14861, new_n14862, new_n14863,
    new_n14864, new_n14865, new_n14866, new_n14867, new_n14868, new_n14869,
    new_n14870, new_n14871, new_n14872, new_n14873, new_n14874, new_n14875,
    new_n14876, new_n14877, new_n14878, new_n14879, new_n14880, new_n14881,
    new_n14882, new_n14883, new_n14884, new_n14885, new_n14886, new_n14887,
    new_n14888, new_n14889, new_n14890, new_n14891, new_n14892, new_n14893,
    new_n14894, new_n14895, new_n14896, new_n14897, new_n14898, new_n14899,
    new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905,
    new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911,
    new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917,
    new_n14918, new_n14919, new_n14920, new_n14921, new_n14922, new_n14923,
    new_n14924, new_n14925, new_n14926, new_n14927, new_n14928, new_n14929,
    new_n14930, new_n14931, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944, new_n14945, new_n14946, new_n14947,
    new_n14948, new_n14949, new_n14950, new_n14951, new_n14952, new_n14953,
    new_n14954, new_n14955, new_n14956, new_n14957, new_n14958, new_n14959,
    new_n14960, new_n14961, new_n14962, new_n14963, new_n14964, new_n14965,
    new_n14966, new_n14967, new_n14968, new_n14969, new_n14970, new_n14971,
    new_n14972, new_n14973, new_n14974, new_n14975, new_n14976, new_n14977,
    new_n14978, new_n14979, new_n14980, new_n14981, new_n14982, new_n14983,
    new_n14984, new_n14985, new_n14986, new_n14987, new_n14988, new_n14989,
    new_n14990, new_n14991, new_n14992, new_n14993, new_n14994, new_n14995,
    new_n14996, new_n14997, new_n14998, new_n14999, new_n15000, new_n15001,
    new_n15002, new_n15003, new_n15004, new_n15005, new_n15006, new_n15007,
    new_n15008, new_n15009, new_n15010, new_n15011, new_n15012, new_n15013,
    new_n15014, new_n15015, new_n15016, new_n15017, new_n15018, new_n15019,
    new_n15020, new_n15021, new_n15022, new_n15023, new_n15024, new_n15025,
    new_n15026, new_n15027, new_n15028, new_n15029, new_n15030, new_n15031,
    new_n15032, new_n15033, new_n15034, new_n15035, new_n15036, new_n15037,
    new_n15038, new_n15039, new_n15041, new_n15042, new_n15043, new_n15044,
    new_n15045, new_n15046, new_n15047, new_n15048, new_n15049, new_n15050,
    new_n15051, new_n15052, new_n15053, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077, new_n15078, new_n15079, new_n15080,
    new_n15081, new_n15082, new_n15083, new_n15084, new_n15085, new_n15086,
    new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094, new_n15095, new_n15096, new_n15097, new_n15098,
    new_n15099, new_n15100, new_n15101, new_n15102, new_n15103, new_n15104,
    new_n15105, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110,
    new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116,
    new_n15117, new_n15118, new_n15119, new_n15120, new_n15121, new_n15122,
    new_n15123, new_n15124, new_n15125, new_n15126, new_n15127, new_n15128,
    new_n15129, new_n15130, new_n15131, new_n15132, new_n15133, new_n15134,
    new_n15135, new_n15136, new_n15137, new_n15138, new_n15139, new_n15140,
    new_n15141, new_n15142, new_n15143, new_n15144, new_n15145, new_n15146,
    new_n15147, new_n15148, new_n15149, new_n15150, new_n15151, new_n15152,
    new_n15153, new_n15154, new_n15155, new_n15156, new_n15157, new_n15158,
    new_n15159, new_n15160, new_n15161, new_n15162, new_n15163, new_n15164,
    new_n15165, new_n15166, new_n15167, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175, new_n15176,
    new_n15177, new_n15178, new_n15179, new_n15180, new_n15181, new_n15182,
    new_n15183, new_n15184, new_n15185, new_n15186, new_n15187, new_n15188,
    new_n15189, new_n15190, new_n15191, new_n15192, new_n15193, new_n15194,
    new_n15195, new_n15196, new_n15197, new_n15198, new_n15199, new_n15200,
    new_n15201, new_n15202, new_n15203, new_n15204, new_n15205, new_n15206,
    new_n15207, new_n15208, new_n15209, new_n15210, new_n15211, new_n15212,
    new_n15213, new_n15214, new_n15215, new_n15216, new_n15217, new_n15218,
    new_n15219, new_n15220, new_n15221, new_n15222, new_n15223, new_n15224,
    new_n15225, new_n15226, new_n15227, new_n15229, new_n15230, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241, new_n15242, new_n15243,
    new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249,
    new_n15250, new_n15251, new_n15252, new_n15253, new_n15254, new_n15255,
    new_n15256, new_n15257, new_n15258, new_n15259, new_n15260, new_n15261,
    new_n15262, new_n15263, new_n15264, new_n15265, new_n15266, new_n15267,
    new_n15268, new_n15269, new_n15270, new_n15271, new_n15272, new_n15273,
    new_n15274, new_n15275, new_n15276, new_n15277, new_n15278, new_n15279,
    new_n15280, new_n15281, new_n15282, new_n15283, new_n15284, new_n15285,
    new_n15286, new_n15287, new_n15288, new_n15289, new_n15290, new_n15291,
    new_n15292, new_n15293, new_n15294, new_n15295, new_n15296, new_n15297,
    new_n15298, new_n15299, new_n15300, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307, new_n15308, new_n15309,
    new_n15310, new_n15311, new_n15312, new_n15313, new_n15314, new_n15315,
    new_n15316, new_n15317, new_n15318, new_n15319, new_n15320, new_n15321,
    new_n15322, new_n15323, new_n15324, new_n15325, new_n15326, new_n15327,
    new_n15328, new_n15329, new_n15330, new_n15331, new_n15332, new_n15333,
    new_n15334, new_n15335, new_n15336, new_n15337, new_n15338, new_n15339,
    new_n15340, new_n15341, new_n15342, new_n15343, new_n15344, new_n15345,
    new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351,
    new_n15352, new_n15353, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366, new_n15367, new_n15368, new_n15369,
    new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378, new_n15379, new_n15380, new_n15381,
    new_n15382, new_n15383, new_n15384, new_n15385, new_n15386, new_n15387,
    new_n15388, new_n15389, new_n15390, new_n15391, new_n15392, new_n15393,
    new_n15394, new_n15395, new_n15397, new_n15398, new_n15399, new_n15400,
    new_n15401, new_n15402, new_n15403, new_n15404, new_n15405, new_n15406,
    new_n15407, new_n15408, new_n15409, new_n15410, new_n15411, new_n15412,
    new_n15413, new_n15414, new_n15415, new_n15416, new_n15417, new_n15418,
    new_n15419, new_n15420, new_n15421, new_n15422, new_n15423, new_n15424,
    new_n15425, new_n15426, new_n15427, new_n15428, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435, new_n15436,
    new_n15437, new_n15438, new_n15439, new_n15440, new_n15441, new_n15442,
    new_n15443, new_n15444, new_n15445, new_n15446, new_n15447, new_n15448,
    new_n15449, new_n15450, new_n15451, new_n15452, new_n15453, new_n15454,
    new_n15455, new_n15456, new_n15457, new_n15458, new_n15459, new_n15460,
    new_n15461, new_n15462, new_n15463, new_n15464, new_n15465, new_n15466,
    new_n15467, new_n15468, new_n15469, new_n15470, new_n15471, new_n15472,
    new_n15473, new_n15474, new_n15475, new_n15476, new_n15477, new_n15478,
    new_n15479, new_n15480, new_n15481, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15490,
    new_n15491, new_n15492, new_n15493, new_n15494, new_n15495, new_n15496,
    new_n15497, new_n15498, new_n15499, new_n15500, new_n15501, new_n15502,
    new_n15503, new_n15504, new_n15505, new_n15506, new_n15507, new_n15508,
    new_n15509, new_n15510, new_n15511, new_n15512, new_n15513, new_n15514,
    new_n15515, new_n15516, new_n15517, new_n15518, new_n15519, new_n15520,
    new_n15521, new_n15522, new_n15523, new_n15524, new_n15525, new_n15526,
    new_n15527, new_n15528, new_n15529, new_n15530, new_n15531, new_n15532,
    new_n15533, new_n15534, new_n15535, new_n15536, new_n15537, new_n15538,
    new_n15539, new_n15540, new_n15541, new_n15542, new_n15543, new_n15544,
    new_n15545, new_n15546, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555, new_n15556,
    new_n15557, new_n15558, new_n15559, new_n15560, new_n15561, new_n15562,
    new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568,
    new_n15569, new_n15570, new_n15571, new_n15572, new_n15573, new_n15574,
    new_n15575, new_n15576, new_n15577, new_n15578, new_n15579, new_n15581,
    new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588, new_n15589, new_n15590, new_n15591, new_n15592, new_n15593,
    new_n15594, new_n15595, new_n15596, new_n15597, new_n15598, new_n15599,
    new_n15600, new_n15601, new_n15602, new_n15603, new_n15604, new_n15605,
    new_n15606, new_n15607, new_n15608, new_n15609, new_n15610, new_n15611,
    new_n15612, new_n15613, new_n15614, new_n15615, new_n15616, new_n15617,
    new_n15618, new_n15619, new_n15620, new_n15621, new_n15622, new_n15623,
    new_n15624, new_n15625, new_n15626, new_n15627, new_n15628, new_n15629,
    new_n15630, new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636, new_n15637, new_n15638, new_n15639, new_n15640, new_n15641,
    new_n15642, new_n15643, new_n15644, new_n15645, new_n15646, new_n15647,
    new_n15648, new_n15649, new_n15650, new_n15651, new_n15652, new_n15653,
    new_n15654, new_n15655, new_n15656, new_n15657, new_n15658, new_n15659,
    new_n15660, new_n15661, new_n15662, new_n15663, new_n15664, new_n15665,
    new_n15666, new_n15667, new_n15668, new_n15669, new_n15670, new_n15671,
    new_n15672, new_n15673, new_n15674, new_n15675, new_n15676, new_n15677,
    new_n15678, new_n15679, new_n15680, new_n15681, new_n15682, new_n15683,
    new_n15684, new_n15685, new_n15686, new_n15687, new_n15688, new_n15689,
    new_n15690, new_n15691, new_n15692, new_n15693, new_n15694, new_n15695,
    new_n15696, new_n15697, new_n15698, new_n15699, new_n15700, new_n15701,
    new_n15702, new_n15703, new_n15704, new_n15705, new_n15706, new_n15707,
    new_n15708, new_n15709, new_n15710, new_n15711, new_n15712, new_n15713,
    new_n15714, new_n15715, new_n15716, new_n15717, new_n15718, new_n15719,
    new_n15720, new_n15721, new_n15722, new_n15723, new_n15724, new_n15725,
    new_n15726, new_n15727, new_n15728, new_n15729, new_n15730, new_n15731,
    new_n15732, new_n15733, new_n15734, new_n15735, new_n15736, new_n15737,
    new_n15738, new_n15739, new_n15740, new_n15741, new_n15742, new_n15743,
    new_n15744, new_n15745, new_n15746, new_n15747, new_n15748, new_n15749,
    new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755,
    new_n15756, new_n15757, new_n15758, new_n15759, new_n15760, new_n15761,
    new_n15762, new_n15763, new_n15764, new_n15765, new_n15766, new_n15767,
    new_n15768, new_n15769, new_n15770, new_n15771, new_n15772, new_n15773,
    new_n15774, new_n15775, new_n15776, new_n15777, new_n15779, new_n15780,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798,
    new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804,
    new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810,
    new_n15811, new_n15812, new_n15813, new_n15814, new_n15815, new_n15816,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845, new_n15846,
    new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859, new_n15860, new_n15861, new_n15862, new_n15863, new_n15864,
    new_n15865, new_n15866, new_n15867, new_n15868, new_n15869, new_n15870,
    new_n15871, new_n15872, new_n15873, new_n15874, new_n15875, new_n15876,
    new_n15877, new_n15878, new_n15879, new_n15880, new_n15881, new_n15882,
    new_n15883, new_n15884, new_n15885, new_n15886, new_n15887, new_n15888,
    new_n15889, new_n15890, new_n15891, new_n15892, new_n15893, new_n15894,
    new_n15895, new_n15896, new_n15897, new_n15898, new_n15899, new_n15900,
    new_n15901, new_n15902, new_n15903, new_n15904, new_n15905, new_n15906,
    new_n15907, new_n15908, new_n15909, new_n15910, new_n15911, new_n15912,
    new_n15913, new_n15914, new_n15915, new_n15916, new_n15917, new_n15918,
    new_n15919, new_n15920, new_n15921, new_n15922, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935, new_n15937,
    new_n15938, new_n15939, new_n15940, new_n15941, new_n15942, new_n15943,
    new_n15944, new_n15945, new_n15946, new_n15947, new_n15948, new_n15949,
    new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955,
    new_n15956, new_n15957, new_n15958, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966, new_n15967,
    new_n15968, new_n15969, new_n15970, new_n15971, new_n15972, new_n15973,
    new_n15974, new_n15975, new_n15976, new_n15977, new_n15978, new_n15979,
    new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985,
    new_n15986, new_n15987, new_n15988, new_n15989, new_n15990, new_n15991,
    new_n15992, new_n15993, new_n15994, new_n15995, new_n15996, new_n15997,
    new_n15998, new_n15999, new_n16000, new_n16001, new_n16002, new_n16003,
    new_n16004, new_n16005, new_n16006, new_n16007, new_n16008, new_n16009,
    new_n16010, new_n16011, new_n16012, new_n16013, new_n16014, new_n16015,
    new_n16016, new_n16017, new_n16018, new_n16019, new_n16020, new_n16021,
    new_n16022, new_n16023, new_n16024, new_n16025, new_n16026, new_n16027,
    new_n16028, new_n16029, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051,
    new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057,
    new_n16058, new_n16059, new_n16060, new_n16061, new_n16062, new_n16063,
    new_n16064, new_n16065, new_n16066, new_n16067, new_n16068, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16078, new_n16079, new_n16080, new_n16081,
    new_n16082, new_n16083, new_n16084, new_n16085, new_n16086, new_n16087,
    new_n16088, new_n16089, new_n16090, new_n16091, new_n16092, new_n16093,
    new_n16094, new_n16095, new_n16096, new_n16097, new_n16098, new_n16099,
    new_n16100, new_n16101, new_n16102, new_n16103, new_n16104, new_n16105,
    new_n16106, new_n16107, new_n16108, new_n16109, new_n16110, new_n16111,
    new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117,
    new_n16118, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124,
    new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220,
    new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16232,
    new_n16233, new_n16234, new_n16235, new_n16236, new_n16237, new_n16238,
    new_n16239, new_n16240, new_n16241, new_n16242, new_n16243, new_n16244,
    new_n16245, new_n16246, new_n16247, new_n16248, new_n16249, new_n16250,
    new_n16251, new_n16252, new_n16253, new_n16254, new_n16255, new_n16256,
    new_n16257, new_n16258, new_n16259, new_n16260, new_n16261, new_n16262,
    new_n16263, new_n16264, new_n16265, new_n16266, new_n16267, new_n16268,
    new_n16269, new_n16270, new_n16271, new_n16272, new_n16273, new_n16274,
    new_n16275, new_n16276, new_n16277, new_n16278, new_n16279, new_n16280,
    new_n16281, new_n16282, new_n16283, new_n16284, new_n16285, new_n16286,
    new_n16287, new_n16288, new_n16289, new_n16290, new_n16291, new_n16292,
    new_n16293, new_n16294, new_n16295, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311,
    new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317,
    new_n16318, new_n16319, new_n16320, new_n16321, new_n16322, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350, new_n16351, new_n16352, new_n16353,
    new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359,
    new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365,
    new_n16366, new_n16367, new_n16368, new_n16369, new_n16370, new_n16371,
    new_n16372, new_n16373, new_n16374, new_n16375, new_n16376, new_n16377,
    new_n16378, new_n16379, new_n16380, new_n16381, new_n16382, new_n16383,
    new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389,
    new_n16390, new_n16391, new_n16392, new_n16393, new_n16394, new_n16395,
    new_n16396, new_n16397, new_n16398, new_n16399, new_n16400, new_n16401,
    new_n16402, new_n16403, new_n16404, new_n16405, new_n16406, new_n16407,
    new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413,
    new_n16414, new_n16415, new_n16416, new_n16417, new_n16418, new_n16419,
    new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425,
    new_n16426, new_n16427, new_n16428, new_n16429, new_n16430, new_n16431,
    new_n16432, new_n16433, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439, new_n16440, new_n16441, new_n16442, new_n16443,
    new_n16444, new_n16445, new_n16446, new_n16447, new_n16448, new_n16449,
    new_n16450, new_n16451, new_n16452, new_n16453, new_n16454, new_n16455,
    new_n16456, new_n16457, new_n16458, new_n16459, new_n16460, new_n16461,
    new_n16462, new_n16463, new_n16464, new_n16465, new_n16467, new_n16468,
    new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474,
    new_n16475, new_n16476, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481, new_n16482, new_n16483, new_n16484, new_n16485, new_n16486,
    new_n16487, new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493, new_n16494, new_n16495, new_n16496, new_n16497, new_n16498,
    new_n16499, new_n16500, new_n16501, new_n16502, new_n16503, new_n16504,
    new_n16505, new_n16506, new_n16507, new_n16508, new_n16509, new_n16510,
    new_n16511, new_n16512, new_n16513, new_n16514, new_n16515, new_n16516,
    new_n16517, new_n16518, new_n16519, new_n16520, new_n16521, new_n16522,
    new_n16523, new_n16524, new_n16525, new_n16526, new_n16527, new_n16528,
    new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534,
    new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540,
    new_n16541, new_n16542, new_n16543, new_n16544, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583, new_n16584, new_n16585, new_n16586, new_n16587, new_n16588,
    new_n16589, new_n16590, new_n16591, new_n16592, new_n16593, new_n16594,
    new_n16595, new_n16596, new_n16597, new_n16598, new_n16599, new_n16600,
    new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606,
    new_n16607, new_n16608, new_n16609, new_n16610, new_n16611, new_n16612,
    new_n16613, new_n16614, new_n16615, new_n16616, new_n16617, new_n16618,
    new_n16619, new_n16620, new_n16621, new_n16622, new_n16623, new_n16624,
    new_n16625, new_n16626, new_n16627, new_n16628, new_n16629, new_n16630,
    new_n16631, new_n16632, new_n16633, new_n16634, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661,
    new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667,
    new_n16668, new_n16669, new_n16670, new_n16671, new_n16672, new_n16673,
    new_n16674, new_n16675, new_n16676, new_n16677, new_n16678, new_n16679,
    new_n16680, new_n16681, new_n16682, new_n16683, new_n16684, new_n16685,
    new_n16686, new_n16687, new_n16688, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722, new_n16723, new_n16724, new_n16725, new_n16726, new_n16727,
    new_n16728, new_n16729, new_n16730, new_n16731, new_n16732, new_n16733,
    new_n16734, new_n16735, new_n16736, new_n16737, new_n16738, new_n16739,
    new_n16740, new_n16741, new_n16742, new_n16743, new_n16744, new_n16745,
    new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751,
    new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16768, new_n16769,
    new_n16770, new_n16771, new_n16772, new_n16773, new_n16774, new_n16775,
    new_n16776, new_n16777, new_n16778, new_n16779, new_n16780, new_n16781,
    new_n16782, new_n16783, new_n16784, new_n16785, new_n16786, new_n16787,
    new_n16788, new_n16789, new_n16790, new_n16791, new_n16792, new_n16793,
    new_n16795, new_n16796, new_n16797, new_n16798, new_n16799, new_n16800,
    new_n16801, new_n16802, new_n16803, new_n16804, new_n16805, new_n16806,
    new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824,
    new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830,
    new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836,
    new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842,
    new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848,
    new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854,
    new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890,
    new_n16891, new_n16892, new_n16893, new_n16894, new_n16895, new_n16896,
    new_n16897, new_n16898, new_n16899, new_n16900, new_n16901, new_n16902,
    new_n16903, new_n16904, new_n16905, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16945,
    new_n16946, new_n16947, new_n16948, new_n16949, new_n16950, new_n16951,
    new_n16952, new_n16953, new_n16954, new_n16955, new_n16956, new_n16957,
    new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963,
    new_n16964, new_n16965, new_n16966, new_n16967, new_n16968, new_n16969,
    new_n16970, new_n16971, new_n16972, new_n16973, new_n16974, new_n16975,
    new_n16976, new_n16977, new_n16978, new_n16979, new_n16980, new_n16981,
    new_n16982, new_n16983, new_n16984, new_n16985, new_n16986, new_n16987,
    new_n16988, new_n16989, new_n16990, new_n16991, new_n16992, new_n16993,
    new_n16994, new_n16995, new_n16996, new_n16997, new_n16998, new_n16999,
    new_n17000, new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006, new_n17007, new_n17008, new_n17009, new_n17010, new_n17011,
    new_n17012, new_n17013, new_n17014, new_n17015, new_n17016, new_n17017,
    new_n17018, new_n17019, new_n17020, new_n17021, new_n17022, new_n17023,
    new_n17024, new_n17025, new_n17026, new_n17027, new_n17028, new_n17029,
    new_n17030, new_n17031, new_n17032, new_n17033, new_n17034, new_n17035,
    new_n17036, new_n17037, new_n17038, new_n17039, new_n17040, new_n17041,
    new_n17042, new_n17043, new_n17044, new_n17045, new_n17046, new_n17047,
    new_n17048, new_n17049, new_n17050, new_n17051, new_n17052, new_n17053,
    new_n17054, new_n17055, new_n17056, new_n17057, new_n17058, new_n17059,
    new_n17060, new_n17061, new_n17062, new_n17063, new_n17064, new_n17065,
    new_n17066, new_n17067, new_n17068, new_n17069, new_n17070, new_n17071,
    new_n17072, new_n17073, new_n17074, new_n17075, new_n17076, new_n17077,
    new_n17078, new_n17079, new_n17080, new_n17081, new_n17082, new_n17083,
    new_n17084, new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090, new_n17091, new_n17092, new_n17093, new_n17094, new_n17095,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104, new_n17105, new_n17106, new_n17107,
    new_n17108, new_n17109, new_n17110, new_n17111, new_n17112, new_n17113,
    new_n17114, new_n17115, new_n17116, new_n17117, new_n17118, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17129, new_n17130, new_n17131, new_n17132,
    new_n17133, new_n17134, new_n17135, new_n17136, new_n17137, new_n17138,
    new_n17139, new_n17140, new_n17141, new_n17142, new_n17143, new_n17144,
    new_n17145, new_n17146, new_n17147, new_n17148, new_n17149, new_n17150,
    new_n17151, new_n17152, new_n17153, new_n17154, new_n17155, new_n17156,
    new_n17157, new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163, new_n17164, new_n17165, new_n17166, new_n17167, new_n17168,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186,
    new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17192,
    new_n17193, new_n17194, new_n17195, new_n17196, new_n17197, new_n17198,
    new_n17199, new_n17200, new_n17201, new_n17202, new_n17203, new_n17204,
    new_n17205, new_n17206, new_n17207, new_n17208, new_n17209, new_n17210,
    new_n17211, new_n17212, new_n17213, new_n17214, new_n17215, new_n17216,
    new_n17217, new_n17218, new_n17219, new_n17220, new_n17221, new_n17222,
    new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228,
    new_n17229, new_n17230, new_n17231, new_n17232, new_n17233, new_n17234,
    new_n17235, new_n17236, new_n17237, new_n17238, new_n17239, new_n17240,
    new_n17241, new_n17242, new_n17243, new_n17244, new_n17245, new_n17246,
    new_n17247, new_n17248, new_n17249, new_n17250, new_n17251, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263, new_n17264,
    new_n17265, new_n17266, new_n17267, new_n17268, new_n17269, new_n17270,
    new_n17271, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277,
    new_n17278, new_n17279, new_n17280, new_n17281, new_n17282, new_n17283,
    new_n17284, new_n17285, new_n17286, new_n17287, new_n17288, new_n17289,
    new_n17290, new_n17291, new_n17292, new_n17293, new_n17294, new_n17295,
    new_n17296, new_n17297, new_n17298, new_n17299, new_n17300, new_n17301,
    new_n17302, new_n17303, new_n17304, new_n17305, new_n17306, new_n17307,
    new_n17308, new_n17309, new_n17310, new_n17311, new_n17312, new_n17313,
    new_n17314, new_n17315, new_n17316, new_n17317, new_n17318, new_n17319,
    new_n17320, new_n17321, new_n17322, new_n17323, new_n17324, new_n17325,
    new_n17326, new_n17327, new_n17328, new_n17329, new_n17330, new_n17331,
    new_n17332, new_n17333, new_n17334, new_n17335, new_n17336, new_n17337,
    new_n17338, new_n17339, new_n17340, new_n17341, new_n17342, new_n17343,
    new_n17344, new_n17345, new_n17346, new_n17347, new_n17348, new_n17349,
    new_n17350, new_n17351, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359, new_n17360, new_n17361,
    new_n17362, new_n17363, new_n17364, new_n17365, new_n17366, new_n17367,
    new_n17368, new_n17369, new_n17370, new_n17371, new_n17372, new_n17373,
    new_n17374, new_n17375, new_n17376, new_n17377, new_n17378, new_n17379,
    new_n17380, new_n17381, new_n17382, new_n17383, new_n17384, new_n17385,
    new_n17386, new_n17387, new_n17388, new_n17389, new_n17390, new_n17391,
    new_n17392, new_n17393, new_n17394, new_n17395, new_n17396, new_n17397,
    new_n17398, new_n17399, new_n17400, new_n17401, new_n17402, new_n17403,
    new_n17404, new_n17405, new_n17406, new_n17407, new_n17408, new_n17409,
    new_n17410, new_n17412, new_n17413, new_n17414, new_n17415, new_n17416,
    new_n17417, new_n17418, new_n17419, new_n17420, new_n17421, new_n17422,
    new_n17423, new_n17424, new_n17425, new_n17426, new_n17427, new_n17428,
    new_n17429, new_n17430, new_n17431, new_n17432, new_n17433, new_n17434,
    new_n17435, new_n17436, new_n17437, new_n17438, new_n17439, new_n17440,
    new_n17441, new_n17442, new_n17443, new_n17444, new_n17445, new_n17446,
    new_n17447, new_n17448, new_n17449, new_n17450, new_n17451, new_n17452,
    new_n17453, new_n17454, new_n17455, new_n17456, new_n17457, new_n17458,
    new_n17459, new_n17460, new_n17461, new_n17462, new_n17463, new_n17464,
    new_n17465, new_n17466, new_n17467, new_n17468, new_n17469, new_n17470,
    new_n17471, new_n17472, new_n17473, new_n17474, new_n17475, new_n17476,
    new_n17477, new_n17478, new_n17479, new_n17480, new_n17481, new_n17482,
    new_n17483, new_n17484, new_n17485, new_n17486, new_n17487, new_n17488,
    new_n17489, new_n17490, new_n17491, new_n17492, new_n17493, new_n17494,
    new_n17495, new_n17496, new_n17497, new_n17498, new_n17499, new_n17500,
    new_n17501, new_n17502, new_n17503, new_n17504, new_n17505, new_n17506,
    new_n17507, new_n17508, new_n17509, new_n17510, new_n17511, new_n17512,
    new_n17513, new_n17514, new_n17515, new_n17516, new_n17517, new_n17518,
    new_n17519, new_n17520, new_n17521, new_n17522, new_n17523, new_n17524,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529, new_n17530,
    new_n17531, new_n17532, new_n17533, new_n17534, new_n17535, new_n17536,
    new_n17537, new_n17538, new_n17539, new_n17540, new_n17541, new_n17542,
    new_n17543, new_n17544, new_n17545, new_n17546, new_n17547, new_n17548,
    new_n17549, new_n17550, new_n17551, new_n17552, new_n17553, new_n17554,
    new_n17555, new_n17556, new_n17557, new_n17558, new_n17559, new_n17560,
    new_n17561, new_n17562, new_n17563, new_n17564, new_n17565, new_n17566,
    new_n17567, new_n17568, new_n17569, new_n17570, new_n17571, new_n17572,
    new_n17573, new_n17574, new_n17575, new_n17577, new_n17578, new_n17579,
    new_n17580, new_n17581, new_n17582, new_n17583, new_n17584, new_n17585,
    new_n17586, new_n17587, new_n17588, new_n17589, new_n17590, new_n17591,
    new_n17592, new_n17593, new_n17594, new_n17595, new_n17596, new_n17597,
    new_n17598, new_n17599, new_n17600, new_n17601, new_n17602, new_n17603,
    new_n17604, new_n17605, new_n17606, new_n17607, new_n17608, new_n17609,
    new_n17610, new_n17611, new_n17612, new_n17613, new_n17614, new_n17615,
    new_n17616, new_n17617, new_n17618, new_n17619, new_n17620, new_n17621,
    new_n17622, new_n17623, new_n17624, new_n17625, new_n17626, new_n17627,
    new_n17628, new_n17629, new_n17630, new_n17631, new_n17632, new_n17633,
    new_n17634, new_n17635, new_n17636, new_n17637, new_n17638, new_n17639,
    new_n17640, new_n17641, new_n17642, new_n17643, new_n17644, new_n17645,
    new_n17646, new_n17647, new_n17648, new_n17649, new_n17650, new_n17651,
    new_n17652, new_n17653, new_n17654, new_n17655, new_n17656, new_n17657,
    new_n17658, new_n17659, new_n17660, new_n17661, new_n17662, new_n17663,
    new_n17664, new_n17665, new_n17666, new_n17667, new_n17668, new_n17669,
    new_n17670, new_n17671, new_n17672, new_n17673, new_n17674, new_n17675,
    new_n17676, new_n17677, new_n17678, new_n17679, new_n17680, new_n17681,
    new_n17682, new_n17683, new_n17684, new_n17685, new_n17686, new_n17687,
    new_n17688, new_n17689, new_n17690, new_n17691, new_n17692, new_n17693,
    new_n17694, new_n17695, new_n17696, new_n17697, new_n17698, new_n17699,
    new_n17700, new_n17701, new_n17702, new_n17703, new_n17704, new_n17705,
    new_n17706, new_n17707, new_n17708, new_n17709, new_n17710, new_n17711,
    new_n17712, new_n17713, new_n17714, new_n17715, new_n17716, new_n17717,
    new_n17718, new_n17719, new_n17720, new_n17721, new_n17722, new_n17723,
    new_n17724, new_n17725, new_n17726, new_n17727, new_n17728, new_n17729,
    new_n17730, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736,
    new_n17737, new_n17738, new_n17739, new_n17740, new_n17741, new_n17742,
    new_n17743, new_n17744, new_n17745, new_n17746, new_n17747, new_n17748,
    new_n17749, new_n17750, new_n17751, new_n17752, new_n17753, new_n17754,
    new_n17755, new_n17756, new_n17757, new_n17758, new_n17759, new_n17760,
    new_n17761, new_n17762, new_n17763, new_n17764, new_n17765, new_n17766,
    new_n17767, new_n17768, new_n17769, new_n17770, new_n17771, new_n17772,
    new_n17773, new_n17774, new_n17775, new_n17776, new_n17777, new_n17778,
    new_n17779, new_n17780, new_n17781, new_n17782, new_n17783, new_n17784,
    new_n17785, new_n17786, new_n17787, new_n17788, new_n17789, new_n17790,
    new_n17791, new_n17792, new_n17793, new_n17794, new_n17795, new_n17796,
    new_n17797, new_n17798, new_n17799, new_n17800, new_n17801, new_n17802,
    new_n17803, new_n17804, new_n17805, new_n17806, new_n17807, new_n17808,
    new_n17809, new_n17810, new_n17811, new_n17812, new_n17813, new_n17814,
    new_n17815, new_n17816, new_n17817, new_n17818, new_n17819, new_n17820,
    new_n17821, new_n17822, new_n17823, new_n17824, new_n17825, new_n17826,
    new_n17827, new_n17828, new_n17829, new_n17830, new_n17831, new_n17832,
    new_n17833, new_n17834, new_n17835, new_n17836, new_n17837, new_n17838,
    new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17844,
    new_n17845, new_n17846, new_n17847, new_n17848, new_n17849, new_n17850,
    new_n17851, new_n17852, new_n17853, new_n17854, new_n17855, new_n17856,
    new_n17857, new_n17858, new_n17859, new_n17860, new_n17861, new_n17862,
    new_n17863, new_n17864, new_n17865, new_n17867, new_n17868, new_n17869,
    new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875,
    new_n17876, new_n17877, new_n17878, new_n17879, new_n17880, new_n17881,
    new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887,
    new_n17888, new_n17889, new_n17890, new_n17891, new_n17892, new_n17893,
    new_n17894, new_n17895, new_n17896, new_n17897, new_n17898, new_n17899,
    new_n17900, new_n17901, new_n17902, new_n17903, new_n17904, new_n17905,
    new_n17906, new_n17907, new_n17908, new_n17909, new_n17910, new_n17911,
    new_n17912, new_n17913, new_n17914, new_n17915, new_n17916, new_n17917,
    new_n17918, new_n17919, new_n17920, new_n17921, new_n17922, new_n17923,
    new_n17924, new_n17925, new_n17926, new_n17927, new_n17928, new_n17929,
    new_n17930, new_n17931, new_n17932, new_n17933, new_n17934, new_n17935,
    new_n17936, new_n17937, new_n17938, new_n17939, new_n17940, new_n17941,
    new_n17942, new_n17943, new_n17944, new_n17945, new_n17946, new_n17947,
    new_n17948, new_n17949, new_n17950, new_n17951, new_n17952, new_n17953,
    new_n17954, new_n17955, new_n17956, new_n17957, new_n17958, new_n17959,
    new_n17960, new_n17961, new_n17962, new_n17963, new_n17964, new_n17965,
    new_n17966, new_n17967, new_n17968, new_n17969, new_n17970, new_n17971,
    new_n17972, new_n17973, new_n17974, new_n17975, new_n17976, new_n17977,
    new_n17978, new_n17979, new_n17980, new_n17981, new_n17982, new_n17983,
    new_n17984, new_n17985, new_n17986, new_n17987, new_n17988, new_n17989,
    new_n17990, new_n17991, new_n17992, new_n17993, new_n17994, new_n17995,
    new_n17996, new_n17997, new_n17998, new_n17999, new_n18000, new_n18001,
    new_n18002, new_n18003, new_n18004, new_n18005, new_n18006, new_n18007,
    new_n18008, new_n18009, new_n18010, new_n18011, new_n18012, new_n18013,
    new_n18014, new_n18015, new_n18016, new_n18017, new_n18018, new_n18019,
    new_n18020, new_n18022, new_n18023, new_n18024, new_n18025, new_n18026,
    new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032,
    new_n18033, new_n18034, new_n18035, new_n18036, new_n18037, new_n18038,
    new_n18039, new_n18040, new_n18041, new_n18042, new_n18043, new_n18044,
    new_n18045, new_n18046, new_n18047, new_n18048, new_n18049, new_n18050,
    new_n18051, new_n18052, new_n18053, new_n18054, new_n18055, new_n18056,
    new_n18057, new_n18058, new_n18059, new_n18060, new_n18061, new_n18062,
    new_n18063, new_n18064, new_n18065, new_n18066, new_n18067, new_n18068,
    new_n18069, new_n18070, new_n18071, new_n18072, new_n18073, new_n18074,
    new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080,
    new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086,
    new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092,
    new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098,
    new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105, new_n18106, new_n18107, new_n18108, new_n18109, new_n18110,
    new_n18111, new_n18112, new_n18113, new_n18114, new_n18115, new_n18116,
    new_n18117, new_n18118, new_n18119, new_n18120, new_n18121, new_n18122,
    new_n18123, new_n18124, new_n18125, new_n18126, new_n18127, new_n18128,
    new_n18129, new_n18130, new_n18131, new_n18132, new_n18133, new_n18134,
    new_n18135, new_n18136, new_n18137, new_n18138, new_n18139, new_n18140,
    new_n18141, new_n18142, new_n18143, new_n18144, new_n18145, new_n18146,
    new_n18147, new_n18148, new_n18149, new_n18150, new_n18151, new_n18152,
    new_n18153, new_n18154, new_n18155, new_n18156, new_n18157, new_n18158,
    new_n18159, new_n18160, new_n18161, new_n18162, new_n18163, new_n18164,
    new_n18165, new_n18166, new_n18168, new_n18169, new_n18170, new_n18171,
    new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177,
    new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183,
    new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189,
    new_n18190, new_n18191, new_n18192, new_n18193, new_n18194, new_n18195,
    new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18210, new_n18211, new_n18212, new_n18213,
    new_n18214, new_n18215, new_n18216, new_n18217, new_n18218, new_n18219,
    new_n18220, new_n18221, new_n18222, new_n18223, new_n18224, new_n18225,
    new_n18226, new_n18227, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232, new_n18233, new_n18234, new_n18235, new_n18236, new_n18237,
    new_n18238, new_n18239, new_n18240, new_n18241, new_n18242, new_n18243,
    new_n18244, new_n18245, new_n18246, new_n18247, new_n18248, new_n18249,
    new_n18250, new_n18251, new_n18252, new_n18253, new_n18254, new_n18255,
    new_n18256, new_n18257, new_n18258, new_n18259, new_n18260, new_n18261,
    new_n18262, new_n18263, new_n18264, new_n18265, new_n18266, new_n18267,
    new_n18268, new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274, new_n18275, new_n18276, new_n18277, new_n18278, new_n18279,
    new_n18280, new_n18281, new_n18282, new_n18283, new_n18284, new_n18285,
    new_n18286, new_n18287, new_n18288, new_n18289, new_n18290, new_n18292,
    new_n18293, new_n18294, new_n18295, new_n18296, new_n18297, new_n18298,
    new_n18299, new_n18300, new_n18301, new_n18302, new_n18303, new_n18304,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309, new_n18310,
    new_n18311, new_n18312, new_n18313, new_n18314, new_n18315, new_n18316,
    new_n18317, new_n18318, new_n18319, new_n18320, new_n18321, new_n18322,
    new_n18323, new_n18324, new_n18325, new_n18326, new_n18327, new_n18328,
    new_n18329, new_n18330, new_n18331, new_n18332, new_n18333, new_n18334,
    new_n18335, new_n18336, new_n18337, new_n18338, new_n18339, new_n18340,
    new_n18341, new_n18342, new_n18343, new_n18344, new_n18345, new_n18346,
    new_n18347, new_n18348, new_n18349, new_n18350, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376,
    new_n18377, new_n18378, new_n18379, new_n18380, new_n18381, new_n18382,
    new_n18383, new_n18384, new_n18385, new_n18386, new_n18387, new_n18388,
    new_n18389, new_n18390, new_n18391, new_n18392, new_n18393, new_n18394,
    new_n18395, new_n18396, new_n18397, new_n18398, new_n18399, new_n18400,
    new_n18401, new_n18402, new_n18403, new_n18404, new_n18405, new_n18406,
    new_n18407, new_n18408, new_n18409, new_n18410, new_n18411, new_n18412,
    new_n18413, new_n18414, new_n18415, new_n18416, new_n18417, new_n18418,
    new_n18419, new_n18420, new_n18421, new_n18422, new_n18423, new_n18424,
    new_n18425, new_n18426, new_n18427, new_n18428, new_n18429, new_n18430,
    new_n18431, new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437, new_n18438, new_n18439, new_n18440, new_n18441, new_n18442,
    new_n18443, new_n18444, new_n18445, new_n18447, new_n18448, new_n18449,
    new_n18450, new_n18451, new_n18452, new_n18453, new_n18454, new_n18455,
    new_n18456, new_n18457, new_n18458, new_n18459, new_n18460, new_n18461,
    new_n18462, new_n18463, new_n18464, new_n18465, new_n18466, new_n18467,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482, new_n18483, new_n18484, new_n18485,
    new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491,
    new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508, new_n18509,
    new_n18510, new_n18511, new_n18512, new_n18513, new_n18514, new_n18515,
    new_n18516, new_n18517, new_n18518, new_n18519, new_n18520, new_n18521,
    new_n18522, new_n18523, new_n18524, new_n18525, new_n18526, new_n18527,
    new_n18528, new_n18529, new_n18530, new_n18531, new_n18532, new_n18533,
    new_n18534, new_n18535, new_n18536, new_n18537, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557,
    new_n18558, new_n18559, new_n18560, new_n18561, new_n18562, new_n18563,
    new_n18564, new_n18565, new_n18566, new_n18567, new_n18568, new_n18569,
    new_n18570, new_n18571, new_n18572, new_n18573, new_n18574, new_n18575,
    new_n18576, new_n18577, new_n18578, new_n18579, new_n18580, new_n18581,
    new_n18582, new_n18583, new_n18584, new_n18585, new_n18586, new_n18588,
    new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594,
    new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600,
    new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18606,
    new_n18607, new_n18608, new_n18609, new_n18610, new_n18611, new_n18612,
    new_n18613, new_n18614, new_n18615, new_n18616, new_n18617, new_n18618,
    new_n18619, new_n18620, new_n18621, new_n18622, new_n18623, new_n18624,
    new_n18625, new_n18626, new_n18627, new_n18628, new_n18629, new_n18630,
    new_n18631, new_n18632, new_n18633, new_n18634, new_n18635, new_n18636,
    new_n18637, new_n18638, new_n18639, new_n18640, new_n18641, new_n18642,
    new_n18643, new_n18644, new_n18645, new_n18646, new_n18647, new_n18648,
    new_n18649, new_n18650, new_n18651, new_n18652, new_n18653, new_n18654,
    new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18715,
    new_n18716, new_n18717, new_n18718, new_n18719, new_n18720, new_n18721,
    new_n18722, new_n18723, new_n18724, new_n18725, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18734, new_n18735, new_n18736, new_n18737, new_n18738, new_n18739,
    new_n18740, new_n18741, new_n18742, new_n18743, new_n18744, new_n18745,
    new_n18746, new_n18747, new_n18748, new_n18749, new_n18750, new_n18751,
    new_n18752, new_n18753, new_n18754, new_n18755, new_n18756, new_n18757,
    new_n18758, new_n18759, new_n18760, new_n18761, new_n18762, new_n18763,
    new_n18764, new_n18765, new_n18766, new_n18767, new_n18768, new_n18769,
    new_n18770, new_n18771, new_n18772, new_n18773, new_n18774, new_n18775,
    new_n18776, new_n18777, new_n18778, new_n18779, new_n18780, new_n18781,
    new_n18782, new_n18783, new_n18784, new_n18785, new_n18786, new_n18787,
    new_n18788, new_n18789, new_n18790, new_n18791, new_n18792, new_n18793,
    new_n18794, new_n18795, new_n18796, new_n18797, new_n18798, new_n18799,
    new_n18800, new_n18801, new_n18802, new_n18803, new_n18804, new_n18805,
    new_n18806, new_n18807, new_n18808, new_n18809, new_n18810, new_n18811,
    new_n18812, new_n18813, new_n18814, new_n18815, new_n18816, new_n18817,
    new_n18818, new_n18819, new_n18820, new_n18821, new_n18822, new_n18823,
    new_n18824, new_n18825, new_n18826, new_n18827, new_n18828, new_n18829,
    new_n18830, new_n18831, new_n18832, new_n18833, new_n18834, new_n18835,
    new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843, new_n18844, new_n18845, new_n18846, new_n18847,
    new_n18848, new_n18849, new_n18850, new_n18851, new_n18852, new_n18853,
    new_n18854, new_n18856, new_n18857, new_n18858, new_n18859, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864, new_n18865, new_n18866,
    new_n18867, new_n18868, new_n18869, new_n18870, new_n18871, new_n18872,
    new_n18873, new_n18874, new_n18875, new_n18876, new_n18877, new_n18878,
    new_n18879, new_n18880, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886, new_n18887, new_n18888, new_n18889, new_n18890,
    new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896,
    new_n18897, new_n18898, new_n18899, new_n18900, new_n18901, new_n18902,
    new_n18903, new_n18904, new_n18905, new_n18906, new_n18907, new_n18908,
    new_n18909, new_n18910, new_n18911, new_n18912, new_n18913, new_n18914,
    new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962,
    new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968,
    new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18985, new_n18986, new_n18987,
    new_n18988, new_n18989, new_n18990, new_n18991, new_n18992, new_n18993,
    new_n18994, new_n18995, new_n18996, new_n18997, new_n18998, new_n18999,
    new_n19000, new_n19001, new_n19002, new_n19003, new_n19004, new_n19005,
    new_n19006, new_n19007, new_n19008, new_n19009, new_n19010, new_n19011,
    new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017,
    new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023,
    new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033, new_n19034, new_n19035,
    new_n19036, new_n19037, new_n19038, new_n19039, new_n19040, new_n19041,
    new_n19042, new_n19043, new_n19044, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077,
    new_n19078, new_n19079, new_n19080, new_n19081, new_n19082, new_n19083,
    new_n19084, new_n19085, new_n19086, new_n19087, new_n19088, new_n19089,
    new_n19090, new_n19092, new_n19093, new_n19094, new_n19095, new_n19096,
    new_n19097, new_n19098, new_n19099, new_n19100, new_n19101, new_n19102,
    new_n19103, new_n19104, new_n19105, new_n19106, new_n19107, new_n19108,
    new_n19109, new_n19110, new_n19111, new_n19112, new_n19113, new_n19114,
    new_n19115, new_n19116, new_n19117, new_n19118, new_n19119, new_n19120,
    new_n19121, new_n19122, new_n19123, new_n19124, new_n19125, new_n19126,
    new_n19127, new_n19128, new_n19129, new_n19130, new_n19131, new_n19132,
    new_n19133, new_n19134, new_n19135, new_n19136, new_n19137, new_n19138,
    new_n19139, new_n19140, new_n19141, new_n19142, new_n19143, new_n19144,
    new_n19145, new_n19146, new_n19147, new_n19148, new_n19149, new_n19150,
    new_n19151, new_n19152, new_n19153, new_n19154, new_n19155, new_n19156,
    new_n19157, new_n19158, new_n19159, new_n19160, new_n19161, new_n19162,
    new_n19163, new_n19164, new_n19165, new_n19166, new_n19167, new_n19168,
    new_n19169, new_n19170, new_n19171, new_n19172, new_n19173, new_n19174,
    new_n19175, new_n19176, new_n19177, new_n19178, new_n19179, new_n19180,
    new_n19181, new_n19182, new_n19183, new_n19184, new_n19185, new_n19186,
    new_n19187, new_n19188, new_n19189, new_n19190, new_n19191, new_n19192,
    new_n19193, new_n19194, new_n19195, new_n19196, new_n19197, new_n19198,
    new_n19199, new_n19200, new_n19201, new_n19202, new_n19203, new_n19204,
    new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210,
    new_n19211, new_n19212, new_n19213, new_n19214, new_n19215, new_n19216,
    new_n19217, new_n19218, new_n19219, new_n19220, new_n19221, new_n19223,
    new_n19224, new_n19225, new_n19226, new_n19227, new_n19228, new_n19229,
    new_n19230, new_n19231, new_n19232, new_n19233, new_n19234, new_n19235,
    new_n19236, new_n19237, new_n19238, new_n19239, new_n19240, new_n19241,
    new_n19242, new_n19243, new_n19244, new_n19245, new_n19246, new_n19247,
    new_n19248, new_n19249, new_n19250, new_n19251, new_n19252, new_n19253,
    new_n19254, new_n19255, new_n19256, new_n19257, new_n19258, new_n19259,
    new_n19260, new_n19261, new_n19262, new_n19263, new_n19264, new_n19265,
    new_n19266, new_n19267, new_n19268, new_n19269, new_n19270, new_n19271,
    new_n19272, new_n19273, new_n19274, new_n19275, new_n19276, new_n19277,
    new_n19278, new_n19279, new_n19280, new_n19281, new_n19282, new_n19283,
    new_n19284, new_n19285, new_n19286, new_n19287, new_n19288, new_n19289,
    new_n19290, new_n19291, new_n19292, new_n19293, new_n19294, new_n19295,
    new_n19296, new_n19297, new_n19298, new_n19299, new_n19300, new_n19301,
    new_n19302, new_n19303, new_n19304, new_n19305, new_n19306, new_n19307,
    new_n19308, new_n19309, new_n19310, new_n19311, new_n19312, new_n19313,
    new_n19314, new_n19315, new_n19316, new_n19317, new_n19318, new_n19319,
    new_n19320, new_n19321, new_n19322, new_n19323, new_n19324, new_n19325,
    new_n19326, new_n19327, new_n19328, new_n19329, new_n19330, new_n19331,
    new_n19332, new_n19333, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19339, new_n19340, new_n19341, new_n19342, new_n19343, new_n19344,
    new_n19345, new_n19346, new_n19347, new_n19348, new_n19349, new_n19350,
    new_n19351, new_n19352, new_n19353, new_n19354, new_n19355, new_n19356,
    new_n19357, new_n19358, new_n19359, new_n19360, new_n19361, new_n19362,
    new_n19363, new_n19364, new_n19365, new_n19366, new_n19367, new_n19368,
    new_n19369, new_n19370, new_n19371, new_n19372, new_n19373, new_n19374,
    new_n19375, new_n19376, new_n19377, new_n19378, new_n19379, new_n19380,
    new_n19381, new_n19382, new_n19383, new_n19384, new_n19385, new_n19386,
    new_n19387, new_n19388, new_n19389, new_n19390, new_n19391, new_n19392,
    new_n19393, new_n19394, new_n19395, new_n19396, new_n19397, new_n19398,
    new_n19399, new_n19400, new_n19401, new_n19402, new_n19403, new_n19404,
    new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410,
    new_n19411, new_n19412, new_n19413, new_n19414, new_n19415, new_n19416,
    new_n19417, new_n19418, new_n19419, new_n19420, new_n19421, new_n19422,
    new_n19423, new_n19424, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19443, new_n19444, new_n19445, new_n19446, new_n19447,
    new_n19448, new_n19449, new_n19450, new_n19451, new_n19452, new_n19453,
    new_n19454, new_n19455, new_n19456, new_n19457, new_n19458, new_n19459,
    new_n19460, new_n19461, new_n19462, new_n19463, new_n19464, new_n19465,
    new_n19466, new_n19467, new_n19468, new_n19469, new_n19470, new_n19471,
    new_n19472, new_n19473, new_n19474, new_n19475, new_n19476, new_n19477,
    new_n19478, new_n19479, new_n19480, new_n19481, new_n19482, new_n19483,
    new_n19484, new_n19485, new_n19486, new_n19487, new_n19488, new_n19489,
    new_n19490, new_n19491, new_n19492, new_n19493, new_n19494, new_n19495,
    new_n19496, new_n19497, new_n19498, new_n19499, new_n19500, new_n19501,
    new_n19502, new_n19503, new_n19504, new_n19505, new_n19506, new_n19507,
    new_n19508, new_n19509, new_n19510, new_n19511, new_n19512, new_n19513,
    new_n19514, new_n19515, new_n19516, new_n19517, new_n19518, new_n19519,
    new_n19520, new_n19521, new_n19522, new_n19523, new_n19524, new_n19525,
    new_n19526, new_n19527, new_n19528, new_n19529, new_n19530, new_n19531,
    new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19537,
    new_n19538, new_n19539, new_n19540, new_n19541, new_n19542, new_n19543,
    new_n19544, new_n19545, new_n19546, new_n19547, new_n19548, new_n19549,
    new_n19550, new_n19552, new_n19553, new_n19554, new_n19555, new_n19556,
    new_n19557, new_n19558, new_n19559, new_n19560, new_n19561, new_n19562,
    new_n19563, new_n19564, new_n19565, new_n19566, new_n19567, new_n19568,
    new_n19569, new_n19570, new_n19571, new_n19572, new_n19573, new_n19574,
    new_n19575, new_n19576, new_n19577, new_n19578, new_n19579, new_n19580,
    new_n19581, new_n19582, new_n19583, new_n19584, new_n19585, new_n19586,
    new_n19587, new_n19588, new_n19589, new_n19590, new_n19591, new_n19592,
    new_n19593, new_n19594, new_n19595, new_n19596, new_n19597, new_n19598,
    new_n19599, new_n19600, new_n19601, new_n19602, new_n19603, new_n19604,
    new_n19605, new_n19606, new_n19607, new_n19608, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617, new_n19618, new_n19619, new_n19620, new_n19621, new_n19622,
    new_n19623, new_n19624, new_n19625, new_n19626, new_n19627, new_n19628,
    new_n19629, new_n19630, new_n19631, new_n19632, new_n19633, new_n19634,
    new_n19635, new_n19636, new_n19637, new_n19638, new_n19639, new_n19640,
    new_n19641, new_n19642, new_n19643, new_n19644, new_n19646, new_n19647,
    new_n19648, new_n19649, new_n19650, new_n19651, new_n19652, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664, new_n19665,
    new_n19666, new_n19667, new_n19668, new_n19669, new_n19670, new_n19671,
    new_n19672, new_n19673, new_n19674, new_n19675, new_n19676, new_n19677,
    new_n19678, new_n19679, new_n19680, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700, new_n19701,
    new_n19702, new_n19703, new_n19704, new_n19705, new_n19706, new_n19707,
    new_n19708, new_n19709, new_n19710, new_n19711, new_n19712, new_n19713,
    new_n19714, new_n19715, new_n19716, new_n19717, new_n19718, new_n19719,
    new_n19720, new_n19721, new_n19722, new_n19723, new_n19724, new_n19725,
    new_n19726, new_n19727, new_n19728, new_n19729, new_n19730, new_n19731,
    new_n19733, new_n19734, new_n19735, new_n19736, new_n19737, new_n19738,
    new_n19739, new_n19740, new_n19741, new_n19742, new_n19743, new_n19744,
    new_n19745, new_n19746, new_n19747, new_n19748, new_n19749, new_n19750,
    new_n19751, new_n19752, new_n19753, new_n19754, new_n19755, new_n19756,
    new_n19757, new_n19758, new_n19759, new_n19760, new_n19761, new_n19762,
    new_n19763, new_n19764, new_n19765, new_n19766, new_n19767, new_n19768,
    new_n19769, new_n19770, new_n19771, new_n19772, new_n19773, new_n19774,
    new_n19775, new_n19776, new_n19777, new_n19778, new_n19779, new_n19780,
    new_n19781, new_n19782, new_n19783, new_n19784, new_n19785, new_n19786,
    new_n19787, new_n19788, new_n19789, new_n19790, new_n19791, new_n19792,
    new_n19793, new_n19794, new_n19795, new_n19796, new_n19797, new_n19798,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803, new_n19804,
    new_n19805, new_n19806, new_n19807, new_n19808, new_n19809, new_n19810,
    new_n19811, new_n19812, new_n19813, new_n19814, new_n19815, new_n19816,
    new_n19817, new_n19818, new_n19819, new_n19820, new_n19821, new_n19822,
    new_n19823, new_n19824, new_n19825, new_n19827, new_n19828, new_n19829,
    new_n19830, new_n19831, new_n19832, new_n19833, new_n19834, new_n19835,
    new_n19836, new_n19837, new_n19838, new_n19839, new_n19840, new_n19841,
    new_n19842, new_n19843, new_n19844, new_n19845, new_n19846, new_n19847,
    new_n19848, new_n19849, new_n19850, new_n19851, new_n19852, new_n19853,
    new_n19854, new_n19855, new_n19856, new_n19857, new_n19858, new_n19859,
    new_n19860, new_n19861, new_n19862, new_n19863, new_n19864, new_n19865,
    new_n19866, new_n19867, new_n19868, new_n19869, new_n19870, new_n19871,
    new_n19872, new_n19873, new_n19874, new_n19875, new_n19876, new_n19877,
    new_n19878, new_n19879, new_n19880, new_n19881, new_n19882, new_n19883,
    new_n19884, new_n19885, new_n19886, new_n19887, new_n19888, new_n19889,
    new_n19890, new_n19891, new_n19892, new_n19893, new_n19894, new_n19895,
    new_n19896, new_n19897, new_n19898, new_n19899, new_n19900, new_n19901,
    new_n19902, new_n19903, new_n19904, new_n19905, new_n19906, new_n19908,
    new_n19909, new_n19910, new_n19911, new_n19912, new_n19913, new_n19914,
    new_n19915, new_n19916, new_n19917, new_n19918, new_n19919, new_n19920,
    new_n19921, new_n19922, new_n19923, new_n19924, new_n19925, new_n19926,
    new_n19927, new_n19928, new_n19929, new_n19930, new_n19931, new_n19932,
    new_n19933, new_n19934, new_n19935, new_n19936, new_n19937, new_n19938,
    new_n19939, new_n19940, new_n19941, new_n19942, new_n19943, new_n19944,
    new_n19945, new_n19946, new_n19947, new_n19948, new_n19949, new_n19950,
    new_n19951, new_n19952, new_n19953, new_n19954, new_n19955, new_n19956,
    new_n19957, new_n19958, new_n19959, new_n19960, new_n19961, new_n19962,
    new_n19963, new_n19964, new_n19965, new_n19966, new_n19967, new_n19968,
    new_n19969, new_n19970, new_n19971, new_n19972, new_n19973, new_n19974,
    new_n19975, new_n19976, new_n19977, new_n19978, new_n19979, new_n19980,
    new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986,
    new_n19987, new_n19988, new_n19989, new_n19990, new_n19992, new_n19993,
    new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999,
    new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005,
    new_n20006, new_n20007, new_n20008, new_n20009, new_n20010, new_n20011,
    new_n20012, new_n20013, new_n20014, new_n20015, new_n20016, new_n20017,
    new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023,
    new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029,
    new_n20030, new_n20031, new_n20032, new_n20033, new_n20034, new_n20035,
    new_n20036, new_n20037, new_n20038, new_n20039, new_n20040, new_n20041,
    new_n20042, new_n20043, new_n20044, new_n20045, new_n20046, new_n20047,
    new_n20048, new_n20049, new_n20050, new_n20051, new_n20052, new_n20053,
    new_n20054, new_n20055, new_n20056, new_n20057, new_n20058, new_n20059,
    new_n20060, new_n20061, new_n20062, new_n20063, new_n20064, new_n20065,
    new_n20066, new_n20067, new_n20068, new_n20069, new_n20070, new_n20071,
    new_n20072, new_n20073, new_n20074, new_n20075, new_n20076, new_n20077,
    new_n20078, new_n20079, new_n20080, new_n20081, new_n20082, new_n20083,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20162, new_n20163,
    new_n20164, new_n20165, new_n20166, new_n20167, new_n20168, new_n20169,
    new_n20170, new_n20171, new_n20172, new_n20173, new_n20174, new_n20175,
    new_n20176, new_n20177, new_n20178, new_n20179, new_n20180, new_n20181,
    new_n20182, new_n20183, new_n20184, new_n20185, new_n20186, new_n20187,
    new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193,
    new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199,
    new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20229, new_n20230,
    new_n20231, new_n20232, new_n20233, new_n20234, new_n20235, new_n20236,
    new_n20237, new_n20238, new_n20239, new_n20240, new_n20241, new_n20242,
    new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248,
    new_n20249, new_n20250, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259, new_n20260,
    new_n20261, new_n20262, new_n20263, new_n20264, new_n20265, new_n20266,
    new_n20267, new_n20268, new_n20269, new_n20270, new_n20271, new_n20272,
    new_n20273, new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279, new_n20280, new_n20281, new_n20282, new_n20283, new_n20284,
    new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20294, new_n20295, new_n20296, new_n20297,
    new_n20298, new_n20299, new_n20300, new_n20301, new_n20302, new_n20303,
    new_n20304, new_n20305, new_n20306, new_n20307, new_n20308, new_n20309,
    new_n20310, new_n20311, new_n20312, new_n20313, new_n20314, new_n20315,
    new_n20316, new_n20317, new_n20318, new_n20319, new_n20320, new_n20321,
    new_n20322, new_n20323, new_n20324, new_n20325, new_n20326, new_n20327,
    new_n20328, new_n20329, new_n20330, new_n20331, new_n20332, new_n20333,
    new_n20334, new_n20335, new_n20336, new_n20337, new_n20338, new_n20339,
    new_n20340, new_n20341, new_n20342, new_n20343, new_n20344, new_n20345,
    new_n20346, new_n20347, new_n20348, new_n20349, new_n20350, new_n20351,
    new_n20352, new_n20353, new_n20354, new_n20355, new_n20356, new_n20357,
    new_n20358, new_n20359, new_n20361, new_n20362, new_n20363, new_n20364,
    new_n20365, new_n20366, new_n20367, new_n20368, new_n20369, new_n20370,
    new_n20371, new_n20372, new_n20373, new_n20374, new_n20375, new_n20376,
    new_n20377, new_n20378, new_n20379, new_n20380, new_n20381, new_n20382,
    new_n20383, new_n20384, new_n20385, new_n20386, new_n20387, new_n20388,
    new_n20389, new_n20390, new_n20391, new_n20392, new_n20393, new_n20394,
    new_n20395, new_n20396, new_n20397, new_n20398, new_n20399, new_n20400,
    new_n20401, new_n20402, new_n20403, new_n20404, new_n20405, new_n20406,
    new_n20407, new_n20408, new_n20409, new_n20410, new_n20411, new_n20412,
    new_n20413, new_n20414, new_n20415, new_n20416, new_n20418, new_n20419,
    new_n20420, new_n20421, new_n20422, new_n20423, new_n20424, new_n20425,
    new_n20426, new_n20427, new_n20428, new_n20429, new_n20430, new_n20431,
    new_n20432, new_n20433, new_n20434, new_n20435, new_n20436, new_n20437,
    new_n20438, new_n20439, new_n20440, new_n20441, new_n20442, new_n20443,
    new_n20444, new_n20445, new_n20446, new_n20447, new_n20448, new_n20449,
    new_n20450, new_n20451, new_n20452, new_n20453, new_n20454, new_n20455,
    new_n20456, new_n20457, new_n20458, new_n20459, new_n20460, new_n20461,
    new_n20462, new_n20463, new_n20464, new_n20465, new_n20466, new_n20467,
    new_n20468, new_n20469, new_n20470, new_n20471, new_n20472, new_n20473,
    new_n20474, new_n20475, new_n20476, new_n20477, new_n20478, new_n20479,
    new_n20480, new_n20481, new_n20482, new_n20483, new_n20485, new_n20486,
    new_n20487, new_n20488, new_n20489, new_n20490, new_n20491, new_n20492,
    new_n20493, new_n20494, new_n20495, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504,
    new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510,
    new_n20511, new_n20512, new_n20513, new_n20514, new_n20515, new_n20516,
    new_n20517, new_n20518, new_n20519, new_n20520, new_n20521, new_n20522,
    new_n20523, new_n20524, new_n20525, new_n20526, new_n20527, new_n20528,
    new_n20529, new_n20530, new_n20531, new_n20532, new_n20533, new_n20534,
    new_n20535, new_n20536, new_n20537, new_n20538, new_n20539, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553,
    new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582, new_n20583,
    new_n20584, new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590, new_n20591, new_n20592, new_n20593, new_n20594, new_n20595,
    new_n20596, new_n20598, new_n20599, new_n20600, new_n20601, new_n20602,
    new_n20603, new_n20604, new_n20605, new_n20606, new_n20607, new_n20608,
    new_n20609, new_n20610, new_n20611, new_n20612, new_n20613, new_n20614,
    new_n20615, new_n20616, new_n20617, new_n20618, new_n20619, new_n20620,
    new_n20621, new_n20622, new_n20623, new_n20624, new_n20625, new_n20626,
    new_n20627, new_n20628, new_n20629, new_n20630, new_n20631, new_n20632,
    new_n20633, new_n20634, new_n20635, new_n20636, new_n20637, new_n20639,
    new_n20640, new_n20641, new_n20642, new_n20643, new_n20644, new_n20645,
    new_n20646, new_n20647, new_n20648, new_n20649, new_n20650, new_n20651,
    new_n20652, new_n20653, new_n20654, new_n20655, new_n20656, new_n20657,
    new_n20658, new_n20659, new_n20660, new_n20661, new_n20662, new_n20663,
    new_n20664, new_n20665, new_n20666, new_n20667, new_n20668, new_n20669,
    new_n20670, new_n20671, new_n20672, new_n20673, new_n20674, new_n20675,
    new_n20676, new_n20677, new_n20678, new_n20679, new_n20680, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685, new_n20687, new_n20688,
    new_n20689, new_n20690, new_n20691, new_n20692, new_n20693, new_n20694,
    new_n20695, new_n20696, new_n20697, new_n20698, new_n20699, new_n20700,
    new_n20701, new_n20702, new_n20703, new_n20704, new_n20705, new_n20706,
    new_n20707, new_n20708, new_n20709, new_n20710, new_n20711, new_n20712,
    new_n20713, new_n20714, new_n20715, new_n20716, new_n20717, new_n20718,
    new_n20719, new_n20720, new_n20721, new_n20722, new_n20723, new_n20724,
    new_n20725, new_n20726, new_n20727, new_n20728, new_n20729, new_n20731,
    new_n20732, new_n20733, new_n20734, new_n20735, new_n20736, new_n20737,
    new_n20738, new_n20739, new_n20740, new_n20741, new_n20742, new_n20743,
    new_n20744, new_n20745, new_n20746, new_n20747, new_n20748, new_n20749,
    new_n20750, new_n20751, new_n20752, new_n20753, new_n20754, new_n20755,
    new_n20756, new_n20757, new_n20758, new_n20759, new_n20760, new_n20761,
    new_n20762, new_n20763, new_n20764, new_n20765, new_n20766, new_n20767,
    new_n20768, new_n20769, new_n20770, new_n20772, new_n20773, new_n20774,
    new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780,
    new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786,
    new_n20787, new_n20788, new_n20789, new_n20790, new_n20791, new_n20792,
    new_n20793, new_n20794, new_n20795, new_n20796, new_n20797, new_n20798,
    new_n20800, new_n20801, new_n20802, new_n20803, new_n20804, new_n20805,
    new_n20806, new_n20807, new_n20808, new_n20809, new_n20810, new_n20811,
    new_n20812, new_n20813, new_n20814, new_n20815, new_n20816, new_n20817,
    new_n20818, new_n20819, new_n20820, new_n20821, new_n20822, new_n20823,
    new_n20824, new_n20825, new_n20826, new_n20827, new_n20828, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836,
    new_n20837, new_n20838, new_n20839, new_n20840, new_n20841, new_n20842,
    new_n20843, new_n20844, new_n20845, new_n20846, new_n20847, new_n20848,
    new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854,
    new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860,
    new_n20862, new_n20863, new_n20864, new_n20865, new_n20866, new_n20867,
    new_n20868, new_n20869, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20878, new_n20879,
    new_n20880, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20894, new_n20895, new_n20896;
  INVx1_ASAP7_75t_L         g00000(.A(\a[0] ), .Y(new_n257));
  INVx1_ASAP7_75t_L         g00001(.A(\b[0] ), .Y(new_n258));
  NOR2xp33_ASAP7_75t_L      g00002(.A(new_n257), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00003(.A(\a[2] ), .B(\f[0] ), .Y(new_n260));
  NAND2xp33_ASAP7_75t_L     g00004(.A(\a[1] ), .B(new_n257), .Y(new_n261));
  NOR2xp33_ASAP7_75t_L      g00005(.A(new_n258), .B(new_n261), .Y(new_n262));
  INVx1_ASAP7_75t_L         g00006(.A(\a[1] ), .Y(new_n263));
  NAND2xp33_ASAP7_75t_L     g00007(.A(\a[2] ), .B(new_n263), .Y(new_n264));
  INVx1_ASAP7_75t_L         g00008(.A(\a[2] ), .Y(new_n265));
  NAND2xp33_ASAP7_75t_L     g00009(.A(\a[1] ), .B(new_n265), .Y(new_n266));
  NAND2xp33_ASAP7_75t_L     g00010(.A(new_n266), .B(new_n264), .Y(new_n267));
  INVx1_ASAP7_75t_L         g00011(.A(new_n267), .Y(new_n268));
  NOR2xp33_ASAP7_75t_L      g00012(.A(new_n257), .B(new_n268), .Y(new_n269));
  XNOR2x2_ASAP7_75t_L       g00013(.A(\b[1] ), .B(\b[0] ), .Y(new_n270));
  INVx1_ASAP7_75t_L         g00014(.A(new_n270), .Y(new_n271));
  NOR2xp33_ASAP7_75t_L      g00015(.A(new_n257), .B(new_n267), .Y(new_n272));
  AOI221xp5_ASAP7_75t_L     g00016(.A1(new_n272), .A2(\b[1] ), .B1(new_n271), .B2(new_n269), .C(new_n262), .Y(new_n273));
  XOR2x2_ASAP7_75t_L        g00017(.A(new_n260), .B(new_n273), .Y(\f[1] ));
  NAND2xp33_ASAP7_75t_L     g00018(.A(\a[2] ), .B(new_n273), .Y(new_n275));
  INVx1_ASAP7_75t_L         g00019(.A(\b[1] ), .Y(new_n276));
  NAND3xp33_ASAP7_75t_L     g00020(.A(new_n257), .B(new_n263), .C(\a[2] ), .Y(new_n277));
  INVx1_ASAP7_75t_L         g00021(.A(\b[2] ), .Y(new_n278));
  NAND3xp33_ASAP7_75t_L     g00022(.A(new_n278), .B(\b[1] ), .C(\b[0] ), .Y(new_n279));
  NAND2xp33_ASAP7_75t_L     g00023(.A(\b[1] ), .B(new_n278), .Y(new_n280));
  NAND2xp33_ASAP7_75t_L     g00024(.A(\b[2] ), .B(new_n276), .Y(new_n281));
  OAI211xp5_ASAP7_75t_L     g00025(.A1(new_n276), .A2(new_n258), .B(new_n280), .C(new_n281), .Y(new_n282));
  NAND2xp33_ASAP7_75t_L     g00026(.A(new_n279), .B(new_n282), .Y(new_n283));
  INVx1_ASAP7_75t_L         g00027(.A(new_n283), .Y(new_n284));
  AOI22xp33_ASAP7_75t_L     g00028(.A1(new_n272), .A2(\b[2] ), .B1(new_n269), .B2(new_n284), .Y(new_n285));
  OAI221xp5_ASAP7_75t_L     g00029(.A1(new_n261), .A2(new_n276), .B1(new_n258), .B2(new_n277), .C(new_n285), .Y(new_n286));
  O2A1O1Ixp33_ASAP7_75t_L   g00030(.A1(\f[0] ), .A2(new_n275), .B(\a[2] ), .C(new_n286), .Y(new_n287));
  O2A1O1Ixp33_ASAP7_75t_L   g00031(.A1(new_n258), .A2(new_n257), .B(new_n273), .C(new_n265), .Y(new_n288));
  AND2x2_ASAP7_75t_L        g00032(.A(new_n286), .B(new_n288), .Y(new_n289));
  NOR2xp33_ASAP7_75t_L      g00033(.A(new_n287), .B(new_n289), .Y(\f[2] ));
  INVx1_ASAP7_75t_L         g00034(.A(new_n277), .Y(new_n291));
  INVx1_ASAP7_75t_L         g00035(.A(new_n269), .Y(new_n292));
  NOR3xp33_ASAP7_75t_L      g00036(.A(new_n258), .B(new_n276), .C(\b[2] ), .Y(new_n293));
  NOR2xp33_ASAP7_75t_L      g00037(.A(\b[2] ), .B(\b[3] ), .Y(new_n294));
  NAND2xp33_ASAP7_75t_L     g00038(.A(\b[3] ), .B(\b[2] ), .Y(new_n295));
  INVx1_ASAP7_75t_L         g00039(.A(new_n295), .Y(new_n296));
  NOR2xp33_ASAP7_75t_L      g00040(.A(new_n294), .B(new_n296), .Y(new_n297));
  A2O1A1Ixp33_ASAP7_75t_L   g00041(.A1(\b[2] ), .A2(\b[1] ), .B(new_n293), .C(new_n297), .Y(new_n298));
  INVx1_ASAP7_75t_L         g00042(.A(\b[3] ), .Y(new_n299));
  NAND2xp33_ASAP7_75t_L     g00043(.A(new_n299), .B(new_n278), .Y(new_n300));
  NAND2xp33_ASAP7_75t_L     g00044(.A(new_n295), .B(new_n300), .Y(new_n301));
  A2O1A1Ixp33_ASAP7_75t_L   g00045(.A1(new_n278), .A2(new_n258), .B(new_n276), .C(new_n301), .Y(new_n302));
  NAND2xp33_ASAP7_75t_L     g00046(.A(new_n302), .B(new_n298), .Y(new_n303));
  NAND2xp33_ASAP7_75t_L     g00047(.A(\b[3] ), .B(new_n272), .Y(new_n304));
  OAI221xp5_ASAP7_75t_L     g00048(.A1(new_n261), .A2(new_n278), .B1(new_n303), .B2(new_n292), .C(new_n304), .Y(new_n305));
  AOI21xp33_ASAP7_75t_L     g00049(.A1(new_n291), .A2(\b[1] ), .B(new_n305), .Y(new_n306));
  NAND2xp33_ASAP7_75t_L     g00050(.A(\a[2] ), .B(new_n306), .Y(new_n307));
  A2O1A1Ixp33_ASAP7_75t_L   g00051(.A1(\b[1] ), .A2(new_n291), .B(new_n305), .C(new_n265), .Y(new_n308));
  NAND2xp33_ASAP7_75t_L     g00052(.A(new_n308), .B(new_n307), .Y(new_n309));
  INVx1_ASAP7_75t_L         g00053(.A(\a[3] ), .Y(new_n310));
  NAND2xp33_ASAP7_75t_L     g00054(.A(\a[2] ), .B(new_n310), .Y(new_n311));
  NAND2xp33_ASAP7_75t_L     g00055(.A(\a[3] ), .B(new_n265), .Y(new_n312));
  NAND2xp33_ASAP7_75t_L     g00056(.A(new_n312), .B(new_n311), .Y(new_n313));
  NAND2xp33_ASAP7_75t_L     g00057(.A(\b[0] ), .B(new_n313), .Y(new_n314));
  INVx1_ASAP7_75t_L         g00058(.A(new_n314), .Y(new_n315));
  XNOR2x2_ASAP7_75t_L       g00059(.A(new_n315), .B(new_n309), .Y(new_n316));
  NOR3xp33_ASAP7_75t_L      g00060(.A(new_n286), .B(new_n275), .C(\f[0] ), .Y(new_n317));
  XNOR2x2_ASAP7_75t_L       g00061(.A(new_n317), .B(new_n316), .Y(\f[3] ));
  OAI21xp33_ASAP7_75t_L     g00062(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n319));
  OAI21xp33_ASAP7_75t_L     g00063(.A1(new_n294), .A2(new_n319), .B(new_n295), .Y(new_n320));
  INVx1_ASAP7_75t_L         g00064(.A(new_n320), .Y(new_n321));
  NOR2xp33_ASAP7_75t_L      g00065(.A(\b[3] ), .B(\b[4] ), .Y(new_n322));
  INVx1_ASAP7_75t_L         g00066(.A(\b[4] ), .Y(new_n323));
  NOR2xp33_ASAP7_75t_L      g00067(.A(new_n299), .B(new_n323), .Y(new_n324));
  NOR3xp33_ASAP7_75t_L      g00068(.A(new_n321), .B(new_n322), .C(new_n324), .Y(new_n325));
  NOR2xp33_ASAP7_75t_L      g00069(.A(new_n322), .B(new_n324), .Y(new_n326));
  NOR2xp33_ASAP7_75t_L      g00070(.A(new_n320), .B(new_n326), .Y(new_n327));
  NOR2xp33_ASAP7_75t_L      g00071(.A(new_n327), .B(new_n325), .Y(new_n328));
  AOI22xp33_ASAP7_75t_L     g00072(.A1(new_n272), .A2(\b[4] ), .B1(new_n269), .B2(new_n328), .Y(new_n329));
  OAI221xp5_ASAP7_75t_L     g00073(.A1(new_n261), .A2(new_n299), .B1(new_n278), .B2(new_n277), .C(new_n329), .Y(new_n330));
  XNOR2x2_ASAP7_75t_L       g00074(.A(\a[2] ), .B(new_n330), .Y(new_n331));
  NAND2xp33_ASAP7_75t_L     g00075(.A(\a[5] ), .B(new_n315), .Y(new_n332));
  XNOR2x2_ASAP7_75t_L       g00076(.A(\a[4] ), .B(\a[3] ), .Y(new_n333));
  NOR2xp33_ASAP7_75t_L      g00077(.A(new_n333), .B(new_n313), .Y(new_n334));
  NAND2xp33_ASAP7_75t_L     g00078(.A(\b[0] ), .B(new_n334), .Y(new_n335));
  AND2x2_ASAP7_75t_L        g00079(.A(new_n311), .B(new_n312), .Y(new_n336));
  INVx1_ASAP7_75t_L         g00080(.A(\a[4] ), .Y(new_n337));
  NAND2xp33_ASAP7_75t_L     g00081(.A(\a[5] ), .B(new_n337), .Y(new_n338));
  INVx1_ASAP7_75t_L         g00082(.A(\a[5] ), .Y(new_n339));
  NAND2xp33_ASAP7_75t_L     g00083(.A(\a[4] ), .B(new_n339), .Y(new_n340));
  AND2x2_ASAP7_75t_L        g00084(.A(new_n338), .B(new_n340), .Y(new_n341));
  NOR2xp33_ASAP7_75t_L      g00085(.A(new_n336), .B(new_n341), .Y(new_n342));
  NAND2xp33_ASAP7_75t_L     g00086(.A(new_n271), .B(new_n342), .Y(new_n343));
  NAND2xp33_ASAP7_75t_L     g00087(.A(new_n340), .B(new_n338), .Y(new_n344));
  NOR2xp33_ASAP7_75t_L      g00088(.A(new_n344), .B(new_n336), .Y(new_n345));
  NAND2xp33_ASAP7_75t_L     g00089(.A(\b[1] ), .B(new_n345), .Y(new_n346));
  AND3x1_ASAP7_75t_L        g00090(.A(new_n343), .B(new_n346), .C(new_n335), .Y(new_n347));
  XNOR2x2_ASAP7_75t_L       g00091(.A(new_n332), .B(new_n347), .Y(new_n348));
  XOR2x2_ASAP7_75t_L        g00092(.A(new_n348), .B(new_n331), .Y(new_n349));
  MAJIxp5_ASAP7_75t_L       g00093(.A(new_n309), .B(new_n315), .C(new_n317), .Y(new_n350));
  XNOR2x2_ASAP7_75t_L       g00094(.A(new_n350), .B(new_n349), .Y(\f[4] ));
  NOR2xp33_ASAP7_75t_L      g00095(.A(\b[4] ), .B(\b[5] ), .Y(new_n352));
  INVx1_ASAP7_75t_L         g00096(.A(\b[5] ), .Y(new_n353));
  NOR2xp33_ASAP7_75t_L      g00097(.A(new_n323), .B(new_n353), .Y(new_n354));
  NOR2xp33_ASAP7_75t_L      g00098(.A(new_n352), .B(new_n354), .Y(new_n355));
  A2O1A1Ixp33_ASAP7_75t_L   g00099(.A1(new_n326), .A2(new_n320), .B(new_n324), .C(new_n355), .Y(new_n356));
  INVx1_ASAP7_75t_L         g00100(.A(new_n324), .Y(new_n357));
  OAI221xp5_ASAP7_75t_L     g00101(.A1(new_n354), .A2(new_n352), .B1(new_n322), .B2(new_n321), .C(new_n357), .Y(new_n358));
  NAND2xp33_ASAP7_75t_L     g00102(.A(new_n356), .B(new_n358), .Y(new_n359));
  INVx1_ASAP7_75t_L         g00103(.A(new_n359), .Y(new_n360));
  AOI22xp33_ASAP7_75t_L     g00104(.A1(new_n272), .A2(\b[5] ), .B1(new_n269), .B2(new_n360), .Y(new_n361));
  OAI221xp5_ASAP7_75t_L     g00105(.A1(new_n261), .A2(new_n323), .B1(new_n299), .B2(new_n277), .C(new_n361), .Y(new_n362));
  XNOR2x2_ASAP7_75t_L       g00106(.A(\a[2] ), .B(new_n362), .Y(new_n363));
  O2A1O1Ixp33_ASAP7_75t_L   g00107(.A1(new_n258), .A2(new_n336), .B(new_n347), .C(new_n339), .Y(new_n364));
  NAND3xp33_ASAP7_75t_L     g00108(.A(new_n336), .B(new_n333), .C(new_n344), .Y(new_n365));
  INVx1_ASAP7_75t_L         g00109(.A(new_n365), .Y(new_n366));
  NAND2xp33_ASAP7_75t_L     g00110(.A(new_n344), .B(new_n313), .Y(new_n367));
  NAND2xp33_ASAP7_75t_L     g00111(.A(new_n313), .B(new_n341), .Y(new_n368));
  NAND2xp33_ASAP7_75t_L     g00112(.A(\b[1] ), .B(new_n334), .Y(new_n369));
  OAI221xp5_ASAP7_75t_L     g00113(.A1(new_n367), .A2(new_n283), .B1(new_n278), .B2(new_n368), .C(new_n369), .Y(new_n370));
  A2O1A1Ixp33_ASAP7_75t_L   g00114(.A1(\b[0] ), .A2(new_n366), .B(new_n370), .C(new_n364), .Y(new_n371));
  AOI21xp33_ASAP7_75t_L     g00115(.A1(new_n366), .A2(\b[0] ), .B(new_n370), .Y(new_n372));
  A2O1A1Ixp33_ASAP7_75t_L   g00116(.A1(new_n314), .A2(new_n347), .B(new_n339), .C(new_n372), .Y(new_n373));
  NAND2xp33_ASAP7_75t_L     g00117(.A(new_n373), .B(new_n371), .Y(new_n374));
  XNOR2x2_ASAP7_75t_L       g00118(.A(new_n374), .B(new_n363), .Y(new_n375));
  MAJx2_ASAP7_75t_L         g00119(.A(new_n350), .B(new_n348), .C(new_n331), .Y(new_n376));
  XOR2x2_ASAP7_75t_L        g00120(.A(new_n376), .B(new_n375), .Y(\f[5] ));
  MAJIxp5_ASAP7_75t_L       g00121(.A(new_n376), .B(new_n363), .C(new_n374), .Y(new_n378));
  NAND2xp33_ASAP7_75t_L     g00122(.A(\b[4] ), .B(new_n291), .Y(new_n379));
  INVx1_ASAP7_75t_L         g00123(.A(new_n261), .Y(new_n380));
  NAND2xp33_ASAP7_75t_L     g00124(.A(\b[5] ), .B(new_n380), .Y(new_n381));
  INVx1_ASAP7_75t_L         g00125(.A(\b[6] ), .Y(new_n382));
  NAND2xp33_ASAP7_75t_L     g00126(.A(new_n382), .B(new_n353), .Y(new_n383));
  NAND2xp33_ASAP7_75t_L     g00127(.A(\b[6] ), .B(\b[5] ), .Y(new_n384));
  NAND2xp33_ASAP7_75t_L     g00128(.A(new_n384), .B(new_n383), .Y(new_n385));
  O2A1O1Ixp33_ASAP7_75t_L   g00129(.A1(new_n323), .A2(new_n353), .B(new_n356), .C(new_n385), .Y(new_n386));
  A2O1A1O1Ixp25_ASAP7_75t_L g00130(.A1(new_n320), .A2(new_n326), .B(new_n324), .C(new_n355), .D(new_n354), .Y(new_n387));
  AND2x2_ASAP7_75t_L        g00131(.A(new_n385), .B(new_n387), .Y(new_n388));
  NOR2xp33_ASAP7_75t_L      g00132(.A(new_n386), .B(new_n388), .Y(new_n389));
  AOI22xp33_ASAP7_75t_L     g00133(.A1(new_n272), .A2(\b[6] ), .B1(new_n269), .B2(new_n389), .Y(new_n390));
  NAND4xp25_ASAP7_75t_L     g00134(.A(new_n390), .B(\a[2] ), .C(new_n379), .D(new_n381), .Y(new_n391));
  NAND2xp33_ASAP7_75t_L     g00135(.A(new_n381), .B(new_n390), .Y(new_n392));
  A2O1A1Ixp33_ASAP7_75t_L   g00136(.A1(\b[4] ), .A2(new_n291), .B(new_n392), .C(new_n265), .Y(new_n393));
  AND2x2_ASAP7_75t_L        g00137(.A(new_n391), .B(new_n393), .Y(new_n394));
  INVx1_ASAP7_75t_L         g00138(.A(\a[6] ), .Y(new_n395));
  NAND2xp33_ASAP7_75t_L     g00139(.A(\a[5] ), .B(new_n395), .Y(new_n396));
  NAND2xp33_ASAP7_75t_L     g00140(.A(\a[6] ), .B(new_n339), .Y(new_n397));
  NAND3xp33_ASAP7_75t_L     g00141(.A(new_n347), .B(new_n314), .C(\a[5] ), .Y(new_n398));
  INVx1_ASAP7_75t_L         g00142(.A(new_n372), .Y(new_n399));
  NOR2xp33_ASAP7_75t_L      g00143(.A(new_n398), .B(new_n399), .Y(new_n400));
  A2O1A1Ixp33_ASAP7_75t_L   g00144(.A1(new_n396), .A2(new_n397), .B(new_n258), .C(new_n400), .Y(new_n401));
  AND2x2_ASAP7_75t_L        g00145(.A(new_n396), .B(new_n397), .Y(new_n402));
  NOR2xp33_ASAP7_75t_L      g00146(.A(new_n258), .B(new_n402), .Y(new_n403));
  OAI21xp33_ASAP7_75t_L     g00147(.A1(new_n399), .A2(new_n398), .B(new_n403), .Y(new_n404));
  NAND2xp33_ASAP7_75t_L     g00148(.A(new_n404), .B(new_n401), .Y(new_n405));
  INVx1_ASAP7_75t_L         g00149(.A(new_n334), .Y(new_n406));
  NAND2xp33_ASAP7_75t_L     g00150(.A(\b[3] ), .B(new_n345), .Y(new_n407));
  OAI221xp5_ASAP7_75t_L     g00151(.A1(new_n278), .A2(new_n406), .B1(new_n367), .B2(new_n303), .C(new_n407), .Y(new_n408));
  AOI21xp33_ASAP7_75t_L     g00152(.A1(new_n366), .A2(\b[1] ), .B(new_n408), .Y(new_n409));
  NAND2xp33_ASAP7_75t_L     g00153(.A(\a[5] ), .B(new_n409), .Y(new_n410));
  A2O1A1Ixp33_ASAP7_75t_L   g00154(.A1(\b[1] ), .A2(new_n366), .B(new_n408), .C(new_n339), .Y(new_n411));
  NAND2xp33_ASAP7_75t_L     g00155(.A(new_n411), .B(new_n410), .Y(new_n412));
  XNOR2x2_ASAP7_75t_L       g00156(.A(new_n412), .B(new_n405), .Y(new_n413));
  NOR2xp33_ASAP7_75t_L      g00157(.A(new_n394), .B(new_n413), .Y(new_n414));
  INVx1_ASAP7_75t_L         g00158(.A(new_n414), .Y(new_n415));
  NAND2xp33_ASAP7_75t_L     g00159(.A(new_n394), .B(new_n413), .Y(new_n416));
  AND3x1_ASAP7_75t_L        g00160(.A(new_n415), .B(new_n416), .C(new_n378), .Y(new_n417));
  AOI21xp33_ASAP7_75t_L     g00161(.A1(new_n415), .A2(new_n416), .B(new_n378), .Y(new_n418));
  NOR2xp33_ASAP7_75t_L      g00162(.A(new_n418), .B(new_n417), .Y(\f[6] ));
  NOR2xp33_ASAP7_75t_L      g00163(.A(\b[6] ), .B(\b[7] ), .Y(new_n420));
  INVx1_ASAP7_75t_L         g00164(.A(\b[7] ), .Y(new_n421));
  NOR2xp33_ASAP7_75t_L      g00165(.A(new_n382), .B(new_n421), .Y(new_n422));
  NOR2xp33_ASAP7_75t_L      g00166(.A(new_n420), .B(new_n422), .Y(new_n423));
  A2O1A1Ixp33_ASAP7_75t_L   g00167(.A1(\b[6] ), .A2(\b[5] ), .B(new_n386), .C(new_n423), .Y(new_n424));
  INVx1_ASAP7_75t_L         g00168(.A(new_n423), .Y(new_n425));
  OAI211xp5_ASAP7_75t_L     g00169(.A1(new_n385), .A2(new_n387), .B(new_n384), .C(new_n425), .Y(new_n426));
  NAND2xp33_ASAP7_75t_L     g00170(.A(new_n426), .B(new_n424), .Y(new_n427));
  NAND2xp33_ASAP7_75t_L     g00171(.A(\b[7] ), .B(new_n272), .Y(new_n428));
  OAI221xp5_ASAP7_75t_L     g00172(.A1(new_n382), .A2(new_n261), .B1(new_n292), .B2(new_n427), .C(new_n428), .Y(new_n429));
  AOI21xp33_ASAP7_75t_L     g00173(.A1(new_n291), .A2(\b[5] ), .B(new_n429), .Y(new_n430));
  NAND2xp33_ASAP7_75t_L     g00174(.A(\a[2] ), .B(new_n430), .Y(new_n431));
  A2O1A1Ixp33_ASAP7_75t_L   g00175(.A1(\b[5] ), .A2(new_n291), .B(new_n429), .C(new_n265), .Y(new_n432));
  NAND2xp33_ASAP7_75t_L     g00176(.A(\b[3] ), .B(new_n334), .Y(new_n433));
  OAI221xp5_ASAP7_75t_L     g00177(.A1(new_n368), .A2(new_n323), .B1(new_n278), .B2(new_n365), .C(new_n433), .Y(new_n434));
  AOI21xp33_ASAP7_75t_L     g00178(.A1(new_n328), .A2(new_n342), .B(new_n434), .Y(new_n435));
  NAND2xp33_ASAP7_75t_L     g00179(.A(\a[5] ), .B(new_n435), .Y(new_n436));
  A2O1A1Ixp33_ASAP7_75t_L   g00180(.A1(new_n328), .A2(new_n342), .B(new_n434), .C(new_n339), .Y(new_n437));
  NAND2xp33_ASAP7_75t_L     g00181(.A(\a[8] ), .B(new_n403), .Y(new_n438));
  NAND2xp33_ASAP7_75t_L     g00182(.A(new_n397), .B(new_n396), .Y(new_n439));
  XNOR2x2_ASAP7_75t_L       g00183(.A(\a[7] ), .B(\a[6] ), .Y(new_n440));
  NOR2xp33_ASAP7_75t_L      g00184(.A(new_n440), .B(new_n439), .Y(new_n441));
  NAND2xp33_ASAP7_75t_L     g00185(.A(\b[0] ), .B(new_n441), .Y(new_n442));
  INVx1_ASAP7_75t_L         g00186(.A(\a[7] ), .Y(new_n443));
  NAND2xp33_ASAP7_75t_L     g00187(.A(\a[8] ), .B(new_n443), .Y(new_n444));
  INVx1_ASAP7_75t_L         g00188(.A(\a[8] ), .Y(new_n445));
  NAND2xp33_ASAP7_75t_L     g00189(.A(\a[7] ), .B(new_n445), .Y(new_n446));
  AND2x2_ASAP7_75t_L        g00190(.A(new_n444), .B(new_n446), .Y(new_n447));
  NOR2xp33_ASAP7_75t_L      g00191(.A(new_n402), .B(new_n447), .Y(new_n448));
  NAND2xp33_ASAP7_75t_L     g00192(.A(new_n271), .B(new_n448), .Y(new_n449));
  NAND2xp33_ASAP7_75t_L     g00193(.A(new_n446), .B(new_n444), .Y(new_n450));
  NOR2xp33_ASAP7_75t_L      g00194(.A(new_n450), .B(new_n402), .Y(new_n451));
  NAND2xp33_ASAP7_75t_L     g00195(.A(\b[1] ), .B(new_n451), .Y(new_n452));
  NAND3xp33_ASAP7_75t_L     g00196(.A(new_n449), .B(new_n452), .C(new_n442), .Y(new_n453));
  XNOR2x2_ASAP7_75t_L       g00197(.A(new_n438), .B(new_n453), .Y(new_n454));
  NAND3xp33_ASAP7_75t_L     g00198(.A(new_n454), .B(new_n437), .C(new_n436), .Y(new_n455));
  INVx1_ASAP7_75t_L         g00199(.A(new_n436), .Y(new_n456));
  INVx1_ASAP7_75t_L         g00200(.A(new_n437), .Y(new_n457));
  INVx1_ASAP7_75t_L         g00201(.A(new_n454), .Y(new_n458));
  OAI21xp33_ASAP7_75t_L     g00202(.A1(new_n456), .A2(new_n457), .B(new_n458), .Y(new_n459));
  MAJIxp5_ASAP7_75t_L       g00203(.A(new_n412), .B(new_n403), .C(new_n400), .Y(new_n460));
  AOI21xp33_ASAP7_75t_L     g00204(.A1(new_n459), .A2(new_n455), .B(new_n460), .Y(new_n461));
  NAND2xp33_ASAP7_75t_L     g00205(.A(new_n455), .B(new_n459), .Y(new_n462));
  INVx1_ASAP7_75t_L         g00206(.A(new_n460), .Y(new_n463));
  NOR2xp33_ASAP7_75t_L      g00207(.A(new_n462), .B(new_n463), .Y(new_n464));
  AOI211xp5_ASAP7_75t_L     g00208(.A1(new_n431), .A2(new_n432), .B(new_n461), .C(new_n464), .Y(new_n465));
  INVx1_ASAP7_75t_L         g00209(.A(new_n465), .Y(new_n466));
  OAI211xp5_ASAP7_75t_L     g00210(.A1(new_n461), .A2(new_n464), .B(new_n431), .C(new_n432), .Y(new_n467));
  NAND2xp33_ASAP7_75t_L     g00211(.A(new_n467), .B(new_n466), .Y(new_n468));
  INVx1_ASAP7_75t_L         g00212(.A(new_n468), .Y(new_n469));
  A2O1A1Ixp33_ASAP7_75t_L   g00213(.A1(new_n416), .A2(new_n378), .B(new_n414), .C(new_n469), .Y(new_n470));
  OR3x1_ASAP7_75t_L         g00214(.A(new_n469), .B(new_n417), .C(new_n414), .Y(new_n471));
  AND2x2_ASAP7_75t_L        g00215(.A(new_n470), .B(new_n471), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g00216(.A(new_n353), .B(new_n368), .Y(new_n473));
  AOI221xp5_ASAP7_75t_L     g00217(.A1(new_n334), .A2(\b[4] ), .B1(new_n366), .B2(\b[3] ), .C(new_n473), .Y(new_n474));
  OAI211xp5_ASAP7_75t_L     g00218(.A1(new_n367), .A2(new_n359), .B(new_n474), .C(\a[5] ), .Y(new_n475));
  INVx1_ASAP7_75t_L         g00219(.A(new_n475), .Y(new_n476));
  O2A1O1Ixp33_ASAP7_75t_L   g00220(.A1(new_n367), .A2(new_n359), .B(new_n474), .C(\a[5] ), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g00221(.A(new_n477), .B(new_n476), .Y(new_n478));
  INVx1_ASAP7_75t_L         g00222(.A(new_n440), .Y(new_n479));
  NOR3xp33_ASAP7_75t_L      g00223(.A(new_n447), .B(new_n479), .C(new_n439), .Y(new_n480));
  INVx1_ASAP7_75t_L         g00224(.A(new_n480), .Y(new_n481));
  NAND2xp33_ASAP7_75t_L     g00225(.A(new_n450), .B(new_n439), .Y(new_n482));
  NOR2xp33_ASAP7_75t_L      g00226(.A(new_n482), .B(new_n283), .Y(new_n483));
  AOI221xp5_ASAP7_75t_L     g00227(.A1(\b[2] ), .A2(new_n451), .B1(new_n441), .B2(\b[1] ), .C(new_n483), .Y(new_n484));
  OAI21xp33_ASAP7_75t_L     g00228(.A1(new_n258), .A2(new_n481), .B(new_n484), .Y(new_n485));
  O2A1O1Ixp33_ASAP7_75t_L   g00229(.A1(new_n403), .A2(new_n453), .B(\a[8] ), .C(new_n485), .Y(new_n486));
  INVx1_ASAP7_75t_L         g00230(.A(new_n486), .Y(new_n487));
  A2O1A1Ixp33_ASAP7_75t_L   g00231(.A1(\b[0] ), .A2(new_n439), .B(new_n453), .C(\a[8] ), .Y(new_n488));
  O2A1O1Ixp33_ASAP7_75t_L   g00232(.A1(new_n481), .A2(new_n258), .B(new_n484), .C(new_n488), .Y(new_n489));
  INVx1_ASAP7_75t_L         g00233(.A(new_n489), .Y(new_n490));
  NAND3xp33_ASAP7_75t_L     g00234(.A(new_n478), .B(new_n490), .C(new_n487), .Y(new_n491));
  INVx1_ASAP7_75t_L         g00235(.A(new_n477), .Y(new_n492));
  NAND2xp33_ASAP7_75t_L     g00236(.A(new_n475), .B(new_n492), .Y(new_n493));
  OAI21xp33_ASAP7_75t_L     g00237(.A1(new_n486), .A2(new_n489), .B(new_n493), .Y(new_n494));
  O2A1O1Ixp33_ASAP7_75t_L   g00238(.A1(new_n456), .A2(new_n457), .B(new_n454), .C(new_n461), .Y(new_n495));
  NAND3xp33_ASAP7_75t_L     g00239(.A(new_n495), .B(new_n494), .C(new_n491), .Y(new_n496));
  NAND2xp33_ASAP7_75t_L     g00240(.A(new_n494), .B(new_n491), .Y(new_n497));
  AOI21xp33_ASAP7_75t_L     g00241(.A1(new_n436), .A2(new_n437), .B(new_n458), .Y(new_n498));
  A2O1A1Ixp33_ASAP7_75t_L   g00242(.A1(new_n462), .A2(new_n463), .B(new_n498), .C(new_n497), .Y(new_n499));
  NAND2xp33_ASAP7_75t_L     g00243(.A(new_n499), .B(new_n496), .Y(new_n500));
  O2A1O1Ixp33_ASAP7_75t_L   g00244(.A1(new_n385), .A2(new_n387), .B(new_n384), .C(new_n425), .Y(new_n501));
  NOR2xp33_ASAP7_75t_L      g00245(.A(\b[7] ), .B(\b[8] ), .Y(new_n502));
  INVx1_ASAP7_75t_L         g00246(.A(\b[8] ), .Y(new_n503));
  NOR2xp33_ASAP7_75t_L      g00247(.A(new_n421), .B(new_n503), .Y(new_n504));
  NOR2xp33_ASAP7_75t_L      g00248(.A(new_n502), .B(new_n504), .Y(new_n505));
  A2O1A1Ixp33_ASAP7_75t_L   g00249(.A1(\b[7] ), .A2(\b[6] ), .B(new_n501), .C(new_n505), .Y(new_n506));
  A2O1A1O1Ixp25_ASAP7_75t_L g00250(.A1(\b[6] ), .A2(\b[5] ), .B(new_n386), .C(new_n423), .D(new_n422), .Y(new_n507));
  OAI21xp33_ASAP7_75t_L     g00251(.A1(new_n502), .A2(new_n504), .B(new_n507), .Y(new_n508));
  NAND2xp33_ASAP7_75t_L     g00252(.A(new_n506), .B(new_n508), .Y(new_n509));
  INVx1_ASAP7_75t_L         g00253(.A(new_n509), .Y(new_n510));
  AOI22xp33_ASAP7_75t_L     g00254(.A1(new_n272), .A2(\b[8] ), .B1(new_n269), .B2(new_n510), .Y(new_n511));
  OAI221xp5_ASAP7_75t_L     g00255(.A1(new_n261), .A2(new_n421), .B1(new_n382), .B2(new_n277), .C(new_n511), .Y(new_n512));
  XNOR2x2_ASAP7_75t_L       g00256(.A(\a[2] ), .B(new_n512), .Y(new_n513));
  XNOR2x2_ASAP7_75t_L       g00257(.A(new_n513), .B(new_n500), .Y(new_n514));
  A2O1A1O1Ixp25_ASAP7_75t_L g00258(.A1(new_n378), .A2(new_n416), .B(new_n414), .C(new_n467), .D(new_n465), .Y(new_n515));
  XOR2x2_ASAP7_75t_L        g00259(.A(new_n515), .B(new_n514), .Y(\f[8] ));
  INVx1_ASAP7_75t_L         g00260(.A(new_n403), .Y(new_n517));
  NAND5xp2_ASAP7_75t_L      g00261(.A(new_n452), .B(new_n449), .C(new_n442), .D(new_n517), .E(\a[8] ), .Y(new_n518));
  INVx1_ASAP7_75t_L         g00262(.A(\a[9] ), .Y(new_n519));
  NAND2xp33_ASAP7_75t_L     g00263(.A(\a[8] ), .B(new_n519), .Y(new_n520));
  NAND2xp33_ASAP7_75t_L     g00264(.A(\a[9] ), .B(new_n445), .Y(new_n521));
  AND2x2_ASAP7_75t_L        g00265(.A(new_n520), .B(new_n521), .Y(new_n522));
  NOR2xp33_ASAP7_75t_L      g00266(.A(new_n258), .B(new_n522), .Y(new_n523));
  OAI21xp33_ASAP7_75t_L     g00267(.A1(new_n518), .A2(new_n485), .B(new_n523), .Y(new_n524));
  INVx1_ASAP7_75t_L         g00268(.A(new_n518), .Y(new_n525));
  NAND2xp33_ASAP7_75t_L     g00269(.A(\b[0] ), .B(new_n480), .Y(new_n526));
  INVx1_ASAP7_75t_L         g00270(.A(new_n523), .Y(new_n527));
  NAND4xp25_ASAP7_75t_L     g00271(.A(new_n525), .B(new_n527), .C(new_n484), .D(new_n526), .Y(new_n528));
  INVx1_ASAP7_75t_L         g00272(.A(new_n441), .Y(new_n529));
  NAND2xp33_ASAP7_75t_L     g00273(.A(\b[3] ), .B(new_n451), .Y(new_n530));
  OAI221xp5_ASAP7_75t_L     g00274(.A1(new_n278), .A2(new_n529), .B1(new_n482), .B2(new_n303), .C(new_n530), .Y(new_n531));
  AOI21xp33_ASAP7_75t_L     g00275(.A1(new_n480), .A2(\b[1] ), .B(new_n531), .Y(new_n532));
  NAND2xp33_ASAP7_75t_L     g00276(.A(\a[8] ), .B(new_n532), .Y(new_n533));
  A2O1A1Ixp33_ASAP7_75t_L   g00277(.A1(\b[1] ), .A2(new_n480), .B(new_n531), .C(new_n445), .Y(new_n534));
  AOI22xp33_ASAP7_75t_L     g00278(.A1(new_n533), .A2(new_n534), .B1(new_n528), .B2(new_n524), .Y(new_n535));
  NAND4xp25_ASAP7_75t_L     g00279(.A(new_n524), .B(new_n528), .C(new_n533), .D(new_n534), .Y(new_n536));
  INVx1_ASAP7_75t_L         g00280(.A(new_n536), .Y(new_n537));
  INVx1_ASAP7_75t_L         g00281(.A(new_n386), .Y(new_n538));
  NAND2xp33_ASAP7_75t_L     g00282(.A(new_n385), .B(new_n387), .Y(new_n539));
  NAND2xp33_ASAP7_75t_L     g00283(.A(new_n539), .B(new_n538), .Y(new_n540));
  NOR2xp33_ASAP7_75t_L      g00284(.A(new_n382), .B(new_n368), .Y(new_n541));
  AOI221xp5_ASAP7_75t_L     g00285(.A1(new_n334), .A2(\b[5] ), .B1(new_n366), .B2(\b[4] ), .C(new_n541), .Y(new_n542));
  OAI211xp5_ASAP7_75t_L     g00286(.A1(new_n367), .A2(new_n540), .B(\a[5] ), .C(new_n542), .Y(new_n543));
  INVx1_ASAP7_75t_L         g00287(.A(new_n542), .Y(new_n544));
  A2O1A1Ixp33_ASAP7_75t_L   g00288(.A1(new_n389), .A2(new_n342), .B(new_n544), .C(new_n339), .Y(new_n545));
  NAND2xp33_ASAP7_75t_L     g00289(.A(new_n545), .B(new_n543), .Y(new_n546));
  NOR3xp33_ASAP7_75t_L      g00290(.A(new_n537), .B(new_n546), .C(new_n535), .Y(new_n547));
  AO22x1_ASAP7_75t_L        g00291(.A1(new_n534), .A2(new_n533), .B1(new_n528), .B2(new_n524), .Y(new_n548));
  AOI22xp33_ASAP7_75t_L     g00292(.A1(new_n543), .A2(new_n545), .B1(new_n536), .B2(new_n548), .Y(new_n549));
  NOR2xp33_ASAP7_75t_L      g00293(.A(new_n549), .B(new_n547), .Y(new_n550));
  NOR3xp33_ASAP7_75t_L      g00294(.A(new_n478), .B(new_n486), .C(new_n489), .Y(new_n551));
  A2O1A1O1Ixp25_ASAP7_75t_L g00295(.A1(new_n462), .A2(new_n463), .B(new_n498), .C(new_n497), .D(new_n551), .Y(new_n552));
  NAND2xp33_ASAP7_75t_L     g00296(.A(new_n550), .B(new_n552), .Y(new_n553));
  INVx1_ASAP7_75t_L         g00297(.A(new_n551), .Y(new_n554));
  AO21x2_ASAP7_75t_L        g00298(.A1(new_n554), .A2(new_n499), .B(new_n550), .Y(new_n555));
  INVx1_ASAP7_75t_L         g00299(.A(new_n422), .Y(new_n556));
  INVx1_ASAP7_75t_L         g00300(.A(new_n504), .Y(new_n557));
  NOR2xp33_ASAP7_75t_L      g00301(.A(\b[8] ), .B(\b[9] ), .Y(new_n558));
  INVx1_ASAP7_75t_L         g00302(.A(\b[9] ), .Y(new_n559));
  NOR2xp33_ASAP7_75t_L      g00303(.A(new_n503), .B(new_n559), .Y(new_n560));
  NOR2xp33_ASAP7_75t_L      g00304(.A(new_n558), .B(new_n560), .Y(new_n561));
  INVx1_ASAP7_75t_L         g00305(.A(new_n561), .Y(new_n562));
  A2O1A1O1Ixp25_ASAP7_75t_L g00306(.A1(new_n556), .A2(new_n424), .B(new_n502), .C(new_n557), .D(new_n562), .Y(new_n563));
  A2O1A1Ixp33_ASAP7_75t_L   g00307(.A1(new_n424), .A2(new_n556), .B(new_n502), .C(new_n557), .Y(new_n564));
  NOR2xp33_ASAP7_75t_L      g00308(.A(new_n561), .B(new_n564), .Y(new_n565));
  NOR2xp33_ASAP7_75t_L      g00309(.A(new_n563), .B(new_n565), .Y(new_n566));
  AOI22xp33_ASAP7_75t_L     g00310(.A1(new_n272), .A2(\b[9] ), .B1(new_n269), .B2(new_n566), .Y(new_n567));
  OAI221xp5_ASAP7_75t_L     g00311(.A1(new_n261), .A2(new_n503), .B1(new_n421), .B2(new_n277), .C(new_n567), .Y(new_n568));
  NOR2xp33_ASAP7_75t_L      g00312(.A(new_n265), .B(new_n568), .Y(new_n569));
  INVx1_ASAP7_75t_L         g00313(.A(new_n569), .Y(new_n570));
  NAND2xp33_ASAP7_75t_L     g00314(.A(new_n265), .B(new_n568), .Y(new_n571));
  NAND4xp25_ASAP7_75t_L     g00315(.A(new_n570), .B(new_n553), .C(new_n555), .D(new_n571), .Y(new_n572));
  AO22x1_ASAP7_75t_L        g00316(.A1(new_n553), .A2(new_n555), .B1(new_n571), .B2(new_n570), .Y(new_n573));
  NAND2xp33_ASAP7_75t_L     g00317(.A(new_n572), .B(new_n573), .Y(new_n574));
  MAJIxp5_ASAP7_75t_L       g00318(.A(new_n515), .B(new_n500), .C(new_n513), .Y(new_n575));
  XOR2x2_ASAP7_75t_L        g00319(.A(new_n575), .B(new_n574), .Y(\f[9] ));
  NAND2xp33_ASAP7_75t_L     g00320(.A(new_n553), .B(new_n555), .Y(new_n577));
  AND2x2_ASAP7_75t_L        g00321(.A(new_n571), .B(new_n570), .Y(new_n578));
  NAND2xp33_ASAP7_75t_L     g00322(.A(new_n575), .B(new_n574), .Y(new_n579));
  NOR3xp33_ASAP7_75t_L      g00323(.A(new_n485), .B(new_n527), .C(new_n518), .Y(new_n580));
  NAND2xp33_ASAP7_75t_L     g00324(.A(\b[2] ), .B(new_n480), .Y(new_n581));
  NAND2xp33_ASAP7_75t_L     g00325(.A(\b[3] ), .B(new_n441), .Y(new_n582));
  AOI22xp33_ASAP7_75t_L     g00326(.A1(new_n451), .A2(\b[4] ), .B1(new_n448), .B2(new_n328), .Y(new_n583));
  NAND4xp25_ASAP7_75t_L     g00327(.A(new_n583), .B(\a[8] ), .C(new_n581), .D(new_n582), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(new_n582), .B(new_n583), .Y(new_n585));
  A2O1A1Ixp33_ASAP7_75t_L   g00329(.A1(\b[2] ), .A2(new_n480), .B(new_n585), .C(new_n445), .Y(new_n586));
  NAND2xp33_ASAP7_75t_L     g00330(.A(\a[11] ), .B(new_n523), .Y(new_n587));
  NAND2xp33_ASAP7_75t_L     g00331(.A(new_n521), .B(new_n520), .Y(new_n588));
  XNOR2x2_ASAP7_75t_L       g00332(.A(\a[10] ), .B(\a[9] ), .Y(new_n589));
  NOR2xp33_ASAP7_75t_L      g00333(.A(new_n589), .B(new_n588), .Y(new_n590));
  NAND2xp33_ASAP7_75t_L     g00334(.A(\b[0] ), .B(new_n590), .Y(new_n591));
  INVx1_ASAP7_75t_L         g00335(.A(\a[10] ), .Y(new_n592));
  NAND2xp33_ASAP7_75t_L     g00336(.A(\a[11] ), .B(new_n592), .Y(new_n593));
  INVx1_ASAP7_75t_L         g00337(.A(\a[11] ), .Y(new_n594));
  NAND2xp33_ASAP7_75t_L     g00338(.A(\a[10] ), .B(new_n594), .Y(new_n595));
  AND2x2_ASAP7_75t_L        g00339(.A(new_n593), .B(new_n595), .Y(new_n596));
  NOR2xp33_ASAP7_75t_L      g00340(.A(new_n522), .B(new_n596), .Y(new_n597));
  NAND2xp33_ASAP7_75t_L     g00341(.A(new_n271), .B(new_n597), .Y(new_n598));
  NAND2xp33_ASAP7_75t_L     g00342(.A(new_n595), .B(new_n593), .Y(new_n599));
  NOR2xp33_ASAP7_75t_L      g00343(.A(new_n599), .B(new_n522), .Y(new_n600));
  NAND2xp33_ASAP7_75t_L     g00344(.A(\b[1] ), .B(new_n600), .Y(new_n601));
  AND3x1_ASAP7_75t_L        g00345(.A(new_n598), .B(new_n601), .C(new_n591), .Y(new_n602));
  XNOR2x2_ASAP7_75t_L       g00346(.A(new_n587), .B(new_n602), .Y(new_n603));
  NAND3xp33_ASAP7_75t_L     g00347(.A(new_n586), .B(new_n584), .C(new_n603), .Y(new_n604));
  AO21x2_ASAP7_75t_L        g00348(.A1(new_n584), .A2(new_n586), .B(new_n603), .Y(new_n605));
  OAI211xp5_ASAP7_75t_L     g00349(.A1(new_n535), .A2(new_n580), .B(new_n605), .C(new_n604), .Y(new_n606));
  NOR2xp33_ASAP7_75t_L      g00350(.A(new_n580), .B(new_n535), .Y(new_n607));
  AND3x1_ASAP7_75t_L        g00351(.A(new_n586), .B(new_n603), .C(new_n584), .Y(new_n608));
  AOI21xp33_ASAP7_75t_L     g00352(.A1(new_n586), .A2(new_n584), .B(new_n603), .Y(new_n609));
  OAI21xp33_ASAP7_75t_L     g00353(.A1(new_n608), .A2(new_n609), .B(new_n607), .Y(new_n610));
  INVx1_ASAP7_75t_L         g00354(.A(new_n427), .Y(new_n611));
  NAND2xp33_ASAP7_75t_L     g00355(.A(\b[6] ), .B(new_n334), .Y(new_n612));
  OAI221xp5_ASAP7_75t_L     g00356(.A1(new_n368), .A2(new_n421), .B1(new_n353), .B2(new_n365), .C(new_n612), .Y(new_n613));
  AOI21xp33_ASAP7_75t_L     g00357(.A1(new_n611), .A2(new_n342), .B(new_n613), .Y(new_n614));
  NAND2xp33_ASAP7_75t_L     g00358(.A(\a[5] ), .B(new_n614), .Y(new_n615));
  A2O1A1Ixp33_ASAP7_75t_L   g00359(.A1(new_n611), .A2(new_n342), .B(new_n613), .C(new_n339), .Y(new_n616));
  AND2x2_ASAP7_75t_L        g00360(.A(new_n616), .B(new_n615), .Y(new_n617));
  NAND3xp33_ASAP7_75t_L     g00361(.A(new_n617), .B(new_n610), .C(new_n606), .Y(new_n618));
  NOR3xp33_ASAP7_75t_L      g00362(.A(new_n607), .B(new_n608), .C(new_n609), .Y(new_n619));
  AOI211xp5_ASAP7_75t_L     g00363(.A1(new_n605), .A2(new_n604), .B(new_n535), .C(new_n580), .Y(new_n620));
  NAND2xp33_ASAP7_75t_L     g00364(.A(new_n616), .B(new_n615), .Y(new_n621));
  OAI21xp33_ASAP7_75t_L     g00365(.A1(new_n620), .A2(new_n619), .B(new_n621), .Y(new_n622));
  NAND2xp33_ASAP7_75t_L     g00366(.A(new_n618), .B(new_n622), .Y(new_n623));
  NAND3xp33_ASAP7_75t_L     g00367(.A(new_n548), .B(new_n536), .C(new_n546), .Y(new_n624));
  A2O1A1Ixp33_ASAP7_75t_L   g00368(.A1(new_n499), .A2(new_n554), .B(new_n550), .C(new_n624), .Y(new_n625));
  NOR2xp33_ASAP7_75t_L      g00369(.A(new_n623), .B(new_n625), .Y(new_n626));
  INVx1_ASAP7_75t_L         g00370(.A(new_n623), .Y(new_n627));
  O2A1O1Ixp33_ASAP7_75t_L   g00371(.A1(new_n552), .A2(new_n550), .B(new_n624), .C(new_n627), .Y(new_n628));
  NOR2xp33_ASAP7_75t_L      g00372(.A(new_n503), .B(new_n277), .Y(new_n629));
  NOR2xp33_ASAP7_75t_L      g00373(.A(new_n559), .B(new_n261), .Y(new_n630));
  INVx1_ASAP7_75t_L         g00374(.A(\b[10] ), .Y(new_n631));
  INVx1_ASAP7_75t_L         g00375(.A(new_n272), .Y(new_n632));
  NOR2xp33_ASAP7_75t_L      g00376(.A(\b[9] ), .B(\b[10] ), .Y(new_n633));
  NOR2xp33_ASAP7_75t_L      g00377(.A(new_n559), .B(new_n631), .Y(new_n634));
  NOR2xp33_ASAP7_75t_L      g00378(.A(new_n633), .B(new_n634), .Y(new_n635));
  A2O1A1Ixp33_ASAP7_75t_L   g00379(.A1(new_n564), .A2(new_n561), .B(new_n560), .C(new_n635), .Y(new_n636));
  INVx1_ASAP7_75t_L         g00380(.A(new_n560), .Y(new_n637));
  A2O1A1Ixp33_ASAP7_75t_L   g00381(.A1(new_n506), .A2(new_n557), .B(new_n558), .C(new_n637), .Y(new_n638));
  NOR2xp33_ASAP7_75t_L      g00382(.A(new_n635), .B(new_n638), .Y(new_n639));
  INVx1_ASAP7_75t_L         g00383(.A(new_n639), .Y(new_n640));
  NAND2xp33_ASAP7_75t_L     g00384(.A(new_n636), .B(new_n640), .Y(new_n641));
  OAI22xp33_ASAP7_75t_L     g00385(.A1(new_n641), .A2(new_n292), .B1(new_n631), .B2(new_n632), .Y(new_n642));
  NOR4xp25_ASAP7_75t_L      g00386(.A(new_n642), .B(new_n265), .C(new_n629), .D(new_n630), .Y(new_n643));
  NOR2xp33_ASAP7_75t_L      g00387(.A(new_n630), .B(new_n642), .Y(new_n644));
  O2A1O1Ixp33_ASAP7_75t_L   g00388(.A1(new_n503), .A2(new_n277), .B(new_n644), .C(\a[2] ), .Y(new_n645));
  NOR2xp33_ASAP7_75t_L      g00389(.A(new_n643), .B(new_n645), .Y(new_n646));
  OAI21xp33_ASAP7_75t_L     g00390(.A1(new_n626), .A2(new_n628), .B(new_n646), .Y(new_n647));
  NOR3xp33_ASAP7_75t_L      g00391(.A(new_n628), .B(new_n646), .C(new_n626), .Y(new_n648));
  INVx1_ASAP7_75t_L         g00392(.A(new_n648), .Y(new_n649));
  NAND2xp33_ASAP7_75t_L     g00393(.A(new_n647), .B(new_n649), .Y(new_n650));
  O2A1O1Ixp33_ASAP7_75t_L   g00394(.A1(new_n577), .A2(new_n578), .B(new_n579), .C(new_n650), .Y(new_n651));
  A2O1A1Ixp33_ASAP7_75t_L   g00395(.A1(new_n570), .A2(new_n571), .B(new_n577), .C(new_n579), .Y(new_n652));
  AOI21xp33_ASAP7_75t_L     g00396(.A1(new_n649), .A2(new_n647), .B(new_n652), .Y(new_n653));
  NOR2xp33_ASAP7_75t_L      g00397(.A(new_n651), .B(new_n653), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g00398(.A(new_n577), .B(new_n578), .Y(new_n655));
  A2O1A1O1Ixp25_ASAP7_75t_L g00399(.A1(new_n575), .A2(new_n574), .B(new_n655), .C(new_n647), .D(new_n648), .Y(new_n656));
  NOR3xp33_ASAP7_75t_L      g00400(.A(new_n620), .B(new_n619), .C(new_n617), .Y(new_n657));
  AOI21xp33_ASAP7_75t_L     g00401(.A1(new_n625), .A2(new_n623), .B(new_n657), .Y(new_n658));
  NAND2xp33_ASAP7_75t_L     g00402(.A(\b[7] ), .B(new_n334), .Y(new_n659));
  OAI221xp5_ASAP7_75t_L     g00403(.A1(new_n368), .A2(new_n503), .B1(new_n382), .B2(new_n365), .C(new_n659), .Y(new_n660));
  AOI21xp33_ASAP7_75t_L     g00404(.A1(new_n510), .A2(new_n342), .B(new_n660), .Y(new_n661));
  NAND2xp33_ASAP7_75t_L     g00405(.A(\a[5] ), .B(new_n661), .Y(new_n662));
  A2O1A1Ixp33_ASAP7_75t_L   g00406(.A1(new_n510), .A2(new_n342), .B(new_n660), .C(new_n339), .Y(new_n663));
  AND2x2_ASAP7_75t_L        g00407(.A(new_n663), .B(new_n662), .Y(new_n664));
  INVx1_ASAP7_75t_L         g00408(.A(new_n580), .Y(new_n665));
  A2O1A1Ixp33_ASAP7_75t_L   g00409(.A1(new_n548), .A2(new_n665), .B(new_n608), .C(new_n605), .Y(new_n666));
  INVx1_ASAP7_75t_L         g00410(.A(new_n451), .Y(new_n667));
  NAND2xp33_ASAP7_75t_L     g00411(.A(\b[4] ), .B(new_n441), .Y(new_n668));
  OAI221xp5_ASAP7_75t_L     g00412(.A1(new_n667), .A2(new_n353), .B1(new_n482), .B2(new_n359), .C(new_n668), .Y(new_n669));
  AOI211xp5_ASAP7_75t_L     g00413(.A1(\b[3] ), .A2(new_n480), .B(new_n445), .C(new_n669), .Y(new_n670));
  INVx1_ASAP7_75t_L         g00414(.A(new_n670), .Y(new_n671));
  A2O1A1Ixp33_ASAP7_75t_L   g00415(.A1(\b[3] ), .A2(new_n480), .B(new_n669), .C(new_n445), .Y(new_n672));
  INVx1_ASAP7_75t_L         g00416(.A(new_n589), .Y(new_n673));
  NOR3xp33_ASAP7_75t_L      g00417(.A(new_n596), .B(new_n673), .C(new_n588), .Y(new_n674));
  NAND2xp33_ASAP7_75t_L     g00418(.A(new_n599), .B(new_n588), .Y(new_n675));
  INVx1_ASAP7_75t_L         g00419(.A(new_n600), .Y(new_n676));
  NAND2xp33_ASAP7_75t_L     g00420(.A(\b[1] ), .B(new_n590), .Y(new_n677));
  OAI221xp5_ASAP7_75t_L     g00421(.A1(new_n675), .A2(new_n283), .B1(new_n278), .B2(new_n676), .C(new_n677), .Y(new_n678));
  AOI21xp33_ASAP7_75t_L     g00422(.A1(new_n674), .A2(\b[0] ), .B(new_n678), .Y(new_n679));
  A2O1A1Ixp33_ASAP7_75t_L   g00423(.A1(new_n527), .A2(new_n602), .B(new_n594), .C(new_n679), .Y(new_n680));
  O2A1O1Ixp33_ASAP7_75t_L   g00424(.A1(new_n258), .A2(new_n522), .B(new_n602), .C(new_n594), .Y(new_n681));
  A2O1A1Ixp33_ASAP7_75t_L   g00425(.A1(\b[0] ), .A2(new_n674), .B(new_n678), .C(new_n681), .Y(new_n682));
  NAND4xp25_ASAP7_75t_L     g00426(.A(new_n682), .B(new_n671), .C(new_n672), .D(new_n680), .Y(new_n683));
  NAND2xp33_ASAP7_75t_L     g00427(.A(new_n672), .B(new_n671), .Y(new_n684));
  NAND2xp33_ASAP7_75t_L     g00428(.A(new_n680), .B(new_n682), .Y(new_n685));
  NAND2xp33_ASAP7_75t_L     g00429(.A(new_n685), .B(new_n684), .Y(new_n686));
  NAND2xp33_ASAP7_75t_L     g00430(.A(new_n683), .B(new_n686), .Y(new_n687));
  NAND2xp33_ASAP7_75t_L     g00431(.A(new_n666), .B(new_n687), .Y(new_n688));
  O2A1O1Ixp33_ASAP7_75t_L   g00432(.A1(new_n580), .A2(new_n535), .B(new_n604), .C(new_n609), .Y(new_n689));
  NAND3xp33_ASAP7_75t_L     g00433(.A(new_n689), .B(new_n683), .C(new_n686), .Y(new_n690));
  NAND2xp33_ASAP7_75t_L     g00434(.A(new_n690), .B(new_n688), .Y(new_n691));
  XNOR2x2_ASAP7_75t_L       g00435(.A(new_n664), .B(new_n691), .Y(new_n692));
  XNOR2x2_ASAP7_75t_L       g00436(.A(new_n658), .B(new_n692), .Y(new_n693));
  NOR2xp33_ASAP7_75t_L      g00437(.A(\b[10] ), .B(\b[11] ), .Y(new_n694));
  INVx1_ASAP7_75t_L         g00438(.A(\b[11] ), .Y(new_n695));
  NOR2xp33_ASAP7_75t_L      g00439(.A(new_n631), .B(new_n695), .Y(new_n696));
  NOR2xp33_ASAP7_75t_L      g00440(.A(new_n694), .B(new_n696), .Y(new_n697));
  A2O1A1Ixp33_ASAP7_75t_L   g00441(.A1(new_n638), .A2(new_n635), .B(new_n634), .C(new_n697), .Y(new_n698));
  A2O1A1O1Ixp25_ASAP7_75t_L g00442(.A1(new_n561), .A2(new_n564), .B(new_n560), .C(new_n635), .D(new_n634), .Y(new_n699));
  OAI21xp33_ASAP7_75t_L     g00443(.A1(new_n694), .A2(new_n696), .B(new_n699), .Y(new_n700));
  NAND2xp33_ASAP7_75t_L     g00444(.A(new_n698), .B(new_n700), .Y(new_n701));
  INVx1_ASAP7_75t_L         g00445(.A(new_n701), .Y(new_n702));
  AOI22xp33_ASAP7_75t_L     g00446(.A1(new_n272), .A2(\b[11] ), .B1(new_n269), .B2(new_n702), .Y(new_n703));
  OAI221xp5_ASAP7_75t_L     g00447(.A1(new_n261), .A2(new_n631), .B1(new_n559), .B2(new_n277), .C(new_n703), .Y(new_n704));
  XNOR2x2_ASAP7_75t_L       g00448(.A(\a[2] ), .B(new_n704), .Y(new_n705));
  NOR2xp33_ASAP7_75t_L      g00449(.A(new_n705), .B(new_n693), .Y(new_n706));
  AND2x2_ASAP7_75t_L        g00450(.A(new_n705), .B(new_n693), .Y(new_n707));
  NOR2xp33_ASAP7_75t_L      g00451(.A(new_n706), .B(new_n707), .Y(new_n708));
  XNOR2x2_ASAP7_75t_L       g00452(.A(new_n656), .B(new_n708), .Y(\f[11] ));
  INVx1_ASAP7_75t_L         g00453(.A(\a[12] ), .Y(new_n710));
  NAND2xp33_ASAP7_75t_L     g00454(.A(\a[11] ), .B(new_n710), .Y(new_n711));
  NAND2xp33_ASAP7_75t_L     g00455(.A(\a[12] ), .B(new_n594), .Y(new_n712));
  AND2x2_ASAP7_75t_L        g00456(.A(new_n711), .B(new_n712), .Y(new_n713));
  NOR2xp33_ASAP7_75t_L      g00457(.A(new_n258), .B(new_n713), .Y(new_n714));
  INVx1_ASAP7_75t_L         g00458(.A(new_n714), .Y(new_n715));
  NAND5xp2_ASAP7_75t_L      g00459(.A(new_n601), .B(new_n598), .C(new_n591), .D(new_n527), .E(\a[11] ), .Y(new_n716));
  AOI211xp5_ASAP7_75t_L     g00460(.A1(new_n674), .A2(\b[0] ), .B(new_n678), .C(new_n716), .Y(new_n717));
  NOR2xp33_ASAP7_75t_L      g00461(.A(new_n715), .B(new_n717), .Y(new_n718));
  AO21x2_ASAP7_75t_L        g00462(.A1(\b[0] ), .A2(new_n674), .B(new_n678), .Y(new_n719));
  NOR3xp33_ASAP7_75t_L      g00463(.A(new_n719), .B(new_n714), .C(new_n716), .Y(new_n720));
  NAND2xp33_ASAP7_75t_L     g00464(.A(new_n673), .B(new_n522), .Y(new_n721));
  NAND2xp33_ASAP7_75t_L     g00465(.A(\b[3] ), .B(new_n600), .Y(new_n722));
  OAI221xp5_ASAP7_75t_L     g00466(.A1(new_n278), .A2(new_n721), .B1(new_n675), .B2(new_n303), .C(new_n722), .Y(new_n723));
  AO211x2_ASAP7_75t_L       g00467(.A1(\b[1] ), .A2(new_n674), .B(new_n594), .C(new_n723), .Y(new_n724));
  A2O1A1Ixp33_ASAP7_75t_L   g00468(.A1(\b[1] ), .A2(new_n674), .B(new_n723), .C(new_n594), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g00469(.A(new_n725), .B(new_n724), .Y(new_n726));
  OAI21xp33_ASAP7_75t_L     g00470(.A1(new_n718), .A2(new_n720), .B(new_n726), .Y(new_n727));
  OAI21xp33_ASAP7_75t_L     g00471(.A1(new_n716), .A2(new_n719), .B(new_n714), .Y(new_n728));
  NAND2xp33_ASAP7_75t_L     g00472(.A(new_n715), .B(new_n717), .Y(new_n729));
  AND2x2_ASAP7_75t_L        g00473(.A(new_n725), .B(new_n724), .Y(new_n730));
  NAND3xp33_ASAP7_75t_L     g00474(.A(new_n730), .B(new_n729), .C(new_n728), .Y(new_n731));
  NAND2xp33_ASAP7_75t_L     g00475(.A(\b[4] ), .B(new_n480), .Y(new_n732));
  NAND2xp33_ASAP7_75t_L     g00476(.A(\b[5] ), .B(new_n441), .Y(new_n733));
  AOI22xp33_ASAP7_75t_L     g00477(.A1(new_n451), .A2(\b[6] ), .B1(new_n448), .B2(new_n389), .Y(new_n734));
  NAND4xp25_ASAP7_75t_L     g00478(.A(new_n734), .B(\a[8] ), .C(new_n732), .D(new_n733), .Y(new_n735));
  AOI31xp33_ASAP7_75t_L     g00479(.A1(new_n734), .A2(new_n733), .A3(new_n732), .B(\a[8] ), .Y(new_n736));
  INVx1_ASAP7_75t_L         g00480(.A(new_n736), .Y(new_n737));
  NAND4xp25_ASAP7_75t_L     g00481(.A(new_n731), .B(new_n737), .C(new_n727), .D(new_n735), .Y(new_n738));
  AOI21xp33_ASAP7_75t_L     g00482(.A1(new_n729), .A2(new_n728), .B(new_n730), .Y(new_n739));
  NOR3xp33_ASAP7_75t_L      g00483(.A(new_n720), .B(new_n718), .C(new_n726), .Y(new_n740));
  INVx1_ASAP7_75t_L         g00484(.A(new_n735), .Y(new_n741));
  OAI22xp33_ASAP7_75t_L     g00485(.A1(new_n739), .A2(new_n740), .B1(new_n736), .B2(new_n741), .Y(new_n742));
  NAND2xp33_ASAP7_75t_L     g00486(.A(new_n738), .B(new_n742), .Y(new_n743));
  AND2x2_ASAP7_75t_L        g00487(.A(new_n680), .B(new_n682), .Y(new_n744));
  NAND2xp33_ASAP7_75t_L     g00488(.A(new_n684), .B(new_n744), .Y(new_n745));
  A2O1A1Ixp33_ASAP7_75t_L   g00489(.A1(new_n683), .A2(new_n686), .B(new_n689), .C(new_n745), .Y(new_n746));
  XNOR2x2_ASAP7_75t_L       g00490(.A(new_n746), .B(new_n743), .Y(new_n747));
  OAI22xp33_ASAP7_75t_L     g00491(.A1(new_n365), .A2(new_n421), .B1(new_n559), .B2(new_n368), .Y(new_n748));
  AOI221xp5_ASAP7_75t_L     g00492(.A1(new_n334), .A2(\b[8] ), .B1(new_n342), .B2(new_n566), .C(new_n748), .Y(new_n749));
  XNOR2x2_ASAP7_75t_L       g00493(.A(new_n339), .B(new_n749), .Y(new_n750));
  NAND2xp33_ASAP7_75t_L     g00494(.A(new_n750), .B(new_n747), .Y(new_n751));
  NOR2xp33_ASAP7_75t_L      g00495(.A(new_n746), .B(new_n743), .Y(new_n752));
  MAJIxp5_ASAP7_75t_L       g00496(.A(new_n666), .B(new_n684), .C(new_n744), .Y(new_n753));
  AOI21xp33_ASAP7_75t_L     g00497(.A1(new_n742), .A2(new_n738), .B(new_n753), .Y(new_n754));
  NOR2xp33_ASAP7_75t_L      g00498(.A(new_n752), .B(new_n754), .Y(new_n755));
  INVx1_ASAP7_75t_L         g00499(.A(new_n750), .Y(new_n756));
  NAND2xp33_ASAP7_75t_L     g00500(.A(new_n756), .B(new_n755), .Y(new_n757));
  NAND2xp33_ASAP7_75t_L     g00501(.A(new_n751), .B(new_n757), .Y(new_n758));
  MAJx2_ASAP7_75t_L         g00502(.A(new_n658), .B(new_n664), .C(new_n691), .Y(new_n759));
  NOR2xp33_ASAP7_75t_L      g00503(.A(new_n758), .B(new_n759), .Y(new_n760));
  MAJIxp5_ASAP7_75t_L       g00504(.A(new_n658), .B(new_n664), .C(new_n691), .Y(new_n761));
  AOI21xp33_ASAP7_75t_L     g00505(.A1(new_n757), .A2(new_n751), .B(new_n761), .Y(new_n762));
  INVx1_ASAP7_75t_L         g00506(.A(\b[12] ), .Y(new_n763));
  A2O1A1Ixp33_ASAP7_75t_L   g00507(.A1(new_n538), .A2(new_n384), .B(new_n425), .C(new_n556), .Y(new_n764));
  A2O1A1Ixp33_ASAP7_75t_L   g00508(.A1(new_n764), .A2(new_n505), .B(new_n504), .C(new_n561), .Y(new_n765));
  INVx1_ASAP7_75t_L         g00509(.A(new_n634), .Y(new_n766));
  A2O1A1Ixp33_ASAP7_75t_L   g00510(.A1(new_n765), .A2(new_n637), .B(new_n633), .C(new_n766), .Y(new_n767));
  NOR2xp33_ASAP7_75t_L      g00511(.A(\b[11] ), .B(\b[12] ), .Y(new_n768));
  NOR2xp33_ASAP7_75t_L      g00512(.A(new_n695), .B(new_n763), .Y(new_n769));
  NOR2xp33_ASAP7_75t_L      g00513(.A(new_n768), .B(new_n769), .Y(new_n770));
  A2O1A1Ixp33_ASAP7_75t_L   g00514(.A1(new_n767), .A2(new_n697), .B(new_n696), .C(new_n770), .Y(new_n771));
  A2O1A1O1Ixp25_ASAP7_75t_L g00515(.A1(new_n635), .A2(new_n638), .B(new_n634), .C(new_n697), .D(new_n696), .Y(new_n772));
  INVx1_ASAP7_75t_L         g00516(.A(new_n770), .Y(new_n773));
  NAND2xp33_ASAP7_75t_L     g00517(.A(new_n773), .B(new_n772), .Y(new_n774));
  NAND2xp33_ASAP7_75t_L     g00518(.A(new_n774), .B(new_n771), .Y(new_n775));
  OAI22xp33_ASAP7_75t_L     g00519(.A1(new_n775), .A2(new_n292), .B1(new_n763), .B2(new_n632), .Y(new_n776));
  AOI221xp5_ASAP7_75t_L     g00520(.A1(\b[10] ), .A2(new_n291), .B1(\b[11] ), .B2(new_n380), .C(new_n776), .Y(new_n777));
  XNOR2x2_ASAP7_75t_L       g00521(.A(\a[2] ), .B(new_n777), .Y(new_n778));
  NOR3xp33_ASAP7_75t_L      g00522(.A(new_n760), .B(new_n762), .C(new_n778), .Y(new_n779));
  OA21x2_ASAP7_75t_L        g00523(.A1(new_n762), .A2(new_n760), .B(new_n778), .Y(new_n780));
  MAJIxp5_ASAP7_75t_L       g00524(.A(new_n656), .B(new_n705), .C(new_n693), .Y(new_n781));
  OAI21xp33_ASAP7_75t_L     g00525(.A1(new_n779), .A2(new_n780), .B(new_n781), .Y(new_n782));
  INVx1_ASAP7_75t_L         g00526(.A(new_n782), .Y(new_n783));
  NOR3xp33_ASAP7_75t_L      g00527(.A(new_n781), .B(new_n780), .C(new_n779), .Y(new_n784));
  NOR2xp33_ASAP7_75t_L      g00528(.A(new_n784), .B(new_n783), .Y(\f[12] ));
  NOR2xp33_ASAP7_75t_L      g00529(.A(new_n762), .B(new_n760), .Y(new_n786));
  NAND2xp33_ASAP7_75t_L     g00530(.A(new_n778), .B(new_n786), .Y(new_n787));
  INVx1_ASAP7_75t_L         g00531(.A(new_n787), .Y(new_n788));
  O2A1O1Ixp33_ASAP7_75t_L   g00532(.A1(new_n779), .A2(new_n780), .B(new_n781), .C(new_n788), .Y(new_n789));
  INVx1_ASAP7_75t_L         g00533(.A(new_n696), .Y(new_n790));
  INVx1_ASAP7_75t_L         g00534(.A(new_n769), .Y(new_n791));
  NOR2xp33_ASAP7_75t_L      g00535(.A(\b[12] ), .B(\b[13] ), .Y(new_n792));
  INVx1_ASAP7_75t_L         g00536(.A(\b[13] ), .Y(new_n793));
  NOR2xp33_ASAP7_75t_L      g00537(.A(new_n763), .B(new_n793), .Y(new_n794));
  NOR2xp33_ASAP7_75t_L      g00538(.A(new_n792), .B(new_n794), .Y(new_n795));
  INVx1_ASAP7_75t_L         g00539(.A(new_n795), .Y(new_n796));
  A2O1A1O1Ixp25_ASAP7_75t_L g00540(.A1(new_n790), .A2(new_n698), .B(new_n768), .C(new_n791), .D(new_n796), .Y(new_n797));
  A2O1A1Ixp33_ASAP7_75t_L   g00541(.A1(new_n698), .A2(new_n790), .B(new_n768), .C(new_n791), .Y(new_n798));
  NOR2xp33_ASAP7_75t_L      g00542(.A(new_n795), .B(new_n798), .Y(new_n799));
  NOR2xp33_ASAP7_75t_L      g00543(.A(new_n797), .B(new_n799), .Y(new_n800));
  AOI22xp33_ASAP7_75t_L     g00544(.A1(new_n272), .A2(\b[13] ), .B1(new_n269), .B2(new_n800), .Y(new_n801));
  OAI221xp5_ASAP7_75t_L     g00545(.A1(new_n261), .A2(new_n763), .B1(new_n695), .B2(new_n277), .C(new_n801), .Y(new_n802));
  XNOR2x2_ASAP7_75t_L       g00546(.A(new_n265), .B(new_n802), .Y(new_n803));
  OAI21xp33_ASAP7_75t_L     g00547(.A1(new_n758), .A2(new_n759), .B(new_n757), .Y(new_n804));
  NAND2xp33_ASAP7_75t_L     g00548(.A(new_n714), .B(new_n717), .Y(new_n805));
  A2O1A1Ixp33_ASAP7_75t_L   g00549(.A1(new_n729), .A2(new_n728), .B(new_n730), .C(new_n805), .Y(new_n806));
  NAND2xp33_ASAP7_75t_L     g00550(.A(\b[2] ), .B(new_n674), .Y(new_n807));
  NAND2xp33_ASAP7_75t_L     g00551(.A(\b[3] ), .B(new_n590), .Y(new_n808));
  AOI22xp33_ASAP7_75t_L     g00552(.A1(new_n600), .A2(\b[4] ), .B1(new_n597), .B2(new_n328), .Y(new_n809));
  NAND4xp25_ASAP7_75t_L     g00553(.A(new_n809), .B(\a[11] ), .C(new_n807), .D(new_n808), .Y(new_n810));
  NAND2xp33_ASAP7_75t_L     g00554(.A(new_n808), .B(new_n809), .Y(new_n811));
  A2O1A1Ixp33_ASAP7_75t_L   g00555(.A1(\b[2] ), .A2(new_n674), .B(new_n811), .C(new_n594), .Y(new_n812));
  INVx1_ASAP7_75t_L         g00556(.A(\a[14] ), .Y(new_n813));
  NOR2xp33_ASAP7_75t_L      g00557(.A(new_n813), .B(new_n715), .Y(new_n814));
  NAND2xp33_ASAP7_75t_L     g00558(.A(new_n712), .B(new_n711), .Y(new_n815));
  XNOR2x2_ASAP7_75t_L       g00559(.A(\a[13] ), .B(\a[12] ), .Y(new_n816));
  NOR2xp33_ASAP7_75t_L      g00560(.A(new_n816), .B(new_n815), .Y(new_n817));
  NAND2xp33_ASAP7_75t_L     g00561(.A(\b[0] ), .B(new_n817), .Y(new_n818));
  INVx1_ASAP7_75t_L         g00562(.A(\a[13] ), .Y(new_n819));
  NAND2xp33_ASAP7_75t_L     g00563(.A(\a[14] ), .B(new_n819), .Y(new_n820));
  NAND2xp33_ASAP7_75t_L     g00564(.A(\a[13] ), .B(new_n813), .Y(new_n821));
  AND2x2_ASAP7_75t_L        g00565(.A(new_n820), .B(new_n821), .Y(new_n822));
  NOR2xp33_ASAP7_75t_L      g00566(.A(new_n713), .B(new_n822), .Y(new_n823));
  NAND2xp33_ASAP7_75t_L     g00567(.A(new_n271), .B(new_n823), .Y(new_n824));
  NAND2xp33_ASAP7_75t_L     g00568(.A(new_n821), .B(new_n820), .Y(new_n825));
  NOR2xp33_ASAP7_75t_L      g00569(.A(new_n825), .B(new_n713), .Y(new_n826));
  NAND2xp33_ASAP7_75t_L     g00570(.A(\b[1] ), .B(new_n826), .Y(new_n827));
  NAND3xp33_ASAP7_75t_L     g00571(.A(new_n824), .B(new_n827), .C(new_n818), .Y(new_n828));
  XNOR2x2_ASAP7_75t_L       g00572(.A(new_n814), .B(new_n828), .Y(new_n829));
  NAND3xp33_ASAP7_75t_L     g00573(.A(new_n812), .B(new_n810), .C(new_n829), .Y(new_n830));
  AO21x2_ASAP7_75t_L        g00574(.A1(new_n810), .A2(new_n812), .B(new_n829), .Y(new_n831));
  NAND3xp33_ASAP7_75t_L     g00575(.A(new_n806), .B(new_n830), .C(new_n831), .Y(new_n832));
  MAJIxp5_ASAP7_75t_L       g00576(.A(new_n726), .B(new_n714), .C(new_n717), .Y(new_n833));
  AND3x1_ASAP7_75t_L        g00577(.A(new_n812), .B(new_n829), .C(new_n810), .Y(new_n834));
  AOI21xp33_ASAP7_75t_L     g00578(.A1(new_n812), .A2(new_n810), .B(new_n829), .Y(new_n835));
  OAI21xp33_ASAP7_75t_L     g00579(.A1(new_n835), .A2(new_n834), .B(new_n833), .Y(new_n836));
  OAI22xp33_ASAP7_75t_L     g00580(.A1(new_n427), .A2(new_n482), .B1(new_n667), .B2(new_n421), .Y(new_n837));
  AOI221xp5_ASAP7_75t_L     g00581(.A1(\b[5] ), .A2(new_n480), .B1(\b[6] ), .B2(new_n441), .C(new_n837), .Y(new_n838));
  NAND2xp33_ASAP7_75t_L     g00582(.A(\a[8] ), .B(new_n838), .Y(new_n839));
  AO21x2_ASAP7_75t_L        g00583(.A1(\b[6] ), .A2(new_n441), .B(new_n837), .Y(new_n840));
  A2O1A1Ixp33_ASAP7_75t_L   g00584(.A1(\b[5] ), .A2(new_n480), .B(new_n840), .C(new_n445), .Y(new_n841));
  NAND4xp25_ASAP7_75t_L     g00585(.A(new_n832), .B(new_n841), .C(new_n839), .D(new_n836), .Y(new_n842));
  AO22x1_ASAP7_75t_L        g00586(.A1(new_n839), .A2(new_n841), .B1(new_n836), .B2(new_n832), .Y(new_n843));
  NOR2xp33_ASAP7_75t_L      g00587(.A(new_n740), .B(new_n739), .Y(new_n844));
  NAND2xp33_ASAP7_75t_L     g00588(.A(new_n735), .B(new_n737), .Y(new_n845));
  MAJIxp5_ASAP7_75t_L       g00589(.A(new_n746), .B(new_n844), .C(new_n845), .Y(new_n846));
  AND3x1_ASAP7_75t_L        g00590(.A(new_n846), .B(new_n843), .C(new_n842), .Y(new_n847));
  AOI21xp33_ASAP7_75t_L     g00591(.A1(new_n843), .A2(new_n842), .B(new_n846), .Y(new_n848));
  O2A1O1Ixp33_ASAP7_75t_L   g00592(.A1(new_n422), .A2(new_n501), .B(new_n505), .C(new_n504), .Y(new_n849));
  INVx1_ASAP7_75t_L         g00593(.A(new_n635), .Y(new_n850));
  O2A1O1Ixp33_ASAP7_75t_L   g00594(.A1(new_n562), .A2(new_n849), .B(new_n637), .C(new_n850), .Y(new_n851));
  NOR2xp33_ASAP7_75t_L      g00595(.A(new_n851), .B(new_n639), .Y(new_n852));
  NOR2xp33_ASAP7_75t_L      g00596(.A(new_n631), .B(new_n368), .Y(new_n853));
  AOI221xp5_ASAP7_75t_L     g00597(.A1(new_n334), .A2(\b[9] ), .B1(new_n342), .B2(new_n852), .C(new_n853), .Y(new_n854));
  OA211x2_ASAP7_75t_L       g00598(.A1(new_n365), .A2(new_n503), .B(new_n854), .C(\a[5] ), .Y(new_n855));
  O2A1O1Ixp33_ASAP7_75t_L   g00599(.A1(new_n503), .A2(new_n365), .B(new_n854), .C(\a[5] ), .Y(new_n856));
  NOR2xp33_ASAP7_75t_L      g00600(.A(new_n856), .B(new_n855), .Y(new_n857));
  OAI21xp33_ASAP7_75t_L     g00601(.A1(new_n848), .A2(new_n847), .B(new_n857), .Y(new_n858));
  NOR3xp33_ASAP7_75t_L      g00602(.A(new_n857), .B(new_n847), .C(new_n848), .Y(new_n859));
  INVx1_ASAP7_75t_L         g00603(.A(new_n859), .Y(new_n860));
  NAND2xp33_ASAP7_75t_L     g00604(.A(new_n858), .B(new_n860), .Y(new_n861));
  NOR2xp33_ASAP7_75t_L      g00605(.A(new_n861), .B(new_n804), .Y(new_n862));
  AND2x2_ASAP7_75t_L        g00606(.A(new_n861), .B(new_n804), .Y(new_n863));
  OAI21xp33_ASAP7_75t_L     g00607(.A1(new_n862), .A2(new_n863), .B(new_n803), .Y(new_n864));
  INVx1_ASAP7_75t_L         g00608(.A(new_n864), .Y(new_n865));
  NOR3xp33_ASAP7_75t_L      g00609(.A(new_n863), .B(new_n862), .C(new_n803), .Y(new_n866));
  NOR2xp33_ASAP7_75t_L      g00610(.A(new_n866), .B(new_n865), .Y(new_n867));
  XNOR2x2_ASAP7_75t_L       g00611(.A(new_n789), .B(new_n867), .Y(\f[13] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00612(.A1(new_n782), .A2(new_n787), .B(new_n866), .C(new_n864), .Y(new_n869));
  NOR2xp33_ASAP7_75t_L      g00613(.A(\b[13] ), .B(\b[14] ), .Y(new_n870));
  INVx1_ASAP7_75t_L         g00614(.A(\b[14] ), .Y(new_n871));
  NOR2xp33_ASAP7_75t_L      g00615(.A(new_n793), .B(new_n871), .Y(new_n872));
  NOR2xp33_ASAP7_75t_L      g00616(.A(new_n870), .B(new_n872), .Y(new_n873));
  A2O1A1Ixp33_ASAP7_75t_L   g00617(.A1(new_n798), .A2(new_n795), .B(new_n794), .C(new_n873), .Y(new_n874));
  A2O1A1Ixp33_ASAP7_75t_L   g00618(.A1(new_n636), .A2(new_n766), .B(new_n694), .C(new_n790), .Y(new_n875));
  A2O1A1O1Ixp25_ASAP7_75t_L g00619(.A1(new_n770), .A2(new_n875), .B(new_n769), .C(new_n795), .D(new_n794), .Y(new_n876));
  OAI21xp33_ASAP7_75t_L     g00620(.A1(new_n870), .A2(new_n872), .B(new_n876), .Y(new_n877));
  NAND2xp33_ASAP7_75t_L     g00621(.A(new_n874), .B(new_n877), .Y(new_n878));
  INVx1_ASAP7_75t_L         g00622(.A(new_n878), .Y(new_n879));
  AOI22xp33_ASAP7_75t_L     g00623(.A1(new_n272), .A2(\b[14] ), .B1(new_n269), .B2(new_n879), .Y(new_n880));
  OAI221xp5_ASAP7_75t_L     g00624(.A1(new_n261), .A2(new_n793), .B1(new_n763), .B2(new_n277), .C(new_n880), .Y(new_n881));
  XNOR2x2_ASAP7_75t_L       g00625(.A(new_n265), .B(new_n881), .Y(new_n882));
  NAND2xp33_ASAP7_75t_L     g00626(.A(\b[9] ), .B(new_n366), .Y(new_n883));
  NAND2xp33_ASAP7_75t_L     g00627(.A(\b[10] ), .B(new_n334), .Y(new_n884));
  AOI22xp33_ASAP7_75t_L     g00628(.A1(new_n345), .A2(\b[11] ), .B1(new_n342), .B2(new_n702), .Y(new_n885));
  NAND4xp25_ASAP7_75t_L     g00629(.A(new_n885), .B(\a[5] ), .C(new_n883), .D(new_n884), .Y(new_n886));
  NAND2xp33_ASAP7_75t_L     g00630(.A(new_n884), .B(new_n885), .Y(new_n887));
  A2O1A1Ixp33_ASAP7_75t_L   g00631(.A1(\b[9] ), .A2(new_n366), .B(new_n887), .C(new_n339), .Y(new_n888));
  AND2x2_ASAP7_75t_L        g00632(.A(new_n886), .B(new_n888), .Y(new_n889));
  NAND2xp33_ASAP7_75t_L     g00633(.A(new_n839), .B(new_n841), .Y(new_n890));
  NAND3xp33_ASAP7_75t_L     g00634(.A(new_n890), .B(new_n836), .C(new_n832), .Y(new_n891));
  A2O1A1Ixp33_ASAP7_75t_L   g00635(.A1(new_n843), .A2(new_n842), .B(new_n846), .C(new_n891), .Y(new_n892));
  NAND2xp33_ASAP7_75t_L     g00636(.A(\b[7] ), .B(new_n441), .Y(new_n893));
  OAI221xp5_ASAP7_75t_L     g00637(.A1(new_n667), .A2(new_n503), .B1(new_n482), .B2(new_n509), .C(new_n893), .Y(new_n894));
  AOI21xp33_ASAP7_75t_L     g00638(.A1(new_n480), .A2(\b[6] ), .B(new_n894), .Y(new_n895));
  NAND2xp33_ASAP7_75t_L     g00639(.A(\a[8] ), .B(new_n895), .Y(new_n896));
  A2O1A1Ixp33_ASAP7_75t_L   g00640(.A1(\b[6] ), .A2(new_n480), .B(new_n894), .C(new_n445), .Y(new_n897));
  NAND2xp33_ASAP7_75t_L     g00641(.A(new_n729), .B(new_n728), .Y(new_n898));
  INVx1_ASAP7_75t_L         g00642(.A(new_n805), .Y(new_n899));
  A2O1A1O1Ixp25_ASAP7_75t_L g00643(.A1(new_n726), .A2(new_n898), .B(new_n899), .C(new_n830), .D(new_n835), .Y(new_n900));
  NAND2xp33_ASAP7_75t_L     g00644(.A(\b[4] ), .B(new_n590), .Y(new_n901));
  OAI221xp5_ASAP7_75t_L     g00645(.A1(new_n676), .A2(new_n353), .B1(new_n675), .B2(new_n359), .C(new_n901), .Y(new_n902));
  AOI211xp5_ASAP7_75t_L     g00646(.A1(\b[3] ), .A2(new_n674), .B(new_n594), .C(new_n902), .Y(new_n903));
  INVx1_ASAP7_75t_L         g00647(.A(new_n903), .Y(new_n904));
  A2O1A1Ixp33_ASAP7_75t_L   g00648(.A1(\b[3] ), .A2(new_n674), .B(new_n902), .C(new_n594), .Y(new_n905));
  AND3x1_ASAP7_75t_L        g00649(.A(new_n824), .B(new_n827), .C(new_n818), .Y(new_n906));
  INVx1_ASAP7_75t_L         g00650(.A(new_n816), .Y(new_n907));
  NOR3xp33_ASAP7_75t_L      g00651(.A(new_n822), .B(new_n907), .C(new_n815), .Y(new_n908));
  INVx1_ASAP7_75t_L         g00652(.A(new_n908), .Y(new_n909));
  NOR2xp33_ASAP7_75t_L      g00653(.A(new_n258), .B(new_n909), .Y(new_n910));
  NAND2xp33_ASAP7_75t_L     g00654(.A(new_n825), .B(new_n815), .Y(new_n911));
  NAND2xp33_ASAP7_75t_L     g00655(.A(new_n815), .B(new_n822), .Y(new_n912));
  NAND2xp33_ASAP7_75t_L     g00656(.A(\b[1] ), .B(new_n817), .Y(new_n913));
  OAI221xp5_ASAP7_75t_L     g00657(.A1(new_n911), .A2(new_n283), .B1(new_n278), .B2(new_n912), .C(new_n913), .Y(new_n914));
  NOR2xp33_ASAP7_75t_L      g00658(.A(new_n914), .B(new_n910), .Y(new_n915));
  A2O1A1Ixp33_ASAP7_75t_L   g00659(.A1(new_n715), .A2(new_n906), .B(new_n813), .C(new_n915), .Y(new_n916));
  INVx1_ASAP7_75t_L         g00660(.A(new_n916), .Y(new_n917));
  A2O1A1Ixp33_ASAP7_75t_L   g00661(.A1(\b[0] ), .A2(new_n815), .B(new_n828), .C(\a[14] ), .Y(new_n918));
  NOR2xp33_ASAP7_75t_L      g00662(.A(new_n911), .B(new_n283), .Y(new_n919));
  AOI221xp5_ASAP7_75t_L     g00663(.A1(\b[2] ), .A2(new_n826), .B1(new_n817), .B2(\b[1] ), .C(new_n919), .Y(new_n920));
  O2A1O1Ixp33_ASAP7_75t_L   g00664(.A1(new_n909), .A2(new_n258), .B(new_n920), .C(new_n918), .Y(new_n921));
  OAI211xp5_ASAP7_75t_L     g00665(.A1(new_n921), .A2(new_n917), .B(new_n905), .C(new_n904), .Y(new_n922));
  INVx1_ASAP7_75t_L         g00666(.A(new_n905), .Y(new_n923));
  O2A1O1Ixp33_ASAP7_75t_L   g00667(.A1(new_n258), .A2(new_n713), .B(new_n906), .C(new_n813), .Y(new_n924));
  A2O1A1Ixp33_ASAP7_75t_L   g00668(.A1(\b[0] ), .A2(new_n908), .B(new_n914), .C(new_n924), .Y(new_n925));
  OAI211xp5_ASAP7_75t_L     g00669(.A1(new_n903), .A2(new_n923), .B(new_n916), .C(new_n925), .Y(new_n926));
  NAND3xp33_ASAP7_75t_L     g00670(.A(new_n900), .B(new_n922), .C(new_n926), .Y(new_n927));
  NAND2xp33_ASAP7_75t_L     g00671(.A(new_n926), .B(new_n922), .Y(new_n928));
  A2O1A1Ixp33_ASAP7_75t_L   g00672(.A1(new_n830), .A2(new_n806), .B(new_n835), .C(new_n928), .Y(new_n929));
  AND4x1_ASAP7_75t_L        g00673(.A(new_n929), .B(new_n927), .C(new_n897), .D(new_n896), .Y(new_n930));
  AOI22xp33_ASAP7_75t_L     g00674(.A1(new_n897), .A2(new_n896), .B1(new_n929), .B2(new_n927), .Y(new_n931));
  NOR2xp33_ASAP7_75t_L      g00675(.A(new_n931), .B(new_n930), .Y(new_n932));
  NAND2xp33_ASAP7_75t_L     g00676(.A(new_n892), .B(new_n932), .Y(new_n933));
  NAND2xp33_ASAP7_75t_L     g00677(.A(new_n842), .B(new_n843), .Y(new_n934));
  A2O1A1Ixp33_ASAP7_75t_L   g00678(.A1(new_n845), .A2(new_n844), .B(new_n754), .C(new_n934), .Y(new_n935));
  OAI211xp5_ASAP7_75t_L     g00679(.A1(new_n930), .A2(new_n931), .B(new_n935), .C(new_n891), .Y(new_n936));
  NAND2xp33_ASAP7_75t_L     g00680(.A(new_n933), .B(new_n936), .Y(new_n937));
  NAND2xp33_ASAP7_75t_L     g00681(.A(new_n889), .B(new_n937), .Y(new_n938));
  NAND2xp33_ASAP7_75t_L     g00682(.A(new_n886), .B(new_n888), .Y(new_n939));
  NAND3xp33_ASAP7_75t_L     g00683(.A(new_n939), .B(new_n933), .C(new_n936), .Y(new_n940));
  NAND2xp33_ASAP7_75t_L     g00684(.A(new_n940), .B(new_n938), .Y(new_n941));
  INVx1_ASAP7_75t_L         g00685(.A(new_n757), .Y(new_n942));
  A2O1A1O1Ixp25_ASAP7_75t_L g00686(.A1(new_n751), .A2(new_n761), .B(new_n942), .C(new_n858), .D(new_n859), .Y(new_n943));
  XOR2x2_ASAP7_75t_L        g00687(.A(new_n943), .B(new_n941), .Y(new_n944));
  XNOR2x2_ASAP7_75t_L       g00688(.A(new_n882), .B(new_n944), .Y(new_n945));
  XNOR2x2_ASAP7_75t_L       g00689(.A(new_n869), .B(new_n945), .Y(\f[14] ));
  MAJIxp5_ASAP7_75t_L       g00690(.A(new_n869), .B(new_n882), .C(new_n944), .Y(new_n947));
  INVx1_ASAP7_75t_L         g00691(.A(new_n794), .Y(new_n948));
  A2O1A1Ixp33_ASAP7_75t_L   g00692(.A1(new_n875), .A2(new_n770), .B(new_n769), .C(new_n795), .Y(new_n949));
  INVx1_ASAP7_75t_L         g00693(.A(new_n872), .Y(new_n950));
  NOR2xp33_ASAP7_75t_L      g00694(.A(\b[14] ), .B(\b[15] ), .Y(new_n951));
  INVx1_ASAP7_75t_L         g00695(.A(\b[15] ), .Y(new_n952));
  NOR2xp33_ASAP7_75t_L      g00696(.A(new_n871), .B(new_n952), .Y(new_n953));
  NOR2xp33_ASAP7_75t_L      g00697(.A(new_n951), .B(new_n953), .Y(new_n954));
  INVx1_ASAP7_75t_L         g00698(.A(new_n954), .Y(new_n955));
  A2O1A1O1Ixp25_ASAP7_75t_L g00699(.A1(new_n948), .A2(new_n949), .B(new_n870), .C(new_n950), .D(new_n955), .Y(new_n956));
  A2O1A1Ixp33_ASAP7_75t_L   g00700(.A1(new_n949), .A2(new_n948), .B(new_n870), .C(new_n950), .Y(new_n957));
  NOR2xp33_ASAP7_75t_L      g00701(.A(new_n954), .B(new_n957), .Y(new_n958));
  NOR2xp33_ASAP7_75t_L      g00702(.A(new_n956), .B(new_n958), .Y(new_n959));
  AOI22xp33_ASAP7_75t_L     g00703(.A1(new_n272), .A2(\b[15] ), .B1(new_n269), .B2(new_n959), .Y(new_n960));
  OAI221xp5_ASAP7_75t_L     g00704(.A1(new_n261), .A2(new_n871), .B1(new_n793), .B2(new_n277), .C(new_n960), .Y(new_n961));
  XNOR2x2_ASAP7_75t_L       g00705(.A(\a[2] ), .B(new_n961), .Y(new_n962));
  INVx1_ASAP7_75t_L         g00706(.A(new_n962), .Y(new_n963));
  NOR2xp33_ASAP7_75t_L      g00707(.A(new_n889), .B(new_n937), .Y(new_n964));
  A2O1A1O1Ixp25_ASAP7_75t_L g00708(.A1(new_n858), .A2(new_n804), .B(new_n859), .C(new_n938), .D(new_n964), .Y(new_n965));
  NAND2xp33_ASAP7_75t_L     g00709(.A(\b[10] ), .B(new_n366), .Y(new_n966));
  NAND2xp33_ASAP7_75t_L     g00710(.A(\b[11] ), .B(new_n334), .Y(new_n967));
  A2O1A1O1Ixp25_ASAP7_75t_L g00711(.A1(new_n766), .A2(new_n636), .B(new_n694), .C(new_n790), .D(new_n773), .Y(new_n968));
  NOR2xp33_ASAP7_75t_L      g00712(.A(new_n770), .B(new_n875), .Y(new_n969));
  NOR2xp33_ASAP7_75t_L      g00713(.A(new_n968), .B(new_n969), .Y(new_n970));
  AOI22xp33_ASAP7_75t_L     g00714(.A1(new_n345), .A2(\b[12] ), .B1(new_n342), .B2(new_n970), .Y(new_n971));
  NAND4xp25_ASAP7_75t_L     g00715(.A(new_n971), .B(\a[5] ), .C(new_n966), .D(new_n967), .Y(new_n972));
  NAND3xp33_ASAP7_75t_L     g00716(.A(new_n971), .B(new_n967), .C(new_n966), .Y(new_n973));
  NAND2xp33_ASAP7_75t_L     g00717(.A(new_n339), .B(new_n973), .Y(new_n974));
  NAND2xp33_ASAP7_75t_L     g00718(.A(new_n972), .B(new_n974), .Y(new_n975));
  NOR2xp33_ASAP7_75t_L      g00719(.A(new_n421), .B(new_n481), .Y(new_n976));
  NAND2xp33_ASAP7_75t_L     g00720(.A(new_n562), .B(new_n849), .Y(new_n977));
  NAND2xp33_ASAP7_75t_L     g00721(.A(new_n977), .B(new_n765), .Y(new_n978));
  NAND2xp33_ASAP7_75t_L     g00722(.A(\b[8] ), .B(new_n441), .Y(new_n979));
  OAI221xp5_ASAP7_75t_L     g00723(.A1(new_n667), .A2(new_n559), .B1(new_n482), .B2(new_n978), .C(new_n979), .Y(new_n980));
  NOR3xp33_ASAP7_75t_L      g00724(.A(new_n980), .B(new_n976), .C(new_n445), .Y(new_n981));
  INVx1_ASAP7_75t_L         g00725(.A(new_n976), .Y(new_n982));
  AOI22xp33_ASAP7_75t_L     g00726(.A1(new_n451), .A2(\b[9] ), .B1(new_n448), .B2(new_n566), .Y(new_n983));
  AOI31xp33_ASAP7_75t_L     g00727(.A1(new_n983), .A2(new_n979), .A3(new_n982), .B(\a[8] ), .Y(new_n984));
  NAND5xp2_ASAP7_75t_L      g00728(.A(new_n827), .B(new_n824), .C(new_n818), .D(new_n715), .E(\a[14] ), .Y(new_n985));
  INVx1_ASAP7_75t_L         g00729(.A(\a[15] ), .Y(new_n986));
  NAND2xp33_ASAP7_75t_L     g00730(.A(\a[14] ), .B(new_n986), .Y(new_n987));
  NAND2xp33_ASAP7_75t_L     g00731(.A(\a[15] ), .B(new_n813), .Y(new_n988));
  AND2x2_ASAP7_75t_L        g00732(.A(new_n987), .B(new_n988), .Y(new_n989));
  NOR2xp33_ASAP7_75t_L      g00733(.A(new_n258), .B(new_n989), .Y(new_n990));
  OAI31xp33_ASAP7_75t_L     g00734(.A1(new_n985), .A2(new_n914), .A3(new_n910), .B(new_n990), .Y(new_n991));
  INVx1_ASAP7_75t_L         g00735(.A(new_n990), .Y(new_n992));
  NAND5xp2_ASAP7_75t_L      g00736(.A(\a[14] ), .B(new_n915), .C(new_n992), .D(new_n906), .E(new_n715), .Y(new_n993));
  NAND2xp33_ASAP7_75t_L     g00737(.A(new_n907), .B(new_n713), .Y(new_n994));
  NAND2xp33_ASAP7_75t_L     g00738(.A(\b[3] ), .B(new_n826), .Y(new_n995));
  OAI221xp5_ASAP7_75t_L     g00739(.A1(new_n278), .A2(new_n994), .B1(new_n911), .B2(new_n303), .C(new_n995), .Y(new_n996));
  AOI211xp5_ASAP7_75t_L     g00740(.A1(\b[1] ), .A2(new_n908), .B(new_n813), .C(new_n996), .Y(new_n997));
  O2A1O1Ixp33_ASAP7_75t_L   g00741(.A1(new_n276), .A2(new_n278), .B(new_n279), .C(new_n301), .Y(new_n998));
  O2A1O1Ixp33_ASAP7_75t_L   g00742(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n297), .Y(new_n999));
  NOR2xp33_ASAP7_75t_L      g00743(.A(new_n998), .B(new_n999), .Y(new_n1000));
  NOR2xp33_ASAP7_75t_L      g00744(.A(new_n278), .B(new_n994), .Y(new_n1001));
  AOI221xp5_ASAP7_75t_L     g00745(.A1(new_n826), .A2(\b[3] ), .B1(new_n823), .B2(new_n1000), .C(new_n1001), .Y(new_n1002));
  O2A1O1Ixp33_ASAP7_75t_L   g00746(.A1(new_n276), .A2(new_n909), .B(new_n1002), .C(\a[14] ), .Y(new_n1003));
  NOR2xp33_ASAP7_75t_L      g00747(.A(new_n997), .B(new_n1003), .Y(new_n1004));
  AO21x2_ASAP7_75t_L        g00748(.A1(new_n991), .A2(new_n993), .B(new_n1004), .Y(new_n1005));
  NAND3xp33_ASAP7_75t_L     g00749(.A(new_n1004), .B(new_n993), .C(new_n991), .Y(new_n1006));
  NAND2xp33_ASAP7_75t_L     g00750(.A(\b[4] ), .B(new_n674), .Y(new_n1007));
  NAND2xp33_ASAP7_75t_L     g00751(.A(\b[5] ), .B(new_n590), .Y(new_n1008));
  AOI22xp33_ASAP7_75t_L     g00752(.A1(new_n600), .A2(\b[6] ), .B1(new_n597), .B2(new_n389), .Y(new_n1009));
  NAND4xp25_ASAP7_75t_L     g00753(.A(new_n1009), .B(\a[11] ), .C(new_n1007), .D(new_n1008), .Y(new_n1010));
  OAI221xp5_ASAP7_75t_L     g00754(.A1(new_n676), .A2(new_n382), .B1(new_n675), .B2(new_n540), .C(new_n1008), .Y(new_n1011));
  A2O1A1Ixp33_ASAP7_75t_L   g00755(.A1(\b[4] ), .A2(new_n674), .B(new_n1011), .C(new_n594), .Y(new_n1012));
  NAND4xp25_ASAP7_75t_L     g00756(.A(new_n1005), .B(new_n1006), .C(new_n1012), .D(new_n1010), .Y(new_n1013));
  AO22x1_ASAP7_75t_L        g00757(.A1(new_n1012), .A2(new_n1010), .B1(new_n1006), .B2(new_n1005), .Y(new_n1014));
  AOI211xp5_ASAP7_75t_L     g00758(.A1(new_n904), .A2(new_n905), .B(new_n917), .C(new_n921), .Y(new_n1015));
  A2O1A1O1Ixp25_ASAP7_75t_L g00759(.A1(new_n830), .A2(new_n806), .B(new_n835), .C(new_n922), .D(new_n1015), .Y(new_n1016));
  AOI21xp33_ASAP7_75t_L     g00760(.A1(new_n1014), .A2(new_n1013), .B(new_n1016), .Y(new_n1017));
  AND4x1_ASAP7_75t_L        g00761(.A(new_n1005), .B(new_n1012), .C(new_n1006), .D(new_n1010), .Y(new_n1018));
  AOI22xp33_ASAP7_75t_L     g00762(.A1(new_n1010), .A2(new_n1012), .B1(new_n1006), .B2(new_n1005), .Y(new_n1019));
  AOI211xp5_ASAP7_75t_L     g00763(.A1(new_n925), .A2(new_n916), .B(new_n903), .C(new_n923), .Y(new_n1020));
  O2A1O1Ixp33_ASAP7_75t_L   g00764(.A1(new_n833), .A2(new_n834), .B(new_n831), .C(new_n1020), .Y(new_n1021));
  NOR4xp25_ASAP7_75t_L      g00765(.A(new_n1021), .B(new_n1018), .C(new_n1015), .D(new_n1019), .Y(new_n1022));
  OAI22xp33_ASAP7_75t_L     g00766(.A1(new_n1017), .A2(new_n1022), .B1(new_n981), .B2(new_n984), .Y(new_n1023));
  NAND4xp25_ASAP7_75t_L     g00767(.A(new_n983), .B(\a[8] ), .C(new_n982), .D(new_n979), .Y(new_n1024));
  A2O1A1Ixp33_ASAP7_75t_L   g00768(.A1(\b[7] ), .A2(new_n480), .B(new_n980), .C(new_n445), .Y(new_n1025));
  OAI22xp33_ASAP7_75t_L     g00769(.A1(new_n1015), .A2(new_n1021), .B1(new_n1019), .B2(new_n1018), .Y(new_n1026));
  NAND3xp33_ASAP7_75t_L     g00770(.A(new_n1016), .B(new_n1014), .C(new_n1013), .Y(new_n1027));
  NAND4xp25_ASAP7_75t_L     g00771(.A(new_n1027), .B(new_n1024), .C(new_n1025), .D(new_n1026), .Y(new_n1028));
  NAND2xp33_ASAP7_75t_L     g00772(.A(new_n1028), .B(new_n1023), .Y(new_n1029));
  A2O1A1Ixp33_ASAP7_75t_L   g00773(.A1(new_n932), .A2(new_n892), .B(new_n931), .C(new_n1029), .Y(new_n1030));
  INVx1_ASAP7_75t_L         g00774(.A(new_n1030), .Y(new_n1031));
  AOI211xp5_ASAP7_75t_L     g00775(.A1(new_n932), .A2(new_n892), .B(new_n931), .C(new_n1029), .Y(new_n1032));
  OAI21xp33_ASAP7_75t_L     g00776(.A1(new_n1032), .A2(new_n1031), .B(new_n975), .Y(new_n1033));
  AND2x2_ASAP7_75t_L        g00777(.A(new_n972), .B(new_n974), .Y(new_n1034));
  INVx1_ASAP7_75t_L         g00778(.A(new_n1032), .Y(new_n1035));
  NAND3xp33_ASAP7_75t_L     g00779(.A(new_n1034), .B(new_n1035), .C(new_n1030), .Y(new_n1036));
  AOI21xp33_ASAP7_75t_L     g00780(.A1(new_n1036), .A2(new_n1033), .B(new_n965), .Y(new_n1037));
  AOI21xp33_ASAP7_75t_L     g00781(.A1(new_n936), .A2(new_n933), .B(new_n939), .Y(new_n1038));
  A2O1A1Ixp33_ASAP7_75t_L   g00782(.A1(new_n761), .A2(new_n751), .B(new_n942), .C(new_n858), .Y(new_n1039));
  A2O1A1Ixp33_ASAP7_75t_L   g00783(.A1(new_n1039), .A2(new_n860), .B(new_n1038), .C(new_n940), .Y(new_n1040));
  NAND2xp33_ASAP7_75t_L     g00784(.A(new_n1033), .B(new_n1036), .Y(new_n1041));
  NOR2xp33_ASAP7_75t_L      g00785(.A(new_n1040), .B(new_n1041), .Y(new_n1042));
  OA21x2_ASAP7_75t_L        g00786(.A1(new_n1042), .A2(new_n1037), .B(new_n963), .Y(new_n1043));
  NOR3xp33_ASAP7_75t_L      g00787(.A(new_n963), .B(new_n1037), .C(new_n1042), .Y(new_n1044));
  NOR2xp33_ASAP7_75t_L      g00788(.A(new_n1044), .B(new_n1043), .Y(new_n1045));
  XOR2x2_ASAP7_75t_L        g00789(.A(new_n1045), .B(new_n947), .Y(\f[15] ));
  NOR2xp33_ASAP7_75t_L      g00790(.A(new_n1042), .B(new_n1037), .Y(new_n1047));
  NAND2xp33_ASAP7_75t_L     g00791(.A(new_n963), .B(new_n1047), .Y(new_n1048));
  INVx1_ASAP7_75t_L         g00792(.A(new_n953), .Y(new_n1049));
  NOR2xp33_ASAP7_75t_L      g00793(.A(\b[15] ), .B(\b[16] ), .Y(new_n1050));
  INVx1_ASAP7_75t_L         g00794(.A(\b[16] ), .Y(new_n1051));
  NOR2xp33_ASAP7_75t_L      g00795(.A(new_n952), .B(new_n1051), .Y(new_n1052));
  NOR2xp33_ASAP7_75t_L      g00796(.A(new_n1050), .B(new_n1052), .Y(new_n1053));
  INVx1_ASAP7_75t_L         g00797(.A(new_n1053), .Y(new_n1054));
  A2O1A1O1Ixp25_ASAP7_75t_L g00798(.A1(new_n950), .A2(new_n874), .B(new_n951), .C(new_n1049), .D(new_n1054), .Y(new_n1055));
  A2O1A1Ixp33_ASAP7_75t_L   g00799(.A1(new_n874), .A2(new_n950), .B(new_n955), .C(new_n1049), .Y(new_n1056));
  NOR2xp33_ASAP7_75t_L      g00800(.A(new_n1053), .B(new_n1056), .Y(new_n1057));
  NOR2xp33_ASAP7_75t_L      g00801(.A(new_n1055), .B(new_n1057), .Y(new_n1058));
  AOI22xp33_ASAP7_75t_L     g00802(.A1(new_n272), .A2(\b[16] ), .B1(new_n269), .B2(new_n1058), .Y(new_n1059));
  OAI221xp5_ASAP7_75t_L     g00803(.A1(new_n261), .A2(new_n952), .B1(new_n871), .B2(new_n277), .C(new_n1059), .Y(new_n1060));
  XNOR2x2_ASAP7_75t_L       g00804(.A(\a[2] ), .B(new_n1060), .Y(new_n1061));
  NOR3xp33_ASAP7_75t_L      g00805(.A(new_n1034), .B(new_n1031), .C(new_n1032), .Y(new_n1062));
  NAND2xp33_ASAP7_75t_L     g00806(.A(new_n342), .B(new_n800), .Y(new_n1063));
  OAI221xp5_ASAP7_75t_L     g00807(.A1(new_n368), .A2(new_n793), .B1(new_n763), .B2(new_n406), .C(new_n1063), .Y(new_n1064));
  AOI21xp33_ASAP7_75t_L     g00808(.A1(new_n366), .A2(\b[11] ), .B(new_n1064), .Y(new_n1065));
  NAND2xp33_ASAP7_75t_L     g00809(.A(\a[5] ), .B(new_n1065), .Y(new_n1066));
  A2O1A1Ixp33_ASAP7_75t_L   g00810(.A1(\b[11] ), .A2(new_n366), .B(new_n1064), .C(new_n339), .Y(new_n1067));
  NAND2xp33_ASAP7_75t_L     g00811(.A(new_n1067), .B(new_n1066), .Y(new_n1068));
  NOR2xp33_ASAP7_75t_L      g00812(.A(new_n981), .B(new_n984), .Y(new_n1069));
  NAND2xp33_ASAP7_75t_L     g00813(.A(new_n1026), .B(new_n1027), .Y(new_n1070));
  NOR2xp33_ASAP7_75t_L      g00814(.A(new_n1069), .B(new_n1070), .Y(new_n1071));
  A2O1A1O1Ixp25_ASAP7_75t_L g00815(.A1(new_n892), .A2(new_n932), .B(new_n931), .C(new_n1029), .D(new_n1071), .Y(new_n1072));
  INVx1_ASAP7_75t_L         g00816(.A(new_n1072), .Y(new_n1073));
  NAND2xp33_ASAP7_75t_L     g00817(.A(\b[8] ), .B(new_n480), .Y(new_n1074));
  NAND2xp33_ASAP7_75t_L     g00818(.A(\b[9] ), .B(new_n441), .Y(new_n1075));
  AOI22xp33_ASAP7_75t_L     g00819(.A1(new_n451), .A2(\b[10] ), .B1(new_n448), .B2(new_n852), .Y(new_n1076));
  NAND4xp25_ASAP7_75t_L     g00820(.A(new_n1076), .B(\a[8] ), .C(new_n1074), .D(new_n1075), .Y(new_n1077));
  NAND2xp33_ASAP7_75t_L     g00821(.A(new_n1075), .B(new_n1076), .Y(new_n1078));
  A2O1A1Ixp33_ASAP7_75t_L   g00822(.A1(\b[8] ), .A2(new_n480), .B(new_n1078), .C(new_n445), .Y(new_n1079));
  NAND2xp33_ASAP7_75t_L     g00823(.A(new_n1077), .B(new_n1079), .Y(new_n1080));
  NAND2xp33_ASAP7_75t_L     g00824(.A(new_n1013), .B(new_n1014), .Y(new_n1081));
  A2O1A1Ixp33_ASAP7_75t_L   g00825(.A1(new_n806), .A2(new_n830), .B(new_n835), .C(new_n922), .Y(new_n1082));
  NAND2xp33_ASAP7_75t_L     g00826(.A(new_n926), .B(new_n1082), .Y(new_n1083));
  NAND2xp33_ASAP7_75t_L     g00827(.A(new_n1006), .B(new_n1005), .Y(new_n1084));
  AOI21xp33_ASAP7_75t_L     g00828(.A1(new_n1012), .A2(new_n1010), .B(new_n1084), .Y(new_n1085));
  NAND2xp33_ASAP7_75t_L     g00829(.A(\b[7] ), .B(new_n600), .Y(new_n1086));
  OAI221xp5_ASAP7_75t_L     g00830(.A1(new_n382), .A2(new_n721), .B1(new_n675), .B2(new_n427), .C(new_n1086), .Y(new_n1087));
  AOI211xp5_ASAP7_75t_L     g00831(.A1(\b[5] ), .A2(new_n674), .B(new_n594), .C(new_n1087), .Y(new_n1088));
  A2O1A1Ixp33_ASAP7_75t_L   g00832(.A1(\b[5] ), .A2(new_n674), .B(new_n1087), .C(new_n594), .Y(new_n1089));
  INVx1_ASAP7_75t_L         g00833(.A(new_n1089), .Y(new_n1090));
  NOR3xp33_ASAP7_75t_L      g00834(.A(new_n985), .B(new_n910), .C(new_n914), .Y(new_n1091));
  NAND2xp33_ASAP7_75t_L     g00835(.A(new_n990), .B(new_n1091), .Y(new_n1092));
  A2O1A1Ixp33_ASAP7_75t_L   g00836(.A1(new_n993), .A2(new_n991), .B(new_n1004), .C(new_n1092), .Y(new_n1093));
  NAND2xp33_ASAP7_75t_L     g00837(.A(\b[2] ), .B(new_n908), .Y(new_n1094));
  NAND2xp33_ASAP7_75t_L     g00838(.A(\b[3] ), .B(new_n817), .Y(new_n1095));
  AOI22xp33_ASAP7_75t_L     g00839(.A1(new_n826), .A2(\b[4] ), .B1(new_n823), .B2(new_n328), .Y(new_n1096));
  NAND4xp25_ASAP7_75t_L     g00840(.A(new_n1096), .B(\a[14] ), .C(new_n1094), .D(new_n1095), .Y(new_n1097));
  AOI31xp33_ASAP7_75t_L     g00841(.A1(new_n1096), .A2(new_n1095), .A3(new_n1094), .B(\a[14] ), .Y(new_n1098));
  INVx1_ASAP7_75t_L         g00842(.A(new_n1098), .Y(new_n1099));
  NAND2xp33_ASAP7_75t_L     g00843(.A(\a[17] ), .B(new_n990), .Y(new_n1100));
  NAND2xp33_ASAP7_75t_L     g00844(.A(new_n988), .B(new_n987), .Y(new_n1101));
  XNOR2x2_ASAP7_75t_L       g00845(.A(\a[16] ), .B(\a[15] ), .Y(new_n1102));
  NOR2xp33_ASAP7_75t_L      g00846(.A(new_n1102), .B(new_n1101), .Y(new_n1103));
  NAND2xp33_ASAP7_75t_L     g00847(.A(\b[0] ), .B(new_n1103), .Y(new_n1104));
  INVx1_ASAP7_75t_L         g00848(.A(\a[16] ), .Y(new_n1105));
  NAND2xp33_ASAP7_75t_L     g00849(.A(\a[17] ), .B(new_n1105), .Y(new_n1106));
  INVx1_ASAP7_75t_L         g00850(.A(\a[17] ), .Y(new_n1107));
  NAND2xp33_ASAP7_75t_L     g00851(.A(\a[16] ), .B(new_n1107), .Y(new_n1108));
  AND2x2_ASAP7_75t_L        g00852(.A(new_n1106), .B(new_n1108), .Y(new_n1109));
  NOR2xp33_ASAP7_75t_L      g00853(.A(new_n989), .B(new_n1109), .Y(new_n1110));
  NAND2xp33_ASAP7_75t_L     g00854(.A(new_n271), .B(new_n1110), .Y(new_n1111));
  NAND2xp33_ASAP7_75t_L     g00855(.A(new_n1108), .B(new_n1106), .Y(new_n1112));
  NOR2xp33_ASAP7_75t_L      g00856(.A(new_n1112), .B(new_n989), .Y(new_n1113));
  NAND2xp33_ASAP7_75t_L     g00857(.A(\b[1] ), .B(new_n1113), .Y(new_n1114));
  NAND3xp33_ASAP7_75t_L     g00858(.A(new_n1111), .B(new_n1114), .C(new_n1104), .Y(new_n1115));
  XOR2x2_ASAP7_75t_L        g00859(.A(new_n1100), .B(new_n1115), .Y(new_n1116));
  NAND3xp33_ASAP7_75t_L     g00860(.A(new_n1099), .B(new_n1097), .C(new_n1116), .Y(new_n1117));
  INVx1_ASAP7_75t_L         g00861(.A(new_n1097), .Y(new_n1118));
  XNOR2x2_ASAP7_75t_L       g00862(.A(new_n1100), .B(new_n1115), .Y(new_n1119));
  OAI21xp33_ASAP7_75t_L     g00863(.A1(new_n1098), .A2(new_n1118), .B(new_n1119), .Y(new_n1120));
  NAND3xp33_ASAP7_75t_L     g00864(.A(new_n1093), .B(new_n1120), .C(new_n1117), .Y(new_n1121));
  OAI211xp5_ASAP7_75t_L     g00865(.A1(new_n276), .A2(new_n909), .B(new_n1002), .C(\a[14] ), .Y(new_n1122));
  A2O1A1Ixp33_ASAP7_75t_L   g00866(.A1(\b[1] ), .A2(new_n908), .B(new_n996), .C(new_n813), .Y(new_n1123));
  NAND2xp33_ASAP7_75t_L     g00867(.A(new_n1123), .B(new_n1122), .Y(new_n1124));
  MAJIxp5_ASAP7_75t_L       g00868(.A(new_n1124), .B(new_n990), .C(new_n1091), .Y(new_n1125));
  NOR3xp33_ASAP7_75t_L      g00869(.A(new_n1118), .B(new_n1098), .C(new_n1119), .Y(new_n1126));
  AOI21xp33_ASAP7_75t_L     g00870(.A1(new_n1099), .A2(new_n1097), .B(new_n1116), .Y(new_n1127));
  OAI21xp33_ASAP7_75t_L     g00871(.A1(new_n1126), .A2(new_n1127), .B(new_n1125), .Y(new_n1128));
  AOI211xp5_ASAP7_75t_L     g00872(.A1(new_n1121), .A2(new_n1128), .B(new_n1090), .C(new_n1088), .Y(new_n1129));
  INVx1_ASAP7_75t_L         g00873(.A(new_n1088), .Y(new_n1130));
  NOR3xp33_ASAP7_75t_L      g00874(.A(new_n1125), .B(new_n1127), .C(new_n1126), .Y(new_n1131));
  AOI21xp33_ASAP7_75t_L     g00875(.A1(new_n1120), .A2(new_n1117), .B(new_n1093), .Y(new_n1132));
  AOI211xp5_ASAP7_75t_L     g00876(.A1(new_n1130), .A2(new_n1089), .B(new_n1131), .C(new_n1132), .Y(new_n1133));
  NOR2xp33_ASAP7_75t_L      g00877(.A(new_n1129), .B(new_n1133), .Y(new_n1134));
  A2O1A1Ixp33_ASAP7_75t_L   g00878(.A1(new_n1083), .A2(new_n1081), .B(new_n1085), .C(new_n1134), .Y(new_n1135));
  O2A1O1Ixp33_ASAP7_75t_L   g00879(.A1(new_n1015), .A2(new_n1021), .B(new_n1081), .C(new_n1085), .Y(new_n1136));
  OAI21xp33_ASAP7_75t_L     g00880(.A1(new_n1129), .A2(new_n1133), .B(new_n1136), .Y(new_n1137));
  AO21x2_ASAP7_75t_L        g00881(.A1(new_n1137), .A2(new_n1135), .B(new_n1080), .Y(new_n1138));
  NAND3xp33_ASAP7_75t_L     g00882(.A(new_n1080), .B(new_n1135), .C(new_n1137), .Y(new_n1139));
  NAND3xp33_ASAP7_75t_L     g00883(.A(new_n1073), .B(new_n1138), .C(new_n1139), .Y(new_n1140));
  NAND2xp33_ASAP7_75t_L     g00884(.A(new_n1139), .B(new_n1138), .Y(new_n1141));
  NAND2xp33_ASAP7_75t_L     g00885(.A(new_n1072), .B(new_n1141), .Y(new_n1142));
  AOI21xp33_ASAP7_75t_L     g00886(.A1(new_n1140), .A2(new_n1142), .B(new_n1068), .Y(new_n1143));
  XNOR2x2_ASAP7_75t_L       g00887(.A(new_n339), .B(new_n1065), .Y(new_n1144));
  O2A1O1Ixp33_ASAP7_75t_L   g00888(.A1(new_n1069), .A2(new_n1070), .B(new_n1030), .C(new_n1141), .Y(new_n1145));
  AOI21xp33_ASAP7_75t_L     g00889(.A1(new_n1139), .A2(new_n1138), .B(new_n1073), .Y(new_n1146));
  NOR3xp33_ASAP7_75t_L      g00890(.A(new_n1144), .B(new_n1146), .C(new_n1145), .Y(new_n1147));
  NOR2xp33_ASAP7_75t_L      g00891(.A(new_n1143), .B(new_n1147), .Y(new_n1148));
  A2O1A1Ixp33_ASAP7_75t_L   g00892(.A1(new_n1041), .A2(new_n1040), .B(new_n1062), .C(new_n1148), .Y(new_n1149));
  NOR2xp33_ASAP7_75t_L      g00893(.A(new_n1032), .B(new_n1031), .Y(new_n1150));
  MAJIxp5_ASAP7_75t_L       g00894(.A(new_n1040), .B(new_n975), .C(new_n1150), .Y(new_n1151));
  OAI21xp33_ASAP7_75t_L     g00895(.A1(new_n1143), .A2(new_n1147), .B(new_n1151), .Y(new_n1152));
  NAND3xp33_ASAP7_75t_L     g00896(.A(new_n1149), .B(new_n1152), .C(new_n1061), .Y(new_n1153));
  AO21x2_ASAP7_75t_L        g00897(.A1(new_n1152), .A2(new_n1149), .B(new_n1061), .Y(new_n1154));
  NAND2xp33_ASAP7_75t_L     g00898(.A(new_n1153), .B(new_n1154), .Y(new_n1155));
  INVx1_ASAP7_75t_L         g00899(.A(new_n1155), .Y(new_n1156));
  O2A1O1Ixp33_ASAP7_75t_L   g00900(.A1(new_n947), .A2(new_n1045), .B(new_n1048), .C(new_n1156), .Y(new_n1157));
  OAI21xp33_ASAP7_75t_L     g00901(.A1(new_n1045), .A2(new_n947), .B(new_n1048), .Y(new_n1158));
  NOR2xp33_ASAP7_75t_L      g00902(.A(new_n1155), .B(new_n1158), .Y(new_n1159));
  NOR2xp33_ASAP7_75t_L      g00903(.A(new_n1159), .B(new_n1157), .Y(\f[16] ));
  INVx1_ASAP7_75t_L         g00904(.A(new_n1062), .Y(new_n1161));
  A2O1A1Ixp33_ASAP7_75t_L   g00905(.A1(new_n1033), .A2(new_n1036), .B(new_n965), .C(new_n1161), .Y(new_n1162));
  OAI21xp33_ASAP7_75t_L     g00906(.A1(new_n1145), .A2(new_n1146), .B(new_n1144), .Y(new_n1163));
  NAND2xp33_ASAP7_75t_L     g00907(.A(\b[13] ), .B(new_n334), .Y(new_n1164));
  OAI221xp5_ASAP7_75t_L     g00908(.A1(new_n368), .A2(new_n871), .B1(new_n367), .B2(new_n878), .C(new_n1164), .Y(new_n1165));
  AOI21xp33_ASAP7_75t_L     g00909(.A1(new_n366), .A2(\b[12] ), .B(new_n1165), .Y(new_n1166));
  NAND2xp33_ASAP7_75t_L     g00910(.A(\a[5] ), .B(new_n1166), .Y(new_n1167));
  A2O1A1Ixp33_ASAP7_75t_L   g00911(.A1(\b[12] ), .A2(new_n366), .B(new_n1165), .C(new_n339), .Y(new_n1168));
  NAND2xp33_ASAP7_75t_L     g00912(.A(new_n1168), .B(new_n1167), .Y(new_n1169));
  AOI21xp33_ASAP7_75t_L     g00913(.A1(new_n1137), .A2(new_n1135), .B(new_n1080), .Y(new_n1170));
  OAI21xp33_ASAP7_75t_L     g00914(.A1(new_n1170), .A2(new_n1072), .B(new_n1139), .Y(new_n1171));
  NAND2xp33_ASAP7_75t_L     g00915(.A(\b[9] ), .B(new_n480), .Y(new_n1172));
  NAND2xp33_ASAP7_75t_L     g00916(.A(\b[10] ), .B(new_n441), .Y(new_n1173));
  AOI32xp33_ASAP7_75t_L     g00917(.A1(new_n700), .A2(new_n698), .A3(new_n448), .B1(new_n451), .B2(\b[11] ), .Y(new_n1174));
  NAND4xp25_ASAP7_75t_L     g00918(.A(new_n1174), .B(\a[8] ), .C(new_n1172), .D(new_n1173), .Y(new_n1175));
  NAND2xp33_ASAP7_75t_L     g00919(.A(new_n1173), .B(new_n1174), .Y(new_n1176));
  A2O1A1Ixp33_ASAP7_75t_L   g00920(.A1(\b[9] ), .A2(new_n480), .B(new_n1176), .C(new_n445), .Y(new_n1177));
  NAND2xp33_ASAP7_75t_L     g00921(.A(new_n1175), .B(new_n1177), .Y(new_n1178));
  AO21x2_ASAP7_75t_L        g00922(.A1(new_n1012), .A2(new_n1010), .B(new_n1084), .Y(new_n1179));
  OAI211xp5_ASAP7_75t_L     g00923(.A1(new_n1088), .A2(new_n1090), .B(new_n1121), .C(new_n1128), .Y(new_n1180));
  A2O1A1Ixp33_ASAP7_75t_L   g00924(.A1(new_n1026), .A2(new_n1179), .B(new_n1129), .C(new_n1180), .Y(new_n1181));
  NAND2xp33_ASAP7_75t_L     g00925(.A(\b[7] ), .B(new_n590), .Y(new_n1182));
  OAI221xp5_ASAP7_75t_L     g00926(.A1(new_n676), .A2(new_n503), .B1(new_n675), .B2(new_n509), .C(new_n1182), .Y(new_n1183));
  AOI211xp5_ASAP7_75t_L     g00927(.A1(\b[6] ), .A2(new_n674), .B(new_n594), .C(new_n1183), .Y(new_n1184));
  INVx1_ASAP7_75t_L         g00928(.A(new_n1184), .Y(new_n1185));
  A2O1A1Ixp33_ASAP7_75t_L   g00929(.A1(\b[6] ), .A2(new_n674), .B(new_n1183), .C(new_n594), .Y(new_n1186));
  NAND2xp33_ASAP7_75t_L     g00930(.A(\b[4] ), .B(new_n817), .Y(new_n1187));
  OAI221xp5_ASAP7_75t_L     g00931(.A1(new_n912), .A2(new_n353), .B1(new_n911), .B2(new_n359), .C(new_n1187), .Y(new_n1188));
  AOI211xp5_ASAP7_75t_L     g00932(.A1(\b[3] ), .A2(new_n908), .B(new_n813), .C(new_n1188), .Y(new_n1189));
  A2O1A1Ixp33_ASAP7_75t_L   g00933(.A1(\b[3] ), .A2(new_n908), .B(new_n1188), .C(new_n813), .Y(new_n1190));
  INVx1_ASAP7_75t_L         g00934(.A(new_n1190), .Y(new_n1191));
  AND3x1_ASAP7_75t_L        g00935(.A(new_n1111), .B(new_n1114), .C(new_n1104), .Y(new_n1192));
  INVx1_ASAP7_75t_L         g00936(.A(new_n1102), .Y(new_n1193));
  NOR3xp33_ASAP7_75t_L      g00937(.A(new_n1109), .B(new_n1193), .C(new_n1101), .Y(new_n1194));
  INVx1_ASAP7_75t_L         g00938(.A(new_n1194), .Y(new_n1195));
  NOR2xp33_ASAP7_75t_L      g00939(.A(new_n258), .B(new_n1195), .Y(new_n1196));
  NAND2xp33_ASAP7_75t_L     g00940(.A(new_n1112), .B(new_n1101), .Y(new_n1197));
  NAND2xp33_ASAP7_75t_L     g00941(.A(new_n1101), .B(new_n1109), .Y(new_n1198));
  NAND2xp33_ASAP7_75t_L     g00942(.A(\b[1] ), .B(new_n1103), .Y(new_n1199));
  OAI221xp5_ASAP7_75t_L     g00943(.A1(new_n1197), .A2(new_n283), .B1(new_n278), .B2(new_n1198), .C(new_n1199), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g00944(.A(new_n1200), .B(new_n1196), .Y(new_n1201));
  A2O1A1Ixp33_ASAP7_75t_L   g00945(.A1(new_n992), .A2(new_n1192), .B(new_n1107), .C(new_n1201), .Y(new_n1202));
  O2A1O1Ixp33_ASAP7_75t_L   g00946(.A1(new_n258), .A2(new_n989), .B(new_n1192), .C(new_n1107), .Y(new_n1203));
  A2O1A1Ixp33_ASAP7_75t_L   g00947(.A1(\b[0] ), .A2(new_n1194), .B(new_n1200), .C(new_n1203), .Y(new_n1204));
  AOI211xp5_ASAP7_75t_L     g00948(.A1(new_n1204), .A2(new_n1202), .B(new_n1189), .C(new_n1191), .Y(new_n1205));
  NAND2xp33_ASAP7_75t_L     g00949(.A(\b[3] ), .B(new_n908), .Y(new_n1206));
  AOI22xp33_ASAP7_75t_L     g00950(.A1(new_n826), .A2(\b[5] ), .B1(new_n823), .B2(new_n360), .Y(new_n1207));
  NAND4xp25_ASAP7_75t_L     g00951(.A(new_n1207), .B(\a[14] ), .C(new_n1206), .D(new_n1187), .Y(new_n1208));
  INVx1_ASAP7_75t_L         g00952(.A(new_n1202), .Y(new_n1209));
  A2O1A1Ixp33_ASAP7_75t_L   g00953(.A1(\b[0] ), .A2(new_n1101), .B(new_n1115), .C(\a[17] ), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g00954(.A(new_n1197), .B(new_n283), .Y(new_n1211));
  AOI221xp5_ASAP7_75t_L     g00955(.A1(\b[2] ), .A2(new_n1113), .B1(new_n1103), .B2(\b[1] ), .C(new_n1211), .Y(new_n1212));
  O2A1O1Ixp33_ASAP7_75t_L   g00956(.A1(new_n1195), .A2(new_n258), .B(new_n1212), .C(new_n1210), .Y(new_n1213));
  AOI211xp5_ASAP7_75t_L     g00957(.A1(new_n1190), .A2(new_n1208), .B(new_n1213), .C(new_n1209), .Y(new_n1214));
  NOR2xp33_ASAP7_75t_L      g00958(.A(new_n1214), .B(new_n1205), .Y(new_n1215));
  NAND3xp33_ASAP7_75t_L     g00959(.A(new_n1215), .B(new_n1121), .C(new_n1120), .Y(new_n1216));
  A2O1A1Ixp33_ASAP7_75t_L   g00960(.A1(new_n1005), .A2(new_n1092), .B(new_n1126), .C(new_n1120), .Y(new_n1217));
  OAI21xp33_ASAP7_75t_L     g00961(.A1(new_n1205), .A2(new_n1214), .B(new_n1217), .Y(new_n1218));
  NAND4xp25_ASAP7_75t_L     g00962(.A(new_n1216), .B(new_n1218), .C(new_n1185), .D(new_n1186), .Y(new_n1219));
  INVx1_ASAP7_75t_L         g00963(.A(new_n1186), .Y(new_n1220));
  NOR3xp33_ASAP7_75t_L      g00964(.A(new_n1217), .B(new_n1205), .C(new_n1214), .Y(new_n1221));
  O2A1O1Ixp33_ASAP7_75t_L   g00965(.A1(new_n1125), .A2(new_n1126), .B(new_n1120), .C(new_n1215), .Y(new_n1222));
  OAI22xp33_ASAP7_75t_L     g00966(.A1(new_n1221), .A2(new_n1222), .B1(new_n1184), .B2(new_n1220), .Y(new_n1223));
  NAND3xp33_ASAP7_75t_L     g00967(.A(new_n1181), .B(new_n1219), .C(new_n1223), .Y(new_n1224));
  OAI211xp5_ASAP7_75t_L     g00968(.A1(new_n1132), .A2(new_n1131), .B(new_n1089), .C(new_n1130), .Y(new_n1225));
  A2O1A1O1Ixp25_ASAP7_75t_L g00969(.A1(new_n1081), .A2(new_n1083), .B(new_n1085), .C(new_n1225), .D(new_n1133), .Y(new_n1226));
  NOR4xp25_ASAP7_75t_L      g00970(.A(new_n1221), .B(new_n1222), .C(new_n1184), .D(new_n1220), .Y(new_n1227));
  AOI22xp33_ASAP7_75t_L     g00971(.A1(new_n1186), .A2(new_n1185), .B1(new_n1218), .B2(new_n1216), .Y(new_n1228));
  OAI21xp33_ASAP7_75t_L     g00972(.A1(new_n1227), .A2(new_n1228), .B(new_n1226), .Y(new_n1229));
  AOI21xp33_ASAP7_75t_L     g00973(.A1(new_n1229), .A2(new_n1224), .B(new_n1178), .Y(new_n1230));
  AND3x1_ASAP7_75t_L        g00974(.A(new_n1229), .B(new_n1178), .C(new_n1224), .Y(new_n1231));
  NOR2xp33_ASAP7_75t_L      g00975(.A(new_n1230), .B(new_n1231), .Y(new_n1232));
  NAND2xp33_ASAP7_75t_L     g00976(.A(new_n1232), .B(new_n1171), .Y(new_n1233));
  OAI221xp5_ASAP7_75t_L     g00977(.A1(new_n1072), .A2(new_n1170), .B1(new_n1230), .B2(new_n1231), .C(new_n1139), .Y(new_n1234));
  AOI21xp33_ASAP7_75t_L     g00978(.A1(new_n1233), .A2(new_n1234), .B(new_n1169), .Y(new_n1235));
  AND3x1_ASAP7_75t_L        g00979(.A(new_n1233), .B(new_n1169), .C(new_n1234), .Y(new_n1236));
  NOR2xp33_ASAP7_75t_L      g00980(.A(new_n1235), .B(new_n1236), .Y(new_n1237));
  A2O1A1Ixp33_ASAP7_75t_L   g00981(.A1(new_n1163), .A2(new_n1162), .B(new_n1147), .C(new_n1237), .Y(new_n1238));
  A2O1A1O1Ixp25_ASAP7_75t_L g00982(.A1(new_n1040), .A2(new_n1041), .B(new_n1062), .C(new_n1163), .D(new_n1147), .Y(new_n1239));
  OAI21xp33_ASAP7_75t_L     g00983(.A1(new_n1235), .A2(new_n1236), .B(new_n1239), .Y(new_n1240));
  NAND2xp33_ASAP7_75t_L     g00984(.A(\b[15] ), .B(new_n291), .Y(new_n1241));
  NAND2xp33_ASAP7_75t_L     g00985(.A(\b[16] ), .B(new_n380), .Y(new_n1242));
  NOR2xp33_ASAP7_75t_L      g00986(.A(\b[16] ), .B(\b[17] ), .Y(new_n1243));
  INVx1_ASAP7_75t_L         g00987(.A(\b[17] ), .Y(new_n1244));
  NOR2xp33_ASAP7_75t_L      g00988(.A(new_n1051), .B(new_n1244), .Y(new_n1245));
  NOR2xp33_ASAP7_75t_L      g00989(.A(new_n1243), .B(new_n1245), .Y(new_n1246));
  A2O1A1Ixp33_ASAP7_75t_L   g00990(.A1(new_n1056), .A2(new_n1053), .B(new_n1052), .C(new_n1246), .Y(new_n1247));
  A2O1A1O1Ixp25_ASAP7_75t_L g00991(.A1(new_n954), .A2(new_n957), .B(new_n953), .C(new_n1053), .D(new_n1052), .Y(new_n1248));
  INVx1_ASAP7_75t_L         g00992(.A(new_n1246), .Y(new_n1249));
  NAND2xp33_ASAP7_75t_L     g00993(.A(new_n1249), .B(new_n1248), .Y(new_n1250));
  NAND2xp33_ASAP7_75t_L     g00994(.A(new_n1247), .B(new_n1250), .Y(new_n1251));
  INVx1_ASAP7_75t_L         g00995(.A(new_n1251), .Y(new_n1252));
  AOI22xp33_ASAP7_75t_L     g00996(.A1(new_n272), .A2(\b[17] ), .B1(new_n269), .B2(new_n1252), .Y(new_n1253));
  NAND4xp25_ASAP7_75t_L     g00997(.A(new_n1253), .B(\a[2] ), .C(new_n1241), .D(new_n1242), .Y(new_n1254));
  NAND2xp33_ASAP7_75t_L     g00998(.A(new_n1242), .B(new_n1253), .Y(new_n1255));
  A2O1A1Ixp33_ASAP7_75t_L   g00999(.A1(\b[15] ), .A2(new_n291), .B(new_n1255), .C(new_n265), .Y(new_n1256));
  NAND4xp25_ASAP7_75t_L     g01000(.A(new_n1238), .B(new_n1256), .C(new_n1254), .D(new_n1240), .Y(new_n1257));
  NOR3xp33_ASAP7_75t_L      g01001(.A(new_n1239), .B(new_n1235), .C(new_n1236), .Y(new_n1258));
  NAND3xp33_ASAP7_75t_L     g01002(.A(new_n1140), .B(new_n1068), .C(new_n1142), .Y(new_n1259));
  OAI21xp33_ASAP7_75t_L     g01003(.A1(new_n1143), .A2(new_n1151), .B(new_n1259), .Y(new_n1260));
  NOR2xp33_ASAP7_75t_L      g01004(.A(new_n1237), .B(new_n1260), .Y(new_n1261));
  NAND2xp33_ASAP7_75t_L     g01005(.A(new_n1254), .B(new_n1256), .Y(new_n1262));
  OAI21xp33_ASAP7_75t_L     g01006(.A1(new_n1258), .A2(new_n1261), .B(new_n1262), .Y(new_n1263));
  NAND2xp33_ASAP7_75t_L     g01007(.A(new_n1257), .B(new_n1263), .Y(new_n1264));
  NAND2xp33_ASAP7_75t_L     g01008(.A(new_n1152), .B(new_n1149), .Y(new_n1265));
  NOR2xp33_ASAP7_75t_L      g01009(.A(new_n1061), .B(new_n1265), .Y(new_n1266));
  A2O1A1Ixp33_ASAP7_75t_L   g01010(.A1(new_n1158), .A2(new_n1155), .B(new_n1266), .C(new_n1264), .Y(new_n1267));
  OR3x1_ASAP7_75t_L         g01011(.A(new_n1157), .B(new_n1264), .C(new_n1266), .Y(new_n1268));
  AND2x2_ASAP7_75t_L        g01012(.A(new_n1267), .B(new_n1268), .Y(\f[17] ));
  NAND3xp33_ASAP7_75t_L     g01013(.A(new_n1233), .B(new_n1169), .C(new_n1234), .Y(new_n1270));
  OAI21xp33_ASAP7_75t_L     g01014(.A1(new_n1235), .A2(new_n1239), .B(new_n1270), .Y(new_n1271));
  NAND2xp33_ASAP7_75t_L     g01015(.A(\b[13] ), .B(new_n366), .Y(new_n1272));
  NAND2xp33_ASAP7_75t_L     g01016(.A(\b[14] ), .B(new_n334), .Y(new_n1273));
  AOI22xp33_ASAP7_75t_L     g01017(.A1(new_n345), .A2(\b[15] ), .B1(new_n342), .B2(new_n959), .Y(new_n1274));
  NAND4xp25_ASAP7_75t_L     g01018(.A(new_n1274), .B(\a[5] ), .C(new_n1272), .D(new_n1273), .Y(new_n1275));
  NAND2xp33_ASAP7_75t_L     g01019(.A(new_n1273), .B(new_n1274), .Y(new_n1276));
  A2O1A1Ixp33_ASAP7_75t_L   g01020(.A1(\b[13] ), .A2(new_n366), .B(new_n1276), .C(new_n339), .Y(new_n1277));
  AND2x2_ASAP7_75t_L        g01021(.A(new_n1275), .B(new_n1277), .Y(new_n1278));
  AOI21xp33_ASAP7_75t_L     g01022(.A1(new_n1171), .A2(new_n1232), .B(new_n1231), .Y(new_n1279));
  NAND2xp33_ASAP7_75t_L     g01023(.A(\b[10] ), .B(new_n480), .Y(new_n1280));
  NAND2xp33_ASAP7_75t_L     g01024(.A(\b[11] ), .B(new_n441), .Y(new_n1281));
  AOI22xp33_ASAP7_75t_L     g01025(.A1(new_n451), .A2(\b[12] ), .B1(new_n448), .B2(new_n970), .Y(new_n1282));
  NAND4xp25_ASAP7_75t_L     g01026(.A(new_n1282), .B(\a[8] ), .C(new_n1280), .D(new_n1281), .Y(new_n1283));
  NAND2xp33_ASAP7_75t_L     g01027(.A(new_n1281), .B(new_n1282), .Y(new_n1284));
  A2O1A1Ixp33_ASAP7_75t_L   g01028(.A1(\b[10] ), .A2(new_n480), .B(new_n1284), .C(new_n445), .Y(new_n1285));
  NAND2xp33_ASAP7_75t_L     g01029(.A(new_n1283), .B(new_n1285), .Y(new_n1286));
  NOR2xp33_ASAP7_75t_L      g01030(.A(new_n1107), .B(new_n1115), .Y(new_n1287));
  INVx1_ASAP7_75t_L         g01031(.A(\a[18] ), .Y(new_n1288));
  NAND2xp33_ASAP7_75t_L     g01032(.A(\a[17] ), .B(new_n1288), .Y(new_n1289));
  NAND2xp33_ASAP7_75t_L     g01033(.A(\a[18] ), .B(new_n1107), .Y(new_n1290));
  AND2x2_ASAP7_75t_L        g01034(.A(new_n1289), .B(new_n1290), .Y(new_n1291));
  NOR2xp33_ASAP7_75t_L      g01035(.A(new_n258), .B(new_n1291), .Y(new_n1292));
  INVx1_ASAP7_75t_L         g01036(.A(new_n1292), .Y(new_n1293));
  AOI31xp33_ASAP7_75t_L     g01037(.A1(new_n1287), .A2(new_n992), .A3(new_n1201), .B(new_n1293), .Y(new_n1294));
  NAND5xp2_ASAP7_75t_L      g01038(.A(new_n1114), .B(new_n1111), .C(new_n1104), .D(new_n992), .E(\a[17] ), .Y(new_n1295));
  OAI21xp33_ASAP7_75t_L     g01039(.A1(new_n258), .A2(new_n1195), .B(new_n1212), .Y(new_n1296));
  NOR3xp33_ASAP7_75t_L      g01040(.A(new_n1296), .B(new_n1292), .C(new_n1295), .Y(new_n1297));
  NAND2xp33_ASAP7_75t_L     g01041(.A(new_n1193), .B(new_n989), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g01042(.A(new_n278), .B(new_n1298), .Y(new_n1299));
  AOI221xp5_ASAP7_75t_L     g01043(.A1(new_n1113), .A2(\b[3] ), .B1(new_n1110), .B2(new_n1000), .C(new_n1299), .Y(new_n1300));
  OAI211xp5_ASAP7_75t_L     g01044(.A1(new_n276), .A2(new_n1195), .B(new_n1300), .C(\a[17] ), .Y(new_n1301));
  NAND2xp33_ASAP7_75t_L     g01045(.A(\b[3] ), .B(new_n1113), .Y(new_n1302));
  OAI221xp5_ASAP7_75t_L     g01046(.A1(new_n278), .A2(new_n1298), .B1(new_n1197), .B2(new_n303), .C(new_n1302), .Y(new_n1303));
  A2O1A1Ixp33_ASAP7_75t_L   g01047(.A1(\b[1] ), .A2(new_n1194), .B(new_n1303), .C(new_n1107), .Y(new_n1304));
  NAND2xp33_ASAP7_75t_L     g01048(.A(new_n1304), .B(new_n1301), .Y(new_n1305));
  OAI21xp33_ASAP7_75t_L     g01049(.A1(new_n1297), .A2(new_n1294), .B(new_n1305), .Y(new_n1306));
  OAI21xp33_ASAP7_75t_L     g01050(.A1(new_n1295), .A2(new_n1296), .B(new_n1292), .Y(new_n1307));
  NAND4xp25_ASAP7_75t_L     g01051(.A(new_n1287), .B(new_n1201), .C(new_n1293), .D(new_n992), .Y(new_n1308));
  NAND4xp25_ASAP7_75t_L     g01052(.A(new_n1307), .B(new_n1308), .C(new_n1304), .D(new_n1301), .Y(new_n1309));
  NAND2xp33_ASAP7_75t_L     g01053(.A(\b[4] ), .B(new_n908), .Y(new_n1310));
  NAND2xp33_ASAP7_75t_L     g01054(.A(\b[5] ), .B(new_n817), .Y(new_n1311));
  AOI22xp33_ASAP7_75t_L     g01055(.A1(new_n826), .A2(\b[6] ), .B1(new_n823), .B2(new_n389), .Y(new_n1312));
  NAND4xp25_ASAP7_75t_L     g01056(.A(new_n1312), .B(\a[14] ), .C(new_n1310), .D(new_n1311), .Y(new_n1313));
  OAI221xp5_ASAP7_75t_L     g01057(.A1(new_n912), .A2(new_n382), .B1(new_n911), .B2(new_n540), .C(new_n1311), .Y(new_n1314));
  A2O1A1Ixp33_ASAP7_75t_L   g01058(.A1(\b[4] ), .A2(new_n908), .B(new_n1314), .C(new_n813), .Y(new_n1315));
  AND4x1_ASAP7_75t_L        g01059(.A(new_n1315), .B(new_n1313), .C(new_n1309), .D(new_n1306), .Y(new_n1316));
  AOI22xp33_ASAP7_75t_L     g01060(.A1(new_n1306), .A2(new_n1309), .B1(new_n1313), .B2(new_n1315), .Y(new_n1317));
  OAI211xp5_ASAP7_75t_L     g01061(.A1(new_n1213), .A2(new_n1209), .B(new_n1190), .C(new_n1208), .Y(new_n1318));
  A2O1A1O1Ixp25_ASAP7_75t_L g01062(.A1(new_n1117), .A2(new_n1093), .B(new_n1127), .C(new_n1318), .D(new_n1214), .Y(new_n1319));
  OR3x1_ASAP7_75t_L         g01063(.A(new_n1319), .B(new_n1316), .C(new_n1317), .Y(new_n1320));
  OAI21xp33_ASAP7_75t_L     g01064(.A1(new_n1316), .A2(new_n1317), .B(new_n1319), .Y(new_n1321));
  NAND2xp33_ASAP7_75t_L     g01065(.A(\b[7] ), .B(new_n674), .Y(new_n1322));
  NAND2xp33_ASAP7_75t_L     g01066(.A(\b[8] ), .B(new_n590), .Y(new_n1323));
  OAI221xp5_ASAP7_75t_L     g01067(.A1(new_n676), .A2(new_n559), .B1(new_n675), .B2(new_n978), .C(new_n1323), .Y(new_n1324));
  INVx1_ASAP7_75t_L         g01068(.A(new_n1324), .Y(new_n1325));
  NAND3xp33_ASAP7_75t_L     g01069(.A(new_n1325), .B(new_n1322), .C(\a[11] ), .Y(new_n1326));
  A2O1A1Ixp33_ASAP7_75t_L   g01070(.A1(\b[7] ), .A2(new_n674), .B(new_n1324), .C(new_n594), .Y(new_n1327));
  AOI22xp33_ASAP7_75t_L     g01071(.A1(new_n1326), .A2(new_n1327), .B1(new_n1321), .B2(new_n1320), .Y(new_n1328));
  AND4x1_ASAP7_75t_L        g01072(.A(new_n1320), .B(new_n1327), .C(new_n1326), .D(new_n1321), .Y(new_n1329));
  NOR2xp33_ASAP7_75t_L      g01073(.A(new_n1328), .B(new_n1329), .Y(new_n1330));
  A2O1A1Ixp33_ASAP7_75t_L   g01074(.A1(new_n1219), .A2(new_n1181), .B(new_n1228), .C(new_n1330), .Y(new_n1331));
  A2O1A1Ixp33_ASAP7_75t_L   g01075(.A1(new_n1014), .A2(new_n1013), .B(new_n1016), .C(new_n1179), .Y(new_n1332));
  A2O1A1O1Ixp25_ASAP7_75t_L g01076(.A1(new_n1225), .A2(new_n1332), .B(new_n1133), .C(new_n1219), .D(new_n1228), .Y(new_n1333));
  OAI21xp33_ASAP7_75t_L     g01077(.A1(new_n1328), .A2(new_n1329), .B(new_n1333), .Y(new_n1334));
  AOI21xp33_ASAP7_75t_L     g01078(.A1(new_n1331), .A2(new_n1334), .B(new_n1286), .Y(new_n1335));
  NOR3xp33_ASAP7_75t_L      g01079(.A(new_n1333), .B(new_n1328), .C(new_n1329), .Y(new_n1336));
  OAI21xp33_ASAP7_75t_L     g01080(.A1(new_n1227), .A2(new_n1226), .B(new_n1223), .Y(new_n1337));
  NOR2xp33_ASAP7_75t_L      g01081(.A(new_n1337), .B(new_n1330), .Y(new_n1338));
  AOI211xp5_ASAP7_75t_L     g01082(.A1(new_n1283), .A2(new_n1285), .B(new_n1336), .C(new_n1338), .Y(new_n1339));
  NOR3xp33_ASAP7_75t_L      g01083(.A(new_n1279), .B(new_n1335), .C(new_n1339), .Y(new_n1340));
  AO21x2_ASAP7_75t_L        g01084(.A1(new_n1232), .A2(new_n1171), .B(new_n1231), .Y(new_n1341));
  NOR2xp33_ASAP7_75t_L      g01085(.A(new_n1339), .B(new_n1335), .Y(new_n1342));
  NOR2xp33_ASAP7_75t_L      g01086(.A(new_n1342), .B(new_n1341), .Y(new_n1343));
  NOR3xp33_ASAP7_75t_L      g01087(.A(new_n1343), .B(new_n1278), .C(new_n1340), .Y(new_n1344));
  INVx1_ASAP7_75t_L         g01088(.A(new_n1344), .Y(new_n1345));
  OAI21xp33_ASAP7_75t_L     g01089(.A1(new_n1340), .A2(new_n1343), .B(new_n1278), .Y(new_n1346));
  NAND3xp33_ASAP7_75t_L     g01090(.A(new_n1271), .B(new_n1345), .C(new_n1346), .Y(new_n1347));
  INVx1_ASAP7_75t_L         g01091(.A(new_n1235), .Y(new_n1348));
  A2O1A1O1Ixp25_ASAP7_75t_L g01092(.A1(new_n1148), .A2(new_n1162), .B(new_n1147), .C(new_n1348), .D(new_n1236), .Y(new_n1349));
  INVx1_ASAP7_75t_L         g01093(.A(new_n1346), .Y(new_n1350));
  OAI21xp33_ASAP7_75t_L     g01094(.A1(new_n1344), .A2(new_n1350), .B(new_n1349), .Y(new_n1351));
  INVx1_ASAP7_75t_L         g01095(.A(new_n1052), .Y(new_n1352));
  A2O1A1Ixp33_ASAP7_75t_L   g01096(.A1(new_n957), .A2(new_n954), .B(new_n953), .C(new_n1053), .Y(new_n1353));
  INVx1_ASAP7_75t_L         g01097(.A(new_n1245), .Y(new_n1354));
  NOR2xp33_ASAP7_75t_L      g01098(.A(\b[17] ), .B(\b[18] ), .Y(new_n1355));
  INVx1_ASAP7_75t_L         g01099(.A(\b[18] ), .Y(new_n1356));
  NOR2xp33_ASAP7_75t_L      g01100(.A(new_n1244), .B(new_n1356), .Y(new_n1357));
  NOR2xp33_ASAP7_75t_L      g01101(.A(new_n1355), .B(new_n1357), .Y(new_n1358));
  INVx1_ASAP7_75t_L         g01102(.A(new_n1358), .Y(new_n1359));
  A2O1A1O1Ixp25_ASAP7_75t_L g01103(.A1(new_n1352), .A2(new_n1353), .B(new_n1243), .C(new_n1354), .D(new_n1359), .Y(new_n1360));
  A2O1A1Ixp33_ASAP7_75t_L   g01104(.A1(new_n1353), .A2(new_n1352), .B(new_n1249), .C(new_n1354), .Y(new_n1361));
  NOR2xp33_ASAP7_75t_L      g01105(.A(new_n1358), .B(new_n1361), .Y(new_n1362));
  NOR2xp33_ASAP7_75t_L      g01106(.A(new_n1360), .B(new_n1362), .Y(new_n1363));
  AOI22xp33_ASAP7_75t_L     g01107(.A1(new_n272), .A2(\b[18] ), .B1(new_n269), .B2(new_n1363), .Y(new_n1364));
  OAI221xp5_ASAP7_75t_L     g01108(.A1(new_n261), .A2(new_n1244), .B1(new_n1051), .B2(new_n277), .C(new_n1364), .Y(new_n1365));
  XNOR2x2_ASAP7_75t_L       g01109(.A(\a[2] ), .B(new_n1365), .Y(new_n1366));
  AND3x1_ASAP7_75t_L        g01110(.A(new_n1351), .B(new_n1347), .C(new_n1366), .Y(new_n1367));
  AOI21xp33_ASAP7_75t_L     g01111(.A1(new_n1351), .A2(new_n1347), .B(new_n1366), .Y(new_n1368));
  NOR2xp33_ASAP7_75t_L      g01112(.A(new_n1368), .B(new_n1367), .Y(new_n1369));
  AND3x1_ASAP7_75t_L        g01113(.A(new_n1238), .B(new_n1262), .C(new_n1240), .Y(new_n1370));
  A2O1A1O1Ixp25_ASAP7_75t_L g01114(.A1(new_n1155), .A2(new_n1158), .B(new_n1266), .C(new_n1264), .D(new_n1370), .Y(new_n1371));
  XOR2x2_ASAP7_75t_L        g01115(.A(new_n1369), .B(new_n1371), .Y(\f[18] ));
  OAI211xp5_ASAP7_75t_L     g01116(.A1(new_n1336), .A2(new_n1338), .B(new_n1285), .C(new_n1283), .Y(new_n1373));
  NAND2xp33_ASAP7_75t_L     g01117(.A(new_n1309), .B(new_n1306), .Y(new_n1374));
  INVx1_ASAP7_75t_L         g01118(.A(new_n1313), .Y(new_n1375));
  AOI31xp33_ASAP7_75t_L     g01119(.A1(new_n1312), .A2(new_n1311), .A3(new_n1310), .B(\a[14] ), .Y(new_n1376));
  NOR2xp33_ASAP7_75t_L      g01120(.A(new_n1376), .B(new_n1375), .Y(new_n1377));
  MAJIxp5_ASAP7_75t_L       g01121(.A(new_n1319), .B(new_n1374), .C(new_n1377), .Y(new_n1378));
  AOI32xp33_ASAP7_75t_L     g01122(.A1(new_n424), .A2(new_n426), .A3(new_n823), .B1(new_n826), .B2(\b[7] ), .Y(new_n1379));
  OAI221xp5_ASAP7_75t_L     g01123(.A1(new_n994), .A2(new_n382), .B1(new_n353), .B2(new_n909), .C(new_n1379), .Y(new_n1380));
  NOR2xp33_ASAP7_75t_L      g01124(.A(new_n813), .B(new_n1380), .Y(new_n1381));
  NAND2xp33_ASAP7_75t_L     g01125(.A(new_n813), .B(new_n1380), .Y(new_n1382));
  INVx1_ASAP7_75t_L         g01126(.A(new_n1382), .Y(new_n1383));
  AOI22xp33_ASAP7_75t_L     g01127(.A1(new_n1301), .A2(new_n1304), .B1(new_n1308), .B2(new_n1307), .Y(new_n1384));
  NOR3xp33_ASAP7_75t_L      g01128(.A(new_n1295), .B(new_n1196), .C(new_n1200), .Y(new_n1385));
  NAND2xp33_ASAP7_75t_L     g01129(.A(new_n1292), .B(new_n1385), .Y(new_n1386));
  INVx1_ASAP7_75t_L         g01130(.A(new_n1386), .Y(new_n1387));
  NAND2xp33_ASAP7_75t_L     g01131(.A(\b[2] ), .B(new_n1194), .Y(new_n1388));
  INVx1_ASAP7_75t_L         g01132(.A(new_n1388), .Y(new_n1389));
  NOR2xp33_ASAP7_75t_L      g01133(.A(new_n299), .B(new_n1298), .Y(new_n1390));
  OAI32xp33_ASAP7_75t_L     g01134(.A1(new_n325), .A2(new_n327), .A3(new_n1197), .B1(new_n323), .B2(new_n1198), .Y(new_n1391));
  NOR4xp25_ASAP7_75t_L      g01135(.A(new_n1389), .B(new_n1391), .C(new_n1107), .D(new_n1390), .Y(new_n1392));
  NOR2xp33_ASAP7_75t_L      g01136(.A(new_n1390), .B(new_n1391), .Y(new_n1393));
  O2A1O1Ixp33_ASAP7_75t_L   g01137(.A1(new_n278), .A2(new_n1195), .B(new_n1393), .C(\a[17] ), .Y(new_n1394));
  NAND2xp33_ASAP7_75t_L     g01138(.A(\a[20] ), .B(new_n1292), .Y(new_n1395));
  XNOR2x2_ASAP7_75t_L       g01139(.A(\a[19] ), .B(\a[18] ), .Y(new_n1396));
  INVx1_ASAP7_75t_L         g01140(.A(new_n1396), .Y(new_n1397));
  NAND2xp33_ASAP7_75t_L     g01141(.A(new_n1397), .B(new_n1291), .Y(new_n1398));
  INVx1_ASAP7_75t_L         g01142(.A(\a[19] ), .Y(new_n1399));
  NAND2xp33_ASAP7_75t_L     g01143(.A(\a[20] ), .B(new_n1399), .Y(new_n1400));
  INVx1_ASAP7_75t_L         g01144(.A(\a[20] ), .Y(new_n1401));
  NAND2xp33_ASAP7_75t_L     g01145(.A(\a[19] ), .B(new_n1401), .Y(new_n1402));
  AND2x2_ASAP7_75t_L        g01146(.A(new_n1400), .B(new_n1402), .Y(new_n1403));
  NOR2xp33_ASAP7_75t_L      g01147(.A(new_n1291), .B(new_n1403), .Y(new_n1404));
  NAND2xp33_ASAP7_75t_L     g01148(.A(new_n1402), .B(new_n1400), .Y(new_n1405));
  NOR2xp33_ASAP7_75t_L      g01149(.A(new_n1405), .B(new_n1291), .Y(new_n1406));
  AOI22xp33_ASAP7_75t_L     g01150(.A1(new_n1406), .A2(\b[1] ), .B1(new_n271), .B2(new_n1404), .Y(new_n1407));
  O2A1O1Ixp33_ASAP7_75t_L   g01151(.A1(new_n1398), .A2(new_n258), .B(new_n1407), .C(new_n1395), .Y(new_n1408));
  NAND2xp33_ASAP7_75t_L     g01152(.A(new_n1290), .B(new_n1289), .Y(new_n1409));
  NOR2xp33_ASAP7_75t_L      g01153(.A(new_n1396), .B(new_n1409), .Y(new_n1410));
  NAND2xp33_ASAP7_75t_L     g01154(.A(new_n1405), .B(new_n1409), .Y(new_n1411));
  NAND2xp33_ASAP7_75t_L     g01155(.A(new_n1409), .B(new_n1403), .Y(new_n1412));
  OAI22xp33_ASAP7_75t_L     g01156(.A1(new_n1412), .A2(new_n276), .B1(new_n270), .B2(new_n1411), .Y(new_n1413));
  A2O1A1O1Ixp25_ASAP7_75t_L g01157(.A1(new_n1409), .A2(\a[20] ), .B(new_n1410), .C(\b[0] ), .D(new_n1413), .Y(new_n1414));
  OR2x4_ASAP7_75t_L         g01158(.A(new_n1414), .B(new_n1408), .Y(new_n1415));
  NOR3xp33_ASAP7_75t_L      g01159(.A(new_n1415), .B(new_n1394), .C(new_n1392), .Y(new_n1416));
  INVx1_ASAP7_75t_L         g01160(.A(new_n1392), .Y(new_n1417));
  OAI31xp33_ASAP7_75t_L     g01161(.A1(new_n1389), .A2(new_n1391), .A3(new_n1390), .B(new_n1107), .Y(new_n1418));
  NOR2xp33_ASAP7_75t_L      g01162(.A(new_n1414), .B(new_n1408), .Y(new_n1419));
  AOI21xp33_ASAP7_75t_L     g01163(.A1(new_n1417), .A2(new_n1418), .B(new_n1419), .Y(new_n1420));
  OAI22xp33_ASAP7_75t_L     g01164(.A1(new_n1384), .A2(new_n1387), .B1(new_n1420), .B2(new_n1416), .Y(new_n1421));
  MAJIxp5_ASAP7_75t_L       g01165(.A(new_n1305), .B(new_n1292), .C(new_n1385), .Y(new_n1422));
  NOR2xp33_ASAP7_75t_L      g01166(.A(new_n1420), .B(new_n1416), .Y(new_n1423));
  NAND2xp33_ASAP7_75t_L     g01167(.A(new_n1422), .B(new_n1423), .Y(new_n1424));
  OAI211xp5_ASAP7_75t_L     g01168(.A1(new_n1381), .A2(new_n1383), .B(new_n1424), .C(new_n1421), .Y(new_n1425));
  INVx1_ASAP7_75t_L         g01169(.A(new_n1381), .Y(new_n1426));
  INVx1_ASAP7_75t_L         g01170(.A(new_n1385), .Y(new_n1427));
  O2A1O1Ixp33_ASAP7_75t_L   g01171(.A1(new_n1293), .A2(new_n1427), .B(new_n1306), .C(new_n1423), .Y(new_n1428));
  AND2x2_ASAP7_75t_L        g01172(.A(new_n1304), .B(new_n1301), .Y(new_n1429));
  A2O1A1Ixp33_ASAP7_75t_L   g01173(.A1(new_n1308), .A2(new_n1307), .B(new_n1429), .C(new_n1386), .Y(new_n1430));
  NAND3xp33_ASAP7_75t_L     g01174(.A(new_n1417), .B(new_n1419), .C(new_n1418), .Y(new_n1431));
  OAI21xp33_ASAP7_75t_L     g01175(.A1(new_n1392), .A2(new_n1394), .B(new_n1415), .Y(new_n1432));
  NAND2xp33_ASAP7_75t_L     g01176(.A(new_n1431), .B(new_n1432), .Y(new_n1433));
  NOR2xp33_ASAP7_75t_L      g01177(.A(new_n1433), .B(new_n1430), .Y(new_n1434));
  OAI211xp5_ASAP7_75t_L     g01178(.A1(new_n1434), .A2(new_n1428), .B(new_n1382), .C(new_n1426), .Y(new_n1435));
  NAND3xp33_ASAP7_75t_L     g01179(.A(new_n1435), .B(new_n1378), .C(new_n1425), .Y(new_n1436));
  OAI211xp5_ASAP7_75t_L     g01180(.A1(new_n1376), .A2(new_n1375), .B(new_n1309), .C(new_n1306), .Y(new_n1437));
  O2A1O1Ixp33_ASAP7_75t_L   g01181(.A1(new_n1125), .A2(new_n1126), .B(new_n1120), .C(new_n1205), .Y(new_n1438));
  OAI22xp33_ASAP7_75t_L     g01182(.A1(new_n1438), .A2(new_n1214), .B1(new_n1316), .B2(new_n1317), .Y(new_n1439));
  AOI211xp5_ASAP7_75t_L     g01183(.A1(new_n1382), .A2(new_n1426), .B(new_n1434), .C(new_n1428), .Y(new_n1440));
  AOI211xp5_ASAP7_75t_L     g01184(.A1(new_n1424), .A2(new_n1421), .B(new_n1381), .C(new_n1383), .Y(new_n1441));
  OAI211xp5_ASAP7_75t_L     g01185(.A1(new_n1441), .A2(new_n1440), .B(new_n1439), .C(new_n1437), .Y(new_n1442));
  NAND2xp33_ASAP7_75t_L     g01186(.A(\b[9] ), .B(new_n590), .Y(new_n1443));
  NAND2xp33_ASAP7_75t_L     g01187(.A(\b[10] ), .B(new_n600), .Y(new_n1444));
  OAI311xp33_ASAP7_75t_L    g01188(.A1(new_n639), .A2(new_n851), .A3(new_n675), .B1(new_n1444), .C1(new_n1443), .Y(new_n1445));
  AOI21xp33_ASAP7_75t_L     g01189(.A1(new_n674), .A2(\b[8] ), .B(new_n1445), .Y(new_n1446));
  NAND2xp33_ASAP7_75t_L     g01190(.A(\a[11] ), .B(new_n1446), .Y(new_n1447));
  A2O1A1Ixp33_ASAP7_75t_L   g01191(.A1(\b[8] ), .A2(new_n674), .B(new_n1445), .C(new_n594), .Y(new_n1448));
  NAND2xp33_ASAP7_75t_L     g01192(.A(new_n1448), .B(new_n1447), .Y(new_n1449));
  INVx1_ASAP7_75t_L         g01193(.A(new_n1449), .Y(new_n1450));
  NAND3xp33_ASAP7_75t_L     g01194(.A(new_n1450), .B(new_n1442), .C(new_n1436), .Y(new_n1451));
  AO22x1_ASAP7_75t_L        g01195(.A1(new_n1448), .A2(new_n1447), .B1(new_n1436), .B2(new_n1442), .Y(new_n1452));
  NAND4xp25_ASAP7_75t_L     g01196(.A(new_n1320), .B(new_n1326), .C(new_n1327), .D(new_n1321), .Y(new_n1453));
  A2O1A1O1Ixp25_ASAP7_75t_L g01197(.A1(new_n1219), .A2(new_n1181), .B(new_n1228), .C(new_n1453), .D(new_n1328), .Y(new_n1454));
  NAND3xp33_ASAP7_75t_L     g01198(.A(new_n1451), .B(new_n1454), .C(new_n1452), .Y(new_n1455));
  AOI21xp33_ASAP7_75t_L     g01199(.A1(new_n1451), .A2(new_n1452), .B(new_n1454), .Y(new_n1456));
  INVx1_ASAP7_75t_L         g01200(.A(new_n1456), .Y(new_n1457));
  NAND2xp33_ASAP7_75t_L     g01201(.A(\b[12] ), .B(new_n441), .Y(new_n1458));
  AOI22xp33_ASAP7_75t_L     g01202(.A1(new_n451), .A2(\b[13] ), .B1(new_n448), .B2(new_n800), .Y(new_n1459));
  AND2x2_ASAP7_75t_L        g01203(.A(new_n1458), .B(new_n1459), .Y(new_n1460));
  OAI211xp5_ASAP7_75t_L     g01204(.A1(new_n695), .A2(new_n481), .B(new_n1460), .C(\a[8] ), .Y(new_n1461));
  NAND2xp33_ASAP7_75t_L     g01205(.A(new_n1458), .B(new_n1459), .Y(new_n1462));
  A2O1A1Ixp33_ASAP7_75t_L   g01206(.A1(\b[11] ), .A2(new_n480), .B(new_n1462), .C(new_n445), .Y(new_n1463));
  NAND2xp33_ASAP7_75t_L     g01207(.A(new_n1463), .B(new_n1461), .Y(new_n1464));
  AOI21xp33_ASAP7_75t_L     g01208(.A1(new_n1455), .A2(new_n1457), .B(new_n1464), .Y(new_n1465));
  INVx1_ASAP7_75t_L         g01209(.A(new_n1455), .Y(new_n1466));
  AOI211xp5_ASAP7_75t_L     g01210(.A1(\b[11] ), .A2(new_n480), .B(new_n445), .C(new_n1462), .Y(new_n1467));
  O2A1O1Ixp33_ASAP7_75t_L   g01211(.A1(new_n695), .A2(new_n481), .B(new_n1460), .C(\a[8] ), .Y(new_n1468));
  NOR2xp33_ASAP7_75t_L      g01212(.A(new_n1467), .B(new_n1468), .Y(new_n1469));
  NOR3xp33_ASAP7_75t_L      g01213(.A(new_n1469), .B(new_n1456), .C(new_n1466), .Y(new_n1470));
  NOR2xp33_ASAP7_75t_L      g01214(.A(new_n1465), .B(new_n1470), .Y(new_n1471));
  A2O1A1Ixp33_ASAP7_75t_L   g01215(.A1(new_n1373), .A2(new_n1341), .B(new_n1339), .C(new_n1471), .Y(new_n1472));
  OAI21xp33_ASAP7_75t_L     g01216(.A1(new_n1466), .A2(new_n1456), .B(new_n1469), .Y(new_n1473));
  NAND3xp33_ASAP7_75t_L     g01217(.A(new_n1464), .B(new_n1457), .C(new_n1455), .Y(new_n1474));
  NAND2xp33_ASAP7_75t_L     g01218(.A(new_n1473), .B(new_n1474), .Y(new_n1475));
  A2O1A1O1Ixp25_ASAP7_75t_L g01219(.A1(new_n1232), .A2(new_n1171), .B(new_n1231), .C(new_n1373), .D(new_n1339), .Y(new_n1476));
  NAND2xp33_ASAP7_75t_L     g01220(.A(new_n1476), .B(new_n1475), .Y(new_n1477));
  AOI22xp33_ASAP7_75t_L     g01221(.A1(new_n345), .A2(\b[16] ), .B1(new_n342), .B2(new_n1058), .Y(new_n1478));
  OAI221xp5_ASAP7_75t_L     g01222(.A1(new_n406), .A2(new_n952), .B1(new_n871), .B2(new_n365), .C(new_n1478), .Y(new_n1479));
  XNOR2x2_ASAP7_75t_L       g01223(.A(\a[5] ), .B(new_n1479), .Y(new_n1480));
  NAND3xp33_ASAP7_75t_L     g01224(.A(new_n1472), .B(new_n1477), .C(new_n1480), .Y(new_n1481));
  INVx1_ASAP7_75t_L         g01225(.A(new_n1339), .Y(new_n1482));
  O2A1O1Ixp33_ASAP7_75t_L   g01226(.A1(new_n1279), .A2(new_n1335), .B(new_n1482), .C(new_n1475), .Y(new_n1483));
  INVx1_ASAP7_75t_L         g01227(.A(new_n1476), .Y(new_n1484));
  NOR2xp33_ASAP7_75t_L      g01228(.A(new_n1484), .B(new_n1471), .Y(new_n1485));
  INVx1_ASAP7_75t_L         g01229(.A(new_n1480), .Y(new_n1486));
  OAI21xp33_ASAP7_75t_L     g01230(.A1(new_n1483), .A2(new_n1485), .B(new_n1486), .Y(new_n1487));
  A2O1A1O1Ixp25_ASAP7_75t_L g01231(.A1(new_n1348), .A2(new_n1260), .B(new_n1236), .C(new_n1346), .D(new_n1344), .Y(new_n1488));
  NAND3xp33_ASAP7_75t_L     g01232(.A(new_n1488), .B(new_n1487), .C(new_n1481), .Y(new_n1489));
  NAND2xp33_ASAP7_75t_L     g01233(.A(new_n1487), .B(new_n1481), .Y(new_n1490));
  A2O1A1Ixp33_ASAP7_75t_L   g01234(.A1(new_n1346), .A2(new_n1271), .B(new_n1344), .C(new_n1490), .Y(new_n1491));
  NOR2xp33_ASAP7_75t_L      g01235(.A(\b[18] ), .B(\b[19] ), .Y(new_n1492));
  INVx1_ASAP7_75t_L         g01236(.A(\b[19] ), .Y(new_n1493));
  NOR2xp33_ASAP7_75t_L      g01237(.A(new_n1356), .B(new_n1493), .Y(new_n1494));
  NOR2xp33_ASAP7_75t_L      g01238(.A(new_n1492), .B(new_n1494), .Y(new_n1495));
  A2O1A1Ixp33_ASAP7_75t_L   g01239(.A1(new_n1361), .A2(new_n1358), .B(new_n1357), .C(new_n1495), .Y(new_n1496));
  INVx1_ASAP7_75t_L         g01240(.A(new_n1496), .Y(new_n1497));
  NOR3xp33_ASAP7_75t_L      g01241(.A(new_n1360), .B(new_n1495), .C(new_n1357), .Y(new_n1498));
  NOR2xp33_ASAP7_75t_L      g01242(.A(new_n1498), .B(new_n1497), .Y(new_n1499));
  AOI22xp33_ASAP7_75t_L     g01243(.A1(new_n272), .A2(\b[19] ), .B1(new_n269), .B2(new_n1499), .Y(new_n1500));
  OAI221xp5_ASAP7_75t_L     g01244(.A1(new_n261), .A2(new_n1356), .B1(new_n1244), .B2(new_n277), .C(new_n1500), .Y(new_n1501));
  XNOR2x2_ASAP7_75t_L       g01245(.A(\a[2] ), .B(new_n1501), .Y(new_n1502));
  NAND3xp33_ASAP7_75t_L     g01246(.A(new_n1491), .B(new_n1489), .C(new_n1502), .Y(new_n1503));
  AO21x2_ASAP7_75t_L        g01247(.A1(new_n1489), .A2(new_n1491), .B(new_n1502), .Y(new_n1504));
  NAND2xp33_ASAP7_75t_L     g01248(.A(new_n1503), .B(new_n1504), .Y(new_n1505));
  INVx1_ASAP7_75t_L         g01249(.A(new_n1505), .Y(new_n1506));
  INVx1_ASAP7_75t_L         g01250(.A(new_n1347), .Y(new_n1507));
  INVx1_ASAP7_75t_L         g01251(.A(new_n1351), .Y(new_n1508));
  OR3x1_ASAP7_75t_L         g01252(.A(new_n1508), .B(new_n1507), .C(new_n1366), .Y(new_n1509));
  O2A1O1Ixp33_ASAP7_75t_L   g01253(.A1(new_n1371), .A2(new_n1369), .B(new_n1509), .C(new_n1506), .Y(new_n1510));
  NAND3xp33_ASAP7_75t_L     g01254(.A(new_n1238), .B(new_n1240), .C(new_n1262), .Y(new_n1511));
  A2O1A1Ixp33_ASAP7_75t_L   g01255(.A1(new_n1511), .A2(new_n1267), .B(new_n1369), .C(new_n1509), .Y(new_n1512));
  NOR2xp33_ASAP7_75t_L      g01256(.A(new_n1505), .B(new_n1512), .Y(new_n1513));
  NOR2xp33_ASAP7_75t_L      g01257(.A(new_n1513), .B(new_n1510), .Y(\f[19] ));
  NAND2xp33_ASAP7_75t_L     g01258(.A(new_n1489), .B(new_n1491), .Y(new_n1515));
  INVx1_ASAP7_75t_L         g01259(.A(new_n1510), .Y(new_n1516));
  NAND3xp33_ASAP7_75t_L     g01260(.A(new_n1472), .B(new_n1477), .C(new_n1486), .Y(new_n1517));
  A2O1A1Ixp33_ASAP7_75t_L   g01261(.A1(new_n1487), .A2(new_n1481), .B(new_n1488), .C(new_n1517), .Y(new_n1518));
  NAND2xp33_ASAP7_75t_L     g01262(.A(\b[16] ), .B(new_n334), .Y(new_n1519));
  OAI221xp5_ASAP7_75t_L     g01263(.A1(new_n368), .A2(new_n1244), .B1(new_n367), .B2(new_n1251), .C(new_n1519), .Y(new_n1520));
  AOI21xp33_ASAP7_75t_L     g01264(.A1(new_n366), .A2(\b[15] ), .B(new_n1520), .Y(new_n1521));
  NAND2xp33_ASAP7_75t_L     g01265(.A(\a[5] ), .B(new_n1521), .Y(new_n1522));
  A2O1A1Ixp33_ASAP7_75t_L   g01266(.A1(\b[15] ), .A2(new_n366), .B(new_n1520), .C(new_n339), .Y(new_n1523));
  NAND2xp33_ASAP7_75t_L     g01267(.A(new_n1523), .B(new_n1522), .Y(new_n1524));
  NAND2xp33_ASAP7_75t_L     g01268(.A(new_n1436), .B(new_n1442), .Y(new_n1525));
  MAJIxp5_ASAP7_75t_L       g01269(.A(new_n1454), .B(new_n1450), .C(new_n1525), .Y(new_n1526));
  NAND2xp33_ASAP7_75t_L     g01270(.A(\b[9] ), .B(new_n674), .Y(new_n1527));
  NAND2xp33_ASAP7_75t_L     g01271(.A(\b[10] ), .B(new_n590), .Y(new_n1528));
  AOI32xp33_ASAP7_75t_L     g01272(.A1(new_n700), .A2(new_n698), .A3(new_n597), .B1(new_n600), .B2(\b[11] ), .Y(new_n1529));
  NAND4xp25_ASAP7_75t_L     g01273(.A(new_n1529), .B(\a[11] ), .C(new_n1527), .D(new_n1528), .Y(new_n1530));
  NAND2xp33_ASAP7_75t_L     g01274(.A(new_n1528), .B(new_n1529), .Y(new_n1531));
  A2O1A1Ixp33_ASAP7_75t_L   g01275(.A1(\b[9] ), .A2(new_n674), .B(new_n1531), .C(new_n594), .Y(new_n1532));
  NAND2xp33_ASAP7_75t_L     g01276(.A(new_n1530), .B(new_n1532), .Y(new_n1533));
  A2O1A1Ixp33_ASAP7_75t_L   g01277(.A1(new_n1439), .A2(new_n1437), .B(new_n1441), .C(new_n1425), .Y(new_n1534));
  NOR2xp33_ASAP7_75t_L      g01278(.A(new_n382), .B(new_n909), .Y(new_n1535));
  NAND2xp33_ASAP7_75t_L     g01279(.A(\b[7] ), .B(new_n817), .Y(new_n1536));
  OAI221xp5_ASAP7_75t_L     g01280(.A1(new_n912), .A2(new_n503), .B1(new_n911), .B2(new_n509), .C(new_n1536), .Y(new_n1537));
  OR3x1_ASAP7_75t_L         g01281(.A(new_n1537), .B(new_n813), .C(new_n1535), .Y(new_n1538));
  A2O1A1Ixp33_ASAP7_75t_L   g01282(.A1(\b[6] ), .A2(new_n908), .B(new_n1537), .C(new_n813), .Y(new_n1539));
  OAI21xp33_ASAP7_75t_L     g01283(.A1(new_n1392), .A2(new_n1394), .B(new_n1419), .Y(new_n1540));
  NAND2xp33_ASAP7_75t_L     g01284(.A(\b[3] ), .B(new_n1194), .Y(new_n1541));
  NAND2xp33_ASAP7_75t_L     g01285(.A(\b[4] ), .B(new_n1103), .Y(new_n1542));
  AOI32xp33_ASAP7_75t_L     g01286(.A1(new_n358), .A2(new_n356), .A3(new_n1110), .B1(\b[5] ), .B2(new_n1113), .Y(new_n1543));
  NAND3xp33_ASAP7_75t_L     g01287(.A(new_n1543), .B(new_n1542), .C(new_n1541), .Y(new_n1544));
  NOR2xp33_ASAP7_75t_L      g01288(.A(new_n1107), .B(new_n1544), .Y(new_n1545));
  AOI31xp33_ASAP7_75t_L     g01289(.A1(new_n1543), .A2(new_n1542), .A3(new_n1541), .B(\a[17] ), .Y(new_n1546));
  A2O1A1O1Ixp25_ASAP7_75t_L g01290(.A1(new_n1396), .A2(new_n1291), .B(new_n258), .C(new_n1407), .D(new_n1401), .Y(new_n1547));
  NOR3xp33_ASAP7_75t_L      g01291(.A(new_n1403), .B(new_n1397), .C(new_n1409), .Y(new_n1548));
  INVx1_ASAP7_75t_L         g01292(.A(new_n1548), .Y(new_n1549));
  NOR2xp33_ASAP7_75t_L      g01293(.A(new_n258), .B(new_n1549), .Y(new_n1550));
  NAND2xp33_ASAP7_75t_L     g01294(.A(\b[1] ), .B(new_n1410), .Y(new_n1551));
  OAI221xp5_ASAP7_75t_L     g01295(.A1(new_n1411), .A2(new_n283), .B1(new_n278), .B2(new_n1412), .C(new_n1551), .Y(new_n1552));
  OR3x1_ASAP7_75t_L         g01296(.A(new_n1547), .B(new_n1550), .C(new_n1552), .Y(new_n1553));
  A2O1A1Ixp33_ASAP7_75t_L   g01297(.A1(\b[0] ), .A2(new_n1548), .B(new_n1552), .C(new_n1547), .Y(new_n1554));
  AOI211xp5_ASAP7_75t_L     g01298(.A1(new_n1553), .A2(new_n1554), .B(new_n1546), .C(new_n1545), .Y(new_n1555));
  INVx1_ASAP7_75t_L         g01299(.A(new_n1555), .Y(new_n1556));
  OAI211xp5_ASAP7_75t_L     g01300(.A1(new_n1546), .A2(new_n1545), .B(new_n1553), .C(new_n1554), .Y(new_n1557));
  NAND4xp25_ASAP7_75t_L     g01301(.A(new_n1421), .B(new_n1557), .C(new_n1556), .D(new_n1540), .Y(new_n1558));
  A2O1A1Ixp33_ASAP7_75t_L   g01302(.A1(new_n1431), .A2(new_n1432), .B(new_n1422), .C(new_n1540), .Y(new_n1559));
  INVx1_ASAP7_75t_L         g01303(.A(new_n1557), .Y(new_n1560));
  OAI21xp33_ASAP7_75t_L     g01304(.A1(new_n1555), .A2(new_n1560), .B(new_n1559), .Y(new_n1561));
  NAND4xp25_ASAP7_75t_L     g01305(.A(new_n1558), .B(new_n1561), .C(new_n1538), .D(new_n1539), .Y(new_n1562));
  AOI22xp33_ASAP7_75t_L     g01306(.A1(new_n1539), .A2(new_n1538), .B1(new_n1561), .B2(new_n1558), .Y(new_n1563));
  INVx1_ASAP7_75t_L         g01307(.A(new_n1563), .Y(new_n1564));
  NAND3xp33_ASAP7_75t_L     g01308(.A(new_n1534), .B(new_n1564), .C(new_n1562), .Y(new_n1565));
  AO21x2_ASAP7_75t_L        g01309(.A1(new_n1564), .A2(new_n1562), .B(new_n1534), .Y(new_n1566));
  AO21x2_ASAP7_75t_L        g01310(.A1(new_n1565), .A2(new_n1566), .B(new_n1533), .Y(new_n1567));
  NAND3xp33_ASAP7_75t_L     g01311(.A(new_n1566), .B(new_n1565), .C(new_n1533), .Y(new_n1568));
  NAND3xp33_ASAP7_75t_L     g01312(.A(new_n1526), .B(new_n1567), .C(new_n1568), .Y(new_n1569));
  AO21x2_ASAP7_75t_L        g01313(.A1(new_n1568), .A2(new_n1567), .B(new_n1526), .Y(new_n1570));
  NOR2xp33_ASAP7_75t_L      g01314(.A(new_n763), .B(new_n481), .Y(new_n1571));
  NAND2xp33_ASAP7_75t_L     g01315(.A(\b[13] ), .B(new_n441), .Y(new_n1572));
  OAI221xp5_ASAP7_75t_L     g01316(.A1(new_n667), .A2(new_n871), .B1(new_n482), .B2(new_n878), .C(new_n1572), .Y(new_n1573));
  OR3x1_ASAP7_75t_L         g01317(.A(new_n1573), .B(new_n445), .C(new_n1571), .Y(new_n1574));
  A2O1A1Ixp33_ASAP7_75t_L   g01318(.A1(\b[12] ), .A2(new_n480), .B(new_n1573), .C(new_n445), .Y(new_n1575));
  NAND4xp25_ASAP7_75t_L     g01319(.A(new_n1570), .B(new_n1569), .C(new_n1574), .D(new_n1575), .Y(new_n1576));
  AND3x1_ASAP7_75t_L        g01320(.A(new_n1526), .B(new_n1568), .C(new_n1567), .Y(new_n1577));
  AOI21xp33_ASAP7_75t_L     g01321(.A1(new_n1568), .A2(new_n1567), .B(new_n1526), .Y(new_n1578));
  NAND2xp33_ASAP7_75t_L     g01322(.A(new_n1575), .B(new_n1574), .Y(new_n1579));
  OAI21xp33_ASAP7_75t_L     g01323(.A1(new_n1578), .A2(new_n1577), .B(new_n1579), .Y(new_n1580));
  AND2x2_ASAP7_75t_L        g01324(.A(new_n1576), .B(new_n1580), .Y(new_n1581));
  O2A1O1Ixp33_ASAP7_75t_L   g01325(.A1(new_n1465), .A2(new_n1476), .B(new_n1474), .C(new_n1581), .Y(new_n1582));
  NAND2xp33_ASAP7_75t_L     g01326(.A(new_n1576), .B(new_n1580), .Y(new_n1583));
  OAI21xp33_ASAP7_75t_L     g01327(.A1(new_n1465), .A2(new_n1476), .B(new_n1474), .Y(new_n1584));
  NOR2xp33_ASAP7_75t_L      g01328(.A(new_n1583), .B(new_n1584), .Y(new_n1585));
  OAI21xp33_ASAP7_75t_L     g01329(.A1(new_n1585), .A2(new_n1582), .B(new_n1524), .Y(new_n1586));
  A2O1A1Ixp33_ASAP7_75t_L   g01330(.A1(new_n1484), .A2(new_n1473), .B(new_n1470), .C(new_n1583), .Y(new_n1587));
  A2O1A1O1Ixp25_ASAP7_75t_L g01331(.A1(new_n1373), .A2(new_n1341), .B(new_n1339), .C(new_n1473), .D(new_n1470), .Y(new_n1588));
  NAND2xp33_ASAP7_75t_L     g01332(.A(new_n1588), .B(new_n1581), .Y(new_n1589));
  NAND4xp25_ASAP7_75t_L     g01333(.A(new_n1589), .B(new_n1587), .C(new_n1522), .D(new_n1523), .Y(new_n1590));
  NAND2xp33_ASAP7_75t_L     g01334(.A(new_n1590), .B(new_n1586), .Y(new_n1591));
  XNOR2x2_ASAP7_75t_L       g01335(.A(new_n1591), .B(new_n1518), .Y(new_n1592));
  NOR2xp33_ASAP7_75t_L      g01336(.A(\b[19] ), .B(\b[20] ), .Y(new_n1593));
  INVx1_ASAP7_75t_L         g01337(.A(\b[20] ), .Y(new_n1594));
  NOR2xp33_ASAP7_75t_L      g01338(.A(new_n1493), .B(new_n1594), .Y(new_n1595));
  NOR2xp33_ASAP7_75t_L      g01339(.A(new_n1593), .B(new_n1595), .Y(new_n1596));
  INVx1_ASAP7_75t_L         g01340(.A(new_n1596), .Y(new_n1597));
  O2A1O1Ixp33_ASAP7_75t_L   g01341(.A1(new_n1356), .A2(new_n1493), .B(new_n1496), .C(new_n1597), .Y(new_n1598));
  NOR3xp33_ASAP7_75t_L      g01342(.A(new_n1497), .B(new_n1596), .C(new_n1494), .Y(new_n1599));
  NOR2xp33_ASAP7_75t_L      g01343(.A(new_n1598), .B(new_n1599), .Y(new_n1600));
  AOI22xp33_ASAP7_75t_L     g01344(.A1(new_n272), .A2(\b[20] ), .B1(new_n269), .B2(new_n1600), .Y(new_n1601));
  OAI221xp5_ASAP7_75t_L     g01345(.A1(new_n261), .A2(new_n1493), .B1(new_n1356), .B2(new_n277), .C(new_n1601), .Y(new_n1602));
  XNOR2x2_ASAP7_75t_L       g01346(.A(\a[2] ), .B(new_n1602), .Y(new_n1603));
  NOR2xp33_ASAP7_75t_L      g01347(.A(new_n1603), .B(new_n1592), .Y(new_n1604));
  INVx1_ASAP7_75t_L         g01348(.A(new_n1604), .Y(new_n1605));
  NAND2xp33_ASAP7_75t_L     g01349(.A(new_n1603), .B(new_n1592), .Y(new_n1606));
  NAND2xp33_ASAP7_75t_L     g01350(.A(new_n1606), .B(new_n1605), .Y(new_n1607));
  O2A1O1Ixp33_ASAP7_75t_L   g01351(.A1(new_n1515), .A2(new_n1502), .B(new_n1516), .C(new_n1607), .Y(new_n1608));
  NOR2xp33_ASAP7_75t_L      g01352(.A(new_n1502), .B(new_n1515), .Y(new_n1609));
  AOI211xp5_ASAP7_75t_L     g01353(.A1(new_n1605), .A2(new_n1606), .B(new_n1609), .C(new_n1510), .Y(new_n1610));
  NOR2xp33_ASAP7_75t_L      g01354(.A(new_n1610), .B(new_n1608), .Y(\f[20] ));
  NAND3xp33_ASAP7_75t_L     g01355(.A(new_n1570), .B(new_n1579), .C(new_n1569), .Y(new_n1612));
  NAND2xp33_ASAP7_75t_L     g01356(.A(\b[13] ), .B(new_n480), .Y(new_n1613));
  NAND2xp33_ASAP7_75t_L     g01357(.A(\b[14] ), .B(new_n441), .Y(new_n1614));
  AOI22xp33_ASAP7_75t_L     g01358(.A1(new_n451), .A2(\b[15] ), .B1(new_n448), .B2(new_n959), .Y(new_n1615));
  AND4x1_ASAP7_75t_L        g01359(.A(new_n1615), .B(new_n1614), .C(new_n1613), .D(\a[8] ), .Y(new_n1616));
  AOI31xp33_ASAP7_75t_L     g01360(.A1(new_n1615), .A2(new_n1614), .A3(new_n1613), .B(\a[8] ), .Y(new_n1617));
  OR2x4_ASAP7_75t_L         g01361(.A(new_n1617), .B(new_n1616), .Y(new_n1618));
  AND3x1_ASAP7_75t_L        g01362(.A(new_n1566), .B(new_n1565), .C(new_n1533), .Y(new_n1619));
  INVx1_ASAP7_75t_L         g01363(.A(new_n674), .Y(new_n1620));
  NOR2xp33_ASAP7_75t_L      g01364(.A(new_n631), .B(new_n1620), .Y(new_n1621));
  NAND2xp33_ASAP7_75t_L     g01365(.A(\b[11] ), .B(new_n590), .Y(new_n1622));
  OAI221xp5_ASAP7_75t_L     g01366(.A1(new_n676), .A2(new_n763), .B1(new_n675), .B2(new_n775), .C(new_n1622), .Y(new_n1623));
  OR3x1_ASAP7_75t_L         g01367(.A(new_n1623), .B(new_n594), .C(new_n1621), .Y(new_n1624));
  A2O1A1Ixp33_ASAP7_75t_L   g01368(.A1(\b[10] ), .A2(new_n674), .B(new_n1623), .C(new_n594), .Y(new_n1625));
  A2O1A1O1Ixp25_ASAP7_75t_L g01369(.A1(new_n1378), .A2(new_n1435), .B(new_n1440), .C(new_n1562), .D(new_n1563), .Y(new_n1626));
  NAND2xp33_ASAP7_75t_L     g01370(.A(\b[0] ), .B(new_n1410), .Y(new_n1627));
  NAND4xp25_ASAP7_75t_L     g01371(.A(new_n1407), .B(\a[20] ), .C(new_n1293), .D(new_n1627), .Y(new_n1628));
  INVx1_ASAP7_75t_L         g01372(.A(\a[21] ), .Y(new_n1629));
  NAND2xp33_ASAP7_75t_L     g01373(.A(\a[20] ), .B(new_n1629), .Y(new_n1630));
  NAND2xp33_ASAP7_75t_L     g01374(.A(\a[21] ), .B(new_n1401), .Y(new_n1631));
  AND2x2_ASAP7_75t_L        g01375(.A(new_n1630), .B(new_n1631), .Y(new_n1632));
  NOR2xp33_ASAP7_75t_L      g01376(.A(new_n258), .B(new_n1632), .Y(new_n1633));
  OAI31xp33_ASAP7_75t_L     g01377(.A1(new_n1628), .A2(new_n1552), .A3(new_n1550), .B(new_n1633), .Y(new_n1634));
  OR4x2_ASAP7_75t_L         g01378(.A(new_n1633), .B(new_n1628), .C(new_n1552), .D(new_n1550), .Y(new_n1635));
  NOR2xp33_ASAP7_75t_L      g01379(.A(new_n278), .B(new_n1398), .Y(new_n1636));
  AOI221xp5_ASAP7_75t_L     g01380(.A1(new_n1406), .A2(\b[3] ), .B1(new_n1404), .B2(new_n1000), .C(new_n1636), .Y(new_n1637));
  OAI211xp5_ASAP7_75t_L     g01381(.A1(new_n276), .A2(new_n1549), .B(new_n1637), .C(\a[20] ), .Y(new_n1638));
  NAND2xp33_ASAP7_75t_L     g01382(.A(\b[3] ), .B(new_n1406), .Y(new_n1639));
  OAI221xp5_ASAP7_75t_L     g01383(.A1(new_n278), .A2(new_n1398), .B1(new_n1411), .B2(new_n303), .C(new_n1639), .Y(new_n1640));
  A2O1A1Ixp33_ASAP7_75t_L   g01384(.A1(\b[1] ), .A2(new_n1548), .B(new_n1640), .C(new_n1401), .Y(new_n1641));
  AO22x1_ASAP7_75t_L        g01385(.A1(new_n1641), .A2(new_n1638), .B1(new_n1634), .B2(new_n1635), .Y(new_n1642));
  AOI211xp5_ASAP7_75t_L     g01386(.A1(\b[1] ), .A2(new_n1548), .B(new_n1401), .C(new_n1640), .Y(new_n1643));
  O2A1O1Ixp33_ASAP7_75t_L   g01387(.A1(new_n276), .A2(new_n1549), .B(new_n1637), .C(\a[20] ), .Y(new_n1644));
  NOR2xp33_ASAP7_75t_L      g01388(.A(new_n1643), .B(new_n1644), .Y(new_n1645));
  NAND3xp33_ASAP7_75t_L     g01389(.A(new_n1645), .B(new_n1635), .C(new_n1634), .Y(new_n1646));
  NAND2xp33_ASAP7_75t_L     g01390(.A(\b[4] ), .B(new_n1194), .Y(new_n1647));
  NAND2xp33_ASAP7_75t_L     g01391(.A(\b[5] ), .B(new_n1103), .Y(new_n1648));
  AOI22xp33_ASAP7_75t_L     g01392(.A1(new_n1113), .A2(\b[6] ), .B1(new_n1110), .B2(new_n389), .Y(new_n1649));
  NAND4xp25_ASAP7_75t_L     g01393(.A(new_n1649), .B(\a[17] ), .C(new_n1647), .D(new_n1648), .Y(new_n1650));
  OAI221xp5_ASAP7_75t_L     g01394(.A1(new_n1198), .A2(new_n382), .B1(new_n1197), .B2(new_n540), .C(new_n1648), .Y(new_n1651));
  A2O1A1Ixp33_ASAP7_75t_L   g01395(.A1(\b[4] ), .A2(new_n1194), .B(new_n1651), .C(new_n1107), .Y(new_n1652));
  NAND4xp25_ASAP7_75t_L     g01396(.A(new_n1646), .B(new_n1652), .C(new_n1642), .D(new_n1650), .Y(new_n1653));
  AO22x1_ASAP7_75t_L        g01397(.A1(new_n1642), .A2(new_n1646), .B1(new_n1652), .B2(new_n1650), .Y(new_n1654));
  A2O1A1O1Ixp25_ASAP7_75t_L g01398(.A1(new_n1431), .A2(new_n1432), .B(new_n1422), .C(new_n1540), .D(new_n1555), .Y(new_n1655));
  OAI211xp5_ASAP7_75t_L     g01399(.A1(new_n1560), .A2(new_n1655), .B(new_n1653), .C(new_n1654), .Y(new_n1656));
  AND4x1_ASAP7_75t_L        g01400(.A(new_n1642), .B(new_n1652), .C(new_n1646), .D(new_n1650), .Y(new_n1657));
  AOI22xp33_ASAP7_75t_L     g01401(.A1(new_n1646), .A2(new_n1642), .B1(new_n1652), .B2(new_n1650), .Y(new_n1658));
  INVx1_ASAP7_75t_L         g01402(.A(new_n1540), .Y(new_n1659));
  A2O1A1O1Ixp25_ASAP7_75t_L g01403(.A1(new_n1433), .A2(new_n1430), .B(new_n1659), .C(new_n1556), .D(new_n1560), .Y(new_n1660));
  OAI21xp33_ASAP7_75t_L     g01404(.A1(new_n1657), .A2(new_n1658), .B(new_n1660), .Y(new_n1661));
  NOR2xp33_ASAP7_75t_L      g01405(.A(new_n421), .B(new_n909), .Y(new_n1662));
  NAND2xp33_ASAP7_75t_L     g01406(.A(\b[8] ), .B(new_n817), .Y(new_n1663));
  OAI221xp5_ASAP7_75t_L     g01407(.A1(new_n912), .A2(new_n559), .B1(new_n911), .B2(new_n978), .C(new_n1663), .Y(new_n1664));
  OR3x1_ASAP7_75t_L         g01408(.A(new_n1664), .B(new_n813), .C(new_n1662), .Y(new_n1665));
  A2O1A1Ixp33_ASAP7_75t_L   g01409(.A1(\b[7] ), .A2(new_n908), .B(new_n1664), .C(new_n813), .Y(new_n1666));
  AOI22xp33_ASAP7_75t_L     g01410(.A1(new_n1661), .A2(new_n1656), .B1(new_n1666), .B2(new_n1665), .Y(new_n1667));
  AND4x1_ASAP7_75t_L        g01411(.A(new_n1661), .B(new_n1665), .C(new_n1656), .D(new_n1666), .Y(new_n1668));
  NOR3xp33_ASAP7_75t_L      g01412(.A(new_n1626), .B(new_n1668), .C(new_n1667), .Y(new_n1669));
  OA21x2_ASAP7_75t_L        g01413(.A1(new_n1667), .A2(new_n1668), .B(new_n1626), .Y(new_n1670));
  OA211x2_ASAP7_75t_L       g01414(.A1(new_n1669), .A2(new_n1670), .B(new_n1624), .C(new_n1625), .Y(new_n1671));
  AOI211xp5_ASAP7_75t_L     g01415(.A1(new_n1624), .A2(new_n1625), .B(new_n1669), .C(new_n1670), .Y(new_n1672));
  NOR2xp33_ASAP7_75t_L      g01416(.A(new_n1672), .B(new_n1671), .Y(new_n1673));
  A2O1A1Ixp33_ASAP7_75t_L   g01417(.A1(new_n1567), .A2(new_n1526), .B(new_n1619), .C(new_n1673), .Y(new_n1674));
  OAI211xp5_ASAP7_75t_L     g01418(.A1(new_n1671), .A2(new_n1672), .B(new_n1569), .C(new_n1568), .Y(new_n1675));
  NAND3xp33_ASAP7_75t_L     g01419(.A(new_n1674), .B(new_n1618), .C(new_n1675), .Y(new_n1676));
  NOR2xp33_ASAP7_75t_L      g01420(.A(new_n1617), .B(new_n1616), .Y(new_n1677));
  AOI211xp5_ASAP7_75t_L     g01421(.A1(new_n1569), .A2(new_n1568), .B(new_n1671), .C(new_n1672), .Y(new_n1678));
  AO21x2_ASAP7_75t_L        g01422(.A1(new_n1567), .A2(new_n1526), .B(new_n1619), .Y(new_n1679));
  NOR2xp33_ASAP7_75t_L      g01423(.A(new_n1679), .B(new_n1673), .Y(new_n1680));
  OAI21xp33_ASAP7_75t_L     g01424(.A1(new_n1678), .A2(new_n1680), .B(new_n1677), .Y(new_n1681));
  NAND2xp33_ASAP7_75t_L     g01425(.A(new_n1681), .B(new_n1676), .Y(new_n1682));
  O2A1O1Ixp33_ASAP7_75t_L   g01426(.A1(new_n1581), .A2(new_n1588), .B(new_n1612), .C(new_n1682), .Y(new_n1683));
  INVx1_ASAP7_75t_L         g01427(.A(new_n1612), .Y(new_n1684));
  AOI221xp5_ASAP7_75t_L     g01428(.A1(new_n1583), .A2(new_n1584), .B1(new_n1681), .B2(new_n1676), .C(new_n1684), .Y(new_n1685));
  AOI22xp33_ASAP7_75t_L     g01429(.A1(new_n345), .A2(\b[18] ), .B1(new_n342), .B2(new_n1363), .Y(new_n1686));
  OAI221xp5_ASAP7_75t_L     g01430(.A1(new_n406), .A2(new_n1244), .B1(new_n1051), .B2(new_n365), .C(new_n1686), .Y(new_n1687));
  XNOR2x2_ASAP7_75t_L       g01431(.A(new_n339), .B(new_n1687), .Y(new_n1688));
  NOR3xp33_ASAP7_75t_L      g01432(.A(new_n1683), .B(new_n1685), .C(new_n1688), .Y(new_n1689));
  NOR3xp33_ASAP7_75t_L      g01433(.A(new_n1680), .B(new_n1678), .C(new_n1677), .Y(new_n1690));
  AOI21xp33_ASAP7_75t_L     g01434(.A1(new_n1674), .A2(new_n1675), .B(new_n1618), .Y(new_n1691));
  NOR2xp33_ASAP7_75t_L      g01435(.A(new_n1690), .B(new_n1691), .Y(new_n1692));
  A2O1A1Ixp33_ASAP7_75t_L   g01436(.A1(new_n1584), .A2(new_n1583), .B(new_n1684), .C(new_n1692), .Y(new_n1693));
  INVx1_ASAP7_75t_L         g01437(.A(new_n1685), .Y(new_n1694));
  XNOR2x2_ASAP7_75t_L       g01438(.A(\a[5] ), .B(new_n1687), .Y(new_n1695));
  AOI21xp33_ASAP7_75t_L     g01439(.A1(new_n1694), .A2(new_n1693), .B(new_n1695), .Y(new_n1696));
  NOR2xp33_ASAP7_75t_L      g01440(.A(new_n1689), .B(new_n1696), .Y(new_n1697));
  AND3x1_ASAP7_75t_L        g01441(.A(new_n1589), .B(new_n1587), .C(new_n1524), .Y(new_n1698));
  AOI21xp33_ASAP7_75t_L     g01442(.A1(new_n1518), .A2(new_n1591), .B(new_n1698), .Y(new_n1699));
  NAND2xp33_ASAP7_75t_L     g01443(.A(new_n1697), .B(new_n1699), .Y(new_n1700));
  NAND3xp33_ASAP7_75t_L     g01444(.A(new_n1694), .B(new_n1693), .C(new_n1695), .Y(new_n1701));
  OAI21xp33_ASAP7_75t_L     g01445(.A1(new_n1685), .A2(new_n1683), .B(new_n1688), .Y(new_n1702));
  NAND2xp33_ASAP7_75t_L     g01446(.A(new_n1702), .B(new_n1701), .Y(new_n1703));
  A2O1A1Ixp33_ASAP7_75t_L   g01447(.A1(new_n1518), .A2(new_n1591), .B(new_n1698), .C(new_n1703), .Y(new_n1704));
  NAND2xp33_ASAP7_75t_L     g01448(.A(new_n1704), .B(new_n1700), .Y(new_n1705));
  A2O1A1O1Ixp25_ASAP7_75t_L g01449(.A1(new_n1358), .A2(new_n1361), .B(new_n1357), .C(new_n1495), .D(new_n1494), .Y(new_n1706));
  INVx1_ASAP7_75t_L         g01450(.A(new_n1595), .Y(new_n1707));
  NOR2xp33_ASAP7_75t_L      g01451(.A(\b[20] ), .B(\b[21] ), .Y(new_n1708));
  INVx1_ASAP7_75t_L         g01452(.A(\b[21] ), .Y(new_n1709));
  NOR2xp33_ASAP7_75t_L      g01453(.A(new_n1594), .B(new_n1709), .Y(new_n1710));
  NOR2xp33_ASAP7_75t_L      g01454(.A(new_n1708), .B(new_n1710), .Y(new_n1711));
  INVx1_ASAP7_75t_L         g01455(.A(new_n1711), .Y(new_n1712));
  O2A1O1Ixp33_ASAP7_75t_L   g01456(.A1(new_n1597), .A2(new_n1706), .B(new_n1707), .C(new_n1712), .Y(new_n1713));
  NOR3xp33_ASAP7_75t_L      g01457(.A(new_n1598), .B(new_n1711), .C(new_n1595), .Y(new_n1714));
  NOR2xp33_ASAP7_75t_L      g01458(.A(new_n1713), .B(new_n1714), .Y(new_n1715));
  AOI22xp33_ASAP7_75t_L     g01459(.A1(new_n272), .A2(\b[21] ), .B1(new_n269), .B2(new_n1715), .Y(new_n1716));
  OAI221xp5_ASAP7_75t_L     g01460(.A1(new_n261), .A2(new_n1594), .B1(new_n1493), .B2(new_n277), .C(new_n1716), .Y(new_n1717));
  XNOR2x2_ASAP7_75t_L       g01461(.A(\a[2] ), .B(new_n1717), .Y(new_n1718));
  XOR2x2_ASAP7_75t_L        g01462(.A(new_n1718), .B(new_n1705), .Y(new_n1719));
  A2O1A1O1Ixp25_ASAP7_75t_L g01463(.A1(new_n1505), .A2(new_n1512), .B(new_n1609), .C(new_n1606), .D(new_n1604), .Y(new_n1720));
  XNOR2x2_ASAP7_75t_L       g01464(.A(new_n1720), .B(new_n1719), .Y(\f[21] ));
  MAJIxp5_ASAP7_75t_L       g01465(.A(new_n1720), .B(new_n1705), .C(new_n1718), .Y(new_n1722));
  A2O1A1O1Ixp25_ASAP7_75t_L g01466(.A1(new_n1583), .A2(new_n1584), .B(new_n1684), .C(new_n1681), .D(new_n1690), .Y(new_n1723));
  NAND2xp33_ASAP7_75t_L     g01467(.A(\b[14] ), .B(new_n480), .Y(new_n1724));
  NAND2xp33_ASAP7_75t_L     g01468(.A(\b[15] ), .B(new_n441), .Y(new_n1725));
  AOI22xp33_ASAP7_75t_L     g01469(.A1(new_n451), .A2(\b[16] ), .B1(new_n448), .B2(new_n1058), .Y(new_n1726));
  NAND4xp25_ASAP7_75t_L     g01470(.A(new_n1726), .B(\a[8] ), .C(new_n1724), .D(new_n1725), .Y(new_n1727));
  NAND2xp33_ASAP7_75t_L     g01471(.A(new_n1725), .B(new_n1726), .Y(new_n1728));
  A2O1A1Ixp33_ASAP7_75t_L   g01472(.A1(\b[14] ), .A2(new_n480), .B(new_n1728), .C(new_n445), .Y(new_n1729));
  AND2x2_ASAP7_75t_L        g01473(.A(new_n1727), .B(new_n1729), .Y(new_n1730));
  OAI211xp5_ASAP7_75t_L     g01474(.A1(new_n1669), .A2(new_n1670), .B(new_n1625), .C(new_n1624), .Y(new_n1731));
  A2O1A1O1Ixp25_ASAP7_75t_L g01475(.A1(new_n1567), .A2(new_n1526), .B(new_n1619), .C(new_n1731), .D(new_n1672), .Y(new_n1732));
  INVx1_ASAP7_75t_L         g01476(.A(new_n1650), .Y(new_n1733));
  INVx1_ASAP7_75t_L         g01477(.A(new_n1652), .Y(new_n1734));
  OAI211xp5_ASAP7_75t_L     g01478(.A1(new_n1733), .A2(new_n1734), .B(new_n1646), .C(new_n1642), .Y(new_n1735));
  A2O1A1Ixp33_ASAP7_75t_L   g01479(.A1(new_n1654), .A2(new_n1653), .B(new_n1660), .C(new_n1735), .Y(new_n1736));
  NAND2xp33_ASAP7_75t_L     g01480(.A(\b[5] ), .B(new_n1194), .Y(new_n1737));
  NAND2xp33_ASAP7_75t_L     g01481(.A(\b[6] ), .B(new_n1103), .Y(new_n1738));
  AOI32xp33_ASAP7_75t_L     g01482(.A1(new_n424), .A2(new_n426), .A3(new_n1110), .B1(new_n1113), .B2(\b[7] ), .Y(new_n1739));
  NAND3xp33_ASAP7_75t_L     g01483(.A(new_n1739), .B(new_n1738), .C(new_n1737), .Y(new_n1740));
  NOR2xp33_ASAP7_75t_L      g01484(.A(new_n1107), .B(new_n1740), .Y(new_n1741));
  NAND2xp33_ASAP7_75t_L     g01485(.A(new_n1107), .B(new_n1740), .Y(new_n1742));
  INVx1_ASAP7_75t_L         g01486(.A(new_n1742), .Y(new_n1743));
  NOR3xp33_ASAP7_75t_L      g01487(.A(new_n1628), .B(new_n1550), .C(new_n1552), .Y(new_n1744));
  NAND2xp33_ASAP7_75t_L     g01488(.A(new_n1633), .B(new_n1744), .Y(new_n1745));
  A2O1A1Ixp33_ASAP7_75t_L   g01489(.A1(new_n1635), .A2(new_n1634), .B(new_n1645), .C(new_n1745), .Y(new_n1746));
  NAND2xp33_ASAP7_75t_L     g01490(.A(\b[2] ), .B(new_n1548), .Y(new_n1747));
  NOR2xp33_ASAP7_75t_L      g01491(.A(new_n299), .B(new_n1398), .Y(new_n1748));
  INVx1_ASAP7_75t_L         g01492(.A(new_n1748), .Y(new_n1749));
  OAI32xp33_ASAP7_75t_L     g01493(.A1(new_n325), .A2(new_n327), .A3(new_n1411), .B1(new_n323), .B2(new_n1412), .Y(new_n1750));
  INVx1_ASAP7_75t_L         g01494(.A(new_n1750), .Y(new_n1751));
  NAND4xp25_ASAP7_75t_L     g01495(.A(new_n1751), .B(\a[20] ), .C(new_n1747), .D(new_n1749), .Y(new_n1752));
  INVx1_ASAP7_75t_L         g01496(.A(new_n1747), .Y(new_n1753));
  OAI31xp33_ASAP7_75t_L     g01497(.A1(new_n1753), .A2(new_n1750), .A3(new_n1748), .B(new_n1401), .Y(new_n1754));
  NAND2xp33_ASAP7_75t_L     g01498(.A(\a[23] ), .B(new_n1633), .Y(new_n1755));
  XNOR2x2_ASAP7_75t_L       g01499(.A(\a[22] ), .B(\a[21] ), .Y(new_n1756));
  INVx1_ASAP7_75t_L         g01500(.A(new_n1756), .Y(new_n1757));
  NAND2xp33_ASAP7_75t_L     g01501(.A(new_n1757), .B(new_n1632), .Y(new_n1758));
  INVx1_ASAP7_75t_L         g01502(.A(\a[22] ), .Y(new_n1759));
  NAND2xp33_ASAP7_75t_L     g01503(.A(\a[23] ), .B(new_n1759), .Y(new_n1760));
  INVx1_ASAP7_75t_L         g01504(.A(\a[23] ), .Y(new_n1761));
  NAND2xp33_ASAP7_75t_L     g01505(.A(\a[22] ), .B(new_n1761), .Y(new_n1762));
  AND2x2_ASAP7_75t_L        g01506(.A(new_n1760), .B(new_n1762), .Y(new_n1763));
  NOR2xp33_ASAP7_75t_L      g01507(.A(new_n1632), .B(new_n1763), .Y(new_n1764));
  NAND2xp33_ASAP7_75t_L     g01508(.A(new_n1762), .B(new_n1760), .Y(new_n1765));
  NOR2xp33_ASAP7_75t_L      g01509(.A(new_n1765), .B(new_n1632), .Y(new_n1766));
  AOI22xp33_ASAP7_75t_L     g01510(.A1(new_n1766), .A2(\b[1] ), .B1(new_n271), .B2(new_n1764), .Y(new_n1767));
  O2A1O1Ixp33_ASAP7_75t_L   g01511(.A1(new_n1758), .A2(new_n258), .B(new_n1767), .C(new_n1755), .Y(new_n1768));
  NAND2xp33_ASAP7_75t_L     g01512(.A(new_n1631), .B(new_n1630), .Y(new_n1769));
  NOR2xp33_ASAP7_75t_L      g01513(.A(new_n1756), .B(new_n1769), .Y(new_n1770));
  NAND2xp33_ASAP7_75t_L     g01514(.A(new_n1765), .B(new_n1769), .Y(new_n1771));
  NAND2xp33_ASAP7_75t_L     g01515(.A(new_n1769), .B(new_n1763), .Y(new_n1772));
  OAI22xp33_ASAP7_75t_L     g01516(.A1(new_n1772), .A2(new_n276), .B1(new_n270), .B2(new_n1771), .Y(new_n1773));
  A2O1A1O1Ixp25_ASAP7_75t_L g01517(.A1(new_n1769), .A2(\a[23] ), .B(new_n1770), .C(\b[0] ), .D(new_n1773), .Y(new_n1774));
  NOR2xp33_ASAP7_75t_L      g01518(.A(new_n1774), .B(new_n1768), .Y(new_n1775));
  NAND3xp33_ASAP7_75t_L     g01519(.A(new_n1752), .B(new_n1775), .C(new_n1754), .Y(new_n1776));
  INVx1_ASAP7_75t_L         g01520(.A(new_n1776), .Y(new_n1777));
  NOR4xp25_ASAP7_75t_L      g01521(.A(new_n1753), .B(new_n1750), .C(new_n1401), .D(new_n1748), .Y(new_n1778));
  AOI31xp33_ASAP7_75t_L     g01522(.A1(new_n1751), .A2(new_n1749), .A3(new_n1747), .B(\a[20] ), .Y(new_n1779));
  NOR2xp33_ASAP7_75t_L      g01523(.A(new_n1778), .B(new_n1779), .Y(new_n1780));
  NOR2xp33_ASAP7_75t_L      g01524(.A(new_n1775), .B(new_n1780), .Y(new_n1781));
  OAI21xp33_ASAP7_75t_L     g01525(.A1(new_n1777), .A2(new_n1781), .B(new_n1746), .Y(new_n1782));
  NAND2xp33_ASAP7_75t_L     g01526(.A(new_n1641), .B(new_n1638), .Y(new_n1783));
  MAJIxp5_ASAP7_75t_L       g01527(.A(new_n1783), .B(new_n1633), .C(new_n1744), .Y(new_n1784));
  OR2x4_ASAP7_75t_L         g01528(.A(new_n1774), .B(new_n1768), .Y(new_n1785));
  OAI21xp33_ASAP7_75t_L     g01529(.A1(new_n1778), .A2(new_n1779), .B(new_n1785), .Y(new_n1786));
  NAND3xp33_ASAP7_75t_L     g01530(.A(new_n1784), .B(new_n1776), .C(new_n1786), .Y(new_n1787));
  OAI211xp5_ASAP7_75t_L     g01531(.A1(new_n1741), .A2(new_n1743), .B(new_n1787), .C(new_n1782), .Y(new_n1788));
  INVx1_ASAP7_75t_L         g01532(.A(new_n1741), .Y(new_n1789));
  AOI21xp33_ASAP7_75t_L     g01533(.A1(new_n1786), .A2(new_n1776), .B(new_n1784), .Y(new_n1790));
  NAND2xp33_ASAP7_75t_L     g01534(.A(new_n1776), .B(new_n1786), .Y(new_n1791));
  NOR2xp33_ASAP7_75t_L      g01535(.A(new_n1746), .B(new_n1791), .Y(new_n1792));
  OAI211xp5_ASAP7_75t_L     g01536(.A1(new_n1790), .A2(new_n1792), .B(new_n1742), .C(new_n1789), .Y(new_n1793));
  NAND3xp33_ASAP7_75t_L     g01537(.A(new_n1736), .B(new_n1788), .C(new_n1793), .Y(new_n1794));
  OAI22xp33_ASAP7_75t_L     g01538(.A1(new_n1658), .A2(new_n1657), .B1(new_n1560), .B2(new_n1655), .Y(new_n1795));
  AOI211xp5_ASAP7_75t_L     g01539(.A1(new_n1789), .A2(new_n1742), .B(new_n1790), .C(new_n1792), .Y(new_n1796));
  AOI211xp5_ASAP7_75t_L     g01540(.A1(new_n1782), .A2(new_n1787), .B(new_n1743), .C(new_n1741), .Y(new_n1797));
  OAI211xp5_ASAP7_75t_L     g01541(.A1(new_n1796), .A2(new_n1797), .B(new_n1795), .C(new_n1735), .Y(new_n1798));
  NOR2xp33_ASAP7_75t_L      g01542(.A(new_n503), .B(new_n909), .Y(new_n1799));
  NAND2xp33_ASAP7_75t_L     g01543(.A(\b[9] ), .B(new_n817), .Y(new_n1800));
  NAND2xp33_ASAP7_75t_L     g01544(.A(\b[10] ), .B(new_n826), .Y(new_n1801));
  OAI311xp33_ASAP7_75t_L    g01545(.A1(new_n639), .A2(new_n851), .A3(new_n911), .B1(new_n1801), .C1(new_n1800), .Y(new_n1802));
  OR3x1_ASAP7_75t_L         g01546(.A(new_n1802), .B(new_n813), .C(new_n1799), .Y(new_n1803));
  A2O1A1Ixp33_ASAP7_75t_L   g01547(.A1(\b[8] ), .A2(new_n908), .B(new_n1802), .C(new_n813), .Y(new_n1804));
  AND2x2_ASAP7_75t_L        g01548(.A(new_n1804), .B(new_n1803), .Y(new_n1805));
  NAND3xp33_ASAP7_75t_L     g01549(.A(new_n1794), .B(new_n1798), .C(new_n1805), .Y(new_n1806));
  AOI211xp5_ASAP7_75t_L     g01550(.A1(new_n1795), .A2(new_n1735), .B(new_n1796), .C(new_n1797), .Y(new_n1807));
  AOI21xp33_ASAP7_75t_L     g01551(.A1(new_n1793), .A2(new_n1788), .B(new_n1736), .Y(new_n1808));
  NAND2xp33_ASAP7_75t_L     g01552(.A(new_n1804), .B(new_n1803), .Y(new_n1809));
  OAI21xp33_ASAP7_75t_L     g01553(.A1(new_n1807), .A2(new_n1808), .B(new_n1809), .Y(new_n1810));
  NAND4xp25_ASAP7_75t_L     g01554(.A(new_n1665), .B(new_n1661), .C(new_n1656), .D(new_n1666), .Y(new_n1811));
  A2O1A1O1Ixp25_ASAP7_75t_L g01555(.A1(new_n1562), .A2(new_n1534), .B(new_n1563), .C(new_n1811), .D(new_n1667), .Y(new_n1812));
  NAND3xp33_ASAP7_75t_L     g01556(.A(new_n1812), .B(new_n1810), .C(new_n1806), .Y(new_n1813));
  NOR3xp33_ASAP7_75t_L      g01557(.A(new_n1808), .B(new_n1807), .C(new_n1809), .Y(new_n1814));
  AOI21xp33_ASAP7_75t_L     g01558(.A1(new_n1794), .A2(new_n1798), .B(new_n1805), .Y(new_n1815));
  AO22x1_ASAP7_75t_L        g01559(.A1(new_n1656), .A2(new_n1661), .B1(new_n1666), .B2(new_n1665), .Y(new_n1816));
  OAI21xp33_ASAP7_75t_L     g01560(.A1(new_n1668), .A2(new_n1626), .B(new_n1816), .Y(new_n1817));
  OAI21xp33_ASAP7_75t_L     g01561(.A1(new_n1814), .A2(new_n1815), .B(new_n1817), .Y(new_n1818));
  NAND2xp33_ASAP7_75t_L     g01562(.A(\b[11] ), .B(new_n674), .Y(new_n1819));
  NAND2xp33_ASAP7_75t_L     g01563(.A(\b[12] ), .B(new_n590), .Y(new_n1820));
  AOI22xp33_ASAP7_75t_L     g01564(.A1(new_n600), .A2(\b[13] ), .B1(new_n597), .B2(new_n800), .Y(new_n1821));
  NAND3xp33_ASAP7_75t_L     g01565(.A(new_n1821), .B(new_n1820), .C(new_n1819), .Y(new_n1822));
  XNOR2x2_ASAP7_75t_L       g01566(.A(new_n594), .B(new_n1822), .Y(new_n1823));
  AOI21xp33_ASAP7_75t_L     g01567(.A1(new_n1818), .A2(new_n1813), .B(new_n1823), .Y(new_n1824));
  NAND2xp33_ASAP7_75t_L     g01568(.A(new_n1806), .B(new_n1810), .Y(new_n1825));
  NOR2xp33_ASAP7_75t_L      g01569(.A(new_n1817), .B(new_n1825), .Y(new_n1826));
  INVx1_ASAP7_75t_L         g01570(.A(new_n1818), .Y(new_n1827));
  XNOR2x2_ASAP7_75t_L       g01571(.A(\a[11] ), .B(new_n1822), .Y(new_n1828));
  NOR3xp33_ASAP7_75t_L      g01572(.A(new_n1828), .B(new_n1827), .C(new_n1826), .Y(new_n1829));
  NOR3xp33_ASAP7_75t_L      g01573(.A(new_n1829), .B(new_n1732), .C(new_n1824), .Y(new_n1830));
  OAI21xp33_ASAP7_75t_L     g01574(.A1(new_n1826), .A2(new_n1827), .B(new_n1828), .Y(new_n1831));
  NAND3xp33_ASAP7_75t_L     g01575(.A(new_n1823), .B(new_n1818), .C(new_n1813), .Y(new_n1832));
  AOI221xp5_ASAP7_75t_L     g01576(.A1(new_n1679), .A2(new_n1731), .B1(new_n1831), .B2(new_n1832), .C(new_n1672), .Y(new_n1833));
  NOR3xp33_ASAP7_75t_L      g01577(.A(new_n1730), .B(new_n1830), .C(new_n1833), .Y(new_n1834));
  OA21x2_ASAP7_75t_L        g01578(.A1(new_n1830), .A2(new_n1833), .B(new_n1730), .Y(new_n1835));
  NOR3xp33_ASAP7_75t_L      g01579(.A(new_n1723), .B(new_n1834), .C(new_n1835), .Y(new_n1836));
  OAI21xp33_ASAP7_75t_L     g01580(.A1(new_n1834), .A2(new_n1835), .B(new_n1723), .Y(new_n1837));
  INVx1_ASAP7_75t_L         g01581(.A(new_n1837), .Y(new_n1838));
  AOI22xp33_ASAP7_75t_L     g01582(.A1(new_n345), .A2(\b[19] ), .B1(new_n342), .B2(new_n1499), .Y(new_n1839));
  OAI221xp5_ASAP7_75t_L     g01583(.A1(new_n406), .A2(new_n1356), .B1(new_n1244), .B2(new_n365), .C(new_n1839), .Y(new_n1840));
  XNOR2x2_ASAP7_75t_L       g01584(.A(new_n339), .B(new_n1840), .Y(new_n1841));
  NOR3xp33_ASAP7_75t_L      g01585(.A(new_n1838), .B(new_n1841), .C(new_n1836), .Y(new_n1842));
  INVx1_ASAP7_75t_L         g01586(.A(new_n1836), .Y(new_n1843));
  XNOR2x2_ASAP7_75t_L       g01587(.A(\a[5] ), .B(new_n1840), .Y(new_n1844));
  AOI21xp33_ASAP7_75t_L     g01588(.A1(new_n1843), .A2(new_n1837), .B(new_n1844), .Y(new_n1845));
  NOR2xp33_ASAP7_75t_L      g01589(.A(new_n1842), .B(new_n1845), .Y(new_n1846));
  NOR3xp33_ASAP7_75t_L      g01590(.A(new_n1683), .B(new_n1685), .C(new_n1695), .Y(new_n1847));
  A2O1A1O1Ixp25_ASAP7_75t_L g01591(.A1(new_n1591), .A2(new_n1518), .B(new_n1698), .C(new_n1703), .D(new_n1847), .Y(new_n1848));
  NAND2xp33_ASAP7_75t_L     g01592(.A(new_n1846), .B(new_n1848), .Y(new_n1849));
  NAND3xp33_ASAP7_75t_L     g01593(.A(new_n1843), .B(new_n1837), .C(new_n1844), .Y(new_n1850));
  OAI21xp33_ASAP7_75t_L     g01594(.A1(new_n1836), .A2(new_n1838), .B(new_n1841), .Y(new_n1851));
  NAND2xp33_ASAP7_75t_L     g01595(.A(new_n1851), .B(new_n1850), .Y(new_n1852));
  INVx1_ASAP7_75t_L         g01596(.A(new_n1847), .Y(new_n1853));
  OAI21xp33_ASAP7_75t_L     g01597(.A1(new_n1697), .A2(new_n1699), .B(new_n1853), .Y(new_n1854));
  NAND2xp33_ASAP7_75t_L     g01598(.A(new_n1852), .B(new_n1854), .Y(new_n1855));
  NOR2xp33_ASAP7_75t_L      g01599(.A(\b[21] ), .B(\b[22] ), .Y(new_n1856));
  INVx1_ASAP7_75t_L         g01600(.A(\b[22] ), .Y(new_n1857));
  NOR2xp33_ASAP7_75t_L      g01601(.A(new_n1709), .B(new_n1857), .Y(new_n1858));
  NOR2xp33_ASAP7_75t_L      g01602(.A(new_n1856), .B(new_n1858), .Y(new_n1859));
  A2O1A1Ixp33_ASAP7_75t_L   g01603(.A1(\b[21] ), .A2(\b[20] ), .B(new_n1713), .C(new_n1859), .Y(new_n1860));
  O2A1O1Ixp33_ASAP7_75t_L   g01604(.A1(new_n1595), .A2(new_n1598), .B(new_n1711), .C(new_n1710), .Y(new_n1861));
  OAI21xp33_ASAP7_75t_L     g01605(.A1(new_n1856), .A2(new_n1858), .B(new_n1861), .Y(new_n1862));
  NAND2xp33_ASAP7_75t_L     g01606(.A(new_n1860), .B(new_n1862), .Y(new_n1863));
  INVx1_ASAP7_75t_L         g01607(.A(new_n1863), .Y(new_n1864));
  NOR2xp33_ASAP7_75t_L      g01608(.A(new_n1857), .B(new_n632), .Y(new_n1865));
  AOI221xp5_ASAP7_75t_L     g01609(.A1(new_n380), .A2(\b[21] ), .B1(new_n269), .B2(new_n1864), .C(new_n1865), .Y(new_n1866));
  OAI21xp33_ASAP7_75t_L     g01610(.A1(new_n1594), .A2(new_n277), .B(new_n1866), .Y(new_n1867));
  XNOR2x2_ASAP7_75t_L       g01611(.A(new_n265), .B(new_n1867), .Y(new_n1868));
  AOI21xp33_ASAP7_75t_L     g01612(.A1(new_n1855), .A2(new_n1849), .B(new_n1868), .Y(new_n1869));
  AND3x1_ASAP7_75t_L        g01613(.A(new_n1855), .B(new_n1849), .C(new_n1868), .Y(new_n1870));
  NOR2xp33_ASAP7_75t_L      g01614(.A(new_n1869), .B(new_n1870), .Y(new_n1871));
  XOR2x2_ASAP7_75t_L        g01615(.A(new_n1871), .B(new_n1722), .Y(\f[22] ));
  NOR3xp33_ASAP7_75t_L      g01616(.A(new_n1838), .B(new_n1844), .C(new_n1836), .Y(new_n1873));
  INVx1_ASAP7_75t_L         g01617(.A(new_n1873), .Y(new_n1874));
  OR3x1_ASAP7_75t_L         g01618(.A(new_n1730), .B(new_n1830), .C(new_n1833), .Y(new_n1875));
  NAND2xp33_ASAP7_75t_L     g01619(.A(\b[15] ), .B(new_n480), .Y(new_n1876));
  NAND2xp33_ASAP7_75t_L     g01620(.A(\b[16] ), .B(new_n441), .Y(new_n1877));
  AOI32xp33_ASAP7_75t_L     g01621(.A1(new_n1250), .A2(new_n1247), .A3(new_n448), .B1(new_n451), .B2(\b[17] ), .Y(new_n1878));
  NAND4xp25_ASAP7_75t_L     g01622(.A(new_n1878), .B(\a[8] ), .C(new_n1876), .D(new_n1877), .Y(new_n1879));
  NAND2xp33_ASAP7_75t_L     g01623(.A(new_n1877), .B(new_n1878), .Y(new_n1880));
  A2O1A1Ixp33_ASAP7_75t_L   g01624(.A1(\b[15] ), .A2(new_n480), .B(new_n1880), .C(new_n445), .Y(new_n1881));
  NAND2xp33_ASAP7_75t_L     g01625(.A(new_n1879), .B(new_n1881), .Y(new_n1882));
  NOR2xp33_ASAP7_75t_L      g01626(.A(new_n1807), .B(new_n1808), .Y(new_n1883));
  MAJIxp5_ASAP7_75t_L       g01627(.A(new_n1817), .B(new_n1809), .C(new_n1883), .Y(new_n1884));
  NOR2xp33_ASAP7_75t_L      g01628(.A(new_n559), .B(new_n909), .Y(new_n1885));
  INVx1_ASAP7_75t_L         g01629(.A(new_n1885), .Y(new_n1886));
  NAND2xp33_ASAP7_75t_L     g01630(.A(\b[10] ), .B(new_n817), .Y(new_n1887));
  AOI32xp33_ASAP7_75t_L     g01631(.A1(new_n700), .A2(new_n698), .A3(new_n823), .B1(\b[11] ), .B2(new_n826), .Y(new_n1888));
  AND4x1_ASAP7_75t_L        g01632(.A(new_n1888), .B(new_n1887), .C(new_n1886), .D(\a[14] ), .Y(new_n1889));
  AOI31xp33_ASAP7_75t_L     g01633(.A1(new_n1888), .A2(new_n1887), .A3(new_n1886), .B(\a[14] ), .Y(new_n1890));
  NOR2xp33_ASAP7_75t_L      g01634(.A(new_n1890), .B(new_n1889), .Y(new_n1891));
  INVx1_ASAP7_75t_L         g01635(.A(new_n1891), .Y(new_n1892));
  A2O1A1Ixp33_ASAP7_75t_L   g01636(.A1(new_n1795), .A2(new_n1735), .B(new_n1797), .C(new_n1788), .Y(new_n1893));
  NAND2xp33_ASAP7_75t_L     g01637(.A(\b[6] ), .B(new_n1194), .Y(new_n1894));
  NAND2xp33_ASAP7_75t_L     g01638(.A(\b[7] ), .B(new_n1103), .Y(new_n1895));
  OAI221xp5_ASAP7_75t_L     g01639(.A1(new_n1198), .A2(new_n503), .B1(new_n1197), .B2(new_n509), .C(new_n1895), .Y(new_n1896));
  INVx1_ASAP7_75t_L         g01640(.A(new_n1896), .Y(new_n1897));
  NAND3xp33_ASAP7_75t_L     g01641(.A(new_n1897), .B(new_n1894), .C(\a[17] ), .Y(new_n1898));
  A2O1A1Ixp33_ASAP7_75t_L   g01642(.A1(\b[6] ), .A2(new_n1194), .B(new_n1896), .C(new_n1107), .Y(new_n1899));
  OAI21xp33_ASAP7_75t_L     g01643(.A1(new_n1778), .A2(new_n1779), .B(new_n1775), .Y(new_n1900));
  NAND2xp33_ASAP7_75t_L     g01644(.A(\b[3] ), .B(new_n1548), .Y(new_n1901));
  NAND2xp33_ASAP7_75t_L     g01645(.A(\b[4] ), .B(new_n1410), .Y(new_n1902));
  AOI32xp33_ASAP7_75t_L     g01646(.A1(new_n358), .A2(new_n356), .A3(new_n1404), .B1(\b[5] ), .B2(new_n1406), .Y(new_n1903));
  NAND3xp33_ASAP7_75t_L     g01647(.A(new_n1903), .B(new_n1902), .C(new_n1901), .Y(new_n1904));
  NOR2xp33_ASAP7_75t_L      g01648(.A(new_n1401), .B(new_n1904), .Y(new_n1905));
  INVx1_ASAP7_75t_L         g01649(.A(new_n1905), .Y(new_n1906));
  AOI31xp33_ASAP7_75t_L     g01650(.A1(new_n1903), .A2(new_n1902), .A3(new_n1901), .B(\a[20] ), .Y(new_n1907));
  INVx1_ASAP7_75t_L         g01651(.A(new_n1907), .Y(new_n1908));
  A2O1A1O1Ixp25_ASAP7_75t_L g01652(.A1(new_n1756), .A2(new_n1632), .B(new_n258), .C(new_n1767), .D(new_n1761), .Y(new_n1909));
  NOR3xp33_ASAP7_75t_L      g01653(.A(new_n1763), .B(new_n1757), .C(new_n1769), .Y(new_n1910));
  INVx1_ASAP7_75t_L         g01654(.A(new_n1910), .Y(new_n1911));
  NOR2xp33_ASAP7_75t_L      g01655(.A(new_n1771), .B(new_n283), .Y(new_n1912));
  AOI221xp5_ASAP7_75t_L     g01656(.A1(\b[2] ), .A2(new_n1766), .B1(new_n1770), .B2(\b[1] ), .C(new_n1912), .Y(new_n1913));
  OAI21xp33_ASAP7_75t_L     g01657(.A1(new_n258), .A2(new_n1911), .B(new_n1913), .Y(new_n1914));
  NOR2xp33_ASAP7_75t_L      g01658(.A(new_n1909), .B(new_n1914), .Y(new_n1915));
  NAND2xp33_ASAP7_75t_L     g01659(.A(\b[1] ), .B(new_n1770), .Y(new_n1916));
  OAI221xp5_ASAP7_75t_L     g01660(.A1(new_n1771), .A2(new_n283), .B1(new_n278), .B2(new_n1772), .C(new_n1916), .Y(new_n1917));
  A2O1A1Ixp33_ASAP7_75t_L   g01661(.A1(\b[0] ), .A2(new_n1910), .B(new_n1917), .C(new_n1909), .Y(new_n1918));
  INVx1_ASAP7_75t_L         g01662(.A(new_n1918), .Y(new_n1919));
  OAI211xp5_ASAP7_75t_L     g01663(.A1(new_n1915), .A2(new_n1919), .B(new_n1906), .C(new_n1908), .Y(new_n1920));
  NOR2xp33_ASAP7_75t_L      g01664(.A(new_n258), .B(new_n1911), .Y(new_n1921));
  OR3x1_ASAP7_75t_L         g01665(.A(new_n1909), .B(new_n1921), .C(new_n1917), .Y(new_n1922));
  OAI211xp5_ASAP7_75t_L     g01666(.A1(new_n1907), .A2(new_n1905), .B(new_n1922), .C(new_n1918), .Y(new_n1923));
  NAND4xp25_ASAP7_75t_L     g01667(.A(new_n1782), .B(new_n1923), .C(new_n1920), .D(new_n1900), .Y(new_n1924));
  INVx1_ASAP7_75t_L         g01668(.A(new_n1900), .Y(new_n1925));
  NAND2xp33_ASAP7_75t_L     g01669(.A(new_n1923), .B(new_n1920), .Y(new_n1926));
  A2O1A1Ixp33_ASAP7_75t_L   g01670(.A1(new_n1791), .A2(new_n1746), .B(new_n1925), .C(new_n1926), .Y(new_n1927));
  NAND4xp25_ASAP7_75t_L     g01671(.A(new_n1924), .B(new_n1927), .C(new_n1898), .D(new_n1899), .Y(new_n1928));
  AOI22xp33_ASAP7_75t_L     g01672(.A1(new_n1898), .A2(new_n1899), .B1(new_n1924), .B2(new_n1927), .Y(new_n1929));
  INVx1_ASAP7_75t_L         g01673(.A(new_n1929), .Y(new_n1930));
  NAND3xp33_ASAP7_75t_L     g01674(.A(new_n1930), .B(new_n1928), .C(new_n1893), .Y(new_n1931));
  AOI21xp33_ASAP7_75t_L     g01675(.A1(new_n1736), .A2(new_n1793), .B(new_n1796), .Y(new_n1932));
  INVx1_ASAP7_75t_L         g01676(.A(new_n1928), .Y(new_n1933));
  OAI21xp33_ASAP7_75t_L     g01677(.A1(new_n1929), .A2(new_n1933), .B(new_n1932), .Y(new_n1934));
  AOI21xp33_ASAP7_75t_L     g01678(.A1(new_n1934), .A2(new_n1931), .B(new_n1892), .Y(new_n1935));
  NOR3xp33_ASAP7_75t_L      g01679(.A(new_n1932), .B(new_n1933), .C(new_n1929), .Y(new_n1936));
  AOI21xp33_ASAP7_75t_L     g01680(.A1(new_n1930), .A2(new_n1928), .B(new_n1893), .Y(new_n1937));
  NOR3xp33_ASAP7_75t_L      g01681(.A(new_n1936), .B(new_n1937), .C(new_n1891), .Y(new_n1938));
  NOR3xp33_ASAP7_75t_L      g01682(.A(new_n1884), .B(new_n1935), .C(new_n1938), .Y(new_n1939));
  NAND2xp33_ASAP7_75t_L     g01683(.A(new_n1798), .B(new_n1794), .Y(new_n1940));
  MAJIxp5_ASAP7_75t_L       g01684(.A(new_n1812), .B(new_n1805), .C(new_n1940), .Y(new_n1941));
  OAI21xp33_ASAP7_75t_L     g01685(.A1(new_n1937), .A2(new_n1936), .B(new_n1891), .Y(new_n1942));
  NAND3xp33_ASAP7_75t_L     g01686(.A(new_n1892), .B(new_n1934), .C(new_n1931), .Y(new_n1943));
  AOI21xp33_ASAP7_75t_L     g01687(.A1(new_n1943), .A2(new_n1942), .B(new_n1941), .Y(new_n1944));
  NOR2xp33_ASAP7_75t_L      g01688(.A(new_n1944), .B(new_n1939), .Y(new_n1945));
  NOR2xp33_ASAP7_75t_L      g01689(.A(new_n763), .B(new_n1620), .Y(new_n1946));
  NAND2xp33_ASAP7_75t_L     g01690(.A(\b[13] ), .B(new_n590), .Y(new_n1947));
  OAI221xp5_ASAP7_75t_L     g01691(.A1(new_n676), .A2(new_n871), .B1(new_n675), .B2(new_n878), .C(new_n1947), .Y(new_n1948));
  OR3x1_ASAP7_75t_L         g01692(.A(new_n1948), .B(new_n594), .C(new_n1946), .Y(new_n1949));
  A2O1A1Ixp33_ASAP7_75t_L   g01693(.A1(\b[12] ), .A2(new_n674), .B(new_n1948), .C(new_n594), .Y(new_n1950));
  AND2x2_ASAP7_75t_L        g01694(.A(new_n1950), .B(new_n1949), .Y(new_n1951));
  NAND2xp33_ASAP7_75t_L     g01695(.A(new_n1951), .B(new_n1945), .Y(new_n1952));
  NAND2xp33_ASAP7_75t_L     g01696(.A(new_n1950), .B(new_n1949), .Y(new_n1953));
  OAI21xp33_ASAP7_75t_L     g01697(.A1(new_n1944), .A2(new_n1939), .B(new_n1953), .Y(new_n1954));
  A2O1A1O1Ixp25_ASAP7_75t_L g01698(.A1(new_n1731), .A2(new_n1679), .B(new_n1672), .C(new_n1831), .D(new_n1829), .Y(new_n1955));
  AOI21xp33_ASAP7_75t_L     g01699(.A1(new_n1952), .A2(new_n1954), .B(new_n1955), .Y(new_n1956));
  NOR3xp33_ASAP7_75t_L      g01700(.A(new_n1953), .B(new_n1944), .C(new_n1939), .Y(new_n1957));
  OA21x2_ASAP7_75t_L        g01701(.A1(new_n1939), .A2(new_n1944), .B(new_n1953), .Y(new_n1958));
  OAI21xp33_ASAP7_75t_L     g01702(.A1(new_n1824), .A2(new_n1732), .B(new_n1832), .Y(new_n1959));
  NOR3xp33_ASAP7_75t_L      g01703(.A(new_n1959), .B(new_n1958), .C(new_n1957), .Y(new_n1960));
  OAI21xp33_ASAP7_75t_L     g01704(.A1(new_n1960), .A2(new_n1956), .B(new_n1882), .Y(new_n1961));
  AND2x2_ASAP7_75t_L        g01705(.A(new_n1879), .B(new_n1881), .Y(new_n1962));
  OAI21xp33_ASAP7_75t_L     g01706(.A1(new_n1957), .A2(new_n1958), .B(new_n1959), .Y(new_n1963));
  NAND3xp33_ASAP7_75t_L     g01707(.A(new_n1955), .B(new_n1952), .C(new_n1954), .Y(new_n1964));
  NAND3xp33_ASAP7_75t_L     g01708(.A(new_n1964), .B(new_n1962), .C(new_n1963), .Y(new_n1965));
  NAND2xp33_ASAP7_75t_L     g01709(.A(new_n1965), .B(new_n1961), .Y(new_n1966));
  O2A1O1Ixp33_ASAP7_75t_L   g01710(.A1(new_n1723), .A2(new_n1835), .B(new_n1875), .C(new_n1966), .Y(new_n1967));
  OAI21xp33_ASAP7_75t_L     g01711(.A1(new_n1835), .A2(new_n1723), .B(new_n1875), .Y(new_n1968));
  AND2x2_ASAP7_75t_L        g01712(.A(new_n1965), .B(new_n1961), .Y(new_n1969));
  NOR2xp33_ASAP7_75t_L      g01713(.A(new_n1968), .B(new_n1969), .Y(new_n1970));
  NAND2xp33_ASAP7_75t_L     g01714(.A(\b[18] ), .B(new_n366), .Y(new_n1971));
  NOR2xp33_ASAP7_75t_L      g01715(.A(new_n1594), .B(new_n368), .Y(new_n1972));
  AOI221xp5_ASAP7_75t_L     g01716(.A1(new_n334), .A2(\b[19] ), .B1(new_n342), .B2(new_n1600), .C(new_n1972), .Y(new_n1973));
  NAND3xp33_ASAP7_75t_L     g01717(.A(new_n1973), .B(new_n1971), .C(\a[5] ), .Y(new_n1974));
  AO21x2_ASAP7_75t_L        g01718(.A1(new_n1971), .A2(new_n1973), .B(\a[5] ), .Y(new_n1975));
  NAND2xp33_ASAP7_75t_L     g01719(.A(new_n1974), .B(new_n1975), .Y(new_n1976));
  OAI21xp33_ASAP7_75t_L     g01720(.A1(new_n1967), .A2(new_n1970), .B(new_n1976), .Y(new_n1977));
  NAND2xp33_ASAP7_75t_L     g01721(.A(new_n1968), .B(new_n1969), .Y(new_n1978));
  A2O1A1Ixp33_ASAP7_75t_L   g01722(.A1(new_n1580), .A2(new_n1576), .B(new_n1588), .C(new_n1612), .Y(new_n1979));
  OAI21xp33_ASAP7_75t_L     g01723(.A1(new_n1830), .A2(new_n1833), .B(new_n1730), .Y(new_n1980));
  A2O1A1O1Ixp25_ASAP7_75t_L g01724(.A1(new_n1681), .A2(new_n1979), .B(new_n1690), .C(new_n1980), .D(new_n1834), .Y(new_n1981));
  NAND2xp33_ASAP7_75t_L     g01725(.A(new_n1966), .B(new_n1981), .Y(new_n1982));
  AND2x2_ASAP7_75t_L        g01726(.A(new_n1974), .B(new_n1975), .Y(new_n1983));
  NAND3xp33_ASAP7_75t_L     g01727(.A(new_n1982), .B(new_n1983), .C(new_n1978), .Y(new_n1984));
  NAND2xp33_ASAP7_75t_L     g01728(.A(new_n1977), .B(new_n1984), .Y(new_n1985));
  OAI211xp5_ASAP7_75t_L     g01729(.A1(new_n1846), .A2(new_n1848), .B(new_n1985), .C(new_n1874), .Y(new_n1986));
  AOI21xp33_ASAP7_75t_L     g01730(.A1(new_n1982), .A2(new_n1978), .B(new_n1983), .Y(new_n1987));
  NOR3xp33_ASAP7_75t_L      g01731(.A(new_n1970), .B(new_n1976), .C(new_n1967), .Y(new_n1988));
  NOR2xp33_ASAP7_75t_L      g01732(.A(new_n1988), .B(new_n1987), .Y(new_n1989));
  A2O1A1Ixp33_ASAP7_75t_L   g01733(.A1(new_n1854), .A2(new_n1852), .B(new_n1873), .C(new_n1989), .Y(new_n1990));
  INVx1_ASAP7_75t_L         g01734(.A(new_n1598), .Y(new_n1991));
  INVx1_ASAP7_75t_L         g01735(.A(new_n1710), .Y(new_n1992));
  A2O1A1Ixp33_ASAP7_75t_L   g01736(.A1(new_n1991), .A2(new_n1707), .B(new_n1708), .C(new_n1992), .Y(new_n1993));
  NOR2xp33_ASAP7_75t_L      g01737(.A(\b[22] ), .B(\b[23] ), .Y(new_n1994));
  INVx1_ASAP7_75t_L         g01738(.A(\b[23] ), .Y(new_n1995));
  NOR2xp33_ASAP7_75t_L      g01739(.A(new_n1857), .B(new_n1995), .Y(new_n1996));
  NOR2xp33_ASAP7_75t_L      g01740(.A(new_n1994), .B(new_n1996), .Y(new_n1997));
  A2O1A1Ixp33_ASAP7_75t_L   g01741(.A1(new_n1993), .A2(new_n1859), .B(new_n1858), .C(new_n1997), .Y(new_n1998));
  O2A1O1Ixp33_ASAP7_75t_L   g01742(.A1(new_n1710), .A2(new_n1713), .B(new_n1859), .C(new_n1858), .Y(new_n1999));
  INVx1_ASAP7_75t_L         g01743(.A(new_n1997), .Y(new_n2000));
  NAND2xp33_ASAP7_75t_L     g01744(.A(new_n2000), .B(new_n1999), .Y(new_n2001));
  AND2x2_ASAP7_75t_L        g01745(.A(new_n2001), .B(new_n1998), .Y(new_n2002));
  AOI22xp33_ASAP7_75t_L     g01746(.A1(new_n272), .A2(\b[23] ), .B1(new_n269), .B2(new_n2002), .Y(new_n2003));
  OAI221xp5_ASAP7_75t_L     g01747(.A1(new_n261), .A2(new_n1857), .B1(new_n1709), .B2(new_n277), .C(new_n2003), .Y(new_n2004));
  XNOR2x2_ASAP7_75t_L       g01748(.A(\a[2] ), .B(new_n2004), .Y(new_n2005));
  NAND3xp33_ASAP7_75t_L     g01749(.A(new_n2005), .B(new_n1990), .C(new_n1986), .Y(new_n2006));
  AOI211xp5_ASAP7_75t_L     g01750(.A1(new_n1852), .A2(new_n1854), .B(new_n1873), .C(new_n1989), .Y(new_n2007));
  O2A1O1Ixp33_ASAP7_75t_L   g01751(.A1(new_n1846), .A2(new_n1848), .B(new_n1874), .C(new_n1985), .Y(new_n2008));
  XNOR2x2_ASAP7_75t_L       g01752(.A(new_n265), .B(new_n2004), .Y(new_n2009));
  OAI21xp33_ASAP7_75t_L     g01753(.A1(new_n2008), .A2(new_n2007), .B(new_n2009), .Y(new_n2010));
  NAND2xp33_ASAP7_75t_L     g01754(.A(new_n2006), .B(new_n2010), .Y(new_n2011));
  AOI21xp33_ASAP7_75t_L     g01755(.A1(new_n1722), .A2(new_n1871), .B(new_n1870), .Y(new_n2012));
  XNOR2x2_ASAP7_75t_L       g01756(.A(new_n2011), .B(new_n2012), .Y(\f[23] ));
  NAND2xp33_ASAP7_75t_L     g01757(.A(new_n1986), .B(new_n1990), .Y(new_n2014));
  A2O1A1Ixp33_ASAP7_75t_L   g01758(.A1(new_n1722), .A2(new_n1871), .B(new_n1870), .C(new_n2011), .Y(new_n2015));
  NAND2xp33_ASAP7_75t_L     g01759(.A(\b[23] ), .B(new_n380), .Y(new_n2016));
  INVx1_ASAP7_75t_L         g01760(.A(new_n1996), .Y(new_n2017));
  NOR2xp33_ASAP7_75t_L      g01761(.A(\b[23] ), .B(\b[24] ), .Y(new_n2018));
  INVx1_ASAP7_75t_L         g01762(.A(\b[24] ), .Y(new_n2019));
  NOR2xp33_ASAP7_75t_L      g01763(.A(new_n1995), .B(new_n2019), .Y(new_n2020));
  NOR2xp33_ASAP7_75t_L      g01764(.A(new_n2018), .B(new_n2020), .Y(new_n2021));
  INVx1_ASAP7_75t_L         g01765(.A(new_n2021), .Y(new_n2022));
  O2A1O1Ixp33_ASAP7_75t_L   g01766(.A1(new_n2000), .A2(new_n1999), .B(new_n2017), .C(new_n2022), .Y(new_n2023));
  INVx1_ASAP7_75t_L         g01767(.A(new_n1858), .Y(new_n2024));
  A2O1A1Ixp33_ASAP7_75t_L   g01768(.A1(new_n1860), .A2(new_n2024), .B(new_n2000), .C(new_n2017), .Y(new_n2025));
  NOR2xp33_ASAP7_75t_L      g01769(.A(new_n2021), .B(new_n2025), .Y(new_n2026));
  NOR2xp33_ASAP7_75t_L      g01770(.A(new_n2023), .B(new_n2026), .Y(new_n2027));
  AOI22xp33_ASAP7_75t_L     g01771(.A1(new_n272), .A2(\b[24] ), .B1(new_n269), .B2(new_n2027), .Y(new_n2028));
  NAND2xp33_ASAP7_75t_L     g01772(.A(new_n2016), .B(new_n2028), .Y(new_n2029));
  AOI21xp33_ASAP7_75t_L     g01773(.A1(new_n291), .A2(\b[22] ), .B(new_n2029), .Y(new_n2030));
  NAND2xp33_ASAP7_75t_L     g01774(.A(\a[2] ), .B(new_n2030), .Y(new_n2031));
  A2O1A1Ixp33_ASAP7_75t_L   g01775(.A1(\b[22] ), .A2(new_n291), .B(new_n2029), .C(new_n265), .Y(new_n2032));
  NAND2xp33_ASAP7_75t_L     g01776(.A(new_n2032), .B(new_n2031), .Y(new_n2033));
  A2O1A1O1Ixp25_ASAP7_75t_L g01777(.A1(new_n1852), .A2(new_n1854), .B(new_n1873), .C(new_n1984), .D(new_n1987), .Y(new_n2034));
  NAND2xp33_ASAP7_75t_L     g01778(.A(\b[20] ), .B(new_n334), .Y(new_n2035));
  AOI22xp33_ASAP7_75t_L     g01779(.A1(new_n345), .A2(\b[21] ), .B1(new_n342), .B2(new_n1715), .Y(new_n2036));
  NAND2xp33_ASAP7_75t_L     g01780(.A(new_n2035), .B(new_n2036), .Y(new_n2037));
  AOI211xp5_ASAP7_75t_L     g01781(.A1(\b[19] ), .A2(new_n366), .B(new_n339), .C(new_n2037), .Y(new_n2038));
  AND2x2_ASAP7_75t_L        g01782(.A(new_n2035), .B(new_n2036), .Y(new_n2039));
  O2A1O1Ixp33_ASAP7_75t_L   g01783(.A1(new_n1493), .A2(new_n365), .B(new_n2039), .C(\a[5] ), .Y(new_n2040));
  NOR2xp33_ASAP7_75t_L      g01784(.A(new_n2038), .B(new_n2040), .Y(new_n2041));
  NOR3xp33_ASAP7_75t_L      g01785(.A(new_n1956), .B(new_n1962), .C(new_n1960), .Y(new_n2042));
  NAND2xp33_ASAP7_75t_L     g01786(.A(new_n1809), .B(new_n1883), .Y(new_n2043));
  A2O1A1Ixp33_ASAP7_75t_L   g01787(.A1(new_n1818), .A2(new_n2043), .B(new_n1935), .C(new_n1943), .Y(new_n2044));
  NOR2xp33_ASAP7_75t_L      g01788(.A(new_n631), .B(new_n909), .Y(new_n2045));
  NAND2xp33_ASAP7_75t_L     g01789(.A(\b[11] ), .B(new_n817), .Y(new_n2046));
  OAI221xp5_ASAP7_75t_L     g01790(.A1(new_n912), .A2(new_n763), .B1(new_n911), .B2(new_n775), .C(new_n2046), .Y(new_n2047));
  OR3x1_ASAP7_75t_L         g01791(.A(new_n2047), .B(new_n813), .C(new_n2045), .Y(new_n2048));
  A2O1A1Ixp33_ASAP7_75t_L   g01792(.A1(\b[10] ), .A2(new_n908), .B(new_n2047), .C(new_n813), .Y(new_n2049));
  A2O1A1O1Ixp25_ASAP7_75t_L g01793(.A1(new_n1793), .A2(new_n1736), .B(new_n1796), .C(new_n1928), .D(new_n1929), .Y(new_n2050));
  INVx1_ASAP7_75t_L         g01794(.A(new_n1923), .Y(new_n2051));
  INVx1_ASAP7_75t_L         g01795(.A(new_n1633), .Y(new_n2052));
  NAND2xp33_ASAP7_75t_L     g01796(.A(\b[0] ), .B(new_n1770), .Y(new_n2053));
  NAND4xp25_ASAP7_75t_L     g01797(.A(new_n1767), .B(\a[23] ), .C(new_n2052), .D(new_n2053), .Y(new_n2054));
  INVx1_ASAP7_75t_L         g01798(.A(\a[24] ), .Y(new_n2055));
  NAND2xp33_ASAP7_75t_L     g01799(.A(\a[23] ), .B(new_n2055), .Y(new_n2056));
  NAND2xp33_ASAP7_75t_L     g01800(.A(\a[24] ), .B(new_n1761), .Y(new_n2057));
  AND2x2_ASAP7_75t_L        g01801(.A(new_n2056), .B(new_n2057), .Y(new_n2058));
  NOR2xp33_ASAP7_75t_L      g01802(.A(new_n258), .B(new_n2058), .Y(new_n2059));
  OA31x2_ASAP7_75t_L        g01803(.A1(new_n1921), .A2(new_n1917), .A3(new_n2054), .B1(new_n2059), .Y(new_n2060));
  NOR3xp33_ASAP7_75t_L      g01804(.A(new_n1914), .B(new_n2059), .C(new_n2054), .Y(new_n2061));
  NOR2xp33_ASAP7_75t_L      g01805(.A(new_n278), .B(new_n1758), .Y(new_n2062));
  AOI221xp5_ASAP7_75t_L     g01806(.A1(new_n1766), .A2(\b[3] ), .B1(new_n1764), .B2(new_n1000), .C(new_n2062), .Y(new_n2063));
  OAI211xp5_ASAP7_75t_L     g01807(.A1(new_n276), .A2(new_n1911), .B(new_n2063), .C(\a[23] ), .Y(new_n2064));
  NAND2xp33_ASAP7_75t_L     g01808(.A(\b[3] ), .B(new_n1766), .Y(new_n2065));
  OAI221xp5_ASAP7_75t_L     g01809(.A1(new_n278), .A2(new_n1758), .B1(new_n1771), .B2(new_n303), .C(new_n2065), .Y(new_n2066));
  A2O1A1Ixp33_ASAP7_75t_L   g01810(.A1(\b[1] ), .A2(new_n1910), .B(new_n2066), .C(new_n1761), .Y(new_n2067));
  NAND2xp33_ASAP7_75t_L     g01811(.A(new_n2067), .B(new_n2064), .Y(new_n2068));
  OAI21xp33_ASAP7_75t_L     g01812(.A1(new_n2060), .A2(new_n2061), .B(new_n2068), .Y(new_n2069));
  OAI21xp33_ASAP7_75t_L     g01813(.A1(new_n2054), .A2(new_n1914), .B(new_n2059), .Y(new_n2070));
  OR4x2_ASAP7_75t_L         g01814(.A(new_n2059), .B(new_n2054), .C(new_n1917), .D(new_n1921), .Y(new_n2071));
  AOI211xp5_ASAP7_75t_L     g01815(.A1(\b[1] ), .A2(new_n1910), .B(new_n1761), .C(new_n2066), .Y(new_n2072));
  O2A1O1Ixp33_ASAP7_75t_L   g01816(.A1(new_n276), .A2(new_n1911), .B(new_n2063), .C(\a[23] ), .Y(new_n2073));
  NOR2xp33_ASAP7_75t_L      g01817(.A(new_n2072), .B(new_n2073), .Y(new_n2074));
  NAND3xp33_ASAP7_75t_L     g01818(.A(new_n2074), .B(new_n2071), .C(new_n2070), .Y(new_n2075));
  NAND2xp33_ASAP7_75t_L     g01819(.A(\b[4] ), .B(new_n1548), .Y(new_n2076));
  NAND2xp33_ASAP7_75t_L     g01820(.A(\b[5] ), .B(new_n1410), .Y(new_n2077));
  AOI22xp33_ASAP7_75t_L     g01821(.A1(new_n1406), .A2(\b[6] ), .B1(new_n1404), .B2(new_n389), .Y(new_n2078));
  NAND4xp25_ASAP7_75t_L     g01822(.A(new_n2078), .B(\a[20] ), .C(new_n2076), .D(new_n2077), .Y(new_n2079));
  OAI221xp5_ASAP7_75t_L     g01823(.A1(new_n1412), .A2(new_n382), .B1(new_n1411), .B2(new_n540), .C(new_n2077), .Y(new_n2080));
  A2O1A1Ixp33_ASAP7_75t_L   g01824(.A1(\b[4] ), .A2(new_n1548), .B(new_n2080), .C(new_n1401), .Y(new_n2081));
  NAND4xp25_ASAP7_75t_L     g01825(.A(new_n2081), .B(new_n2075), .C(new_n2069), .D(new_n2079), .Y(new_n2082));
  AOI21xp33_ASAP7_75t_L     g01826(.A1(new_n2071), .A2(new_n2070), .B(new_n2074), .Y(new_n2083));
  NOR3xp33_ASAP7_75t_L      g01827(.A(new_n2068), .B(new_n2061), .C(new_n2060), .Y(new_n2084));
  AOI211xp5_ASAP7_75t_L     g01828(.A1(\b[4] ), .A2(new_n1548), .B(new_n1401), .C(new_n2080), .Y(new_n2085));
  AOI31xp33_ASAP7_75t_L     g01829(.A1(new_n2078), .A2(new_n2077), .A3(new_n2076), .B(\a[20] ), .Y(new_n2086));
  OAI22xp33_ASAP7_75t_L     g01830(.A1(new_n2085), .A2(new_n2086), .B1(new_n2083), .B2(new_n2084), .Y(new_n2087));
  AOI211xp5_ASAP7_75t_L     g01831(.A1(new_n1922), .A2(new_n1918), .B(new_n1907), .C(new_n1905), .Y(new_n2088));
  A2O1A1O1Ixp25_ASAP7_75t_L g01832(.A1(new_n1776), .A2(new_n1786), .B(new_n1784), .C(new_n1900), .D(new_n2088), .Y(new_n2089));
  OAI211xp5_ASAP7_75t_L     g01833(.A1(new_n2051), .A2(new_n2089), .B(new_n2082), .C(new_n2087), .Y(new_n2090));
  NAND2xp33_ASAP7_75t_L     g01834(.A(new_n2082), .B(new_n2087), .Y(new_n2091));
  A2O1A1O1Ixp25_ASAP7_75t_L g01835(.A1(new_n1746), .A2(new_n1791), .B(new_n1925), .C(new_n1920), .D(new_n2051), .Y(new_n2092));
  NAND2xp33_ASAP7_75t_L     g01836(.A(new_n2092), .B(new_n2091), .Y(new_n2093));
  NAND2xp33_ASAP7_75t_L     g01837(.A(\b[7] ), .B(new_n1194), .Y(new_n2094));
  NAND2xp33_ASAP7_75t_L     g01838(.A(\b[8] ), .B(new_n1103), .Y(new_n2095));
  AOI22xp33_ASAP7_75t_L     g01839(.A1(new_n1113), .A2(\b[9] ), .B1(new_n1110), .B2(new_n566), .Y(new_n2096));
  NAND4xp25_ASAP7_75t_L     g01840(.A(new_n2096), .B(\a[17] ), .C(new_n2094), .D(new_n2095), .Y(new_n2097));
  OAI221xp5_ASAP7_75t_L     g01841(.A1(new_n1198), .A2(new_n559), .B1(new_n1197), .B2(new_n978), .C(new_n2095), .Y(new_n2098));
  A2O1A1Ixp33_ASAP7_75t_L   g01842(.A1(\b[7] ), .A2(new_n1194), .B(new_n2098), .C(new_n1107), .Y(new_n2099));
  AOI22xp33_ASAP7_75t_L     g01843(.A1(new_n2097), .A2(new_n2099), .B1(new_n2090), .B2(new_n2093), .Y(new_n2100));
  O2A1O1Ixp33_ASAP7_75t_L   g01844(.A1(new_n1777), .A2(new_n1781), .B(new_n1746), .C(new_n1925), .Y(new_n2101));
  O2A1O1Ixp33_ASAP7_75t_L   g01845(.A1(new_n2101), .A2(new_n2088), .B(new_n1923), .C(new_n2091), .Y(new_n2102));
  AOI211xp5_ASAP7_75t_L     g01846(.A1(new_n2082), .A2(new_n2087), .B(new_n2051), .C(new_n2089), .Y(new_n2103));
  NAND2xp33_ASAP7_75t_L     g01847(.A(new_n2097), .B(new_n2099), .Y(new_n2104));
  NOR3xp33_ASAP7_75t_L      g01848(.A(new_n2104), .B(new_n2103), .C(new_n2102), .Y(new_n2105));
  NOR3xp33_ASAP7_75t_L      g01849(.A(new_n2050), .B(new_n2100), .C(new_n2105), .Y(new_n2106));
  OAI21xp33_ASAP7_75t_L     g01850(.A1(new_n2102), .A2(new_n2103), .B(new_n2104), .Y(new_n2107));
  NAND4xp25_ASAP7_75t_L     g01851(.A(new_n2093), .B(new_n2097), .C(new_n2099), .D(new_n2090), .Y(new_n2108));
  AOI221xp5_ASAP7_75t_L     g01852(.A1(new_n1893), .A2(new_n1928), .B1(new_n2108), .B2(new_n2107), .C(new_n1929), .Y(new_n2109));
  OAI211xp5_ASAP7_75t_L     g01853(.A1(new_n2109), .A2(new_n2106), .B(new_n2049), .C(new_n2048), .Y(new_n2110));
  AOI211xp5_ASAP7_75t_L     g01854(.A1(new_n2048), .A2(new_n2049), .B(new_n2109), .C(new_n2106), .Y(new_n2111));
  INVx1_ASAP7_75t_L         g01855(.A(new_n2111), .Y(new_n2112));
  NAND3xp33_ASAP7_75t_L     g01856(.A(new_n2044), .B(new_n2112), .C(new_n2110), .Y(new_n2113));
  NOR2xp33_ASAP7_75t_L      g01857(.A(new_n1805), .B(new_n1940), .Y(new_n2114));
  A2O1A1O1Ixp25_ASAP7_75t_L g01858(.A1(new_n1817), .A2(new_n1825), .B(new_n2114), .C(new_n1942), .D(new_n1938), .Y(new_n2115));
  NAND2xp33_ASAP7_75t_L     g01859(.A(new_n2049), .B(new_n2048), .Y(new_n2116));
  INVx1_ASAP7_75t_L         g01860(.A(new_n2106), .Y(new_n2117));
  INVx1_ASAP7_75t_L         g01861(.A(new_n2109), .Y(new_n2118));
  AOI21xp33_ASAP7_75t_L     g01862(.A1(new_n2117), .A2(new_n2118), .B(new_n2116), .Y(new_n2119));
  OAI21xp33_ASAP7_75t_L     g01863(.A1(new_n2111), .A2(new_n2119), .B(new_n2115), .Y(new_n2120));
  NAND2xp33_ASAP7_75t_L     g01864(.A(\b[13] ), .B(new_n674), .Y(new_n2121));
  NAND2xp33_ASAP7_75t_L     g01865(.A(\b[14] ), .B(new_n590), .Y(new_n2122));
  AOI22xp33_ASAP7_75t_L     g01866(.A1(new_n600), .A2(\b[15] ), .B1(new_n597), .B2(new_n959), .Y(new_n2123));
  AND4x1_ASAP7_75t_L        g01867(.A(new_n2123), .B(new_n2122), .C(new_n2121), .D(\a[11] ), .Y(new_n2124));
  AOI31xp33_ASAP7_75t_L     g01868(.A1(new_n2123), .A2(new_n2122), .A3(new_n2121), .B(\a[11] ), .Y(new_n2125));
  NOR2xp33_ASAP7_75t_L      g01869(.A(new_n2125), .B(new_n2124), .Y(new_n2126));
  NAND3xp33_ASAP7_75t_L     g01870(.A(new_n2113), .B(new_n2126), .C(new_n2120), .Y(new_n2127));
  NAND2xp33_ASAP7_75t_L     g01871(.A(new_n2120), .B(new_n2113), .Y(new_n2128));
  OAI21xp33_ASAP7_75t_L     g01872(.A1(new_n2124), .A2(new_n2125), .B(new_n2128), .Y(new_n2129));
  NOR3xp33_ASAP7_75t_L      g01873(.A(new_n1951), .B(new_n1944), .C(new_n1939), .Y(new_n2130));
  O2A1O1Ixp33_ASAP7_75t_L   g01874(.A1(new_n1957), .A2(new_n1958), .B(new_n1959), .C(new_n2130), .Y(new_n2131));
  NAND3xp33_ASAP7_75t_L     g01875(.A(new_n2129), .B(new_n2131), .C(new_n2127), .Y(new_n2132));
  AO21x2_ASAP7_75t_L        g01876(.A1(new_n2127), .A2(new_n2129), .B(new_n2131), .Y(new_n2133));
  NAND2xp33_ASAP7_75t_L     g01877(.A(\b[16] ), .B(new_n480), .Y(new_n2134));
  NOR2xp33_ASAP7_75t_L      g01878(.A(new_n1356), .B(new_n667), .Y(new_n2135));
  AOI221xp5_ASAP7_75t_L     g01879(.A1(new_n441), .A2(\b[17] ), .B1(new_n448), .B2(new_n1363), .C(new_n2135), .Y(new_n2136));
  AND3x1_ASAP7_75t_L        g01880(.A(new_n2136), .B(new_n2134), .C(\a[8] ), .Y(new_n2137));
  O2A1O1Ixp33_ASAP7_75t_L   g01881(.A1(new_n1051), .A2(new_n481), .B(new_n2136), .C(\a[8] ), .Y(new_n2138));
  OR2x4_ASAP7_75t_L         g01882(.A(new_n2138), .B(new_n2137), .Y(new_n2139));
  AOI21xp33_ASAP7_75t_L     g01883(.A1(new_n2133), .A2(new_n2132), .B(new_n2139), .Y(new_n2140));
  AND3x1_ASAP7_75t_L        g01884(.A(new_n2129), .B(new_n2131), .C(new_n2127), .Y(new_n2141));
  AOI21xp33_ASAP7_75t_L     g01885(.A1(new_n2129), .A2(new_n2127), .B(new_n2131), .Y(new_n2142));
  NOR2xp33_ASAP7_75t_L      g01886(.A(new_n2138), .B(new_n2137), .Y(new_n2143));
  NOR3xp33_ASAP7_75t_L      g01887(.A(new_n2141), .B(new_n2142), .C(new_n2143), .Y(new_n2144));
  NOR2xp33_ASAP7_75t_L      g01888(.A(new_n2140), .B(new_n2144), .Y(new_n2145));
  A2O1A1Ixp33_ASAP7_75t_L   g01889(.A1(new_n1966), .A2(new_n1968), .B(new_n2042), .C(new_n2145), .Y(new_n2146));
  O2A1O1Ixp33_ASAP7_75t_L   g01890(.A1(new_n1834), .A2(new_n1836), .B(new_n1966), .C(new_n2042), .Y(new_n2147));
  OAI21xp33_ASAP7_75t_L     g01891(.A1(new_n2142), .A2(new_n2141), .B(new_n2143), .Y(new_n2148));
  NAND3xp33_ASAP7_75t_L     g01892(.A(new_n2139), .B(new_n2133), .C(new_n2132), .Y(new_n2149));
  NAND2xp33_ASAP7_75t_L     g01893(.A(new_n2148), .B(new_n2149), .Y(new_n2150));
  NAND2xp33_ASAP7_75t_L     g01894(.A(new_n2150), .B(new_n2147), .Y(new_n2151));
  AOI21xp33_ASAP7_75t_L     g01895(.A1(new_n2146), .A2(new_n2151), .B(new_n2041), .Y(new_n2152));
  OAI211xp5_ASAP7_75t_L     g01896(.A1(new_n1493), .A2(new_n365), .B(new_n2039), .C(\a[5] ), .Y(new_n2153));
  A2O1A1Ixp33_ASAP7_75t_L   g01897(.A1(\b[19] ), .A2(new_n366), .B(new_n2037), .C(new_n339), .Y(new_n2154));
  NAND2xp33_ASAP7_75t_L     g01898(.A(new_n2154), .B(new_n2153), .Y(new_n2155));
  INVx1_ASAP7_75t_L         g01899(.A(new_n2042), .Y(new_n2156));
  O2A1O1Ixp33_ASAP7_75t_L   g01900(.A1(new_n1981), .A2(new_n1969), .B(new_n2156), .C(new_n2150), .Y(new_n2157));
  A2O1A1Ixp33_ASAP7_75t_L   g01901(.A1(new_n1961), .A2(new_n1965), .B(new_n1981), .C(new_n2156), .Y(new_n2158));
  NOR2xp33_ASAP7_75t_L      g01902(.A(new_n2145), .B(new_n2158), .Y(new_n2159));
  NOR3xp33_ASAP7_75t_L      g01903(.A(new_n2159), .B(new_n2157), .C(new_n2155), .Y(new_n2160));
  NOR2xp33_ASAP7_75t_L      g01904(.A(new_n2152), .B(new_n2160), .Y(new_n2161));
  NOR2xp33_ASAP7_75t_L      g01905(.A(new_n2161), .B(new_n2034), .Y(new_n2162));
  OAI21xp33_ASAP7_75t_L     g01906(.A1(new_n2157), .A2(new_n2159), .B(new_n2155), .Y(new_n2163));
  NAND3xp33_ASAP7_75t_L     g01907(.A(new_n2146), .B(new_n2151), .C(new_n2041), .Y(new_n2164));
  NAND2xp33_ASAP7_75t_L     g01908(.A(new_n2164), .B(new_n2163), .Y(new_n2165));
  NOR3xp33_ASAP7_75t_L      g01909(.A(new_n2165), .B(new_n2008), .C(new_n1987), .Y(new_n2166));
  NOR3xp33_ASAP7_75t_L      g01910(.A(new_n2166), .B(new_n2162), .C(new_n2033), .Y(new_n2167));
  NAND2xp33_ASAP7_75t_L     g01911(.A(new_n1978), .B(new_n1982), .Y(new_n2168));
  A2O1A1Ixp33_ASAP7_75t_L   g01912(.A1(new_n1976), .A2(new_n2168), .B(new_n2008), .C(new_n2165), .Y(new_n2169));
  NAND2xp33_ASAP7_75t_L     g01913(.A(new_n2161), .B(new_n2034), .Y(new_n2170));
  AOI22xp33_ASAP7_75t_L     g01914(.A1(new_n2031), .A2(new_n2032), .B1(new_n2169), .B2(new_n2170), .Y(new_n2171));
  NOR2xp33_ASAP7_75t_L      g01915(.A(new_n2171), .B(new_n2167), .Y(new_n2172));
  O2A1O1Ixp33_ASAP7_75t_L   g01916(.A1(new_n2014), .A2(new_n2005), .B(new_n2015), .C(new_n2172), .Y(new_n2173));
  NOR2xp33_ASAP7_75t_L      g01917(.A(new_n2005), .B(new_n2014), .Y(new_n2174));
  A2O1A1O1Ixp25_ASAP7_75t_L g01918(.A1(new_n1871), .A2(new_n1722), .B(new_n1870), .C(new_n2011), .D(new_n2174), .Y(new_n2175));
  AND2x2_ASAP7_75t_L        g01919(.A(new_n2172), .B(new_n2175), .Y(new_n2176));
  NOR2xp33_ASAP7_75t_L      g01920(.A(new_n2173), .B(new_n2176), .Y(\f[24] ));
  NAND3xp33_ASAP7_75t_L     g01921(.A(new_n2169), .B(new_n2170), .C(new_n2033), .Y(new_n2178));
  NOR2xp33_ASAP7_75t_L      g01922(.A(\b[24] ), .B(\b[25] ), .Y(new_n2179));
  INVx1_ASAP7_75t_L         g01923(.A(\b[25] ), .Y(new_n2180));
  NOR2xp33_ASAP7_75t_L      g01924(.A(new_n2019), .B(new_n2180), .Y(new_n2181));
  NOR2xp33_ASAP7_75t_L      g01925(.A(new_n2179), .B(new_n2181), .Y(new_n2182));
  A2O1A1Ixp33_ASAP7_75t_L   g01926(.A1(new_n2025), .A2(new_n2021), .B(new_n2020), .C(new_n2182), .Y(new_n2183));
  O2A1O1Ixp33_ASAP7_75t_L   g01927(.A1(new_n1856), .A2(new_n1861), .B(new_n2024), .C(new_n2000), .Y(new_n2184));
  O2A1O1Ixp33_ASAP7_75t_L   g01928(.A1(new_n1996), .A2(new_n2184), .B(new_n2021), .C(new_n2020), .Y(new_n2185));
  OAI21xp33_ASAP7_75t_L     g01929(.A1(new_n2179), .A2(new_n2181), .B(new_n2185), .Y(new_n2186));
  NAND2xp33_ASAP7_75t_L     g01930(.A(new_n2183), .B(new_n2186), .Y(new_n2187));
  INVx1_ASAP7_75t_L         g01931(.A(new_n2187), .Y(new_n2188));
  NOR2xp33_ASAP7_75t_L      g01932(.A(new_n2180), .B(new_n632), .Y(new_n2189));
  AOI221xp5_ASAP7_75t_L     g01933(.A1(new_n380), .A2(\b[24] ), .B1(new_n269), .B2(new_n2188), .C(new_n2189), .Y(new_n2190));
  OAI21xp33_ASAP7_75t_L     g01934(.A1(new_n1995), .A2(new_n277), .B(new_n2190), .Y(new_n2191));
  NOR2xp33_ASAP7_75t_L      g01935(.A(new_n265), .B(new_n2191), .Y(new_n2192));
  O2A1O1Ixp33_ASAP7_75t_L   g01936(.A1(new_n1995), .A2(new_n277), .B(new_n2190), .C(\a[2] ), .Y(new_n2193));
  NOR2xp33_ASAP7_75t_L      g01937(.A(new_n2193), .B(new_n2192), .Y(new_n2194));
  NOR3xp33_ASAP7_75t_L      g01938(.A(new_n2159), .B(new_n2157), .C(new_n2041), .Y(new_n2195));
  INVx1_ASAP7_75t_L         g01939(.A(new_n2195), .Y(new_n2196));
  OAI211xp5_ASAP7_75t_L     g01940(.A1(new_n2086), .A2(new_n2085), .B(new_n2075), .C(new_n2069), .Y(new_n2197));
  NOR4xp25_ASAP7_75t_L      g01941(.A(new_n2085), .B(new_n2084), .C(new_n2083), .D(new_n2086), .Y(new_n2198));
  AOI22xp33_ASAP7_75t_L     g01942(.A1(new_n2075), .A2(new_n2069), .B1(new_n2081), .B2(new_n2079), .Y(new_n2199));
  OAI22xp33_ASAP7_75t_L     g01943(.A1(new_n2089), .A2(new_n2051), .B1(new_n2198), .B2(new_n2199), .Y(new_n2200));
  NAND2xp33_ASAP7_75t_L     g01944(.A(\b[6] ), .B(new_n1410), .Y(new_n2201));
  AOI32xp33_ASAP7_75t_L     g01945(.A1(new_n424), .A2(new_n426), .A3(new_n1404), .B1(new_n1406), .B2(\b[7] ), .Y(new_n2202));
  NAND2xp33_ASAP7_75t_L     g01946(.A(new_n2201), .B(new_n2202), .Y(new_n2203));
  AOI211xp5_ASAP7_75t_L     g01947(.A1(\b[5] ), .A2(new_n1548), .B(new_n1401), .C(new_n2203), .Y(new_n2204));
  INVx1_ASAP7_75t_L         g01948(.A(new_n2204), .Y(new_n2205));
  A2O1A1Ixp33_ASAP7_75t_L   g01949(.A1(\b[5] ), .A2(new_n1548), .B(new_n2203), .C(new_n1401), .Y(new_n2206));
  NOR3xp33_ASAP7_75t_L      g01950(.A(new_n2054), .B(new_n1921), .C(new_n1917), .Y(new_n2207));
  MAJIxp5_ASAP7_75t_L       g01951(.A(new_n2068), .B(new_n2059), .C(new_n2207), .Y(new_n2208));
  NAND2xp33_ASAP7_75t_L     g01952(.A(\b[2] ), .B(new_n1910), .Y(new_n2209));
  NOR2xp33_ASAP7_75t_L      g01953(.A(new_n299), .B(new_n1758), .Y(new_n2210));
  INVx1_ASAP7_75t_L         g01954(.A(new_n2210), .Y(new_n2211));
  OAI32xp33_ASAP7_75t_L     g01955(.A1(new_n325), .A2(new_n327), .A3(new_n1771), .B1(new_n323), .B2(new_n1772), .Y(new_n2212));
  INVx1_ASAP7_75t_L         g01956(.A(new_n2212), .Y(new_n2213));
  NAND4xp25_ASAP7_75t_L     g01957(.A(new_n2213), .B(\a[23] ), .C(new_n2209), .D(new_n2211), .Y(new_n2214));
  INVx1_ASAP7_75t_L         g01958(.A(new_n2209), .Y(new_n2215));
  OAI31xp33_ASAP7_75t_L     g01959(.A1(new_n2215), .A2(new_n2212), .A3(new_n2210), .B(new_n1761), .Y(new_n2216));
  NAND2xp33_ASAP7_75t_L     g01960(.A(\a[26] ), .B(new_n2059), .Y(new_n2217));
  XNOR2x2_ASAP7_75t_L       g01961(.A(\a[25] ), .B(\a[24] ), .Y(new_n2218));
  INVx1_ASAP7_75t_L         g01962(.A(new_n2218), .Y(new_n2219));
  NAND2xp33_ASAP7_75t_L     g01963(.A(new_n2219), .B(new_n2058), .Y(new_n2220));
  INVx1_ASAP7_75t_L         g01964(.A(\a[25] ), .Y(new_n2221));
  NAND2xp33_ASAP7_75t_L     g01965(.A(\a[26] ), .B(new_n2221), .Y(new_n2222));
  INVx1_ASAP7_75t_L         g01966(.A(\a[26] ), .Y(new_n2223));
  NAND2xp33_ASAP7_75t_L     g01967(.A(\a[25] ), .B(new_n2223), .Y(new_n2224));
  AND2x2_ASAP7_75t_L        g01968(.A(new_n2222), .B(new_n2224), .Y(new_n2225));
  NOR2xp33_ASAP7_75t_L      g01969(.A(new_n2058), .B(new_n2225), .Y(new_n2226));
  NAND2xp33_ASAP7_75t_L     g01970(.A(new_n2224), .B(new_n2222), .Y(new_n2227));
  NOR2xp33_ASAP7_75t_L      g01971(.A(new_n2227), .B(new_n2058), .Y(new_n2228));
  AOI22xp33_ASAP7_75t_L     g01972(.A1(new_n2228), .A2(\b[1] ), .B1(new_n271), .B2(new_n2226), .Y(new_n2229));
  O2A1O1Ixp33_ASAP7_75t_L   g01973(.A1(new_n2220), .A2(new_n258), .B(new_n2229), .C(new_n2217), .Y(new_n2230));
  NAND2xp33_ASAP7_75t_L     g01974(.A(new_n2057), .B(new_n2056), .Y(new_n2231));
  NOR2xp33_ASAP7_75t_L      g01975(.A(new_n2218), .B(new_n2231), .Y(new_n2232));
  NAND2xp33_ASAP7_75t_L     g01976(.A(new_n2227), .B(new_n2231), .Y(new_n2233));
  NAND2xp33_ASAP7_75t_L     g01977(.A(new_n2231), .B(new_n2225), .Y(new_n2234));
  OAI22xp33_ASAP7_75t_L     g01978(.A1(new_n2234), .A2(new_n276), .B1(new_n270), .B2(new_n2233), .Y(new_n2235));
  A2O1A1O1Ixp25_ASAP7_75t_L g01979(.A1(new_n2231), .A2(\a[26] ), .B(new_n2232), .C(\b[0] ), .D(new_n2235), .Y(new_n2236));
  NOR2xp33_ASAP7_75t_L      g01980(.A(new_n2236), .B(new_n2230), .Y(new_n2237));
  NAND3xp33_ASAP7_75t_L     g01981(.A(new_n2214), .B(new_n2237), .C(new_n2216), .Y(new_n2238));
  NOR4xp25_ASAP7_75t_L      g01982(.A(new_n2215), .B(new_n2212), .C(new_n1761), .D(new_n2210), .Y(new_n2239));
  AOI31xp33_ASAP7_75t_L     g01983(.A1(new_n2213), .A2(new_n2211), .A3(new_n2209), .B(\a[23] ), .Y(new_n2240));
  OR2x4_ASAP7_75t_L         g01984(.A(new_n2236), .B(new_n2230), .Y(new_n2241));
  OAI21xp33_ASAP7_75t_L     g01985(.A1(new_n2239), .A2(new_n2240), .B(new_n2241), .Y(new_n2242));
  AOI21xp33_ASAP7_75t_L     g01986(.A1(new_n2242), .A2(new_n2238), .B(new_n2208), .Y(new_n2243));
  NAND2xp33_ASAP7_75t_L     g01987(.A(new_n2059), .B(new_n2207), .Y(new_n2244));
  A2O1A1Ixp33_ASAP7_75t_L   g01988(.A1(new_n2071), .A2(new_n2070), .B(new_n2074), .C(new_n2244), .Y(new_n2245));
  NAND2xp33_ASAP7_75t_L     g01989(.A(new_n2238), .B(new_n2242), .Y(new_n2246));
  NOR2xp33_ASAP7_75t_L      g01990(.A(new_n2245), .B(new_n2246), .Y(new_n2247));
  AOI211xp5_ASAP7_75t_L     g01991(.A1(new_n2205), .A2(new_n2206), .B(new_n2243), .C(new_n2247), .Y(new_n2248));
  INVx1_ASAP7_75t_L         g01992(.A(new_n2206), .Y(new_n2249));
  INVx1_ASAP7_75t_L         g01993(.A(new_n2238), .Y(new_n2250));
  AOI21xp33_ASAP7_75t_L     g01994(.A1(new_n2214), .A2(new_n2216), .B(new_n2237), .Y(new_n2251));
  OAI21xp33_ASAP7_75t_L     g01995(.A1(new_n2250), .A2(new_n2251), .B(new_n2245), .Y(new_n2252));
  NAND3xp33_ASAP7_75t_L     g01996(.A(new_n2208), .B(new_n2238), .C(new_n2242), .Y(new_n2253));
  AOI211xp5_ASAP7_75t_L     g01997(.A1(new_n2253), .A2(new_n2252), .B(new_n2204), .C(new_n2249), .Y(new_n2254));
  AOI211xp5_ASAP7_75t_L     g01998(.A1(new_n2200), .A2(new_n2197), .B(new_n2248), .C(new_n2254), .Y(new_n2255));
  A2O1A1Ixp33_ASAP7_75t_L   g01999(.A1(new_n2087), .A2(new_n2082), .B(new_n2092), .C(new_n2197), .Y(new_n2256));
  OAI211xp5_ASAP7_75t_L     g02000(.A1(new_n2204), .A2(new_n2249), .B(new_n2252), .C(new_n2253), .Y(new_n2257));
  OAI211xp5_ASAP7_75t_L     g02001(.A1(new_n2243), .A2(new_n2247), .B(new_n2206), .C(new_n2205), .Y(new_n2258));
  AOI21xp33_ASAP7_75t_L     g02002(.A1(new_n2258), .A2(new_n2257), .B(new_n2256), .Y(new_n2259));
  NOR2xp33_ASAP7_75t_L      g02003(.A(new_n503), .B(new_n1195), .Y(new_n2260));
  NAND2xp33_ASAP7_75t_L     g02004(.A(\b[9] ), .B(new_n1103), .Y(new_n2261));
  NAND2xp33_ASAP7_75t_L     g02005(.A(\b[10] ), .B(new_n1113), .Y(new_n2262));
  OAI311xp33_ASAP7_75t_L    g02006(.A1(new_n639), .A2(new_n851), .A3(new_n1197), .B1(new_n2262), .C1(new_n2261), .Y(new_n2263));
  OR3x1_ASAP7_75t_L         g02007(.A(new_n2263), .B(new_n1107), .C(new_n2260), .Y(new_n2264));
  A2O1A1Ixp33_ASAP7_75t_L   g02008(.A1(\b[8] ), .A2(new_n1194), .B(new_n2263), .C(new_n1107), .Y(new_n2265));
  NAND2xp33_ASAP7_75t_L     g02009(.A(new_n2265), .B(new_n2264), .Y(new_n2266));
  NOR3xp33_ASAP7_75t_L      g02010(.A(new_n2259), .B(new_n2255), .C(new_n2266), .Y(new_n2267));
  NAND3xp33_ASAP7_75t_L     g02011(.A(new_n2256), .B(new_n2257), .C(new_n2258), .Y(new_n2268));
  OAI211xp5_ASAP7_75t_L     g02012(.A1(new_n2254), .A2(new_n2248), .B(new_n2200), .C(new_n2197), .Y(new_n2269));
  AND2x2_ASAP7_75t_L        g02013(.A(new_n2265), .B(new_n2264), .Y(new_n2270));
  AOI21xp33_ASAP7_75t_L     g02014(.A1(new_n2268), .A2(new_n2269), .B(new_n2270), .Y(new_n2271));
  NOR2xp33_ASAP7_75t_L      g02015(.A(new_n2271), .B(new_n2267), .Y(new_n2272));
  A2O1A1O1Ixp25_ASAP7_75t_L g02016(.A1(new_n1928), .A2(new_n1893), .B(new_n1929), .C(new_n2108), .D(new_n2100), .Y(new_n2273));
  NAND2xp33_ASAP7_75t_L     g02017(.A(new_n2273), .B(new_n2272), .Y(new_n2274));
  NAND3xp33_ASAP7_75t_L     g02018(.A(new_n2268), .B(new_n2270), .C(new_n2269), .Y(new_n2275));
  OAI21xp33_ASAP7_75t_L     g02019(.A1(new_n2255), .A2(new_n2259), .B(new_n2266), .Y(new_n2276));
  AOI21xp33_ASAP7_75t_L     g02020(.A1(new_n2276), .A2(new_n2275), .B(new_n2273), .Y(new_n2277));
  INVx1_ASAP7_75t_L         g02021(.A(new_n2277), .Y(new_n2278));
  NOR2xp33_ASAP7_75t_L      g02022(.A(new_n695), .B(new_n909), .Y(new_n2279));
  INVx1_ASAP7_75t_L         g02023(.A(new_n2279), .Y(new_n2280));
  NAND2xp33_ASAP7_75t_L     g02024(.A(\b[12] ), .B(new_n817), .Y(new_n2281));
  AOI22xp33_ASAP7_75t_L     g02025(.A1(new_n826), .A2(\b[13] ), .B1(new_n823), .B2(new_n800), .Y(new_n2282));
  AND4x1_ASAP7_75t_L        g02026(.A(new_n2282), .B(new_n2281), .C(new_n2280), .D(\a[14] ), .Y(new_n2283));
  AOI31xp33_ASAP7_75t_L     g02027(.A1(new_n2282), .A2(new_n2281), .A3(new_n2280), .B(\a[14] ), .Y(new_n2284));
  OR2x4_ASAP7_75t_L         g02028(.A(new_n2284), .B(new_n2283), .Y(new_n2285));
  AOI21xp33_ASAP7_75t_L     g02029(.A1(new_n2278), .A2(new_n2274), .B(new_n2285), .Y(new_n2286));
  NAND2xp33_ASAP7_75t_L     g02030(.A(new_n2276), .B(new_n2275), .Y(new_n2287));
  OAI21xp33_ASAP7_75t_L     g02031(.A1(new_n2105), .A2(new_n2050), .B(new_n2107), .Y(new_n2288));
  NOR2xp33_ASAP7_75t_L      g02032(.A(new_n2288), .B(new_n2287), .Y(new_n2289));
  NOR2xp33_ASAP7_75t_L      g02033(.A(new_n2284), .B(new_n2283), .Y(new_n2290));
  NOR3xp33_ASAP7_75t_L      g02034(.A(new_n2289), .B(new_n2277), .C(new_n2290), .Y(new_n2291));
  A2O1A1O1Ixp25_ASAP7_75t_L g02035(.A1(new_n1942), .A2(new_n1941), .B(new_n1938), .C(new_n2110), .D(new_n2111), .Y(new_n2292));
  OR3x1_ASAP7_75t_L         g02036(.A(new_n2292), .B(new_n2286), .C(new_n2291), .Y(new_n2293));
  OAI21xp33_ASAP7_75t_L     g02037(.A1(new_n2291), .A2(new_n2286), .B(new_n2292), .Y(new_n2294));
  NAND2xp33_ASAP7_75t_L     g02038(.A(\b[14] ), .B(new_n674), .Y(new_n2295));
  NAND2xp33_ASAP7_75t_L     g02039(.A(\b[15] ), .B(new_n590), .Y(new_n2296));
  AOI22xp33_ASAP7_75t_L     g02040(.A1(new_n600), .A2(\b[16] ), .B1(new_n597), .B2(new_n1058), .Y(new_n2297));
  AND4x1_ASAP7_75t_L        g02041(.A(new_n2297), .B(new_n2296), .C(new_n2295), .D(\a[11] ), .Y(new_n2298));
  AOI31xp33_ASAP7_75t_L     g02042(.A1(new_n2297), .A2(new_n2296), .A3(new_n2295), .B(\a[11] ), .Y(new_n2299));
  NOR2xp33_ASAP7_75t_L      g02043(.A(new_n2299), .B(new_n2298), .Y(new_n2300));
  NAND3xp33_ASAP7_75t_L     g02044(.A(new_n2293), .B(new_n2294), .C(new_n2300), .Y(new_n2301));
  NOR3xp33_ASAP7_75t_L      g02045(.A(new_n2292), .B(new_n2286), .C(new_n2291), .Y(new_n2302));
  OA21x2_ASAP7_75t_L        g02046(.A1(new_n2291), .A2(new_n2286), .B(new_n2292), .Y(new_n2303));
  OR2x4_ASAP7_75t_L         g02047(.A(new_n2299), .B(new_n2298), .Y(new_n2304));
  OAI21xp33_ASAP7_75t_L     g02048(.A1(new_n2302), .A2(new_n2303), .B(new_n2304), .Y(new_n2305));
  AND2x2_ASAP7_75t_L        g02049(.A(new_n2305), .B(new_n2301), .Y(new_n2306));
  MAJx2_ASAP7_75t_L         g02050(.A(new_n2131), .B(new_n2126), .C(new_n2128), .Y(new_n2307));
  NAND2xp33_ASAP7_75t_L     g02051(.A(new_n2306), .B(new_n2307), .Y(new_n2308));
  NAND2xp33_ASAP7_75t_L     g02052(.A(new_n2305), .B(new_n2301), .Y(new_n2309));
  MAJIxp5_ASAP7_75t_L       g02053(.A(new_n2131), .B(new_n2128), .C(new_n2126), .Y(new_n2310));
  NAND2xp33_ASAP7_75t_L     g02054(.A(new_n2310), .B(new_n2309), .Y(new_n2311));
  AOI22xp33_ASAP7_75t_L     g02055(.A1(new_n451), .A2(\b[19] ), .B1(new_n448), .B2(new_n1499), .Y(new_n2312));
  OAI221xp5_ASAP7_75t_L     g02056(.A1(new_n529), .A2(new_n1356), .B1(new_n1244), .B2(new_n481), .C(new_n2312), .Y(new_n2313));
  XNOR2x2_ASAP7_75t_L       g02057(.A(\a[8] ), .B(new_n2313), .Y(new_n2314));
  AND3x1_ASAP7_75t_L        g02058(.A(new_n2314), .B(new_n2308), .C(new_n2311), .Y(new_n2315));
  AOI21xp33_ASAP7_75t_L     g02059(.A1(new_n2308), .A2(new_n2311), .B(new_n2314), .Y(new_n2316));
  A2O1A1O1Ixp25_ASAP7_75t_L g02060(.A1(new_n1966), .A2(new_n1968), .B(new_n2042), .C(new_n2148), .D(new_n2144), .Y(new_n2317));
  OA21x2_ASAP7_75t_L        g02061(.A1(new_n2316), .A2(new_n2315), .B(new_n2317), .Y(new_n2318));
  NOR3xp33_ASAP7_75t_L      g02062(.A(new_n2315), .B(new_n2317), .C(new_n2316), .Y(new_n2319));
  NAND2xp33_ASAP7_75t_L     g02063(.A(\b[21] ), .B(new_n334), .Y(new_n2320));
  OAI221xp5_ASAP7_75t_L     g02064(.A1(new_n368), .A2(new_n1857), .B1(new_n367), .B2(new_n1863), .C(new_n2320), .Y(new_n2321));
  INVx1_ASAP7_75t_L         g02065(.A(new_n2321), .Y(new_n2322));
  OAI211xp5_ASAP7_75t_L     g02066(.A1(new_n1594), .A2(new_n365), .B(new_n2322), .C(\a[5] ), .Y(new_n2323));
  A2O1A1Ixp33_ASAP7_75t_L   g02067(.A1(\b[20] ), .A2(new_n366), .B(new_n2321), .C(new_n339), .Y(new_n2324));
  NAND2xp33_ASAP7_75t_L     g02068(.A(new_n2324), .B(new_n2323), .Y(new_n2325));
  OAI21xp33_ASAP7_75t_L     g02069(.A1(new_n2319), .A2(new_n2318), .B(new_n2325), .Y(new_n2326));
  OR3x1_ASAP7_75t_L         g02070(.A(new_n2318), .B(new_n2325), .C(new_n2319), .Y(new_n2327));
  NAND2xp33_ASAP7_75t_L     g02071(.A(new_n2326), .B(new_n2327), .Y(new_n2328));
  O2A1O1Ixp33_ASAP7_75t_L   g02072(.A1(new_n2034), .A2(new_n2161), .B(new_n2196), .C(new_n2328), .Y(new_n2329));
  OA21x2_ASAP7_75t_L        g02073(.A1(new_n2319), .A2(new_n2318), .B(new_n2325), .Y(new_n2330));
  NOR3xp33_ASAP7_75t_L      g02074(.A(new_n2318), .B(new_n2325), .C(new_n2319), .Y(new_n2331));
  NOR2xp33_ASAP7_75t_L      g02075(.A(new_n2331), .B(new_n2330), .Y(new_n2332));
  NOR3xp33_ASAP7_75t_L      g02076(.A(new_n2162), .B(new_n2332), .C(new_n2195), .Y(new_n2333));
  NOR3xp33_ASAP7_75t_L      g02077(.A(new_n2333), .B(new_n2329), .C(new_n2194), .Y(new_n2334));
  XNOR2x2_ASAP7_75t_L       g02078(.A(new_n265), .B(new_n2191), .Y(new_n2335));
  INVx1_ASAP7_75t_L         g02079(.A(new_n2034), .Y(new_n2336));
  A2O1A1Ixp33_ASAP7_75t_L   g02080(.A1(new_n2336), .A2(new_n2165), .B(new_n2195), .C(new_n2332), .Y(new_n2337));
  O2A1O1Ixp33_ASAP7_75t_L   g02081(.A1(new_n1987), .A2(new_n2008), .B(new_n2165), .C(new_n2195), .Y(new_n2338));
  NAND2xp33_ASAP7_75t_L     g02082(.A(new_n2328), .B(new_n2338), .Y(new_n2339));
  AOI21xp33_ASAP7_75t_L     g02083(.A1(new_n2339), .A2(new_n2337), .B(new_n2335), .Y(new_n2340));
  NOR2xp33_ASAP7_75t_L      g02084(.A(new_n2340), .B(new_n2334), .Y(new_n2341));
  INVx1_ASAP7_75t_L         g02085(.A(new_n2341), .Y(new_n2342));
  O2A1O1Ixp33_ASAP7_75t_L   g02086(.A1(new_n2172), .A2(new_n2175), .B(new_n2178), .C(new_n2342), .Y(new_n2343));
  OAI21xp33_ASAP7_75t_L     g02087(.A1(new_n2172), .A2(new_n2175), .B(new_n2178), .Y(new_n2344));
  NOR2xp33_ASAP7_75t_L      g02088(.A(new_n2341), .B(new_n2344), .Y(new_n2345));
  NOR2xp33_ASAP7_75t_L      g02089(.A(new_n2345), .B(new_n2343), .Y(\f[25] ));
  INVx1_ASAP7_75t_L         g02090(.A(new_n2178), .Y(new_n2347));
  O2A1O1Ixp33_ASAP7_75t_L   g02091(.A1(new_n2347), .A2(new_n2173), .B(new_n2341), .C(new_n2334), .Y(new_n2348));
  A2O1A1Ixp33_ASAP7_75t_L   g02092(.A1(new_n2169), .A2(new_n2196), .B(new_n2331), .C(new_n2326), .Y(new_n2349));
  NOR3xp33_ASAP7_75t_L      g02093(.A(new_n2303), .B(new_n2300), .C(new_n2302), .Y(new_n2350));
  INVx1_ASAP7_75t_L         g02094(.A(new_n2350), .Y(new_n2351));
  NAND2xp33_ASAP7_75t_L     g02095(.A(\b[15] ), .B(new_n674), .Y(new_n2352));
  NAND2xp33_ASAP7_75t_L     g02096(.A(\b[16] ), .B(new_n590), .Y(new_n2353));
  AOI32xp33_ASAP7_75t_L     g02097(.A1(new_n1250), .A2(new_n1247), .A3(new_n597), .B1(new_n600), .B2(\b[17] ), .Y(new_n2354));
  NAND4xp25_ASAP7_75t_L     g02098(.A(new_n2354), .B(\a[11] ), .C(new_n2352), .D(new_n2353), .Y(new_n2355));
  AOI31xp33_ASAP7_75t_L     g02099(.A1(new_n2354), .A2(new_n2353), .A3(new_n2352), .B(\a[11] ), .Y(new_n2356));
  INVx1_ASAP7_75t_L         g02100(.A(new_n2356), .Y(new_n2357));
  NAND2xp33_ASAP7_75t_L     g02101(.A(new_n2355), .B(new_n2357), .Y(new_n2358));
  NAND3xp33_ASAP7_75t_L     g02102(.A(new_n2278), .B(new_n2285), .C(new_n2274), .Y(new_n2359));
  OAI21xp33_ASAP7_75t_L     g02103(.A1(new_n2286), .A2(new_n2292), .B(new_n2359), .Y(new_n2360));
  NAND3xp33_ASAP7_75t_L     g02104(.A(new_n2268), .B(new_n2269), .C(new_n2266), .Y(new_n2361));
  INVx1_ASAP7_75t_L         g02105(.A(new_n2361), .Y(new_n2362));
  O2A1O1Ixp33_ASAP7_75t_L   g02106(.A1(new_n2267), .A2(new_n2271), .B(new_n2288), .C(new_n2362), .Y(new_n2363));
  NAND2xp33_ASAP7_75t_L     g02107(.A(\b[9] ), .B(new_n1194), .Y(new_n2364));
  NAND2xp33_ASAP7_75t_L     g02108(.A(\b[10] ), .B(new_n1103), .Y(new_n2365));
  AOI32xp33_ASAP7_75t_L     g02109(.A1(new_n700), .A2(new_n698), .A3(new_n1110), .B1(\b[11] ), .B2(new_n1113), .Y(new_n2366));
  NAND4xp25_ASAP7_75t_L     g02110(.A(new_n2366), .B(\a[17] ), .C(new_n2364), .D(new_n2365), .Y(new_n2367));
  NAND2xp33_ASAP7_75t_L     g02111(.A(new_n2365), .B(new_n2366), .Y(new_n2368));
  A2O1A1Ixp33_ASAP7_75t_L   g02112(.A1(\b[9] ), .A2(new_n1194), .B(new_n2368), .C(new_n1107), .Y(new_n2369));
  NAND2xp33_ASAP7_75t_L     g02113(.A(new_n2367), .B(new_n2369), .Y(new_n2370));
  A2O1A1Ixp33_ASAP7_75t_L   g02114(.A1(new_n2200), .A2(new_n2197), .B(new_n2254), .C(new_n2257), .Y(new_n2371));
  NOR2xp33_ASAP7_75t_L      g02115(.A(new_n382), .B(new_n1549), .Y(new_n2372));
  NAND2xp33_ASAP7_75t_L     g02116(.A(\b[7] ), .B(new_n1410), .Y(new_n2373));
  OAI221xp5_ASAP7_75t_L     g02117(.A1(new_n1412), .A2(new_n503), .B1(new_n1411), .B2(new_n509), .C(new_n2373), .Y(new_n2374));
  OR3x1_ASAP7_75t_L         g02118(.A(new_n2374), .B(new_n1401), .C(new_n2372), .Y(new_n2375));
  A2O1A1Ixp33_ASAP7_75t_L   g02119(.A1(\b[6] ), .A2(new_n1548), .B(new_n2374), .C(new_n1401), .Y(new_n2376));
  AOI21xp33_ASAP7_75t_L     g02120(.A1(new_n2216), .A2(new_n2214), .B(new_n2241), .Y(new_n2377));
  INVx1_ASAP7_75t_L         g02121(.A(new_n2377), .Y(new_n2378));
  NAND2xp33_ASAP7_75t_L     g02122(.A(\b[3] ), .B(new_n1910), .Y(new_n2379));
  NAND2xp33_ASAP7_75t_L     g02123(.A(\b[4] ), .B(new_n1770), .Y(new_n2380));
  AOI32xp33_ASAP7_75t_L     g02124(.A1(new_n358), .A2(new_n356), .A3(new_n1764), .B1(\b[5] ), .B2(new_n1766), .Y(new_n2381));
  NAND4xp25_ASAP7_75t_L     g02125(.A(new_n2381), .B(\a[23] ), .C(new_n2379), .D(new_n2380), .Y(new_n2382));
  AOI31xp33_ASAP7_75t_L     g02126(.A1(new_n2381), .A2(new_n2380), .A3(new_n2379), .B(\a[23] ), .Y(new_n2383));
  INVx1_ASAP7_75t_L         g02127(.A(new_n2383), .Y(new_n2384));
  A2O1A1O1Ixp25_ASAP7_75t_L g02128(.A1(new_n2218), .A2(new_n2058), .B(new_n258), .C(new_n2229), .D(new_n2223), .Y(new_n2385));
  NOR3xp33_ASAP7_75t_L      g02129(.A(new_n2225), .B(new_n2219), .C(new_n2231), .Y(new_n2386));
  INVx1_ASAP7_75t_L         g02130(.A(new_n2386), .Y(new_n2387));
  NOR2xp33_ASAP7_75t_L      g02131(.A(new_n258), .B(new_n2387), .Y(new_n2388));
  NAND2xp33_ASAP7_75t_L     g02132(.A(\b[1] ), .B(new_n2232), .Y(new_n2389));
  OAI221xp5_ASAP7_75t_L     g02133(.A1(new_n2233), .A2(new_n283), .B1(new_n278), .B2(new_n2234), .C(new_n2389), .Y(new_n2390));
  NOR3xp33_ASAP7_75t_L      g02134(.A(new_n2385), .B(new_n2388), .C(new_n2390), .Y(new_n2391));
  A2O1A1Ixp33_ASAP7_75t_L   g02135(.A1(\b[0] ), .A2(new_n2386), .B(new_n2390), .C(new_n2385), .Y(new_n2392));
  INVx1_ASAP7_75t_L         g02136(.A(new_n2392), .Y(new_n2393));
  OAI211xp5_ASAP7_75t_L     g02137(.A1(new_n2391), .A2(new_n2393), .B(new_n2384), .C(new_n2382), .Y(new_n2394));
  INVx1_ASAP7_75t_L         g02138(.A(new_n2382), .Y(new_n2395));
  INVx1_ASAP7_75t_L         g02139(.A(new_n2391), .Y(new_n2396));
  OAI211xp5_ASAP7_75t_L     g02140(.A1(new_n2383), .A2(new_n2395), .B(new_n2396), .C(new_n2392), .Y(new_n2397));
  NAND4xp25_ASAP7_75t_L     g02141(.A(new_n2252), .B(new_n2397), .C(new_n2394), .D(new_n2378), .Y(new_n2398));
  NAND2xp33_ASAP7_75t_L     g02142(.A(new_n2397), .B(new_n2394), .Y(new_n2399));
  A2O1A1Ixp33_ASAP7_75t_L   g02143(.A1(new_n2246), .A2(new_n2245), .B(new_n2377), .C(new_n2399), .Y(new_n2400));
  NAND4xp25_ASAP7_75t_L     g02144(.A(new_n2400), .B(new_n2398), .C(new_n2375), .D(new_n2376), .Y(new_n2401));
  AOI22xp33_ASAP7_75t_L     g02145(.A1(new_n2376), .A2(new_n2375), .B1(new_n2398), .B2(new_n2400), .Y(new_n2402));
  INVx1_ASAP7_75t_L         g02146(.A(new_n2402), .Y(new_n2403));
  NAND3xp33_ASAP7_75t_L     g02147(.A(new_n2403), .B(new_n2401), .C(new_n2371), .Y(new_n2404));
  AOI21xp33_ASAP7_75t_L     g02148(.A1(new_n2256), .A2(new_n2258), .B(new_n2248), .Y(new_n2405));
  INVx1_ASAP7_75t_L         g02149(.A(new_n2401), .Y(new_n2406));
  OAI21xp33_ASAP7_75t_L     g02150(.A1(new_n2402), .A2(new_n2406), .B(new_n2405), .Y(new_n2407));
  AOI21xp33_ASAP7_75t_L     g02151(.A1(new_n2404), .A2(new_n2407), .B(new_n2370), .Y(new_n2408));
  NOR3xp33_ASAP7_75t_L      g02152(.A(new_n2405), .B(new_n2406), .C(new_n2402), .Y(new_n2409));
  AOI21xp33_ASAP7_75t_L     g02153(.A1(new_n2403), .A2(new_n2401), .B(new_n2371), .Y(new_n2410));
  AOI211xp5_ASAP7_75t_L     g02154(.A1(new_n2369), .A2(new_n2367), .B(new_n2410), .C(new_n2409), .Y(new_n2411));
  NOR3xp33_ASAP7_75t_L      g02155(.A(new_n2363), .B(new_n2408), .C(new_n2411), .Y(new_n2412));
  A2O1A1Ixp33_ASAP7_75t_L   g02156(.A1(new_n2276), .A2(new_n2275), .B(new_n2273), .C(new_n2361), .Y(new_n2413));
  OAI211xp5_ASAP7_75t_L     g02157(.A1(new_n2410), .A2(new_n2409), .B(new_n2369), .C(new_n2367), .Y(new_n2414));
  NAND3xp33_ASAP7_75t_L     g02158(.A(new_n2370), .B(new_n2404), .C(new_n2407), .Y(new_n2415));
  AOI21xp33_ASAP7_75t_L     g02159(.A1(new_n2415), .A2(new_n2414), .B(new_n2413), .Y(new_n2416));
  NAND2xp33_ASAP7_75t_L     g02160(.A(\b[12] ), .B(new_n908), .Y(new_n2417));
  NAND2xp33_ASAP7_75t_L     g02161(.A(\b[13] ), .B(new_n817), .Y(new_n2418));
  AOI32xp33_ASAP7_75t_L     g02162(.A1(new_n877), .A2(new_n874), .A3(new_n823), .B1(new_n826), .B2(\b[14] ), .Y(new_n2419));
  NAND4xp25_ASAP7_75t_L     g02163(.A(new_n2419), .B(\a[14] ), .C(new_n2417), .D(new_n2418), .Y(new_n2420));
  NAND2xp33_ASAP7_75t_L     g02164(.A(new_n2418), .B(new_n2419), .Y(new_n2421));
  A2O1A1Ixp33_ASAP7_75t_L   g02165(.A1(\b[12] ), .A2(new_n908), .B(new_n2421), .C(new_n813), .Y(new_n2422));
  NAND2xp33_ASAP7_75t_L     g02166(.A(new_n2420), .B(new_n2422), .Y(new_n2423));
  NOR3xp33_ASAP7_75t_L      g02167(.A(new_n2412), .B(new_n2416), .C(new_n2423), .Y(new_n2424));
  NAND3xp33_ASAP7_75t_L     g02168(.A(new_n2413), .B(new_n2414), .C(new_n2415), .Y(new_n2425));
  OAI21xp33_ASAP7_75t_L     g02169(.A1(new_n2408), .A2(new_n2411), .B(new_n2363), .Y(new_n2426));
  AND2x2_ASAP7_75t_L        g02170(.A(new_n2420), .B(new_n2422), .Y(new_n2427));
  AOI21xp33_ASAP7_75t_L     g02171(.A1(new_n2426), .A2(new_n2425), .B(new_n2427), .Y(new_n2428));
  OAI21xp33_ASAP7_75t_L     g02172(.A1(new_n2424), .A2(new_n2428), .B(new_n2360), .Y(new_n2429));
  OAI21xp33_ASAP7_75t_L     g02173(.A1(new_n2277), .A2(new_n2289), .B(new_n2290), .Y(new_n2430));
  A2O1A1O1Ixp25_ASAP7_75t_L g02174(.A1(new_n2110), .A2(new_n2044), .B(new_n2111), .C(new_n2430), .D(new_n2291), .Y(new_n2431));
  NAND3xp33_ASAP7_75t_L     g02175(.A(new_n2427), .B(new_n2426), .C(new_n2425), .Y(new_n2432));
  OAI21xp33_ASAP7_75t_L     g02176(.A1(new_n2416), .A2(new_n2412), .B(new_n2423), .Y(new_n2433));
  NAND3xp33_ASAP7_75t_L     g02177(.A(new_n2431), .B(new_n2432), .C(new_n2433), .Y(new_n2434));
  NAND3xp33_ASAP7_75t_L     g02178(.A(new_n2434), .B(new_n2429), .C(new_n2358), .Y(new_n2435));
  INVx1_ASAP7_75t_L         g02179(.A(new_n2355), .Y(new_n2436));
  NOR2xp33_ASAP7_75t_L      g02180(.A(new_n2356), .B(new_n2436), .Y(new_n2437));
  AOI21xp33_ASAP7_75t_L     g02181(.A1(new_n2433), .A2(new_n2432), .B(new_n2431), .Y(new_n2438));
  NOR3xp33_ASAP7_75t_L      g02182(.A(new_n2360), .B(new_n2428), .C(new_n2424), .Y(new_n2439));
  OAI21xp33_ASAP7_75t_L     g02183(.A1(new_n2438), .A2(new_n2439), .B(new_n2437), .Y(new_n2440));
  NAND2xp33_ASAP7_75t_L     g02184(.A(new_n2435), .B(new_n2440), .Y(new_n2441));
  OAI211xp5_ASAP7_75t_L     g02185(.A1(new_n2306), .A2(new_n2307), .B(new_n2441), .C(new_n2351), .Y(new_n2442));
  NOR3xp33_ASAP7_75t_L      g02186(.A(new_n2439), .B(new_n2437), .C(new_n2438), .Y(new_n2443));
  AOI21xp33_ASAP7_75t_L     g02187(.A1(new_n2434), .A2(new_n2429), .B(new_n2358), .Y(new_n2444));
  NOR2xp33_ASAP7_75t_L      g02188(.A(new_n2444), .B(new_n2443), .Y(new_n2445));
  A2O1A1Ixp33_ASAP7_75t_L   g02189(.A1(new_n2310), .A2(new_n2309), .B(new_n2350), .C(new_n2445), .Y(new_n2446));
  NOR2xp33_ASAP7_75t_L      g02190(.A(new_n1356), .B(new_n481), .Y(new_n2447));
  NAND2xp33_ASAP7_75t_L     g02191(.A(\b[19] ), .B(new_n441), .Y(new_n2448));
  NAND2xp33_ASAP7_75t_L     g02192(.A(\b[20] ), .B(new_n451), .Y(new_n2449));
  OAI311xp33_ASAP7_75t_L    g02193(.A1(new_n1599), .A2(new_n1598), .A3(new_n482), .B1(new_n2449), .C1(new_n2448), .Y(new_n2450));
  OR3x1_ASAP7_75t_L         g02194(.A(new_n2450), .B(new_n445), .C(new_n2447), .Y(new_n2451));
  A2O1A1Ixp33_ASAP7_75t_L   g02195(.A1(\b[18] ), .A2(new_n480), .B(new_n2450), .C(new_n445), .Y(new_n2452));
  AND2x2_ASAP7_75t_L        g02196(.A(new_n2452), .B(new_n2451), .Y(new_n2453));
  NAND3xp33_ASAP7_75t_L     g02197(.A(new_n2446), .B(new_n2442), .C(new_n2453), .Y(new_n2454));
  AOI221xp5_ASAP7_75t_L     g02198(.A1(new_n2440), .A2(new_n2435), .B1(new_n2310), .B2(new_n2309), .C(new_n2350), .Y(new_n2455));
  O2A1O1Ixp33_ASAP7_75t_L   g02199(.A1(new_n2306), .A2(new_n2307), .B(new_n2351), .C(new_n2441), .Y(new_n2456));
  NAND2xp33_ASAP7_75t_L     g02200(.A(new_n2452), .B(new_n2451), .Y(new_n2457));
  OAI21xp33_ASAP7_75t_L     g02201(.A1(new_n2455), .A2(new_n2456), .B(new_n2457), .Y(new_n2458));
  NAND2xp33_ASAP7_75t_L     g02202(.A(new_n2458), .B(new_n2454), .Y(new_n2459));
  XNOR2x2_ASAP7_75t_L       g02203(.A(new_n2310), .B(new_n2309), .Y(new_n2460));
  MAJIxp5_ASAP7_75t_L       g02204(.A(new_n2317), .B(new_n2460), .C(new_n2314), .Y(new_n2461));
  NOR2xp33_ASAP7_75t_L      g02205(.A(new_n2461), .B(new_n2459), .Y(new_n2462));
  AND2x2_ASAP7_75t_L        g02206(.A(new_n2461), .B(new_n2459), .Y(new_n2463));
  NAND2xp33_ASAP7_75t_L     g02207(.A(\b[21] ), .B(new_n366), .Y(new_n2464));
  NAND2xp33_ASAP7_75t_L     g02208(.A(\b[22] ), .B(new_n334), .Y(new_n2465));
  AOI22xp33_ASAP7_75t_L     g02209(.A1(new_n345), .A2(\b[23] ), .B1(new_n342), .B2(new_n2002), .Y(new_n2466));
  NAND4xp25_ASAP7_75t_L     g02210(.A(new_n2466), .B(\a[5] ), .C(new_n2464), .D(new_n2465), .Y(new_n2467));
  NAND2xp33_ASAP7_75t_L     g02211(.A(new_n2465), .B(new_n2466), .Y(new_n2468));
  A2O1A1Ixp33_ASAP7_75t_L   g02212(.A1(\b[21] ), .A2(new_n366), .B(new_n2468), .C(new_n339), .Y(new_n2469));
  NAND2xp33_ASAP7_75t_L     g02213(.A(new_n2467), .B(new_n2469), .Y(new_n2470));
  OR3x1_ASAP7_75t_L         g02214(.A(new_n2470), .B(new_n2462), .C(new_n2463), .Y(new_n2471));
  OAI21xp33_ASAP7_75t_L     g02215(.A1(new_n2462), .A2(new_n2463), .B(new_n2470), .Y(new_n2472));
  NAND3xp33_ASAP7_75t_L     g02216(.A(new_n2349), .B(new_n2471), .C(new_n2472), .Y(new_n2473));
  A2O1A1O1Ixp25_ASAP7_75t_L g02217(.A1(new_n2165), .A2(new_n2336), .B(new_n2195), .C(new_n2332), .D(new_n2330), .Y(new_n2474));
  NAND2xp33_ASAP7_75t_L     g02218(.A(new_n2472), .B(new_n2471), .Y(new_n2475));
  NAND2xp33_ASAP7_75t_L     g02219(.A(new_n2475), .B(new_n2474), .Y(new_n2476));
  INVx1_ASAP7_75t_L         g02220(.A(\b[26] ), .Y(new_n2477));
  INVx1_ASAP7_75t_L         g02221(.A(new_n2020), .Y(new_n2478));
  A2O1A1Ixp33_ASAP7_75t_L   g02222(.A1(new_n1998), .A2(new_n2017), .B(new_n2018), .C(new_n2478), .Y(new_n2479));
  NOR2xp33_ASAP7_75t_L      g02223(.A(\b[25] ), .B(\b[26] ), .Y(new_n2480));
  NOR2xp33_ASAP7_75t_L      g02224(.A(new_n2180), .B(new_n2477), .Y(new_n2481));
  NOR2xp33_ASAP7_75t_L      g02225(.A(new_n2480), .B(new_n2481), .Y(new_n2482));
  A2O1A1Ixp33_ASAP7_75t_L   g02226(.A1(new_n2479), .A2(new_n2182), .B(new_n2181), .C(new_n2482), .Y(new_n2483));
  A2O1A1O1Ixp25_ASAP7_75t_L g02227(.A1(new_n2021), .A2(new_n2025), .B(new_n2020), .C(new_n2182), .D(new_n2181), .Y(new_n2484));
  INVx1_ASAP7_75t_L         g02228(.A(new_n2482), .Y(new_n2485));
  NAND2xp33_ASAP7_75t_L     g02229(.A(new_n2485), .B(new_n2484), .Y(new_n2486));
  NAND2xp33_ASAP7_75t_L     g02230(.A(new_n2486), .B(new_n2483), .Y(new_n2487));
  OAI22xp33_ASAP7_75t_L     g02231(.A1(new_n2487), .A2(new_n292), .B1(new_n2477), .B2(new_n632), .Y(new_n2488));
  AOI221xp5_ASAP7_75t_L     g02232(.A1(\b[24] ), .A2(new_n291), .B1(\b[25] ), .B2(new_n380), .C(new_n2488), .Y(new_n2489));
  XNOR2x2_ASAP7_75t_L       g02233(.A(new_n265), .B(new_n2489), .Y(new_n2490));
  AOI21xp33_ASAP7_75t_L     g02234(.A1(new_n2473), .A2(new_n2476), .B(new_n2490), .Y(new_n2491));
  INVx1_ASAP7_75t_L         g02235(.A(new_n2491), .Y(new_n2492));
  NAND3xp33_ASAP7_75t_L     g02236(.A(new_n2473), .B(new_n2476), .C(new_n2490), .Y(new_n2493));
  NAND2xp33_ASAP7_75t_L     g02237(.A(new_n2493), .B(new_n2492), .Y(new_n2494));
  XOR2x2_ASAP7_75t_L        g02238(.A(new_n2348), .B(new_n2494), .Y(\f[26] ));
  OAI21xp33_ASAP7_75t_L     g02239(.A1(new_n2408), .A2(new_n2363), .B(new_n2415), .Y(new_n2496));
  NOR2xp33_ASAP7_75t_L      g02240(.A(new_n763), .B(new_n1198), .Y(new_n2497));
  AOI221xp5_ASAP7_75t_L     g02241(.A1(new_n1103), .A2(\b[11] ), .B1(new_n1110), .B2(new_n970), .C(new_n2497), .Y(new_n2498));
  OAI211xp5_ASAP7_75t_L     g02242(.A1(new_n631), .A2(new_n1195), .B(new_n2498), .C(\a[17] ), .Y(new_n2499));
  NAND2xp33_ASAP7_75t_L     g02243(.A(\b[11] ), .B(new_n1103), .Y(new_n2500));
  OAI221xp5_ASAP7_75t_L     g02244(.A1(new_n1198), .A2(new_n763), .B1(new_n1197), .B2(new_n775), .C(new_n2500), .Y(new_n2501));
  A2O1A1Ixp33_ASAP7_75t_L   g02245(.A1(\b[10] ), .A2(new_n1194), .B(new_n2501), .C(new_n1107), .Y(new_n2502));
  A2O1A1O1Ixp25_ASAP7_75t_L g02246(.A1(new_n2258), .A2(new_n2256), .B(new_n2248), .C(new_n2401), .D(new_n2402), .Y(new_n2503));
  AOI211xp5_ASAP7_75t_L     g02247(.A1(new_n2382), .A2(new_n2384), .B(new_n2391), .C(new_n2393), .Y(new_n2504));
  INVx1_ASAP7_75t_L         g02248(.A(new_n2059), .Y(new_n2505));
  NAND2xp33_ASAP7_75t_L     g02249(.A(\b[0] ), .B(new_n2232), .Y(new_n2506));
  NAND4xp25_ASAP7_75t_L     g02250(.A(new_n2229), .B(\a[26] ), .C(new_n2505), .D(new_n2506), .Y(new_n2507));
  INVx1_ASAP7_75t_L         g02251(.A(\a[27] ), .Y(new_n2508));
  NAND2xp33_ASAP7_75t_L     g02252(.A(\a[26] ), .B(new_n2508), .Y(new_n2509));
  NAND2xp33_ASAP7_75t_L     g02253(.A(\a[27] ), .B(new_n2223), .Y(new_n2510));
  AND2x2_ASAP7_75t_L        g02254(.A(new_n2509), .B(new_n2510), .Y(new_n2511));
  NOR2xp33_ASAP7_75t_L      g02255(.A(new_n258), .B(new_n2511), .Y(new_n2512));
  OA31x2_ASAP7_75t_L        g02256(.A1(new_n2388), .A2(new_n2390), .A3(new_n2507), .B1(new_n2512), .Y(new_n2513));
  NOR4xp25_ASAP7_75t_L      g02257(.A(new_n2507), .B(new_n2512), .C(new_n2390), .D(new_n2388), .Y(new_n2514));
  NAND2xp33_ASAP7_75t_L     g02258(.A(\b[3] ), .B(new_n2228), .Y(new_n2515));
  OAI221xp5_ASAP7_75t_L     g02259(.A1(new_n278), .A2(new_n2220), .B1(new_n2233), .B2(new_n303), .C(new_n2515), .Y(new_n2516));
  AOI211xp5_ASAP7_75t_L     g02260(.A1(\b[1] ), .A2(new_n2386), .B(new_n2223), .C(new_n2516), .Y(new_n2517));
  NOR2xp33_ASAP7_75t_L      g02261(.A(new_n278), .B(new_n2220), .Y(new_n2518));
  AOI221xp5_ASAP7_75t_L     g02262(.A1(new_n2228), .A2(\b[3] ), .B1(new_n2226), .B2(new_n1000), .C(new_n2518), .Y(new_n2519));
  O2A1O1Ixp33_ASAP7_75t_L   g02263(.A1(new_n276), .A2(new_n2387), .B(new_n2519), .C(\a[26] ), .Y(new_n2520));
  OAI22xp33_ASAP7_75t_L     g02264(.A1(new_n2513), .A2(new_n2514), .B1(new_n2520), .B2(new_n2517), .Y(new_n2521));
  OAI31xp33_ASAP7_75t_L     g02265(.A1(new_n2507), .A2(new_n2390), .A3(new_n2388), .B(new_n2512), .Y(new_n2522));
  OR4x2_ASAP7_75t_L         g02266(.A(new_n2512), .B(new_n2507), .C(new_n2390), .D(new_n2388), .Y(new_n2523));
  NOR2xp33_ASAP7_75t_L      g02267(.A(new_n2517), .B(new_n2520), .Y(new_n2524));
  NAND3xp33_ASAP7_75t_L     g02268(.A(new_n2524), .B(new_n2523), .C(new_n2522), .Y(new_n2525));
  NAND2xp33_ASAP7_75t_L     g02269(.A(\b[5] ), .B(new_n1770), .Y(new_n2526));
  NAND2xp33_ASAP7_75t_L     g02270(.A(\b[6] ), .B(new_n1766), .Y(new_n2527));
  OAI311xp33_ASAP7_75t_L    g02271(.A1(new_n388), .A2(new_n386), .A3(new_n1771), .B1(new_n2527), .C1(new_n2526), .Y(new_n2528));
  AOI211xp5_ASAP7_75t_L     g02272(.A1(\b[4] ), .A2(new_n1910), .B(new_n1761), .C(new_n2528), .Y(new_n2529));
  INVx1_ASAP7_75t_L         g02273(.A(new_n2529), .Y(new_n2530));
  A2O1A1Ixp33_ASAP7_75t_L   g02274(.A1(\b[4] ), .A2(new_n1910), .B(new_n2528), .C(new_n1761), .Y(new_n2531));
  NAND4xp25_ASAP7_75t_L     g02275(.A(new_n2525), .B(new_n2531), .C(new_n2521), .D(new_n2530), .Y(new_n2532));
  OAI211xp5_ASAP7_75t_L     g02276(.A1(new_n276), .A2(new_n2387), .B(new_n2519), .C(\a[26] ), .Y(new_n2533));
  A2O1A1Ixp33_ASAP7_75t_L   g02277(.A1(\b[1] ), .A2(new_n2386), .B(new_n2516), .C(new_n2223), .Y(new_n2534));
  AOI22xp33_ASAP7_75t_L     g02278(.A1(new_n2533), .A2(new_n2534), .B1(new_n2522), .B2(new_n2523), .Y(new_n2535));
  NOR4xp25_ASAP7_75t_L      g02279(.A(new_n2513), .B(new_n2520), .C(new_n2517), .D(new_n2514), .Y(new_n2536));
  INVx1_ASAP7_75t_L         g02280(.A(new_n2531), .Y(new_n2537));
  OAI22xp33_ASAP7_75t_L     g02281(.A1(new_n2535), .A2(new_n2536), .B1(new_n2537), .B2(new_n2529), .Y(new_n2538));
  AOI211xp5_ASAP7_75t_L     g02282(.A1(new_n2396), .A2(new_n2392), .B(new_n2383), .C(new_n2395), .Y(new_n2539));
  A2O1A1O1Ixp25_ASAP7_75t_L g02283(.A1(new_n2238), .A2(new_n2242), .B(new_n2208), .C(new_n2378), .D(new_n2539), .Y(new_n2540));
  OAI211xp5_ASAP7_75t_L     g02284(.A1(new_n2504), .A2(new_n2540), .B(new_n2532), .C(new_n2538), .Y(new_n2541));
  NAND2xp33_ASAP7_75t_L     g02285(.A(new_n2538), .B(new_n2532), .Y(new_n2542));
  A2O1A1O1Ixp25_ASAP7_75t_L g02286(.A1(new_n2245), .A2(new_n2246), .B(new_n2377), .C(new_n2394), .D(new_n2504), .Y(new_n2543));
  NAND2xp33_ASAP7_75t_L     g02287(.A(new_n2543), .B(new_n2542), .Y(new_n2544));
  NOR2xp33_ASAP7_75t_L      g02288(.A(new_n421), .B(new_n1549), .Y(new_n2545));
  INVx1_ASAP7_75t_L         g02289(.A(new_n2545), .Y(new_n2546));
  NAND2xp33_ASAP7_75t_L     g02290(.A(\b[8] ), .B(new_n1410), .Y(new_n2547));
  AOI22xp33_ASAP7_75t_L     g02291(.A1(new_n1406), .A2(\b[9] ), .B1(new_n1404), .B2(new_n566), .Y(new_n2548));
  NAND4xp25_ASAP7_75t_L     g02292(.A(new_n2548), .B(\a[20] ), .C(new_n2546), .D(new_n2547), .Y(new_n2549));
  OAI221xp5_ASAP7_75t_L     g02293(.A1(new_n1412), .A2(new_n559), .B1(new_n1411), .B2(new_n978), .C(new_n2547), .Y(new_n2550));
  A2O1A1Ixp33_ASAP7_75t_L   g02294(.A1(\b[7] ), .A2(new_n1548), .B(new_n2550), .C(new_n1401), .Y(new_n2551));
  AOI22xp33_ASAP7_75t_L     g02295(.A1(new_n2549), .A2(new_n2551), .B1(new_n2544), .B2(new_n2541), .Y(new_n2552));
  NOR2xp33_ASAP7_75t_L      g02296(.A(new_n2543), .B(new_n2542), .Y(new_n2553));
  AOI211xp5_ASAP7_75t_L     g02297(.A1(new_n2532), .A2(new_n2538), .B(new_n2504), .C(new_n2540), .Y(new_n2554));
  NOR3xp33_ASAP7_75t_L      g02298(.A(new_n2550), .B(new_n2545), .C(new_n1401), .Y(new_n2555));
  AOI31xp33_ASAP7_75t_L     g02299(.A1(new_n2548), .A2(new_n2547), .A3(new_n2546), .B(\a[20] ), .Y(new_n2556));
  NOR4xp25_ASAP7_75t_L      g02300(.A(new_n2553), .B(new_n2554), .C(new_n2556), .D(new_n2555), .Y(new_n2557));
  NOR3xp33_ASAP7_75t_L      g02301(.A(new_n2503), .B(new_n2552), .C(new_n2557), .Y(new_n2558));
  OAI22xp33_ASAP7_75t_L     g02302(.A1(new_n2553), .A2(new_n2554), .B1(new_n2556), .B2(new_n2555), .Y(new_n2559));
  NAND4xp25_ASAP7_75t_L     g02303(.A(new_n2541), .B(new_n2544), .C(new_n2551), .D(new_n2549), .Y(new_n2560));
  AOI221xp5_ASAP7_75t_L     g02304(.A1(new_n2371), .A2(new_n2401), .B1(new_n2560), .B2(new_n2559), .C(new_n2402), .Y(new_n2561));
  OAI211xp5_ASAP7_75t_L     g02305(.A1(new_n2561), .A2(new_n2558), .B(new_n2502), .C(new_n2499), .Y(new_n2562));
  AO211x2_ASAP7_75t_L       g02306(.A1(new_n2499), .A2(new_n2502), .B(new_n2561), .C(new_n2558), .Y(new_n2563));
  NAND3xp33_ASAP7_75t_L     g02307(.A(new_n2496), .B(new_n2562), .C(new_n2563), .Y(new_n2564));
  A2O1A1O1Ixp25_ASAP7_75t_L g02308(.A1(new_n2288), .A2(new_n2287), .B(new_n2362), .C(new_n2414), .D(new_n2411), .Y(new_n2565));
  INVx1_ASAP7_75t_L         g02309(.A(new_n2562), .Y(new_n2566));
  AOI211xp5_ASAP7_75t_L     g02310(.A1(new_n2502), .A2(new_n2499), .B(new_n2561), .C(new_n2558), .Y(new_n2567));
  OAI21xp33_ASAP7_75t_L     g02311(.A1(new_n2567), .A2(new_n2566), .B(new_n2565), .Y(new_n2568));
  A2O1A1Ixp33_ASAP7_75t_L   g02312(.A1(new_n771), .A2(new_n791), .B(new_n796), .C(new_n948), .Y(new_n2569));
  A2O1A1Ixp33_ASAP7_75t_L   g02313(.A1(new_n2569), .A2(new_n873), .B(new_n872), .C(new_n954), .Y(new_n2570));
  A2O1A1O1Ixp25_ASAP7_75t_L g02314(.A1(new_n795), .A2(new_n798), .B(new_n794), .C(new_n873), .D(new_n872), .Y(new_n2571));
  NAND2xp33_ASAP7_75t_L     g02315(.A(new_n955), .B(new_n2571), .Y(new_n2572));
  NAND2xp33_ASAP7_75t_L     g02316(.A(new_n2572), .B(new_n2570), .Y(new_n2573));
  NAND2xp33_ASAP7_75t_L     g02317(.A(\b[14] ), .B(new_n817), .Y(new_n2574));
  OAI221xp5_ASAP7_75t_L     g02318(.A1(new_n912), .A2(new_n952), .B1(new_n911), .B2(new_n2573), .C(new_n2574), .Y(new_n2575));
  AOI211xp5_ASAP7_75t_L     g02319(.A1(\b[13] ), .A2(new_n908), .B(new_n813), .C(new_n2575), .Y(new_n2576));
  NAND2xp33_ASAP7_75t_L     g02320(.A(\b[13] ), .B(new_n908), .Y(new_n2577));
  AOI22xp33_ASAP7_75t_L     g02321(.A1(new_n826), .A2(\b[15] ), .B1(new_n823), .B2(new_n959), .Y(new_n2578));
  AOI31xp33_ASAP7_75t_L     g02322(.A1(new_n2578), .A2(new_n2574), .A3(new_n2577), .B(\a[14] ), .Y(new_n2579));
  NOR2xp33_ASAP7_75t_L      g02323(.A(new_n2579), .B(new_n2576), .Y(new_n2580));
  NAND3xp33_ASAP7_75t_L     g02324(.A(new_n2564), .B(new_n2568), .C(new_n2580), .Y(new_n2581));
  NOR3xp33_ASAP7_75t_L      g02325(.A(new_n2565), .B(new_n2566), .C(new_n2567), .Y(new_n2582));
  AOI221xp5_ASAP7_75t_L     g02326(.A1(new_n2413), .A2(new_n2414), .B1(new_n2562), .B2(new_n2563), .C(new_n2411), .Y(new_n2583));
  NAND4xp25_ASAP7_75t_L     g02327(.A(new_n2578), .B(\a[14] ), .C(new_n2577), .D(new_n2574), .Y(new_n2584));
  A2O1A1Ixp33_ASAP7_75t_L   g02328(.A1(\b[13] ), .A2(new_n908), .B(new_n2575), .C(new_n813), .Y(new_n2585));
  NAND2xp33_ASAP7_75t_L     g02329(.A(new_n2584), .B(new_n2585), .Y(new_n2586));
  OAI21xp33_ASAP7_75t_L     g02330(.A1(new_n2583), .A2(new_n2582), .B(new_n2586), .Y(new_n2587));
  NOR2xp33_ASAP7_75t_L      g02331(.A(new_n2416), .B(new_n2412), .Y(new_n2588));
  MAJIxp5_ASAP7_75t_L       g02332(.A(new_n2360), .B(new_n2423), .C(new_n2588), .Y(new_n2589));
  NAND3xp33_ASAP7_75t_L     g02333(.A(new_n2589), .B(new_n2587), .C(new_n2581), .Y(new_n2590));
  NAND2xp33_ASAP7_75t_L     g02334(.A(new_n2587), .B(new_n2581), .Y(new_n2591));
  A2O1A1Ixp33_ASAP7_75t_L   g02335(.A1(new_n2423), .A2(new_n2588), .B(new_n2438), .C(new_n2591), .Y(new_n2592));
  NOR2xp33_ASAP7_75t_L      g02336(.A(new_n1356), .B(new_n676), .Y(new_n2593));
  AOI221xp5_ASAP7_75t_L     g02337(.A1(new_n590), .A2(\b[17] ), .B1(new_n597), .B2(new_n1363), .C(new_n2593), .Y(new_n2594));
  OAI21xp33_ASAP7_75t_L     g02338(.A1(new_n1051), .A2(new_n1620), .B(new_n2594), .Y(new_n2595));
  NOR2xp33_ASAP7_75t_L      g02339(.A(new_n594), .B(new_n2595), .Y(new_n2596));
  O2A1O1Ixp33_ASAP7_75t_L   g02340(.A1(new_n1051), .A2(new_n1620), .B(new_n2594), .C(\a[11] ), .Y(new_n2597));
  NOR2xp33_ASAP7_75t_L      g02341(.A(new_n2597), .B(new_n2596), .Y(new_n2598));
  NAND3xp33_ASAP7_75t_L     g02342(.A(new_n2598), .B(new_n2592), .C(new_n2590), .Y(new_n2599));
  NAND2xp33_ASAP7_75t_L     g02343(.A(new_n2425), .B(new_n2426), .Y(new_n2600));
  MAJIxp5_ASAP7_75t_L       g02344(.A(new_n2431), .B(new_n2427), .C(new_n2600), .Y(new_n2601));
  NOR2xp33_ASAP7_75t_L      g02345(.A(new_n2601), .B(new_n2591), .Y(new_n2602));
  AOI21xp33_ASAP7_75t_L     g02346(.A1(new_n2587), .A2(new_n2581), .B(new_n2589), .Y(new_n2603));
  XNOR2x2_ASAP7_75t_L       g02347(.A(new_n594), .B(new_n2595), .Y(new_n2604));
  OAI21xp33_ASAP7_75t_L     g02348(.A1(new_n2602), .A2(new_n2603), .B(new_n2604), .Y(new_n2605));
  A2O1A1O1Ixp25_ASAP7_75t_L g02349(.A1(new_n2310), .A2(new_n2309), .B(new_n2350), .C(new_n2440), .D(new_n2443), .Y(new_n2606));
  NAND3xp33_ASAP7_75t_L     g02350(.A(new_n2606), .B(new_n2605), .C(new_n2599), .Y(new_n2607));
  AO21x2_ASAP7_75t_L        g02351(.A1(new_n2599), .A2(new_n2605), .B(new_n2606), .Y(new_n2608));
  NOR2xp33_ASAP7_75t_L      g02352(.A(new_n1493), .B(new_n481), .Y(new_n2609));
  INVx1_ASAP7_75t_L         g02353(.A(new_n2609), .Y(new_n2610));
  NOR2xp33_ASAP7_75t_L      g02354(.A(new_n1594), .B(new_n529), .Y(new_n2611));
  INVx1_ASAP7_75t_L         g02355(.A(new_n2611), .Y(new_n2612));
  AOI22xp33_ASAP7_75t_L     g02356(.A1(new_n451), .A2(\b[21] ), .B1(new_n448), .B2(new_n1715), .Y(new_n2613));
  AND4x1_ASAP7_75t_L        g02357(.A(new_n2613), .B(new_n2612), .C(new_n2610), .D(\a[8] ), .Y(new_n2614));
  AOI31xp33_ASAP7_75t_L     g02358(.A1(new_n2613), .A2(new_n2612), .A3(new_n2610), .B(\a[8] ), .Y(new_n2615));
  NOR2xp33_ASAP7_75t_L      g02359(.A(new_n2615), .B(new_n2614), .Y(new_n2616));
  INVx1_ASAP7_75t_L         g02360(.A(new_n2616), .Y(new_n2617));
  AOI21xp33_ASAP7_75t_L     g02361(.A1(new_n2608), .A2(new_n2607), .B(new_n2617), .Y(new_n2618));
  AND3x1_ASAP7_75t_L        g02362(.A(new_n2606), .B(new_n2605), .C(new_n2599), .Y(new_n2619));
  AOI21xp33_ASAP7_75t_L     g02363(.A1(new_n2605), .A2(new_n2599), .B(new_n2606), .Y(new_n2620));
  NOR3xp33_ASAP7_75t_L      g02364(.A(new_n2619), .B(new_n2616), .C(new_n2620), .Y(new_n2621));
  NOR2xp33_ASAP7_75t_L      g02365(.A(new_n2618), .B(new_n2621), .Y(new_n2622));
  NOR3xp33_ASAP7_75t_L      g02366(.A(new_n2456), .B(new_n2453), .C(new_n2455), .Y(new_n2623));
  A2O1A1Ixp33_ASAP7_75t_L   g02367(.A1(new_n2459), .A2(new_n2461), .B(new_n2623), .C(new_n2622), .Y(new_n2624));
  AOI21xp33_ASAP7_75t_L     g02368(.A1(new_n2459), .A2(new_n2461), .B(new_n2623), .Y(new_n2625));
  OAI21xp33_ASAP7_75t_L     g02369(.A1(new_n2618), .A2(new_n2621), .B(new_n2625), .Y(new_n2626));
  NAND2xp33_ASAP7_75t_L     g02370(.A(\b[22] ), .B(new_n366), .Y(new_n2627));
  NAND2xp33_ASAP7_75t_L     g02371(.A(\b[23] ), .B(new_n334), .Y(new_n2628));
  AOI22xp33_ASAP7_75t_L     g02372(.A1(new_n345), .A2(\b[24] ), .B1(new_n342), .B2(new_n2027), .Y(new_n2629));
  NAND4xp25_ASAP7_75t_L     g02373(.A(new_n2629), .B(\a[5] ), .C(new_n2627), .D(new_n2628), .Y(new_n2630));
  NAND2xp33_ASAP7_75t_L     g02374(.A(new_n2628), .B(new_n2629), .Y(new_n2631));
  A2O1A1Ixp33_ASAP7_75t_L   g02375(.A1(\b[22] ), .A2(new_n366), .B(new_n2631), .C(new_n339), .Y(new_n2632));
  AND2x2_ASAP7_75t_L        g02376(.A(new_n2630), .B(new_n2632), .Y(new_n2633));
  NAND3xp33_ASAP7_75t_L     g02377(.A(new_n2624), .B(new_n2633), .C(new_n2626), .Y(new_n2634));
  NOR3xp33_ASAP7_75t_L      g02378(.A(new_n2625), .B(new_n2621), .C(new_n2618), .Y(new_n2635));
  OAI21xp33_ASAP7_75t_L     g02379(.A1(new_n2620), .A2(new_n2619), .B(new_n2616), .Y(new_n2636));
  INVx1_ASAP7_75t_L         g02380(.A(new_n2621), .Y(new_n2637));
  AOI221xp5_ASAP7_75t_L     g02381(.A1(new_n2461), .A2(new_n2459), .B1(new_n2636), .B2(new_n2637), .C(new_n2623), .Y(new_n2638));
  NAND2xp33_ASAP7_75t_L     g02382(.A(new_n2630), .B(new_n2632), .Y(new_n2639));
  OAI21xp33_ASAP7_75t_L     g02383(.A1(new_n2635), .A2(new_n2638), .B(new_n2639), .Y(new_n2640));
  NOR2xp33_ASAP7_75t_L      g02384(.A(new_n2462), .B(new_n2463), .Y(new_n2641));
  NAND2xp33_ASAP7_75t_L     g02385(.A(new_n2470), .B(new_n2641), .Y(new_n2642));
  INVx1_ASAP7_75t_L         g02386(.A(new_n2642), .Y(new_n2643));
  O2A1O1Ixp33_ASAP7_75t_L   g02387(.A1(new_n2330), .A2(new_n2329), .B(new_n2475), .C(new_n2643), .Y(new_n2644));
  NAND3xp33_ASAP7_75t_L     g02388(.A(new_n2644), .B(new_n2640), .C(new_n2634), .Y(new_n2645));
  NAND2xp33_ASAP7_75t_L     g02389(.A(new_n2634), .B(new_n2640), .Y(new_n2646));
  A2O1A1Ixp33_ASAP7_75t_L   g02390(.A1(new_n2349), .A2(new_n2475), .B(new_n2643), .C(new_n2646), .Y(new_n2647));
  INVx1_ASAP7_75t_L         g02391(.A(new_n2481), .Y(new_n2648));
  NOR2xp33_ASAP7_75t_L      g02392(.A(\b[26] ), .B(\b[27] ), .Y(new_n2649));
  INVx1_ASAP7_75t_L         g02393(.A(\b[27] ), .Y(new_n2650));
  NOR2xp33_ASAP7_75t_L      g02394(.A(new_n2477), .B(new_n2650), .Y(new_n2651));
  NOR2xp33_ASAP7_75t_L      g02395(.A(new_n2649), .B(new_n2651), .Y(new_n2652));
  INVx1_ASAP7_75t_L         g02396(.A(new_n2652), .Y(new_n2653));
  O2A1O1Ixp33_ASAP7_75t_L   g02397(.A1(new_n2485), .A2(new_n2484), .B(new_n2648), .C(new_n2653), .Y(new_n2654));
  O2A1O1Ixp33_ASAP7_75t_L   g02398(.A1(new_n2019), .A2(new_n2180), .B(new_n2183), .C(new_n2485), .Y(new_n2655));
  NOR3xp33_ASAP7_75t_L      g02399(.A(new_n2655), .B(new_n2652), .C(new_n2481), .Y(new_n2656));
  NOR2xp33_ASAP7_75t_L      g02400(.A(new_n2654), .B(new_n2656), .Y(new_n2657));
  AOI22xp33_ASAP7_75t_L     g02401(.A1(new_n272), .A2(\b[27] ), .B1(new_n269), .B2(new_n2657), .Y(new_n2658));
  OAI221xp5_ASAP7_75t_L     g02402(.A1(new_n261), .A2(new_n2477), .B1(new_n2180), .B2(new_n277), .C(new_n2658), .Y(new_n2659));
  XNOR2x2_ASAP7_75t_L       g02403(.A(new_n265), .B(new_n2659), .Y(new_n2660));
  AOI21xp33_ASAP7_75t_L     g02404(.A1(new_n2645), .A2(new_n2647), .B(new_n2660), .Y(new_n2661));
  NAND3xp33_ASAP7_75t_L     g02405(.A(new_n2645), .B(new_n2647), .C(new_n2660), .Y(new_n2662));
  INVx1_ASAP7_75t_L         g02406(.A(new_n2662), .Y(new_n2663));
  NOR2xp33_ASAP7_75t_L      g02407(.A(new_n2661), .B(new_n2663), .Y(new_n2664));
  INVx1_ASAP7_75t_L         g02408(.A(new_n2664), .Y(new_n2665));
  O2A1O1Ixp33_ASAP7_75t_L   g02409(.A1(new_n2348), .A2(new_n2494), .B(new_n2492), .C(new_n2665), .Y(new_n2666));
  A2O1A1O1Ixp25_ASAP7_75t_L g02410(.A1(new_n2341), .A2(new_n2344), .B(new_n2334), .C(new_n2493), .D(new_n2491), .Y(new_n2667));
  INVx1_ASAP7_75t_L         g02411(.A(new_n2667), .Y(new_n2668));
  NOR2xp33_ASAP7_75t_L      g02412(.A(new_n2668), .B(new_n2664), .Y(new_n2669));
  NOR2xp33_ASAP7_75t_L      g02413(.A(new_n2669), .B(new_n2666), .Y(\f[27] ));
  NOR3xp33_ASAP7_75t_L      g02414(.A(new_n2582), .B(new_n2583), .C(new_n2580), .Y(new_n2671));
  NAND2xp33_ASAP7_75t_L     g02415(.A(new_n2521), .B(new_n2525), .Y(new_n2672));
  NOR2xp33_ASAP7_75t_L      g02416(.A(new_n2529), .B(new_n2537), .Y(new_n2673));
  MAJIxp5_ASAP7_75t_L       g02417(.A(new_n2543), .B(new_n2672), .C(new_n2673), .Y(new_n2674));
  NAND2xp33_ASAP7_75t_L     g02418(.A(\b[5] ), .B(new_n1910), .Y(new_n2675));
  NAND2xp33_ASAP7_75t_L     g02419(.A(\b[6] ), .B(new_n1770), .Y(new_n2676));
  AOI32xp33_ASAP7_75t_L     g02420(.A1(new_n424), .A2(new_n426), .A3(new_n1764), .B1(new_n1766), .B2(\b[7] ), .Y(new_n2677));
  NAND4xp25_ASAP7_75t_L     g02421(.A(new_n2677), .B(\a[23] ), .C(new_n2675), .D(new_n2676), .Y(new_n2678));
  INVx1_ASAP7_75t_L         g02422(.A(new_n2678), .Y(new_n2679));
  AOI31xp33_ASAP7_75t_L     g02423(.A1(new_n2677), .A2(new_n2676), .A3(new_n2675), .B(\a[23] ), .Y(new_n2680));
  NOR3xp33_ASAP7_75t_L      g02424(.A(new_n2507), .B(new_n2388), .C(new_n2390), .Y(new_n2681));
  NAND2xp33_ASAP7_75t_L     g02425(.A(new_n2512), .B(new_n2681), .Y(new_n2682));
  NAND2xp33_ASAP7_75t_L     g02426(.A(\b[2] ), .B(new_n2386), .Y(new_n2683));
  NOR2xp33_ASAP7_75t_L      g02427(.A(new_n299), .B(new_n2220), .Y(new_n2684));
  INVx1_ASAP7_75t_L         g02428(.A(new_n2684), .Y(new_n2685));
  OAI32xp33_ASAP7_75t_L     g02429(.A1(new_n325), .A2(new_n327), .A3(new_n2233), .B1(new_n323), .B2(new_n2234), .Y(new_n2686));
  INVx1_ASAP7_75t_L         g02430(.A(new_n2686), .Y(new_n2687));
  NAND4xp25_ASAP7_75t_L     g02431(.A(new_n2687), .B(\a[26] ), .C(new_n2683), .D(new_n2685), .Y(new_n2688));
  INVx1_ASAP7_75t_L         g02432(.A(new_n2683), .Y(new_n2689));
  OAI31xp33_ASAP7_75t_L     g02433(.A1(new_n2689), .A2(new_n2686), .A3(new_n2684), .B(new_n2223), .Y(new_n2690));
  NAND2xp33_ASAP7_75t_L     g02434(.A(\a[29] ), .B(new_n2512), .Y(new_n2691));
  XNOR2x2_ASAP7_75t_L       g02435(.A(\a[28] ), .B(\a[27] ), .Y(new_n2692));
  INVx1_ASAP7_75t_L         g02436(.A(new_n2692), .Y(new_n2693));
  NAND2xp33_ASAP7_75t_L     g02437(.A(new_n2693), .B(new_n2511), .Y(new_n2694));
  INVx1_ASAP7_75t_L         g02438(.A(\a[28] ), .Y(new_n2695));
  NAND2xp33_ASAP7_75t_L     g02439(.A(\a[29] ), .B(new_n2695), .Y(new_n2696));
  INVx1_ASAP7_75t_L         g02440(.A(\a[29] ), .Y(new_n2697));
  NAND2xp33_ASAP7_75t_L     g02441(.A(\a[28] ), .B(new_n2697), .Y(new_n2698));
  AND2x2_ASAP7_75t_L        g02442(.A(new_n2696), .B(new_n2698), .Y(new_n2699));
  NOR2xp33_ASAP7_75t_L      g02443(.A(new_n2511), .B(new_n2699), .Y(new_n2700));
  NAND2xp33_ASAP7_75t_L     g02444(.A(new_n2698), .B(new_n2696), .Y(new_n2701));
  NOR2xp33_ASAP7_75t_L      g02445(.A(new_n2701), .B(new_n2511), .Y(new_n2702));
  AOI22xp33_ASAP7_75t_L     g02446(.A1(new_n2702), .A2(\b[1] ), .B1(new_n271), .B2(new_n2700), .Y(new_n2703));
  O2A1O1Ixp33_ASAP7_75t_L   g02447(.A1(new_n2694), .A2(new_n258), .B(new_n2703), .C(new_n2691), .Y(new_n2704));
  NAND2xp33_ASAP7_75t_L     g02448(.A(new_n2510), .B(new_n2509), .Y(new_n2705));
  NOR2xp33_ASAP7_75t_L      g02449(.A(new_n2692), .B(new_n2705), .Y(new_n2706));
  NAND2xp33_ASAP7_75t_L     g02450(.A(new_n2701), .B(new_n2705), .Y(new_n2707));
  NAND2xp33_ASAP7_75t_L     g02451(.A(new_n2705), .B(new_n2699), .Y(new_n2708));
  OAI22xp33_ASAP7_75t_L     g02452(.A1(new_n2708), .A2(new_n276), .B1(new_n270), .B2(new_n2707), .Y(new_n2709));
  A2O1A1O1Ixp25_ASAP7_75t_L g02453(.A1(new_n2705), .A2(\a[29] ), .B(new_n2706), .C(\b[0] ), .D(new_n2709), .Y(new_n2710));
  NOR2xp33_ASAP7_75t_L      g02454(.A(new_n2710), .B(new_n2704), .Y(new_n2711));
  NAND3xp33_ASAP7_75t_L     g02455(.A(new_n2688), .B(new_n2711), .C(new_n2690), .Y(new_n2712));
  NOR4xp25_ASAP7_75t_L      g02456(.A(new_n2689), .B(new_n2686), .C(new_n2223), .D(new_n2684), .Y(new_n2713));
  AOI31xp33_ASAP7_75t_L     g02457(.A1(new_n2687), .A2(new_n2685), .A3(new_n2683), .B(\a[26] ), .Y(new_n2714));
  OR2x4_ASAP7_75t_L         g02458(.A(new_n2710), .B(new_n2704), .Y(new_n2715));
  OAI21xp33_ASAP7_75t_L     g02459(.A1(new_n2713), .A2(new_n2714), .B(new_n2715), .Y(new_n2716));
  AO22x1_ASAP7_75t_L        g02460(.A1(new_n2716), .A2(new_n2712), .B1(new_n2682), .B2(new_n2521), .Y(new_n2717));
  NAND2xp33_ASAP7_75t_L     g02461(.A(new_n2534), .B(new_n2533), .Y(new_n2718));
  INVx1_ASAP7_75t_L         g02462(.A(new_n2512), .Y(new_n2719));
  NOR4xp25_ASAP7_75t_L      g02463(.A(new_n2507), .B(new_n2719), .C(new_n2390), .D(new_n2388), .Y(new_n2720));
  O2A1O1Ixp33_ASAP7_75t_L   g02464(.A1(new_n2513), .A2(new_n2514), .B(new_n2718), .C(new_n2720), .Y(new_n2721));
  NAND3xp33_ASAP7_75t_L     g02465(.A(new_n2721), .B(new_n2712), .C(new_n2716), .Y(new_n2722));
  OAI211xp5_ASAP7_75t_L     g02466(.A1(new_n2680), .A2(new_n2679), .B(new_n2722), .C(new_n2717), .Y(new_n2723));
  INVx1_ASAP7_75t_L         g02467(.A(new_n2680), .Y(new_n2724));
  AOI22xp33_ASAP7_75t_L     g02468(.A1(new_n2712), .A2(new_n2716), .B1(new_n2682), .B2(new_n2521), .Y(new_n2725));
  AND4x1_ASAP7_75t_L        g02469(.A(new_n2521), .B(new_n2716), .C(new_n2682), .D(new_n2712), .Y(new_n2726));
  OAI211xp5_ASAP7_75t_L     g02470(.A1(new_n2725), .A2(new_n2726), .B(new_n2724), .C(new_n2678), .Y(new_n2727));
  NAND3xp33_ASAP7_75t_L     g02471(.A(new_n2674), .B(new_n2723), .C(new_n2727), .Y(new_n2728));
  NOR2xp33_ASAP7_75t_L      g02472(.A(new_n2673), .B(new_n2672), .Y(new_n2729));
  O2A1O1Ixp33_ASAP7_75t_L   g02473(.A1(new_n2504), .A2(new_n2540), .B(new_n2542), .C(new_n2729), .Y(new_n2730));
  AOI211xp5_ASAP7_75t_L     g02474(.A1(new_n2724), .A2(new_n2678), .B(new_n2725), .C(new_n2726), .Y(new_n2731));
  AOI211xp5_ASAP7_75t_L     g02475(.A1(new_n2722), .A2(new_n2717), .B(new_n2679), .C(new_n2680), .Y(new_n2732));
  OAI21xp33_ASAP7_75t_L     g02476(.A1(new_n2731), .A2(new_n2732), .B(new_n2730), .Y(new_n2733));
  NAND2xp33_ASAP7_75t_L     g02477(.A(\b[9] ), .B(new_n1410), .Y(new_n2734));
  NAND2xp33_ASAP7_75t_L     g02478(.A(\b[10] ), .B(new_n1406), .Y(new_n2735));
  OAI311xp33_ASAP7_75t_L    g02479(.A1(new_n639), .A2(new_n851), .A3(new_n1411), .B1(new_n2735), .C1(new_n2734), .Y(new_n2736));
  AOI21xp33_ASAP7_75t_L     g02480(.A1(new_n1548), .A2(\b[8] ), .B(new_n2736), .Y(new_n2737));
  NAND2xp33_ASAP7_75t_L     g02481(.A(\a[20] ), .B(new_n2737), .Y(new_n2738));
  A2O1A1Ixp33_ASAP7_75t_L   g02482(.A1(\b[8] ), .A2(new_n1548), .B(new_n2736), .C(new_n1401), .Y(new_n2739));
  NAND4xp25_ASAP7_75t_L     g02483(.A(new_n2733), .B(new_n2728), .C(new_n2738), .D(new_n2739), .Y(new_n2740));
  NOR3xp33_ASAP7_75t_L      g02484(.A(new_n2730), .B(new_n2731), .C(new_n2732), .Y(new_n2741));
  AOI21xp33_ASAP7_75t_L     g02485(.A1(new_n2727), .A2(new_n2723), .B(new_n2674), .Y(new_n2742));
  NAND2xp33_ASAP7_75t_L     g02486(.A(new_n2739), .B(new_n2738), .Y(new_n2743));
  OAI21xp33_ASAP7_75t_L     g02487(.A1(new_n2742), .A2(new_n2741), .B(new_n2743), .Y(new_n2744));
  A2O1A1O1Ixp25_ASAP7_75t_L g02488(.A1(new_n2401), .A2(new_n2371), .B(new_n2402), .C(new_n2560), .D(new_n2552), .Y(new_n2745));
  NAND3xp33_ASAP7_75t_L     g02489(.A(new_n2745), .B(new_n2744), .C(new_n2740), .Y(new_n2746));
  NOR3xp33_ASAP7_75t_L      g02490(.A(new_n2741), .B(new_n2742), .C(new_n2743), .Y(new_n2747));
  AND2x2_ASAP7_75t_L        g02491(.A(new_n2739), .B(new_n2738), .Y(new_n2748));
  AOI21xp33_ASAP7_75t_L     g02492(.A1(new_n2733), .A2(new_n2728), .B(new_n2748), .Y(new_n2749));
  OAI21xp33_ASAP7_75t_L     g02493(.A1(new_n2557), .A2(new_n2503), .B(new_n2559), .Y(new_n2750));
  OAI21xp33_ASAP7_75t_L     g02494(.A1(new_n2747), .A2(new_n2749), .B(new_n2750), .Y(new_n2751));
  NAND2xp33_ASAP7_75t_L     g02495(.A(\b[12] ), .B(new_n1103), .Y(new_n2752));
  NAND2xp33_ASAP7_75t_L     g02496(.A(\b[13] ), .B(new_n1113), .Y(new_n2753));
  OAI311xp33_ASAP7_75t_L    g02497(.A1(new_n799), .A2(new_n797), .A3(new_n1197), .B1(new_n2753), .C1(new_n2752), .Y(new_n2754));
  AOI21xp33_ASAP7_75t_L     g02498(.A1(new_n1194), .A2(\b[11] ), .B(new_n2754), .Y(new_n2755));
  NAND2xp33_ASAP7_75t_L     g02499(.A(\a[17] ), .B(new_n2755), .Y(new_n2756));
  A2O1A1Ixp33_ASAP7_75t_L   g02500(.A1(\b[11] ), .A2(new_n1194), .B(new_n2754), .C(new_n1107), .Y(new_n2757));
  NAND4xp25_ASAP7_75t_L     g02501(.A(new_n2751), .B(new_n2746), .C(new_n2756), .D(new_n2757), .Y(new_n2758));
  NOR3xp33_ASAP7_75t_L      g02502(.A(new_n2750), .B(new_n2749), .C(new_n2747), .Y(new_n2759));
  AOI21xp33_ASAP7_75t_L     g02503(.A1(new_n2744), .A2(new_n2740), .B(new_n2745), .Y(new_n2760));
  NAND2xp33_ASAP7_75t_L     g02504(.A(new_n2757), .B(new_n2756), .Y(new_n2761));
  OAI21xp33_ASAP7_75t_L     g02505(.A1(new_n2760), .A2(new_n2759), .B(new_n2761), .Y(new_n2762));
  AOI221xp5_ASAP7_75t_L     g02506(.A1(new_n2762), .A2(new_n2758), .B1(new_n2562), .B2(new_n2496), .C(new_n2567), .Y(new_n2763));
  NOR3xp33_ASAP7_75t_L      g02507(.A(new_n2759), .B(new_n2760), .C(new_n2761), .Y(new_n2764));
  AOI22xp33_ASAP7_75t_L     g02508(.A1(new_n2756), .A2(new_n2757), .B1(new_n2746), .B2(new_n2751), .Y(new_n2765));
  A2O1A1O1Ixp25_ASAP7_75t_L g02509(.A1(new_n2414), .A2(new_n2413), .B(new_n2411), .C(new_n2562), .D(new_n2567), .Y(new_n2766));
  NOR3xp33_ASAP7_75t_L      g02510(.A(new_n2766), .B(new_n2765), .C(new_n2764), .Y(new_n2767));
  NAND2xp33_ASAP7_75t_L     g02511(.A(\b[15] ), .B(new_n817), .Y(new_n2768));
  NAND2xp33_ASAP7_75t_L     g02512(.A(\b[16] ), .B(new_n826), .Y(new_n2769));
  OAI311xp33_ASAP7_75t_L    g02513(.A1(new_n1057), .A2(new_n1055), .A3(new_n911), .B1(new_n2769), .C1(new_n2768), .Y(new_n2770));
  AOI21xp33_ASAP7_75t_L     g02514(.A1(new_n908), .A2(\b[14] ), .B(new_n2770), .Y(new_n2771));
  NAND2xp33_ASAP7_75t_L     g02515(.A(\a[14] ), .B(new_n2771), .Y(new_n2772));
  A2O1A1Ixp33_ASAP7_75t_L   g02516(.A1(\b[14] ), .A2(new_n908), .B(new_n2770), .C(new_n813), .Y(new_n2773));
  NAND2xp33_ASAP7_75t_L     g02517(.A(new_n2773), .B(new_n2772), .Y(new_n2774));
  OAI21xp33_ASAP7_75t_L     g02518(.A1(new_n2767), .A2(new_n2763), .B(new_n2774), .Y(new_n2775));
  OAI21xp33_ASAP7_75t_L     g02519(.A1(new_n2764), .A2(new_n2765), .B(new_n2766), .Y(new_n2776));
  OR3x1_ASAP7_75t_L         g02520(.A(new_n2766), .B(new_n2764), .C(new_n2765), .Y(new_n2777));
  NAND4xp25_ASAP7_75t_L     g02521(.A(new_n2777), .B(new_n2772), .C(new_n2773), .D(new_n2776), .Y(new_n2778));
  AOI221xp5_ASAP7_75t_L     g02522(.A1(new_n2778), .A2(new_n2775), .B1(new_n2601), .B2(new_n2591), .C(new_n2671), .Y(new_n2779));
  NOR2xp33_ASAP7_75t_L      g02523(.A(new_n2583), .B(new_n2582), .Y(new_n2780));
  MAJIxp5_ASAP7_75t_L       g02524(.A(new_n2601), .B(new_n2780), .C(new_n2586), .Y(new_n2781));
  OA21x2_ASAP7_75t_L        g02525(.A1(new_n2767), .A2(new_n2763), .B(new_n2774), .Y(new_n2782));
  NOR3xp33_ASAP7_75t_L      g02526(.A(new_n2763), .B(new_n2767), .C(new_n2774), .Y(new_n2783));
  NOR3xp33_ASAP7_75t_L      g02527(.A(new_n2781), .B(new_n2782), .C(new_n2783), .Y(new_n2784));
  NOR2xp33_ASAP7_75t_L      g02528(.A(new_n1244), .B(new_n1620), .Y(new_n2785));
  INVx1_ASAP7_75t_L         g02529(.A(new_n2785), .Y(new_n2786));
  NAND2xp33_ASAP7_75t_L     g02530(.A(\b[18] ), .B(new_n590), .Y(new_n2787));
  AOI22xp33_ASAP7_75t_L     g02531(.A1(new_n600), .A2(\b[19] ), .B1(new_n597), .B2(new_n1499), .Y(new_n2788));
  NAND4xp25_ASAP7_75t_L     g02532(.A(new_n2788), .B(\a[11] ), .C(new_n2786), .D(new_n2787), .Y(new_n2789));
  A2O1A1Ixp33_ASAP7_75t_L   g02533(.A1(new_n2570), .A2(new_n1049), .B(new_n1050), .C(new_n1352), .Y(new_n2790));
  A2O1A1O1Ixp25_ASAP7_75t_L g02534(.A1(new_n1246), .A2(new_n2790), .B(new_n1245), .C(new_n1358), .D(new_n1357), .Y(new_n2791));
  OAI21xp33_ASAP7_75t_L     g02535(.A1(new_n1492), .A2(new_n1494), .B(new_n2791), .Y(new_n2792));
  NAND2xp33_ASAP7_75t_L     g02536(.A(new_n1496), .B(new_n2792), .Y(new_n2793));
  OAI221xp5_ASAP7_75t_L     g02537(.A1(new_n676), .A2(new_n1493), .B1(new_n675), .B2(new_n2793), .C(new_n2787), .Y(new_n2794));
  A2O1A1Ixp33_ASAP7_75t_L   g02538(.A1(\b[17] ), .A2(new_n674), .B(new_n2794), .C(new_n594), .Y(new_n2795));
  NAND2xp33_ASAP7_75t_L     g02539(.A(new_n2789), .B(new_n2795), .Y(new_n2796));
  NOR3xp33_ASAP7_75t_L      g02540(.A(new_n2784), .B(new_n2796), .C(new_n2779), .Y(new_n2797));
  OAI21xp33_ASAP7_75t_L     g02541(.A1(new_n2782), .A2(new_n2783), .B(new_n2781), .Y(new_n2798));
  INVx1_ASAP7_75t_L         g02542(.A(new_n2671), .Y(new_n2799));
  A2O1A1Ixp33_ASAP7_75t_L   g02543(.A1(new_n2587), .A2(new_n2581), .B(new_n2589), .C(new_n2799), .Y(new_n2800));
  NOR2xp33_ASAP7_75t_L      g02544(.A(new_n2783), .B(new_n2782), .Y(new_n2801));
  NAND2xp33_ASAP7_75t_L     g02545(.A(new_n2801), .B(new_n2800), .Y(new_n2802));
  NOR3xp33_ASAP7_75t_L      g02546(.A(new_n2794), .B(new_n2785), .C(new_n594), .Y(new_n2803));
  AOI31xp33_ASAP7_75t_L     g02547(.A1(new_n2788), .A2(new_n2787), .A3(new_n2786), .B(\a[11] ), .Y(new_n2804));
  NOR2xp33_ASAP7_75t_L      g02548(.A(new_n2804), .B(new_n2803), .Y(new_n2805));
  AOI21xp33_ASAP7_75t_L     g02549(.A1(new_n2802), .A2(new_n2798), .B(new_n2805), .Y(new_n2806));
  NOR2xp33_ASAP7_75t_L      g02550(.A(new_n2806), .B(new_n2797), .Y(new_n2807));
  NAND2xp33_ASAP7_75t_L     g02551(.A(new_n2590), .B(new_n2592), .Y(new_n2808));
  INVx1_ASAP7_75t_L         g02552(.A(new_n2808), .Y(new_n2809));
  NAND2xp33_ASAP7_75t_L     g02553(.A(new_n2604), .B(new_n2809), .Y(new_n2810));
  NAND3xp33_ASAP7_75t_L     g02554(.A(new_n2807), .B(new_n2608), .C(new_n2810), .Y(new_n2811));
  NAND3xp33_ASAP7_75t_L     g02555(.A(new_n2802), .B(new_n2805), .C(new_n2798), .Y(new_n2812));
  OAI21xp33_ASAP7_75t_L     g02556(.A1(new_n2779), .A2(new_n2784), .B(new_n2796), .Y(new_n2813));
  NAND2xp33_ASAP7_75t_L     g02557(.A(new_n2812), .B(new_n2813), .Y(new_n2814));
  A2O1A1Ixp33_ASAP7_75t_L   g02558(.A1(new_n2604), .A2(new_n2809), .B(new_n2620), .C(new_n2814), .Y(new_n2815));
  NAND2xp33_ASAP7_75t_L     g02559(.A(\b[21] ), .B(new_n441), .Y(new_n2816));
  OAI221xp5_ASAP7_75t_L     g02560(.A1(new_n667), .A2(new_n1857), .B1(new_n482), .B2(new_n1863), .C(new_n2816), .Y(new_n2817));
  INVx1_ASAP7_75t_L         g02561(.A(new_n2817), .Y(new_n2818));
  OAI211xp5_ASAP7_75t_L     g02562(.A1(new_n1594), .A2(new_n481), .B(new_n2818), .C(\a[8] ), .Y(new_n2819));
  A2O1A1Ixp33_ASAP7_75t_L   g02563(.A1(\b[20] ), .A2(new_n480), .B(new_n2817), .C(new_n445), .Y(new_n2820));
  NAND2xp33_ASAP7_75t_L     g02564(.A(new_n2820), .B(new_n2819), .Y(new_n2821));
  AO21x2_ASAP7_75t_L        g02565(.A1(new_n2815), .A2(new_n2811), .B(new_n2821), .Y(new_n2822));
  NAND3xp33_ASAP7_75t_L     g02566(.A(new_n2811), .B(new_n2815), .C(new_n2821), .Y(new_n2823));
  A2O1A1O1Ixp25_ASAP7_75t_L g02567(.A1(new_n2461), .A2(new_n2459), .B(new_n2623), .C(new_n2636), .D(new_n2621), .Y(new_n2824));
  INVx1_ASAP7_75t_L         g02568(.A(new_n2824), .Y(new_n2825));
  NAND3xp33_ASAP7_75t_L     g02569(.A(new_n2825), .B(new_n2823), .C(new_n2822), .Y(new_n2826));
  NAND2xp33_ASAP7_75t_L     g02570(.A(new_n2823), .B(new_n2822), .Y(new_n2827));
  NAND2xp33_ASAP7_75t_L     g02571(.A(new_n2824), .B(new_n2827), .Y(new_n2828));
  NOR2xp33_ASAP7_75t_L      g02572(.A(new_n1995), .B(new_n365), .Y(new_n2829));
  NOR2xp33_ASAP7_75t_L      g02573(.A(new_n2180), .B(new_n368), .Y(new_n2830));
  INVx1_ASAP7_75t_L         g02574(.A(new_n2830), .Y(new_n2831));
  OAI221xp5_ASAP7_75t_L     g02575(.A1(new_n2019), .A2(new_n406), .B1(new_n367), .B2(new_n2187), .C(new_n2831), .Y(new_n2832));
  NOR3xp33_ASAP7_75t_L      g02576(.A(new_n2832), .B(new_n2829), .C(new_n339), .Y(new_n2833));
  INVx1_ASAP7_75t_L         g02577(.A(new_n2833), .Y(new_n2834));
  A2O1A1Ixp33_ASAP7_75t_L   g02578(.A1(\b[23] ), .A2(new_n366), .B(new_n2832), .C(new_n339), .Y(new_n2835));
  NAND2xp33_ASAP7_75t_L     g02579(.A(new_n2835), .B(new_n2834), .Y(new_n2836));
  INVx1_ASAP7_75t_L         g02580(.A(new_n2836), .Y(new_n2837));
  NAND3xp33_ASAP7_75t_L     g02581(.A(new_n2837), .B(new_n2828), .C(new_n2826), .Y(new_n2838));
  NOR2xp33_ASAP7_75t_L      g02582(.A(new_n2824), .B(new_n2827), .Y(new_n2839));
  AOI21xp33_ASAP7_75t_L     g02583(.A1(new_n2823), .A2(new_n2822), .B(new_n2825), .Y(new_n2840));
  OAI21xp33_ASAP7_75t_L     g02584(.A1(new_n2840), .A2(new_n2839), .B(new_n2836), .Y(new_n2841));
  NAND2xp33_ASAP7_75t_L     g02585(.A(new_n2841), .B(new_n2838), .Y(new_n2842));
  NAND2xp33_ASAP7_75t_L     g02586(.A(new_n2626), .B(new_n2624), .Y(new_n2843));
  NOR2xp33_ASAP7_75t_L      g02587(.A(new_n2633), .B(new_n2843), .Y(new_n2844));
  A2O1A1O1Ixp25_ASAP7_75t_L g02588(.A1(new_n2475), .A2(new_n2349), .B(new_n2643), .C(new_n2646), .D(new_n2844), .Y(new_n2845));
  INVx1_ASAP7_75t_L         g02589(.A(new_n2845), .Y(new_n2846));
  NOR2xp33_ASAP7_75t_L      g02590(.A(new_n2842), .B(new_n2846), .Y(new_n2847));
  A2O1A1Ixp33_ASAP7_75t_L   g02591(.A1(new_n2471), .A2(new_n2472), .B(new_n2474), .C(new_n2642), .Y(new_n2848));
  A2O1A1Ixp33_ASAP7_75t_L   g02592(.A1(new_n2848), .A2(new_n2646), .B(new_n2844), .C(new_n2842), .Y(new_n2849));
  INVx1_ASAP7_75t_L         g02593(.A(new_n2849), .Y(new_n2850));
  NOR2xp33_ASAP7_75t_L      g02594(.A(\b[27] ), .B(\b[28] ), .Y(new_n2851));
  INVx1_ASAP7_75t_L         g02595(.A(\b[28] ), .Y(new_n2852));
  NOR2xp33_ASAP7_75t_L      g02596(.A(new_n2650), .B(new_n2852), .Y(new_n2853));
  NOR2xp33_ASAP7_75t_L      g02597(.A(new_n2851), .B(new_n2853), .Y(new_n2854));
  A2O1A1Ixp33_ASAP7_75t_L   g02598(.A1(\b[27] ), .A2(\b[26] ), .B(new_n2654), .C(new_n2854), .Y(new_n2855));
  O2A1O1Ixp33_ASAP7_75t_L   g02599(.A1(new_n2481), .A2(new_n2655), .B(new_n2652), .C(new_n2651), .Y(new_n2856));
  OAI21xp33_ASAP7_75t_L     g02600(.A1(new_n2851), .A2(new_n2853), .B(new_n2856), .Y(new_n2857));
  AND2x2_ASAP7_75t_L        g02601(.A(new_n2855), .B(new_n2857), .Y(new_n2858));
  AOI22xp33_ASAP7_75t_L     g02602(.A1(new_n272), .A2(\b[28] ), .B1(new_n269), .B2(new_n2858), .Y(new_n2859));
  OAI221xp5_ASAP7_75t_L     g02603(.A1(new_n261), .A2(new_n2650), .B1(new_n2477), .B2(new_n277), .C(new_n2859), .Y(new_n2860));
  XNOR2x2_ASAP7_75t_L       g02604(.A(\a[2] ), .B(new_n2860), .Y(new_n2861));
  OAI21xp33_ASAP7_75t_L     g02605(.A1(new_n2850), .A2(new_n2847), .B(new_n2861), .Y(new_n2862));
  NOR3xp33_ASAP7_75t_L      g02606(.A(new_n2847), .B(new_n2850), .C(new_n2861), .Y(new_n2863));
  INVx1_ASAP7_75t_L         g02607(.A(new_n2863), .Y(new_n2864));
  NAND2xp33_ASAP7_75t_L     g02608(.A(new_n2862), .B(new_n2864), .Y(new_n2865));
  O2A1O1Ixp33_ASAP7_75t_L   g02609(.A1(new_n2667), .A2(new_n2661), .B(new_n2662), .C(new_n2865), .Y(new_n2866));
  OAI21xp33_ASAP7_75t_L     g02610(.A1(new_n2661), .A2(new_n2667), .B(new_n2662), .Y(new_n2867));
  AOI21xp33_ASAP7_75t_L     g02611(.A1(new_n2864), .A2(new_n2862), .B(new_n2867), .Y(new_n2868));
  NOR2xp33_ASAP7_75t_L      g02612(.A(new_n2868), .B(new_n2866), .Y(\f[28] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02613(.A1(new_n2668), .A2(new_n2664), .B(new_n2663), .C(new_n2862), .D(new_n2863), .Y(new_n2870));
  INVx1_ASAP7_75t_L         g02614(.A(\b[29] ), .Y(new_n2871));
  INVx1_ASAP7_75t_L         g02615(.A(new_n2651), .Y(new_n2872));
  A2O1A1Ixp33_ASAP7_75t_L   g02616(.A1(new_n2483), .A2(new_n2648), .B(new_n2649), .C(new_n2872), .Y(new_n2873));
  NOR2xp33_ASAP7_75t_L      g02617(.A(\b[28] ), .B(\b[29] ), .Y(new_n2874));
  NOR2xp33_ASAP7_75t_L      g02618(.A(new_n2852), .B(new_n2871), .Y(new_n2875));
  NOR2xp33_ASAP7_75t_L      g02619(.A(new_n2874), .B(new_n2875), .Y(new_n2876));
  A2O1A1Ixp33_ASAP7_75t_L   g02620(.A1(new_n2873), .A2(new_n2854), .B(new_n2853), .C(new_n2876), .Y(new_n2877));
  O2A1O1Ixp33_ASAP7_75t_L   g02621(.A1(new_n2651), .A2(new_n2654), .B(new_n2854), .C(new_n2853), .Y(new_n2878));
  INVx1_ASAP7_75t_L         g02622(.A(new_n2876), .Y(new_n2879));
  NAND2xp33_ASAP7_75t_L     g02623(.A(new_n2879), .B(new_n2878), .Y(new_n2880));
  NAND2xp33_ASAP7_75t_L     g02624(.A(new_n2880), .B(new_n2877), .Y(new_n2881));
  OAI22xp33_ASAP7_75t_L     g02625(.A1(new_n2881), .A2(new_n292), .B1(new_n2871), .B2(new_n632), .Y(new_n2882));
  AOI221xp5_ASAP7_75t_L     g02626(.A1(\b[27] ), .A2(new_n291), .B1(\b[28] ), .B2(new_n380), .C(new_n2882), .Y(new_n2883));
  XNOR2x2_ASAP7_75t_L       g02627(.A(new_n265), .B(new_n2883), .Y(new_n2884));
  NAND2xp33_ASAP7_75t_L     g02628(.A(new_n2828), .B(new_n2826), .Y(new_n2885));
  NAND2xp33_ASAP7_75t_L     g02629(.A(\b[24] ), .B(new_n366), .Y(new_n2886));
  NAND2xp33_ASAP7_75t_L     g02630(.A(\b[25] ), .B(new_n334), .Y(new_n2887));
  AND2x2_ASAP7_75t_L        g02631(.A(new_n2486), .B(new_n2483), .Y(new_n2888));
  AOI22xp33_ASAP7_75t_L     g02632(.A1(new_n345), .A2(\b[26] ), .B1(new_n342), .B2(new_n2888), .Y(new_n2889));
  AND4x1_ASAP7_75t_L        g02633(.A(new_n2889), .B(new_n2887), .C(new_n2886), .D(\a[5] ), .Y(new_n2890));
  AOI31xp33_ASAP7_75t_L     g02634(.A1(new_n2889), .A2(new_n2887), .A3(new_n2886), .B(\a[5] ), .Y(new_n2891));
  NOR2xp33_ASAP7_75t_L      g02635(.A(new_n2891), .B(new_n2890), .Y(new_n2892));
  AOI21xp33_ASAP7_75t_L     g02636(.A1(new_n2811), .A2(new_n2815), .B(new_n2821), .Y(new_n2893));
  OAI21xp33_ASAP7_75t_L     g02637(.A1(new_n2893), .A2(new_n2824), .B(new_n2823), .Y(new_n2894));
  AOI32xp33_ASAP7_75t_L     g02638(.A1(new_n1998), .A2(new_n2001), .A3(new_n448), .B1(new_n451), .B2(\b[23] ), .Y(new_n2895));
  OAI221xp5_ASAP7_75t_L     g02639(.A1(new_n529), .A2(new_n1857), .B1(new_n1709), .B2(new_n481), .C(new_n2895), .Y(new_n2896));
  XNOR2x2_ASAP7_75t_L       g02640(.A(\a[8] ), .B(new_n2896), .Y(new_n2897));
  INVx1_ASAP7_75t_L         g02641(.A(new_n2897), .Y(new_n2898));
  O2A1O1Ixp33_ASAP7_75t_L   g02642(.A1(new_n2808), .A2(new_n2598), .B(new_n2608), .C(new_n2807), .Y(new_n2899));
  NOR3xp33_ASAP7_75t_L      g02643(.A(new_n2784), .B(new_n2805), .C(new_n2779), .Y(new_n2900));
  NOR2xp33_ASAP7_75t_L      g02644(.A(new_n2742), .B(new_n2741), .Y(new_n2901));
  MAJIxp5_ASAP7_75t_L       g02645(.A(new_n2750), .B(new_n2743), .C(new_n2901), .Y(new_n2902));
  NOR2xp33_ASAP7_75t_L      g02646(.A(new_n559), .B(new_n1549), .Y(new_n2903));
  INVx1_ASAP7_75t_L         g02647(.A(new_n2903), .Y(new_n2904));
  NAND2xp33_ASAP7_75t_L     g02648(.A(\b[10] ), .B(new_n1410), .Y(new_n2905));
  AOI32xp33_ASAP7_75t_L     g02649(.A1(new_n700), .A2(new_n698), .A3(new_n1404), .B1(\b[11] ), .B2(new_n1406), .Y(new_n2906));
  AND4x1_ASAP7_75t_L        g02650(.A(new_n2906), .B(new_n2905), .C(new_n2904), .D(\a[20] ), .Y(new_n2907));
  AOI31xp33_ASAP7_75t_L     g02651(.A1(new_n2906), .A2(new_n2905), .A3(new_n2904), .B(\a[20] ), .Y(new_n2908));
  NOR2xp33_ASAP7_75t_L      g02652(.A(new_n2908), .B(new_n2907), .Y(new_n2909));
  INVx1_ASAP7_75t_L         g02653(.A(new_n2909), .Y(new_n2910));
  INVx1_ASAP7_75t_L         g02654(.A(new_n2729), .Y(new_n2911));
  NOR4xp25_ASAP7_75t_L      g02655(.A(new_n2535), .B(new_n2536), .C(new_n2537), .D(new_n2529), .Y(new_n2912));
  AOI22xp33_ASAP7_75t_L     g02656(.A1(new_n2530), .A2(new_n2531), .B1(new_n2521), .B2(new_n2525), .Y(new_n2913));
  OAI22xp33_ASAP7_75t_L     g02657(.A1(new_n2540), .A2(new_n2504), .B1(new_n2912), .B2(new_n2913), .Y(new_n2914));
  A2O1A1Ixp33_ASAP7_75t_L   g02658(.A1(new_n2914), .A2(new_n2911), .B(new_n2732), .C(new_n2723), .Y(new_n2915));
  NAND2xp33_ASAP7_75t_L     g02659(.A(\b[6] ), .B(new_n1910), .Y(new_n2916));
  NAND2xp33_ASAP7_75t_L     g02660(.A(\b[7] ), .B(new_n1770), .Y(new_n2917));
  AOI22xp33_ASAP7_75t_L     g02661(.A1(new_n1766), .A2(\b[8] ), .B1(new_n1764), .B2(new_n510), .Y(new_n2918));
  NAND4xp25_ASAP7_75t_L     g02662(.A(new_n2918), .B(\a[23] ), .C(new_n2916), .D(new_n2917), .Y(new_n2919));
  OAI221xp5_ASAP7_75t_L     g02663(.A1(new_n1772), .A2(new_n503), .B1(new_n1771), .B2(new_n509), .C(new_n2917), .Y(new_n2920));
  A2O1A1Ixp33_ASAP7_75t_L   g02664(.A1(\b[6] ), .A2(new_n1910), .B(new_n2920), .C(new_n1761), .Y(new_n2921));
  OAI21xp33_ASAP7_75t_L     g02665(.A1(new_n2713), .A2(new_n2714), .B(new_n2711), .Y(new_n2922));
  NAND2xp33_ASAP7_75t_L     g02666(.A(\b[3] ), .B(new_n2386), .Y(new_n2923));
  NAND2xp33_ASAP7_75t_L     g02667(.A(\b[4] ), .B(new_n2232), .Y(new_n2924));
  AOI32xp33_ASAP7_75t_L     g02668(.A1(new_n358), .A2(new_n356), .A3(new_n2226), .B1(\b[5] ), .B2(new_n2228), .Y(new_n2925));
  NAND3xp33_ASAP7_75t_L     g02669(.A(new_n2925), .B(new_n2924), .C(new_n2923), .Y(new_n2926));
  NOR2xp33_ASAP7_75t_L      g02670(.A(new_n2223), .B(new_n2926), .Y(new_n2927));
  INVx1_ASAP7_75t_L         g02671(.A(new_n2927), .Y(new_n2928));
  NAND2xp33_ASAP7_75t_L     g02672(.A(new_n2223), .B(new_n2926), .Y(new_n2929));
  A2O1A1O1Ixp25_ASAP7_75t_L g02673(.A1(new_n2692), .A2(new_n2511), .B(new_n258), .C(new_n2703), .D(new_n2697), .Y(new_n2930));
  NOR3xp33_ASAP7_75t_L      g02674(.A(new_n2699), .B(new_n2693), .C(new_n2705), .Y(new_n2931));
  INVx1_ASAP7_75t_L         g02675(.A(new_n2931), .Y(new_n2932));
  NOR2xp33_ASAP7_75t_L      g02676(.A(new_n258), .B(new_n2932), .Y(new_n2933));
  NAND2xp33_ASAP7_75t_L     g02677(.A(\b[1] ), .B(new_n2706), .Y(new_n2934));
  OAI221xp5_ASAP7_75t_L     g02678(.A1(new_n2707), .A2(new_n283), .B1(new_n278), .B2(new_n2708), .C(new_n2934), .Y(new_n2935));
  NOR3xp33_ASAP7_75t_L      g02679(.A(new_n2930), .B(new_n2933), .C(new_n2935), .Y(new_n2936));
  A2O1A1Ixp33_ASAP7_75t_L   g02680(.A1(\b[0] ), .A2(new_n2931), .B(new_n2935), .C(new_n2930), .Y(new_n2937));
  INVx1_ASAP7_75t_L         g02681(.A(new_n2937), .Y(new_n2938));
  OAI211xp5_ASAP7_75t_L     g02682(.A1(new_n2936), .A2(new_n2938), .B(new_n2928), .C(new_n2929), .Y(new_n2939));
  INVx1_ASAP7_75t_L         g02683(.A(new_n2929), .Y(new_n2940));
  INVx1_ASAP7_75t_L         g02684(.A(new_n2936), .Y(new_n2941));
  OAI211xp5_ASAP7_75t_L     g02685(.A1(new_n2927), .A2(new_n2940), .B(new_n2941), .C(new_n2937), .Y(new_n2942));
  NAND4xp25_ASAP7_75t_L     g02686(.A(new_n2717), .B(new_n2942), .C(new_n2939), .D(new_n2922), .Y(new_n2943));
  INVx1_ASAP7_75t_L         g02687(.A(new_n2922), .Y(new_n2944));
  AOI211xp5_ASAP7_75t_L     g02688(.A1(new_n2941), .A2(new_n2937), .B(new_n2927), .C(new_n2940), .Y(new_n2945));
  AOI211xp5_ASAP7_75t_L     g02689(.A1(new_n2928), .A2(new_n2929), .B(new_n2936), .C(new_n2938), .Y(new_n2946));
  OAI22xp33_ASAP7_75t_L     g02690(.A1(new_n2725), .A2(new_n2944), .B1(new_n2946), .B2(new_n2945), .Y(new_n2947));
  NAND4xp25_ASAP7_75t_L     g02691(.A(new_n2943), .B(new_n2919), .C(new_n2947), .D(new_n2921), .Y(new_n2948));
  AOI22xp33_ASAP7_75t_L     g02692(.A1(new_n2919), .A2(new_n2921), .B1(new_n2947), .B2(new_n2943), .Y(new_n2949));
  INVx1_ASAP7_75t_L         g02693(.A(new_n2949), .Y(new_n2950));
  NAND3xp33_ASAP7_75t_L     g02694(.A(new_n2915), .B(new_n2950), .C(new_n2948), .Y(new_n2951));
  INVx1_ASAP7_75t_L         g02695(.A(new_n2543), .Y(new_n2952));
  A2O1A1O1Ixp25_ASAP7_75t_L g02696(.A1(new_n2542), .A2(new_n2952), .B(new_n2729), .C(new_n2727), .D(new_n2731), .Y(new_n2953));
  INVx1_ASAP7_75t_L         g02697(.A(new_n2948), .Y(new_n2954));
  OAI21xp33_ASAP7_75t_L     g02698(.A1(new_n2949), .A2(new_n2954), .B(new_n2953), .Y(new_n2955));
  AOI21xp33_ASAP7_75t_L     g02699(.A1(new_n2955), .A2(new_n2951), .B(new_n2910), .Y(new_n2956));
  NOR3xp33_ASAP7_75t_L      g02700(.A(new_n2953), .B(new_n2954), .C(new_n2949), .Y(new_n2957));
  AOI21xp33_ASAP7_75t_L     g02701(.A1(new_n2950), .A2(new_n2948), .B(new_n2915), .Y(new_n2958));
  NOR3xp33_ASAP7_75t_L      g02702(.A(new_n2957), .B(new_n2958), .C(new_n2909), .Y(new_n2959));
  NOR3xp33_ASAP7_75t_L      g02703(.A(new_n2902), .B(new_n2956), .C(new_n2959), .Y(new_n2960));
  NAND2xp33_ASAP7_75t_L     g02704(.A(new_n2728), .B(new_n2733), .Y(new_n2961));
  MAJIxp5_ASAP7_75t_L       g02705(.A(new_n2745), .B(new_n2748), .C(new_n2961), .Y(new_n2962));
  OAI21xp33_ASAP7_75t_L     g02706(.A1(new_n2958), .A2(new_n2957), .B(new_n2909), .Y(new_n2963));
  NAND3xp33_ASAP7_75t_L     g02707(.A(new_n2910), .B(new_n2951), .C(new_n2955), .Y(new_n2964));
  AOI21xp33_ASAP7_75t_L     g02708(.A1(new_n2964), .A2(new_n2963), .B(new_n2962), .Y(new_n2965));
  NAND2xp33_ASAP7_75t_L     g02709(.A(\b[12] ), .B(new_n1194), .Y(new_n2966));
  NAND2xp33_ASAP7_75t_L     g02710(.A(\b[13] ), .B(new_n1103), .Y(new_n2967));
  AOI32xp33_ASAP7_75t_L     g02711(.A1(new_n877), .A2(new_n874), .A3(new_n1110), .B1(\b[14] ), .B2(new_n1113), .Y(new_n2968));
  NAND4xp25_ASAP7_75t_L     g02712(.A(new_n2968), .B(\a[17] ), .C(new_n2966), .D(new_n2967), .Y(new_n2969));
  NAND2xp33_ASAP7_75t_L     g02713(.A(new_n2967), .B(new_n2968), .Y(new_n2970));
  A2O1A1Ixp33_ASAP7_75t_L   g02714(.A1(\b[12] ), .A2(new_n1194), .B(new_n2970), .C(new_n1107), .Y(new_n2971));
  NAND2xp33_ASAP7_75t_L     g02715(.A(new_n2969), .B(new_n2971), .Y(new_n2972));
  OR3x1_ASAP7_75t_L         g02716(.A(new_n2960), .B(new_n2965), .C(new_n2972), .Y(new_n2973));
  OAI21xp33_ASAP7_75t_L     g02717(.A1(new_n2965), .A2(new_n2960), .B(new_n2972), .Y(new_n2974));
  NAND3xp33_ASAP7_75t_L     g02718(.A(new_n2761), .B(new_n2751), .C(new_n2746), .Y(new_n2975));
  AO21x2_ASAP7_75t_L        g02719(.A1(new_n2758), .A2(new_n2762), .B(new_n2766), .Y(new_n2976));
  NAND4xp25_ASAP7_75t_L     g02720(.A(new_n2976), .B(new_n2973), .C(new_n2974), .D(new_n2975), .Y(new_n2977));
  NOR3xp33_ASAP7_75t_L      g02721(.A(new_n2960), .B(new_n2965), .C(new_n2972), .Y(new_n2978));
  OA21x2_ASAP7_75t_L        g02722(.A1(new_n2965), .A2(new_n2960), .B(new_n2972), .Y(new_n2979));
  A2O1A1Ixp33_ASAP7_75t_L   g02723(.A1(new_n2762), .A2(new_n2758), .B(new_n2766), .C(new_n2975), .Y(new_n2980));
  OAI21xp33_ASAP7_75t_L     g02724(.A1(new_n2978), .A2(new_n2979), .B(new_n2980), .Y(new_n2981));
  NAND2xp33_ASAP7_75t_L     g02725(.A(\b[15] ), .B(new_n908), .Y(new_n2982));
  NAND2xp33_ASAP7_75t_L     g02726(.A(\b[16] ), .B(new_n817), .Y(new_n2983));
  AOI32xp33_ASAP7_75t_L     g02727(.A1(new_n1250), .A2(new_n1247), .A3(new_n823), .B1(new_n826), .B2(\b[17] ), .Y(new_n2984));
  NAND4xp25_ASAP7_75t_L     g02728(.A(new_n2984), .B(\a[14] ), .C(new_n2982), .D(new_n2983), .Y(new_n2985));
  OAI221xp5_ASAP7_75t_L     g02729(.A1(new_n912), .A2(new_n1244), .B1(new_n911), .B2(new_n1251), .C(new_n2983), .Y(new_n2986));
  A2O1A1Ixp33_ASAP7_75t_L   g02730(.A1(\b[15] ), .A2(new_n908), .B(new_n2986), .C(new_n813), .Y(new_n2987));
  AND2x2_ASAP7_75t_L        g02731(.A(new_n2985), .B(new_n2987), .Y(new_n2988));
  NAND3xp33_ASAP7_75t_L     g02732(.A(new_n2977), .B(new_n2988), .C(new_n2981), .Y(new_n2989));
  NOR3xp33_ASAP7_75t_L      g02733(.A(new_n2980), .B(new_n2979), .C(new_n2978), .Y(new_n2990));
  AOI22xp33_ASAP7_75t_L     g02734(.A1(new_n2973), .A2(new_n2974), .B1(new_n2975), .B2(new_n2976), .Y(new_n2991));
  NAND2xp33_ASAP7_75t_L     g02735(.A(new_n2985), .B(new_n2987), .Y(new_n2992));
  OAI21xp33_ASAP7_75t_L     g02736(.A1(new_n2990), .A2(new_n2991), .B(new_n2992), .Y(new_n2993));
  NAND2xp33_ASAP7_75t_L     g02737(.A(new_n2989), .B(new_n2993), .Y(new_n2994));
  OAI21xp33_ASAP7_75t_L     g02738(.A1(new_n2783), .A2(new_n2781), .B(new_n2775), .Y(new_n2995));
  NOR2xp33_ASAP7_75t_L      g02739(.A(new_n2995), .B(new_n2994), .Y(new_n2996));
  A2O1A1O1Ixp25_ASAP7_75t_L g02740(.A1(new_n2601), .A2(new_n2591), .B(new_n2671), .C(new_n2778), .D(new_n2782), .Y(new_n2997));
  AOI21xp33_ASAP7_75t_L     g02741(.A1(new_n2993), .A2(new_n2989), .B(new_n2997), .Y(new_n2998));
  NOR2xp33_ASAP7_75t_L      g02742(.A(new_n1356), .B(new_n1620), .Y(new_n2999));
  NAND2xp33_ASAP7_75t_L     g02743(.A(new_n1597), .B(new_n1706), .Y(new_n3000));
  NAND2xp33_ASAP7_75t_L     g02744(.A(new_n3000), .B(new_n1991), .Y(new_n3001));
  NAND2xp33_ASAP7_75t_L     g02745(.A(\b[19] ), .B(new_n590), .Y(new_n3002));
  OAI221xp5_ASAP7_75t_L     g02746(.A1(new_n676), .A2(new_n1594), .B1(new_n675), .B2(new_n3001), .C(new_n3002), .Y(new_n3003));
  NOR3xp33_ASAP7_75t_L      g02747(.A(new_n3003), .B(new_n2999), .C(new_n594), .Y(new_n3004));
  INVx1_ASAP7_75t_L         g02748(.A(new_n2999), .Y(new_n3005));
  AOI22xp33_ASAP7_75t_L     g02749(.A1(new_n600), .A2(\b[20] ), .B1(new_n597), .B2(new_n1600), .Y(new_n3006));
  AOI31xp33_ASAP7_75t_L     g02750(.A1(new_n3006), .A2(new_n3002), .A3(new_n3005), .B(\a[11] ), .Y(new_n3007));
  NOR2xp33_ASAP7_75t_L      g02751(.A(new_n3007), .B(new_n3004), .Y(new_n3008));
  OAI21xp33_ASAP7_75t_L     g02752(.A1(new_n2998), .A2(new_n2996), .B(new_n3008), .Y(new_n3009));
  NAND3xp33_ASAP7_75t_L     g02753(.A(new_n2997), .B(new_n2993), .C(new_n2989), .Y(new_n3010));
  A2O1A1Ixp33_ASAP7_75t_L   g02754(.A1(new_n2778), .A2(new_n2800), .B(new_n2782), .C(new_n2994), .Y(new_n3011));
  OR2x4_ASAP7_75t_L         g02755(.A(new_n3007), .B(new_n3004), .Y(new_n3012));
  NAND3xp33_ASAP7_75t_L     g02756(.A(new_n3012), .B(new_n3011), .C(new_n3010), .Y(new_n3013));
  NAND2xp33_ASAP7_75t_L     g02757(.A(new_n3009), .B(new_n3013), .Y(new_n3014));
  NOR3xp33_ASAP7_75t_L      g02758(.A(new_n2899), .B(new_n2900), .C(new_n3014), .Y(new_n3015));
  INVx1_ASAP7_75t_L         g02759(.A(new_n2900), .Y(new_n3016));
  AOI21xp33_ASAP7_75t_L     g02760(.A1(new_n3011), .A2(new_n3010), .B(new_n3012), .Y(new_n3017));
  NOR3xp33_ASAP7_75t_L      g02761(.A(new_n2996), .B(new_n2998), .C(new_n3008), .Y(new_n3018));
  NOR2xp33_ASAP7_75t_L      g02762(.A(new_n3018), .B(new_n3017), .Y(new_n3019));
  A2O1A1O1Ixp25_ASAP7_75t_L g02763(.A1(new_n2608), .A2(new_n2810), .B(new_n2807), .C(new_n3016), .D(new_n3019), .Y(new_n3020));
  OAI21xp33_ASAP7_75t_L     g02764(.A1(new_n3015), .A2(new_n3020), .B(new_n2898), .Y(new_n3021));
  MAJIxp5_ASAP7_75t_L       g02765(.A(new_n2606), .B(new_n2598), .C(new_n2808), .Y(new_n3022));
  O2A1O1Ixp33_ASAP7_75t_L   g02766(.A1(new_n2797), .A2(new_n2806), .B(new_n3022), .C(new_n2900), .Y(new_n3023));
  NAND2xp33_ASAP7_75t_L     g02767(.A(new_n3023), .B(new_n3019), .Y(new_n3024));
  A2O1A1Ixp33_ASAP7_75t_L   g02768(.A1(new_n3022), .A2(new_n2814), .B(new_n2900), .C(new_n3014), .Y(new_n3025));
  NAND3xp33_ASAP7_75t_L     g02769(.A(new_n3025), .B(new_n3024), .C(new_n2897), .Y(new_n3026));
  NAND3xp33_ASAP7_75t_L     g02770(.A(new_n2894), .B(new_n3021), .C(new_n3026), .Y(new_n3027));
  OA21x2_ASAP7_75t_L        g02771(.A1(new_n2893), .A2(new_n2824), .B(new_n2823), .Y(new_n3028));
  AOI21xp33_ASAP7_75t_L     g02772(.A1(new_n3025), .A2(new_n3024), .B(new_n2897), .Y(new_n3029));
  NOR3xp33_ASAP7_75t_L      g02773(.A(new_n3020), .B(new_n3015), .C(new_n2898), .Y(new_n3030));
  OAI21xp33_ASAP7_75t_L     g02774(.A1(new_n3029), .A2(new_n3030), .B(new_n3028), .Y(new_n3031));
  AOI21xp33_ASAP7_75t_L     g02775(.A1(new_n3031), .A2(new_n3027), .B(new_n2892), .Y(new_n3032));
  NAND3xp33_ASAP7_75t_L     g02776(.A(new_n3031), .B(new_n3027), .C(new_n2892), .Y(new_n3033));
  INVx1_ASAP7_75t_L         g02777(.A(new_n3033), .Y(new_n3034));
  NOR2xp33_ASAP7_75t_L      g02778(.A(new_n3032), .B(new_n3034), .Y(new_n3035));
  O2A1O1Ixp33_ASAP7_75t_L   g02779(.A1(new_n2885), .A2(new_n2837), .B(new_n2849), .C(new_n3035), .Y(new_n3036));
  MAJIxp5_ASAP7_75t_L       g02780(.A(new_n2845), .B(new_n2885), .C(new_n2837), .Y(new_n3037));
  INVx1_ASAP7_75t_L         g02781(.A(new_n3032), .Y(new_n3038));
  NAND2xp33_ASAP7_75t_L     g02782(.A(new_n3033), .B(new_n3038), .Y(new_n3039));
  NOR2xp33_ASAP7_75t_L      g02783(.A(new_n3039), .B(new_n3037), .Y(new_n3040));
  NOR3xp33_ASAP7_75t_L      g02784(.A(new_n3036), .B(new_n3040), .C(new_n2884), .Y(new_n3041));
  INVx1_ASAP7_75t_L         g02785(.A(new_n3041), .Y(new_n3042));
  OAI21xp33_ASAP7_75t_L     g02786(.A1(new_n3040), .A2(new_n3036), .B(new_n2884), .Y(new_n3043));
  NAND2xp33_ASAP7_75t_L     g02787(.A(new_n3043), .B(new_n3042), .Y(new_n3044));
  XOR2x2_ASAP7_75t_L        g02788(.A(new_n2870), .B(new_n3044), .Y(\f[29] ));
  NAND3xp33_ASAP7_75t_L     g02789(.A(new_n2826), .B(new_n2828), .C(new_n2836), .Y(new_n3046));
  INVx1_ASAP7_75t_L         g02790(.A(new_n3046), .Y(new_n3047));
  A2O1A1Ixp33_ASAP7_75t_L   g02791(.A1(new_n2846), .A2(new_n2842), .B(new_n3047), .C(new_n3039), .Y(new_n3048));
  AOI21xp33_ASAP7_75t_L     g02792(.A1(new_n2894), .A2(new_n3026), .B(new_n3029), .Y(new_n3049));
  NAND2xp33_ASAP7_75t_L     g02793(.A(new_n2743), .B(new_n2901), .Y(new_n3050));
  A2O1A1Ixp33_ASAP7_75t_L   g02794(.A1(new_n2751), .A2(new_n3050), .B(new_n2956), .C(new_n2964), .Y(new_n3051));
  NOR2xp33_ASAP7_75t_L      g02795(.A(new_n631), .B(new_n1549), .Y(new_n3052));
  INVx1_ASAP7_75t_L         g02796(.A(new_n3052), .Y(new_n3053));
  NAND2xp33_ASAP7_75t_L     g02797(.A(\b[11] ), .B(new_n1410), .Y(new_n3054));
  AOI32xp33_ASAP7_75t_L     g02798(.A1(new_n771), .A2(new_n774), .A3(new_n1404), .B1(new_n1406), .B2(\b[12] ), .Y(new_n3055));
  NAND4xp25_ASAP7_75t_L     g02799(.A(new_n3055), .B(\a[20] ), .C(new_n3053), .D(new_n3054), .Y(new_n3056));
  NAND2xp33_ASAP7_75t_L     g02800(.A(new_n3054), .B(new_n3055), .Y(new_n3057));
  A2O1A1Ixp33_ASAP7_75t_L   g02801(.A1(\b[10] ), .A2(new_n1548), .B(new_n3057), .C(new_n1401), .Y(new_n3058));
  A2O1A1O1Ixp25_ASAP7_75t_L g02802(.A1(new_n2727), .A2(new_n2674), .B(new_n2731), .C(new_n2948), .D(new_n2949), .Y(new_n3059));
  NAND2xp33_ASAP7_75t_L     g02803(.A(\b[0] ), .B(new_n2706), .Y(new_n3060));
  NAND4xp25_ASAP7_75t_L     g02804(.A(new_n2703), .B(\a[29] ), .C(new_n2719), .D(new_n3060), .Y(new_n3061));
  INVx1_ASAP7_75t_L         g02805(.A(\a[30] ), .Y(new_n3062));
  NAND2xp33_ASAP7_75t_L     g02806(.A(\a[29] ), .B(new_n3062), .Y(new_n3063));
  NAND2xp33_ASAP7_75t_L     g02807(.A(\a[30] ), .B(new_n2697), .Y(new_n3064));
  AND2x2_ASAP7_75t_L        g02808(.A(new_n3063), .B(new_n3064), .Y(new_n3065));
  NOR2xp33_ASAP7_75t_L      g02809(.A(new_n258), .B(new_n3065), .Y(new_n3066));
  OAI31xp33_ASAP7_75t_L     g02810(.A1(new_n3061), .A2(new_n2935), .A3(new_n2933), .B(new_n3066), .Y(new_n3067));
  OR4x2_ASAP7_75t_L         g02811(.A(new_n3066), .B(new_n3061), .C(new_n2935), .D(new_n2933), .Y(new_n3068));
  NOR2xp33_ASAP7_75t_L      g02812(.A(new_n278), .B(new_n2694), .Y(new_n3069));
  AOI221xp5_ASAP7_75t_L     g02813(.A1(new_n2702), .A2(\b[3] ), .B1(new_n2700), .B2(new_n1000), .C(new_n3069), .Y(new_n3070));
  OAI211xp5_ASAP7_75t_L     g02814(.A1(new_n276), .A2(new_n2932), .B(new_n3070), .C(\a[29] ), .Y(new_n3071));
  NAND2xp33_ASAP7_75t_L     g02815(.A(\b[3] ), .B(new_n2702), .Y(new_n3072));
  OAI221xp5_ASAP7_75t_L     g02816(.A1(new_n278), .A2(new_n2694), .B1(new_n2707), .B2(new_n303), .C(new_n3072), .Y(new_n3073));
  A2O1A1Ixp33_ASAP7_75t_L   g02817(.A1(\b[1] ), .A2(new_n2931), .B(new_n3073), .C(new_n2697), .Y(new_n3074));
  AO22x1_ASAP7_75t_L        g02818(.A1(new_n3074), .A2(new_n3071), .B1(new_n3067), .B2(new_n3068), .Y(new_n3075));
  NAND4xp25_ASAP7_75t_L     g02819(.A(new_n3068), .B(new_n3067), .C(new_n3071), .D(new_n3074), .Y(new_n3076));
  NAND2xp33_ASAP7_75t_L     g02820(.A(\b[4] ), .B(new_n2386), .Y(new_n3077));
  NAND2xp33_ASAP7_75t_L     g02821(.A(\b[5] ), .B(new_n2232), .Y(new_n3078));
  AOI22xp33_ASAP7_75t_L     g02822(.A1(new_n2228), .A2(\b[6] ), .B1(new_n2226), .B2(new_n389), .Y(new_n3079));
  NAND4xp25_ASAP7_75t_L     g02823(.A(new_n3079), .B(\a[26] ), .C(new_n3077), .D(new_n3078), .Y(new_n3080));
  OAI221xp5_ASAP7_75t_L     g02824(.A1(new_n2234), .A2(new_n382), .B1(new_n2233), .B2(new_n540), .C(new_n3078), .Y(new_n3081));
  A2O1A1Ixp33_ASAP7_75t_L   g02825(.A1(\b[4] ), .A2(new_n2386), .B(new_n3081), .C(new_n2223), .Y(new_n3082));
  NAND4xp25_ASAP7_75t_L     g02826(.A(new_n3082), .B(new_n3075), .C(new_n3076), .D(new_n3080), .Y(new_n3083));
  AOI22xp33_ASAP7_75t_L     g02827(.A1(new_n3071), .A2(new_n3074), .B1(new_n3067), .B2(new_n3068), .Y(new_n3084));
  AND4x1_ASAP7_75t_L        g02828(.A(new_n3068), .B(new_n3067), .C(new_n3074), .D(new_n3071), .Y(new_n3085));
  INVx1_ASAP7_75t_L         g02829(.A(new_n3080), .Y(new_n3086));
  AOI31xp33_ASAP7_75t_L     g02830(.A1(new_n3079), .A2(new_n3078), .A3(new_n3077), .B(\a[26] ), .Y(new_n3087));
  OAI22xp33_ASAP7_75t_L     g02831(.A1(new_n3086), .A2(new_n3087), .B1(new_n3084), .B2(new_n3085), .Y(new_n3088));
  A2O1A1O1Ixp25_ASAP7_75t_L g02832(.A1(new_n2712), .A2(new_n2716), .B(new_n2721), .C(new_n2922), .D(new_n2945), .Y(new_n3089));
  OAI211xp5_ASAP7_75t_L     g02833(.A1(new_n2946), .A2(new_n3089), .B(new_n3083), .C(new_n3088), .Y(new_n3090));
  NAND2xp33_ASAP7_75t_L     g02834(.A(new_n3083), .B(new_n3088), .Y(new_n3091));
  A2O1A1Ixp33_ASAP7_75t_L   g02835(.A1(new_n2523), .A2(new_n2522), .B(new_n2524), .C(new_n2682), .Y(new_n3092));
  NAND2xp33_ASAP7_75t_L     g02836(.A(new_n2712), .B(new_n2716), .Y(new_n3093));
  A2O1A1O1Ixp25_ASAP7_75t_L g02837(.A1(new_n3092), .A2(new_n3093), .B(new_n2944), .C(new_n2939), .D(new_n2946), .Y(new_n3094));
  NAND2xp33_ASAP7_75t_L     g02838(.A(new_n3094), .B(new_n3091), .Y(new_n3095));
  NOR2xp33_ASAP7_75t_L      g02839(.A(new_n421), .B(new_n1911), .Y(new_n3096));
  NAND2xp33_ASAP7_75t_L     g02840(.A(\b[8] ), .B(new_n1770), .Y(new_n3097));
  OAI221xp5_ASAP7_75t_L     g02841(.A1(new_n1772), .A2(new_n559), .B1(new_n1771), .B2(new_n978), .C(new_n3097), .Y(new_n3098));
  OR3x1_ASAP7_75t_L         g02842(.A(new_n3098), .B(new_n1761), .C(new_n3096), .Y(new_n3099));
  A2O1A1Ixp33_ASAP7_75t_L   g02843(.A1(\b[7] ), .A2(new_n1910), .B(new_n3098), .C(new_n1761), .Y(new_n3100));
  AOI22xp33_ASAP7_75t_L     g02844(.A1(new_n3099), .A2(new_n3100), .B1(new_n3090), .B2(new_n3095), .Y(new_n3101));
  AND4x1_ASAP7_75t_L        g02845(.A(new_n3095), .B(new_n3090), .C(new_n3100), .D(new_n3099), .Y(new_n3102));
  NOR3xp33_ASAP7_75t_L      g02846(.A(new_n3059), .B(new_n3102), .C(new_n3101), .Y(new_n3103));
  OA21x2_ASAP7_75t_L        g02847(.A1(new_n3101), .A2(new_n3102), .B(new_n3059), .Y(new_n3104));
  OAI211xp5_ASAP7_75t_L     g02848(.A1(new_n3103), .A2(new_n3104), .B(new_n3058), .C(new_n3056), .Y(new_n3105));
  INVx1_ASAP7_75t_L         g02849(.A(new_n3056), .Y(new_n3106));
  INVx1_ASAP7_75t_L         g02850(.A(new_n3058), .Y(new_n3107));
  INVx1_ASAP7_75t_L         g02851(.A(new_n3103), .Y(new_n3108));
  OAI21xp33_ASAP7_75t_L     g02852(.A1(new_n3101), .A2(new_n3102), .B(new_n3059), .Y(new_n3109));
  OAI211xp5_ASAP7_75t_L     g02853(.A1(new_n3107), .A2(new_n3106), .B(new_n3108), .C(new_n3109), .Y(new_n3110));
  NAND3xp33_ASAP7_75t_L     g02854(.A(new_n3051), .B(new_n3105), .C(new_n3110), .Y(new_n3111));
  NOR2xp33_ASAP7_75t_L      g02855(.A(new_n2748), .B(new_n2961), .Y(new_n3112));
  O2A1O1Ixp33_ASAP7_75t_L   g02856(.A1(new_n3112), .A2(new_n2760), .B(new_n2963), .C(new_n2959), .Y(new_n3113));
  AOI211xp5_ASAP7_75t_L     g02857(.A1(new_n3108), .A2(new_n3109), .B(new_n3107), .C(new_n3106), .Y(new_n3114));
  AOI211xp5_ASAP7_75t_L     g02858(.A1(new_n3056), .A2(new_n3058), .B(new_n3103), .C(new_n3104), .Y(new_n3115));
  OAI21xp33_ASAP7_75t_L     g02859(.A1(new_n3115), .A2(new_n3114), .B(new_n3113), .Y(new_n3116));
  NOR2xp33_ASAP7_75t_L      g02860(.A(new_n793), .B(new_n1195), .Y(new_n3117));
  NAND2xp33_ASAP7_75t_L     g02861(.A(\b[14] ), .B(new_n1103), .Y(new_n3118));
  OAI221xp5_ASAP7_75t_L     g02862(.A1(new_n1198), .A2(new_n952), .B1(new_n1197), .B2(new_n2573), .C(new_n3118), .Y(new_n3119));
  NOR3xp33_ASAP7_75t_L      g02863(.A(new_n3119), .B(new_n3117), .C(new_n1107), .Y(new_n3120));
  INVx1_ASAP7_75t_L         g02864(.A(new_n3117), .Y(new_n3121));
  AOI22xp33_ASAP7_75t_L     g02865(.A1(new_n1113), .A2(\b[15] ), .B1(new_n1110), .B2(new_n959), .Y(new_n3122));
  AOI31xp33_ASAP7_75t_L     g02866(.A1(new_n3122), .A2(new_n3118), .A3(new_n3121), .B(\a[17] ), .Y(new_n3123));
  NOR2xp33_ASAP7_75t_L      g02867(.A(new_n3120), .B(new_n3123), .Y(new_n3124));
  NAND3xp33_ASAP7_75t_L     g02868(.A(new_n3111), .B(new_n3116), .C(new_n3124), .Y(new_n3125));
  AO21x2_ASAP7_75t_L        g02869(.A1(new_n3116), .A2(new_n3111), .B(new_n3124), .Y(new_n3126));
  NOR2xp33_ASAP7_75t_L      g02870(.A(new_n2965), .B(new_n2960), .Y(new_n3127));
  NAND2xp33_ASAP7_75t_L     g02871(.A(new_n2972), .B(new_n3127), .Y(new_n3128));
  AND4x1_ASAP7_75t_L        g02872(.A(new_n2981), .B(new_n3128), .C(new_n3126), .D(new_n3125), .Y(new_n3129));
  MAJIxp5_ASAP7_75t_L       g02873(.A(new_n2980), .B(new_n2972), .C(new_n3127), .Y(new_n3130));
  AOI21xp33_ASAP7_75t_L     g02874(.A1(new_n3126), .A2(new_n3125), .B(new_n3130), .Y(new_n3131));
  NOR2xp33_ASAP7_75t_L      g02875(.A(new_n1356), .B(new_n912), .Y(new_n3132));
  AOI221xp5_ASAP7_75t_L     g02876(.A1(new_n817), .A2(\b[17] ), .B1(new_n823), .B2(new_n1363), .C(new_n3132), .Y(new_n3133));
  OAI211xp5_ASAP7_75t_L     g02877(.A1(new_n1051), .A2(new_n909), .B(new_n3133), .C(\a[14] ), .Y(new_n3134));
  A2O1A1Ixp33_ASAP7_75t_L   g02878(.A1(new_n2790), .A2(new_n1246), .B(new_n1245), .C(new_n1358), .Y(new_n3135));
  A2O1A1O1Ixp25_ASAP7_75t_L g02879(.A1(new_n1053), .A2(new_n1056), .B(new_n1052), .C(new_n1246), .D(new_n1245), .Y(new_n3136));
  NAND2xp33_ASAP7_75t_L     g02880(.A(new_n1359), .B(new_n3136), .Y(new_n3137));
  NAND2xp33_ASAP7_75t_L     g02881(.A(new_n3137), .B(new_n3135), .Y(new_n3138));
  INVx1_ASAP7_75t_L         g02882(.A(new_n3132), .Y(new_n3139));
  OAI221xp5_ASAP7_75t_L     g02883(.A1(new_n1244), .A2(new_n994), .B1(new_n911), .B2(new_n3138), .C(new_n3139), .Y(new_n3140));
  A2O1A1Ixp33_ASAP7_75t_L   g02884(.A1(\b[16] ), .A2(new_n908), .B(new_n3140), .C(new_n813), .Y(new_n3141));
  NAND2xp33_ASAP7_75t_L     g02885(.A(new_n3141), .B(new_n3134), .Y(new_n3142));
  NOR3xp33_ASAP7_75t_L      g02886(.A(new_n3129), .B(new_n3131), .C(new_n3142), .Y(new_n3143));
  NAND3xp33_ASAP7_75t_L     g02887(.A(new_n3130), .B(new_n3126), .C(new_n3125), .Y(new_n3144));
  AO22x1_ASAP7_75t_L        g02888(.A1(new_n3125), .A2(new_n3126), .B1(new_n3128), .B2(new_n2981), .Y(new_n3145));
  AND2x2_ASAP7_75t_L        g02889(.A(new_n3141), .B(new_n3134), .Y(new_n3146));
  AOI21xp33_ASAP7_75t_L     g02890(.A1(new_n3145), .A2(new_n3144), .B(new_n3146), .Y(new_n3147));
  NOR2xp33_ASAP7_75t_L      g02891(.A(new_n3143), .B(new_n3147), .Y(new_n3148));
  NAND3xp33_ASAP7_75t_L     g02892(.A(new_n2977), .B(new_n2981), .C(new_n2992), .Y(new_n3149));
  INVx1_ASAP7_75t_L         g02893(.A(new_n3149), .Y(new_n3150));
  AOI21xp33_ASAP7_75t_L     g02894(.A1(new_n2994), .A2(new_n2995), .B(new_n3150), .Y(new_n3151));
  NAND2xp33_ASAP7_75t_L     g02895(.A(new_n3148), .B(new_n3151), .Y(new_n3152));
  NAND3xp33_ASAP7_75t_L     g02896(.A(new_n3145), .B(new_n3146), .C(new_n3144), .Y(new_n3153));
  OAI21xp33_ASAP7_75t_L     g02897(.A1(new_n3131), .A2(new_n3129), .B(new_n3142), .Y(new_n3154));
  NAND2xp33_ASAP7_75t_L     g02898(.A(new_n3154), .B(new_n3153), .Y(new_n3155));
  A2O1A1Ixp33_ASAP7_75t_L   g02899(.A1(new_n2994), .A2(new_n2995), .B(new_n3150), .C(new_n3155), .Y(new_n3156));
  NAND2xp33_ASAP7_75t_L     g02900(.A(\b[19] ), .B(new_n674), .Y(new_n3157));
  NAND2xp33_ASAP7_75t_L     g02901(.A(\b[20] ), .B(new_n590), .Y(new_n3158));
  AOI22xp33_ASAP7_75t_L     g02902(.A1(new_n600), .A2(\b[21] ), .B1(new_n597), .B2(new_n1715), .Y(new_n3159));
  NAND4xp25_ASAP7_75t_L     g02903(.A(new_n3159), .B(\a[11] ), .C(new_n3157), .D(new_n3158), .Y(new_n3160));
  NAND2xp33_ASAP7_75t_L     g02904(.A(new_n3158), .B(new_n3159), .Y(new_n3161));
  A2O1A1Ixp33_ASAP7_75t_L   g02905(.A1(\b[19] ), .A2(new_n674), .B(new_n3161), .C(new_n594), .Y(new_n3162));
  AND2x2_ASAP7_75t_L        g02906(.A(new_n3160), .B(new_n3162), .Y(new_n3163));
  NAND3xp33_ASAP7_75t_L     g02907(.A(new_n3163), .B(new_n3152), .C(new_n3156), .Y(new_n3164));
  A2O1A1Ixp33_ASAP7_75t_L   g02908(.A1(new_n2993), .A2(new_n2989), .B(new_n2997), .C(new_n3149), .Y(new_n3165));
  NOR2xp33_ASAP7_75t_L      g02909(.A(new_n3165), .B(new_n3155), .Y(new_n3166));
  A2O1A1O1Ixp25_ASAP7_75t_L g02910(.A1(new_n2993), .A2(new_n2989), .B(new_n2997), .C(new_n3149), .D(new_n3148), .Y(new_n3167));
  NAND2xp33_ASAP7_75t_L     g02911(.A(new_n3160), .B(new_n3162), .Y(new_n3168));
  OAI21xp33_ASAP7_75t_L     g02912(.A1(new_n3166), .A2(new_n3167), .B(new_n3168), .Y(new_n3169));
  A2O1A1O1Ixp25_ASAP7_75t_L g02913(.A1(new_n2810), .A2(new_n2608), .B(new_n2807), .C(new_n3016), .D(new_n3017), .Y(new_n3170));
  OAI211xp5_ASAP7_75t_L     g02914(.A1(new_n3018), .A2(new_n3170), .B(new_n3164), .C(new_n3169), .Y(new_n3171));
  NOR3xp33_ASAP7_75t_L      g02915(.A(new_n3167), .B(new_n3168), .C(new_n3166), .Y(new_n3172));
  AOI21xp33_ASAP7_75t_L     g02916(.A1(new_n3152), .A2(new_n3156), .B(new_n3163), .Y(new_n3173));
  A2O1A1O1Ixp25_ASAP7_75t_L g02917(.A1(new_n3022), .A2(new_n2814), .B(new_n2900), .C(new_n3009), .D(new_n3018), .Y(new_n3174));
  OAI21xp33_ASAP7_75t_L     g02918(.A1(new_n3173), .A2(new_n3172), .B(new_n3174), .Y(new_n3175));
  NAND2xp33_ASAP7_75t_L     g02919(.A(\b[22] ), .B(new_n480), .Y(new_n3176));
  NAND2xp33_ASAP7_75t_L     g02920(.A(\b[23] ), .B(new_n441), .Y(new_n3177));
  AOI22xp33_ASAP7_75t_L     g02921(.A1(new_n451), .A2(\b[24] ), .B1(new_n448), .B2(new_n2027), .Y(new_n3178));
  AND4x1_ASAP7_75t_L        g02922(.A(new_n3178), .B(new_n3177), .C(new_n3176), .D(\a[8] ), .Y(new_n3179));
  AOI31xp33_ASAP7_75t_L     g02923(.A1(new_n3178), .A2(new_n3177), .A3(new_n3176), .B(\a[8] ), .Y(new_n3180));
  NOR2xp33_ASAP7_75t_L      g02924(.A(new_n3180), .B(new_n3179), .Y(new_n3181));
  AOI21xp33_ASAP7_75t_L     g02925(.A1(new_n3171), .A2(new_n3175), .B(new_n3181), .Y(new_n3182));
  NAND3xp33_ASAP7_75t_L     g02926(.A(new_n3171), .B(new_n3175), .C(new_n3181), .Y(new_n3183));
  INVx1_ASAP7_75t_L         g02927(.A(new_n3183), .Y(new_n3184));
  OAI21xp33_ASAP7_75t_L     g02928(.A1(new_n3182), .A2(new_n3184), .B(new_n3049), .Y(new_n3185));
  OAI21xp33_ASAP7_75t_L     g02929(.A1(new_n3030), .A2(new_n3028), .B(new_n3021), .Y(new_n3186));
  NOR3xp33_ASAP7_75t_L      g02930(.A(new_n3174), .B(new_n3173), .C(new_n3172), .Y(new_n3187));
  INVx1_ASAP7_75t_L         g02931(.A(new_n3175), .Y(new_n3188));
  INVx1_ASAP7_75t_L         g02932(.A(new_n3181), .Y(new_n3189));
  OAI21xp33_ASAP7_75t_L     g02933(.A1(new_n3187), .A2(new_n3188), .B(new_n3189), .Y(new_n3190));
  NAND3xp33_ASAP7_75t_L     g02934(.A(new_n3186), .B(new_n3190), .C(new_n3183), .Y(new_n3191));
  NAND2xp33_ASAP7_75t_L     g02935(.A(\b[25] ), .B(new_n366), .Y(new_n3192));
  NAND2xp33_ASAP7_75t_L     g02936(.A(\b[26] ), .B(new_n334), .Y(new_n3193));
  AOI22xp33_ASAP7_75t_L     g02937(.A1(new_n345), .A2(\b[27] ), .B1(new_n342), .B2(new_n2657), .Y(new_n3194));
  AND4x1_ASAP7_75t_L        g02938(.A(new_n3194), .B(new_n3193), .C(new_n3192), .D(\a[5] ), .Y(new_n3195));
  AOI31xp33_ASAP7_75t_L     g02939(.A1(new_n3194), .A2(new_n3193), .A3(new_n3192), .B(\a[5] ), .Y(new_n3196));
  NOR2xp33_ASAP7_75t_L      g02940(.A(new_n3196), .B(new_n3195), .Y(new_n3197));
  NAND3xp33_ASAP7_75t_L     g02941(.A(new_n3191), .B(new_n3185), .C(new_n3197), .Y(new_n3198));
  AOI221xp5_ASAP7_75t_L     g02942(.A1(new_n3026), .A2(new_n2894), .B1(new_n3183), .B2(new_n3190), .C(new_n3029), .Y(new_n3199));
  NOR3xp33_ASAP7_75t_L      g02943(.A(new_n3049), .B(new_n3184), .C(new_n3182), .Y(new_n3200));
  OAI22xp33_ASAP7_75t_L     g02944(.A1(new_n3200), .A2(new_n3199), .B1(new_n3196), .B2(new_n3195), .Y(new_n3201));
  AND2x2_ASAP7_75t_L        g02945(.A(new_n3201), .B(new_n3198), .Y(new_n3202));
  INVx1_ASAP7_75t_L         g02946(.A(new_n2892), .Y(new_n3203));
  NAND3xp33_ASAP7_75t_L     g02947(.A(new_n3203), .B(new_n3027), .C(new_n3031), .Y(new_n3204));
  NAND3xp33_ASAP7_75t_L     g02948(.A(new_n3048), .B(new_n3202), .C(new_n3204), .Y(new_n3205));
  NAND2xp33_ASAP7_75t_L     g02949(.A(new_n3201), .B(new_n3198), .Y(new_n3206));
  INVx1_ASAP7_75t_L         g02950(.A(new_n3204), .Y(new_n3207));
  A2O1A1Ixp33_ASAP7_75t_L   g02951(.A1(new_n3037), .A2(new_n3039), .B(new_n3207), .C(new_n3206), .Y(new_n3208));
  NAND2xp33_ASAP7_75t_L     g02952(.A(new_n3208), .B(new_n3205), .Y(new_n3209));
  INVx1_ASAP7_75t_L         g02953(.A(new_n2875), .Y(new_n3210));
  NOR2xp33_ASAP7_75t_L      g02954(.A(\b[29] ), .B(\b[30] ), .Y(new_n3211));
  INVx1_ASAP7_75t_L         g02955(.A(\b[30] ), .Y(new_n3212));
  NOR2xp33_ASAP7_75t_L      g02956(.A(new_n2871), .B(new_n3212), .Y(new_n3213));
  NOR2xp33_ASAP7_75t_L      g02957(.A(new_n3211), .B(new_n3213), .Y(new_n3214));
  INVx1_ASAP7_75t_L         g02958(.A(new_n3214), .Y(new_n3215));
  O2A1O1Ixp33_ASAP7_75t_L   g02959(.A1(new_n2879), .A2(new_n2878), .B(new_n3210), .C(new_n3215), .Y(new_n3216));
  O2A1O1Ixp33_ASAP7_75t_L   g02960(.A1(new_n2650), .A2(new_n2852), .B(new_n2855), .C(new_n2879), .Y(new_n3217));
  NOR3xp33_ASAP7_75t_L      g02961(.A(new_n3217), .B(new_n3214), .C(new_n2875), .Y(new_n3218));
  NOR2xp33_ASAP7_75t_L      g02962(.A(new_n3216), .B(new_n3218), .Y(new_n3219));
  AOI22xp33_ASAP7_75t_L     g02963(.A1(new_n272), .A2(\b[30] ), .B1(new_n269), .B2(new_n3219), .Y(new_n3220));
  OAI221xp5_ASAP7_75t_L     g02964(.A1(new_n261), .A2(new_n2871), .B1(new_n2852), .B2(new_n277), .C(new_n3220), .Y(new_n3221));
  XNOR2x2_ASAP7_75t_L       g02965(.A(\a[2] ), .B(new_n3221), .Y(new_n3222));
  XNOR2x2_ASAP7_75t_L       g02966(.A(new_n3222), .B(new_n3209), .Y(new_n3223));
  O2A1O1Ixp33_ASAP7_75t_L   g02967(.A1(new_n2870), .A2(new_n3044), .B(new_n3042), .C(new_n3223), .Y(new_n3224));
  A2O1A1O1Ixp25_ASAP7_75t_L g02968(.A1(new_n2862), .A2(new_n2867), .B(new_n2863), .C(new_n3043), .D(new_n3041), .Y(new_n3225));
  AND2x2_ASAP7_75t_L        g02969(.A(new_n3225), .B(new_n3223), .Y(new_n3226));
  NOR2xp33_ASAP7_75t_L      g02970(.A(new_n3224), .B(new_n3226), .Y(\f[30] ));
  OAI211xp5_ASAP7_75t_L     g02971(.A1(new_n3087), .A2(new_n3086), .B(new_n3076), .C(new_n3075), .Y(new_n3228));
  A2O1A1Ixp33_ASAP7_75t_L   g02972(.A1(new_n3088), .A2(new_n3083), .B(new_n3094), .C(new_n3228), .Y(new_n3229));
  NAND2xp33_ASAP7_75t_L     g02973(.A(\b[5] ), .B(new_n2386), .Y(new_n3230));
  NAND2xp33_ASAP7_75t_L     g02974(.A(\b[6] ), .B(new_n2232), .Y(new_n3231));
  AOI32xp33_ASAP7_75t_L     g02975(.A1(new_n424), .A2(new_n426), .A3(new_n2226), .B1(new_n2228), .B2(\b[7] ), .Y(new_n3232));
  AND4x1_ASAP7_75t_L        g02976(.A(new_n3232), .B(new_n3231), .C(new_n3230), .D(\a[26] ), .Y(new_n3233));
  AOI31xp33_ASAP7_75t_L     g02977(.A1(new_n3232), .A2(new_n3231), .A3(new_n3230), .B(\a[26] ), .Y(new_n3234));
  NOR3xp33_ASAP7_75t_L      g02978(.A(new_n3061), .B(new_n2933), .C(new_n2935), .Y(new_n3235));
  NAND2xp33_ASAP7_75t_L     g02979(.A(new_n3066), .B(new_n3235), .Y(new_n3236));
  INVx1_ASAP7_75t_L         g02980(.A(new_n3236), .Y(new_n3237));
  NAND2xp33_ASAP7_75t_L     g02981(.A(\b[2] ), .B(new_n2931), .Y(new_n3238));
  INVx1_ASAP7_75t_L         g02982(.A(new_n3238), .Y(new_n3239));
  NOR2xp33_ASAP7_75t_L      g02983(.A(new_n299), .B(new_n2694), .Y(new_n3240));
  OAI32xp33_ASAP7_75t_L     g02984(.A1(new_n325), .A2(new_n327), .A3(new_n2707), .B1(new_n323), .B2(new_n2708), .Y(new_n3241));
  NOR4xp25_ASAP7_75t_L      g02985(.A(new_n3239), .B(new_n3241), .C(new_n2697), .D(new_n3240), .Y(new_n3242));
  OAI31xp33_ASAP7_75t_L     g02986(.A1(new_n3239), .A2(new_n3241), .A3(new_n3240), .B(new_n2697), .Y(new_n3243));
  INVx1_ASAP7_75t_L         g02987(.A(new_n3243), .Y(new_n3244));
  NAND2xp33_ASAP7_75t_L     g02988(.A(\a[32] ), .B(new_n3066), .Y(new_n3245));
  XNOR2x2_ASAP7_75t_L       g02989(.A(\a[31] ), .B(\a[30] ), .Y(new_n3246));
  INVx1_ASAP7_75t_L         g02990(.A(new_n3246), .Y(new_n3247));
  NAND2xp33_ASAP7_75t_L     g02991(.A(new_n3247), .B(new_n3065), .Y(new_n3248));
  INVx1_ASAP7_75t_L         g02992(.A(\a[31] ), .Y(new_n3249));
  NAND2xp33_ASAP7_75t_L     g02993(.A(\a[32] ), .B(new_n3249), .Y(new_n3250));
  INVx1_ASAP7_75t_L         g02994(.A(\a[32] ), .Y(new_n3251));
  NAND2xp33_ASAP7_75t_L     g02995(.A(\a[31] ), .B(new_n3251), .Y(new_n3252));
  AND2x2_ASAP7_75t_L        g02996(.A(new_n3250), .B(new_n3252), .Y(new_n3253));
  NOR2xp33_ASAP7_75t_L      g02997(.A(new_n3065), .B(new_n3253), .Y(new_n3254));
  NAND2xp33_ASAP7_75t_L     g02998(.A(new_n3252), .B(new_n3250), .Y(new_n3255));
  NOR2xp33_ASAP7_75t_L      g02999(.A(new_n3255), .B(new_n3065), .Y(new_n3256));
  AOI22xp33_ASAP7_75t_L     g03000(.A1(new_n3256), .A2(\b[1] ), .B1(new_n271), .B2(new_n3254), .Y(new_n3257));
  O2A1O1Ixp33_ASAP7_75t_L   g03001(.A1(new_n3248), .A2(new_n258), .B(new_n3257), .C(new_n3245), .Y(new_n3258));
  NAND2xp33_ASAP7_75t_L     g03002(.A(new_n3064), .B(new_n3063), .Y(new_n3259));
  NOR2xp33_ASAP7_75t_L      g03003(.A(new_n3246), .B(new_n3259), .Y(new_n3260));
  NAND2xp33_ASAP7_75t_L     g03004(.A(new_n3255), .B(new_n3259), .Y(new_n3261));
  NAND2xp33_ASAP7_75t_L     g03005(.A(new_n3259), .B(new_n3253), .Y(new_n3262));
  OAI22xp33_ASAP7_75t_L     g03006(.A1(new_n3262), .A2(new_n276), .B1(new_n270), .B2(new_n3261), .Y(new_n3263));
  A2O1A1O1Ixp25_ASAP7_75t_L g03007(.A1(new_n3259), .A2(\a[32] ), .B(new_n3260), .C(\b[0] ), .D(new_n3263), .Y(new_n3264));
  OR2x4_ASAP7_75t_L         g03008(.A(new_n3264), .B(new_n3258), .Y(new_n3265));
  NOR3xp33_ASAP7_75t_L      g03009(.A(new_n3265), .B(new_n3244), .C(new_n3242), .Y(new_n3266));
  INVx1_ASAP7_75t_L         g03010(.A(new_n3242), .Y(new_n3267));
  NOR2xp33_ASAP7_75t_L      g03011(.A(new_n3264), .B(new_n3258), .Y(new_n3268));
  AOI21xp33_ASAP7_75t_L     g03012(.A1(new_n3267), .A2(new_n3243), .B(new_n3268), .Y(new_n3269));
  OAI22xp33_ASAP7_75t_L     g03013(.A1(new_n3084), .A2(new_n3237), .B1(new_n3269), .B2(new_n3266), .Y(new_n3270));
  NAND2xp33_ASAP7_75t_L     g03014(.A(new_n3074), .B(new_n3071), .Y(new_n3271));
  MAJIxp5_ASAP7_75t_L       g03015(.A(new_n3271), .B(new_n3066), .C(new_n3235), .Y(new_n3272));
  NAND3xp33_ASAP7_75t_L     g03016(.A(new_n3267), .B(new_n3268), .C(new_n3243), .Y(new_n3273));
  OAI21xp33_ASAP7_75t_L     g03017(.A1(new_n3242), .A2(new_n3244), .B(new_n3265), .Y(new_n3274));
  NAND3xp33_ASAP7_75t_L     g03018(.A(new_n3272), .B(new_n3273), .C(new_n3274), .Y(new_n3275));
  OAI211xp5_ASAP7_75t_L     g03019(.A1(new_n3233), .A2(new_n3234), .B(new_n3275), .C(new_n3270), .Y(new_n3276));
  NOR2xp33_ASAP7_75t_L      g03020(.A(new_n3234), .B(new_n3233), .Y(new_n3277));
  AOI21xp33_ASAP7_75t_L     g03021(.A1(new_n3274), .A2(new_n3273), .B(new_n3272), .Y(new_n3278));
  NOR4xp25_ASAP7_75t_L      g03022(.A(new_n3084), .B(new_n3237), .C(new_n3266), .D(new_n3269), .Y(new_n3279));
  OAI21xp33_ASAP7_75t_L     g03023(.A1(new_n3279), .A2(new_n3278), .B(new_n3277), .Y(new_n3280));
  NAND3xp33_ASAP7_75t_L     g03024(.A(new_n3229), .B(new_n3276), .C(new_n3280), .Y(new_n3281));
  NOR4xp25_ASAP7_75t_L      g03025(.A(new_n3086), .B(new_n3087), .C(new_n3085), .D(new_n3084), .Y(new_n3282));
  AOI22xp33_ASAP7_75t_L     g03026(.A1(new_n3075), .A2(new_n3076), .B1(new_n3080), .B2(new_n3082), .Y(new_n3283));
  OAI22xp33_ASAP7_75t_L     g03027(.A1(new_n3089), .A2(new_n2946), .B1(new_n3282), .B2(new_n3283), .Y(new_n3284));
  NOR3xp33_ASAP7_75t_L      g03028(.A(new_n3278), .B(new_n3279), .C(new_n3277), .Y(new_n3285));
  AOI211xp5_ASAP7_75t_L     g03029(.A1(new_n3275), .A2(new_n3270), .B(new_n3233), .C(new_n3234), .Y(new_n3286));
  OAI211xp5_ASAP7_75t_L     g03030(.A1(new_n3286), .A2(new_n3285), .B(new_n3284), .C(new_n3228), .Y(new_n3287));
  NOR2xp33_ASAP7_75t_L      g03031(.A(new_n503), .B(new_n1911), .Y(new_n3288));
  NAND2xp33_ASAP7_75t_L     g03032(.A(\b[9] ), .B(new_n1770), .Y(new_n3289));
  NAND2xp33_ASAP7_75t_L     g03033(.A(\b[10] ), .B(new_n1766), .Y(new_n3290));
  OAI311xp33_ASAP7_75t_L    g03034(.A1(new_n639), .A2(new_n851), .A3(new_n1771), .B1(new_n3290), .C1(new_n3289), .Y(new_n3291));
  OR3x1_ASAP7_75t_L         g03035(.A(new_n3291), .B(new_n1761), .C(new_n3288), .Y(new_n3292));
  A2O1A1Ixp33_ASAP7_75t_L   g03036(.A1(\b[8] ), .A2(new_n1910), .B(new_n3291), .C(new_n1761), .Y(new_n3293));
  AND2x2_ASAP7_75t_L        g03037(.A(new_n3293), .B(new_n3292), .Y(new_n3294));
  NAND3xp33_ASAP7_75t_L     g03038(.A(new_n3281), .B(new_n3294), .C(new_n3287), .Y(new_n3295));
  AOI211xp5_ASAP7_75t_L     g03039(.A1(new_n3284), .A2(new_n3228), .B(new_n3285), .C(new_n3286), .Y(new_n3296));
  AOI21xp33_ASAP7_75t_L     g03040(.A1(new_n3280), .A2(new_n3276), .B(new_n3229), .Y(new_n3297));
  NAND2xp33_ASAP7_75t_L     g03041(.A(new_n3293), .B(new_n3292), .Y(new_n3298));
  OAI21xp33_ASAP7_75t_L     g03042(.A1(new_n3297), .A2(new_n3296), .B(new_n3298), .Y(new_n3299));
  NAND4xp25_ASAP7_75t_L     g03043(.A(new_n3095), .B(new_n3099), .C(new_n3100), .D(new_n3090), .Y(new_n3300));
  A2O1A1O1Ixp25_ASAP7_75t_L g03044(.A1(new_n2948), .A2(new_n2915), .B(new_n2949), .C(new_n3300), .D(new_n3101), .Y(new_n3301));
  NAND3xp33_ASAP7_75t_L     g03045(.A(new_n3301), .B(new_n3299), .C(new_n3295), .Y(new_n3302));
  NOR3xp33_ASAP7_75t_L      g03046(.A(new_n3296), .B(new_n3297), .C(new_n3298), .Y(new_n3303));
  AOI21xp33_ASAP7_75t_L     g03047(.A1(new_n3281), .A2(new_n3287), .B(new_n3294), .Y(new_n3304));
  AO22x1_ASAP7_75t_L        g03048(.A1(new_n3100), .A2(new_n3099), .B1(new_n3090), .B2(new_n3095), .Y(new_n3305));
  OAI21xp33_ASAP7_75t_L     g03049(.A1(new_n3102), .A2(new_n3059), .B(new_n3305), .Y(new_n3306));
  OAI21xp33_ASAP7_75t_L     g03050(.A1(new_n3303), .A2(new_n3304), .B(new_n3306), .Y(new_n3307));
  NAND2xp33_ASAP7_75t_L     g03051(.A(\b[12] ), .B(new_n1410), .Y(new_n3308));
  NAND2xp33_ASAP7_75t_L     g03052(.A(\b[13] ), .B(new_n1406), .Y(new_n3309));
  OAI311xp33_ASAP7_75t_L    g03053(.A1(new_n799), .A2(new_n797), .A3(new_n1411), .B1(new_n3309), .C1(new_n3308), .Y(new_n3310));
  AOI21xp33_ASAP7_75t_L     g03054(.A1(new_n1548), .A2(\b[11] ), .B(new_n3310), .Y(new_n3311));
  NAND2xp33_ASAP7_75t_L     g03055(.A(\a[20] ), .B(new_n3311), .Y(new_n3312));
  A2O1A1Ixp33_ASAP7_75t_L   g03056(.A1(\b[11] ), .A2(new_n1548), .B(new_n3310), .C(new_n1401), .Y(new_n3313));
  NAND2xp33_ASAP7_75t_L     g03057(.A(new_n3313), .B(new_n3312), .Y(new_n3314));
  AOI21xp33_ASAP7_75t_L     g03058(.A1(new_n3302), .A2(new_n3307), .B(new_n3314), .Y(new_n3315));
  AND3x1_ASAP7_75t_L        g03059(.A(new_n3302), .B(new_n3314), .C(new_n3307), .Y(new_n3316));
  A2O1A1O1Ixp25_ASAP7_75t_L g03060(.A1(new_n2963), .A2(new_n2962), .B(new_n2959), .C(new_n3105), .D(new_n3115), .Y(new_n3317));
  NOR3xp33_ASAP7_75t_L      g03061(.A(new_n3317), .B(new_n3316), .C(new_n3315), .Y(new_n3318));
  AO21x2_ASAP7_75t_L        g03062(.A1(new_n3307), .A2(new_n3302), .B(new_n3314), .Y(new_n3319));
  NAND3xp33_ASAP7_75t_L     g03063(.A(new_n3302), .B(new_n3314), .C(new_n3307), .Y(new_n3320));
  AOI221xp5_ASAP7_75t_L     g03064(.A1(new_n3051), .A2(new_n3105), .B1(new_n3319), .B2(new_n3320), .C(new_n3115), .Y(new_n3321));
  NAND2xp33_ASAP7_75t_L     g03065(.A(\b[15] ), .B(new_n1103), .Y(new_n3322));
  NAND2xp33_ASAP7_75t_L     g03066(.A(\b[16] ), .B(new_n1113), .Y(new_n3323));
  OAI311xp33_ASAP7_75t_L    g03067(.A1(new_n1057), .A2(new_n1055), .A3(new_n1197), .B1(new_n3323), .C1(new_n3322), .Y(new_n3324));
  AOI21xp33_ASAP7_75t_L     g03068(.A1(new_n1194), .A2(\b[14] ), .B(new_n3324), .Y(new_n3325));
  NAND2xp33_ASAP7_75t_L     g03069(.A(\a[17] ), .B(new_n3325), .Y(new_n3326));
  A2O1A1Ixp33_ASAP7_75t_L   g03070(.A1(\b[14] ), .A2(new_n1194), .B(new_n3324), .C(new_n1107), .Y(new_n3327));
  NAND2xp33_ASAP7_75t_L     g03071(.A(new_n3327), .B(new_n3326), .Y(new_n3328));
  NOR3xp33_ASAP7_75t_L      g03072(.A(new_n3318), .B(new_n3321), .C(new_n3328), .Y(new_n3329));
  OA21x2_ASAP7_75t_L        g03073(.A1(new_n3321), .A2(new_n3318), .B(new_n3328), .Y(new_n3330));
  NOR2xp33_ASAP7_75t_L      g03074(.A(new_n3329), .B(new_n3330), .Y(new_n3331));
  OAI211xp5_ASAP7_75t_L     g03075(.A1(new_n3120), .A2(new_n3123), .B(new_n3111), .C(new_n3116), .Y(new_n3332));
  NAND3xp33_ASAP7_75t_L     g03076(.A(new_n3331), .B(new_n3145), .C(new_n3332), .Y(new_n3333));
  OAI21xp33_ASAP7_75t_L     g03077(.A1(new_n3114), .A2(new_n3113), .B(new_n3110), .Y(new_n3334));
  NAND3xp33_ASAP7_75t_L     g03078(.A(new_n3334), .B(new_n3320), .C(new_n3319), .Y(new_n3335));
  OAI21xp33_ASAP7_75t_L     g03079(.A1(new_n3315), .A2(new_n3316), .B(new_n3317), .Y(new_n3336));
  NAND4xp25_ASAP7_75t_L     g03080(.A(new_n3335), .B(new_n3327), .C(new_n3326), .D(new_n3336), .Y(new_n3337));
  OAI21xp33_ASAP7_75t_L     g03081(.A1(new_n3321), .A2(new_n3318), .B(new_n3328), .Y(new_n3338));
  NAND2xp33_ASAP7_75t_L     g03082(.A(new_n3338), .B(new_n3337), .Y(new_n3339));
  A2O1A1Ixp33_ASAP7_75t_L   g03083(.A1(new_n3126), .A2(new_n3125), .B(new_n3130), .C(new_n3332), .Y(new_n3340));
  NAND2xp33_ASAP7_75t_L     g03084(.A(new_n3340), .B(new_n3339), .Y(new_n3341));
  NAND2xp33_ASAP7_75t_L     g03085(.A(\b[18] ), .B(new_n817), .Y(new_n3342));
  OAI221xp5_ASAP7_75t_L     g03086(.A1(new_n912), .A2(new_n1493), .B1(new_n911), .B2(new_n2793), .C(new_n3342), .Y(new_n3343));
  AOI211xp5_ASAP7_75t_L     g03087(.A1(\b[17] ), .A2(new_n908), .B(new_n813), .C(new_n3343), .Y(new_n3344));
  NOR2xp33_ASAP7_75t_L      g03088(.A(new_n1493), .B(new_n912), .Y(new_n3345));
  AOI221xp5_ASAP7_75t_L     g03089(.A1(new_n817), .A2(\b[18] ), .B1(new_n823), .B2(new_n1499), .C(new_n3345), .Y(new_n3346));
  O2A1O1Ixp33_ASAP7_75t_L   g03090(.A1(new_n1244), .A2(new_n909), .B(new_n3346), .C(\a[14] ), .Y(new_n3347));
  NOR2xp33_ASAP7_75t_L      g03091(.A(new_n3347), .B(new_n3344), .Y(new_n3348));
  NAND3xp33_ASAP7_75t_L     g03092(.A(new_n3333), .B(new_n3341), .C(new_n3348), .Y(new_n3349));
  NOR2xp33_ASAP7_75t_L      g03093(.A(new_n3340), .B(new_n3339), .Y(new_n3350));
  AOI21xp33_ASAP7_75t_L     g03094(.A1(new_n3145), .A2(new_n3332), .B(new_n3331), .Y(new_n3351));
  OR2x4_ASAP7_75t_L         g03095(.A(new_n3347), .B(new_n3344), .Y(new_n3352));
  OAI21xp33_ASAP7_75t_L     g03096(.A1(new_n3350), .A2(new_n3351), .B(new_n3352), .Y(new_n3353));
  NOR3xp33_ASAP7_75t_L      g03097(.A(new_n3146), .B(new_n3129), .C(new_n3131), .Y(new_n3354));
  O2A1O1Ixp33_ASAP7_75t_L   g03098(.A1(new_n3143), .A2(new_n3147), .B(new_n3165), .C(new_n3354), .Y(new_n3355));
  NAND3xp33_ASAP7_75t_L     g03099(.A(new_n3355), .B(new_n3353), .C(new_n3349), .Y(new_n3356));
  NAND2xp33_ASAP7_75t_L     g03100(.A(new_n3349), .B(new_n3353), .Y(new_n3357));
  A2O1A1Ixp33_ASAP7_75t_L   g03101(.A1(new_n3155), .A2(new_n3165), .B(new_n3354), .C(new_n3357), .Y(new_n3358));
  NAND2xp33_ASAP7_75t_L     g03102(.A(\b[21] ), .B(new_n590), .Y(new_n3359));
  OAI221xp5_ASAP7_75t_L     g03103(.A1(new_n676), .A2(new_n1857), .B1(new_n675), .B2(new_n1863), .C(new_n3359), .Y(new_n3360));
  AOI21xp33_ASAP7_75t_L     g03104(.A1(new_n674), .A2(\b[20] ), .B(new_n3360), .Y(new_n3361));
  NAND2xp33_ASAP7_75t_L     g03105(.A(\a[11] ), .B(new_n3361), .Y(new_n3362));
  A2O1A1Ixp33_ASAP7_75t_L   g03106(.A1(\b[20] ), .A2(new_n674), .B(new_n3360), .C(new_n594), .Y(new_n3363));
  NAND4xp25_ASAP7_75t_L     g03107(.A(new_n3358), .B(new_n3356), .C(new_n3362), .D(new_n3363), .Y(new_n3364));
  INVx1_ASAP7_75t_L         g03108(.A(new_n3354), .Y(new_n3365));
  OAI21xp33_ASAP7_75t_L     g03109(.A1(new_n3148), .A2(new_n3151), .B(new_n3365), .Y(new_n3366));
  NOR2xp33_ASAP7_75t_L      g03110(.A(new_n3357), .B(new_n3366), .Y(new_n3367));
  AOI21xp33_ASAP7_75t_L     g03111(.A1(new_n3353), .A2(new_n3349), .B(new_n3355), .Y(new_n3368));
  NAND2xp33_ASAP7_75t_L     g03112(.A(new_n3363), .B(new_n3362), .Y(new_n3369));
  OAI21xp33_ASAP7_75t_L     g03113(.A1(new_n3368), .A2(new_n3367), .B(new_n3369), .Y(new_n3370));
  NAND3xp33_ASAP7_75t_L     g03114(.A(new_n3156), .B(new_n3152), .C(new_n3168), .Y(new_n3371));
  OAI22xp33_ASAP7_75t_L     g03115(.A1(new_n3170), .A2(new_n3018), .B1(new_n3172), .B2(new_n3173), .Y(new_n3372));
  NAND4xp25_ASAP7_75t_L     g03116(.A(new_n3372), .B(new_n3364), .C(new_n3370), .D(new_n3371), .Y(new_n3373));
  NOR3xp33_ASAP7_75t_L      g03117(.A(new_n3367), .B(new_n3368), .C(new_n3369), .Y(new_n3374));
  AOI22xp33_ASAP7_75t_L     g03118(.A1(new_n3362), .A2(new_n3363), .B1(new_n3356), .B2(new_n3358), .Y(new_n3375));
  A2O1A1Ixp33_ASAP7_75t_L   g03119(.A1(new_n3169), .A2(new_n3164), .B(new_n3174), .C(new_n3371), .Y(new_n3376));
  OAI21xp33_ASAP7_75t_L     g03120(.A1(new_n3374), .A2(new_n3375), .B(new_n3376), .Y(new_n3377));
  NAND2xp33_ASAP7_75t_L     g03121(.A(new_n3377), .B(new_n3373), .Y(new_n3378));
  NOR2xp33_ASAP7_75t_L      g03122(.A(new_n2180), .B(new_n667), .Y(new_n3379));
  AOI221xp5_ASAP7_75t_L     g03123(.A1(new_n441), .A2(\b[24] ), .B1(new_n448), .B2(new_n2188), .C(new_n3379), .Y(new_n3380));
  OAI211xp5_ASAP7_75t_L     g03124(.A1(new_n1995), .A2(new_n481), .B(new_n3380), .C(\a[8] ), .Y(new_n3381));
  O2A1O1Ixp33_ASAP7_75t_L   g03125(.A1(new_n1995), .A2(new_n481), .B(new_n3380), .C(\a[8] ), .Y(new_n3382));
  INVx1_ASAP7_75t_L         g03126(.A(new_n3382), .Y(new_n3383));
  NAND2xp33_ASAP7_75t_L     g03127(.A(new_n3381), .B(new_n3383), .Y(new_n3384));
  NOR2xp33_ASAP7_75t_L      g03128(.A(new_n3384), .B(new_n3378), .Y(new_n3385));
  INVx1_ASAP7_75t_L         g03129(.A(new_n3381), .Y(new_n3386));
  NOR2xp33_ASAP7_75t_L      g03130(.A(new_n3382), .B(new_n3386), .Y(new_n3387));
  AOI21xp33_ASAP7_75t_L     g03131(.A1(new_n3377), .A2(new_n3373), .B(new_n3387), .Y(new_n3388));
  OAI21xp33_ASAP7_75t_L     g03132(.A1(new_n3184), .A2(new_n3049), .B(new_n3190), .Y(new_n3389));
  NOR3xp33_ASAP7_75t_L      g03133(.A(new_n3389), .B(new_n3385), .C(new_n3388), .Y(new_n3390));
  NAND3xp33_ASAP7_75t_L     g03134(.A(new_n3387), .B(new_n3377), .C(new_n3373), .Y(new_n3391));
  NAND2xp33_ASAP7_75t_L     g03135(.A(new_n3384), .B(new_n3378), .Y(new_n3392));
  A2O1A1O1Ixp25_ASAP7_75t_L g03136(.A1(new_n3026), .A2(new_n2894), .B(new_n3029), .C(new_n3183), .D(new_n3182), .Y(new_n3393));
  AOI21xp33_ASAP7_75t_L     g03137(.A1(new_n3392), .A2(new_n3391), .B(new_n3393), .Y(new_n3394));
  NAND2xp33_ASAP7_75t_L     g03138(.A(\b[26] ), .B(new_n366), .Y(new_n3395));
  NOR2xp33_ASAP7_75t_L      g03139(.A(new_n2852), .B(new_n368), .Y(new_n3396));
  AOI221xp5_ASAP7_75t_L     g03140(.A1(new_n334), .A2(\b[27] ), .B1(new_n342), .B2(new_n2858), .C(new_n3396), .Y(new_n3397));
  AND3x1_ASAP7_75t_L        g03141(.A(new_n3397), .B(new_n3395), .C(\a[5] ), .Y(new_n3398));
  O2A1O1Ixp33_ASAP7_75t_L   g03142(.A1(new_n2477), .A2(new_n365), .B(new_n3397), .C(\a[5] ), .Y(new_n3399));
  NOR2xp33_ASAP7_75t_L      g03143(.A(new_n3399), .B(new_n3398), .Y(new_n3400));
  INVx1_ASAP7_75t_L         g03144(.A(new_n3400), .Y(new_n3401));
  NOR3xp33_ASAP7_75t_L      g03145(.A(new_n3401), .B(new_n3390), .C(new_n3394), .Y(new_n3402));
  NAND3xp33_ASAP7_75t_L     g03146(.A(new_n3392), .B(new_n3391), .C(new_n3393), .Y(new_n3403));
  OAI21xp33_ASAP7_75t_L     g03147(.A1(new_n3388), .A2(new_n3385), .B(new_n3389), .Y(new_n3404));
  AOI21xp33_ASAP7_75t_L     g03148(.A1(new_n3404), .A2(new_n3403), .B(new_n3400), .Y(new_n3405));
  NOR2xp33_ASAP7_75t_L      g03149(.A(new_n3405), .B(new_n3402), .Y(new_n3406));
  NAND2xp33_ASAP7_75t_L     g03150(.A(new_n3185), .B(new_n3191), .Y(new_n3407));
  NOR2xp33_ASAP7_75t_L      g03151(.A(new_n3197), .B(new_n3407), .Y(new_n3408));
  A2O1A1O1Ixp25_ASAP7_75t_L g03152(.A1(new_n3039), .A2(new_n3037), .B(new_n3207), .C(new_n3206), .D(new_n3408), .Y(new_n3409));
  NAND2xp33_ASAP7_75t_L     g03153(.A(new_n3406), .B(new_n3409), .Y(new_n3410));
  A2O1A1Ixp33_ASAP7_75t_L   g03154(.A1(new_n2849), .A2(new_n3046), .B(new_n3035), .C(new_n3204), .Y(new_n3411));
  NAND3xp33_ASAP7_75t_L     g03155(.A(new_n3404), .B(new_n3403), .C(new_n3400), .Y(new_n3412));
  OAI21xp33_ASAP7_75t_L     g03156(.A1(new_n3394), .A2(new_n3390), .B(new_n3401), .Y(new_n3413));
  NAND2xp33_ASAP7_75t_L     g03157(.A(new_n3412), .B(new_n3413), .Y(new_n3414));
  A2O1A1Ixp33_ASAP7_75t_L   g03158(.A1(new_n3411), .A2(new_n3206), .B(new_n3408), .C(new_n3414), .Y(new_n3415));
  NAND2xp33_ASAP7_75t_L     g03159(.A(\b[29] ), .B(new_n291), .Y(new_n3416));
  NAND2xp33_ASAP7_75t_L     g03160(.A(\b[30] ), .B(new_n380), .Y(new_n3417));
  NOR2xp33_ASAP7_75t_L      g03161(.A(\b[30] ), .B(\b[31] ), .Y(new_n3418));
  INVx1_ASAP7_75t_L         g03162(.A(\b[31] ), .Y(new_n3419));
  NOR2xp33_ASAP7_75t_L      g03163(.A(new_n3212), .B(new_n3419), .Y(new_n3420));
  NOR2xp33_ASAP7_75t_L      g03164(.A(new_n3418), .B(new_n3420), .Y(new_n3421));
  A2O1A1Ixp33_ASAP7_75t_L   g03165(.A1(\b[30] ), .A2(\b[29] ), .B(new_n3216), .C(new_n3421), .Y(new_n3422));
  O2A1O1Ixp33_ASAP7_75t_L   g03166(.A1(new_n2875), .A2(new_n3217), .B(new_n3214), .C(new_n3213), .Y(new_n3423));
  INVx1_ASAP7_75t_L         g03167(.A(new_n3421), .Y(new_n3424));
  NAND2xp33_ASAP7_75t_L     g03168(.A(new_n3424), .B(new_n3423), .Y(new_n3425));
  AND2x2_ASAP7_75t_L        g03169(.A(new_n3422), .B(new_n3425), .Y(new_n3426));
  AOI22xp33_ASAP7_75t_L     g03170(.A1(new_n272), .A2(\b[31] ), .B1(new_n269), .B2(new_n3426), .Y(new_n3427));
  NAND4xp25_ASAP7_75t_L     g03171(.A(new_n3427), .B(\a[2] ), .C(new_n3416), .D(new_n3417), .Y(new_n3428));
  NAND2xp33_ASAP7_75t_L     g03172(.A(new_n3417), .B(new_n3427), .Y(new_n3429));
  A2O1A1Ixp33_ASAP7_75t_L   g03173(.A1(\b[29] ), .A2(new_n291), .B(new_n3429), .C(new_n265), .Y(new_n3430));
  AND2x2_ASAP7_75t_L        g03174(.A(new_n3428), .B(new_n3430), .Y(new_n3431));
  NAND3xp33_ASAP7_75t_L     g03175(.A(new_n3410), .B(new_n3415), .C(new_n3431), .Y(new_n3432));
  AO21x2_ASAP7_75t_L        g03176(.A1(new_n3415), .A2(new_n3410), .B(new_n3431), .Y(new_n3433));
  NAND2xp33_ASAP7_75t_L     g03177(.A(new_n3432), .B(new_n3433), .Y(new_n3434));
  MAJIxp5_ASAP7_75t_L       g03178(.A(new_n3225), .B(new_n3209), .C(new_n3222), .Y(new_n3435));
  XOR2x2_ASAP7_75t_L        g03179(.A(new_n3434), .B(new_n3435), .Y(\f[31] ));
  NAND2xp33_ASAP7_75t_L     g03180(.A(new_n3415), .B(new_n3410), .Y(new_n3437));
  NAND2xp33_ASAP7_75t_L     g03181(.A(new_n3434), .B(new_n3435), .Y(new_n3438));
  A2O1A1Ixp33_ASAP7_75t_L   g03182(.A1(new_n3428), .A2(new_n3430), .B(new_n3437), .C(new_n3438), .Y(new_n3439));
  NAND2xp33_ASAP7_75t_L     g03183(.A(\b[30] ), .B(new_n291), .Y(new_n3440));
  NAND2xp33_ASAP7_75t_L     g03184(.A(\b[31] ), .B(new_n380), .Y(new_n3441));
  NOR2xp33_ASAP7_75t_L      g03185(.A(\b[31] ), .B(\b[32] ), .Y(new_n3442));
  INVx1_ASAP7_75t_L         g03186(.A(\b[32] ), .Y(new_n3443));
  NOR2xp33_ASAP7_75t_L      g03187(.A(new_n3419), .B(new_n3443), .Y(new_n3444));
  NOR2xp33_ASAP7_75t_L      g03188(.A(new_n3442), .B(new_n3444), .Y(new_n3445));
  INVx1_ASAP7_75t_L         g03189(.A(new_n3445), .Y(new_n3446));
  O2A1O1Ixp33_ASAP7_75t_L   g03190(.A1(new_n3212), .A2(new_n3419), .B(new_n3422), .C(new_n3446), .Y(new_n3447));
  OAI21xp33_ASAP7_75t_L     g03191(.A1(new_n3212), .A2(new_n3419), .B(new_n3422), .Y(new_n3448));
  NOR2xp33_ASAP7_75t_L      g03192(.A(new_n3445), .B(new_n3448), .Y(new_n3449));
  NOR2xp33_ASAP7_75t_L      g03193(.A(new_n3447), .B(new_n3449), .Y(new_n3450));
  AOI22xp33_ASAP7_75t_L     g03194(.A1(new_n272), .A2(\b[32] ), .B1(new_n269), .B2(new_n3450), .Y(new_n3451));
  NAND4xp25_ASAP7_75t_L     g03195(.A(new_n3451), .B(\a[2] ), .C(new_n3440), .D(new_n3441), .Y(new_n3452));
  NAND2xp33_ASAP7_75t_L     g03196(.A(new_n3441), .B(new_n3451), .Y(new_n3453));
  A2O1A1Ixp33_ASAP7_75t_L   g03197(.A1(\b[30] ), .A2(new_n291), .B(new_n3453), .C(new_n265), .Y(new_n3454));
  AND2x2_ASAP7_75t_L        g03198(.A(new_n3452), .B(new_n3454), .Y(new_n3455));
  NOR3xp33_ASAP7_75t_L      g03199(.A(new_n3390), .B(new_n3394), .C(new_n3400), .Y(new_n3456));
  A2O1A1O1Ixp25_ASAP7_75t_L g03200(.A1(new_n3206), .A2(new_n3411), .B(new_n3408), .C(new_n3414), .D(new_n3456), .Y(new_n3457));
  XNOR2x2_ASAP7_75t_L       g03201(.A(new_n3355), .B(new_n3357), .Y(new_n3458));
  MAJIxp5_ASAP7_75t_L       g03202(.A(new_n3376), .B(new_n3458), .C(new_n3369), .Y(new_n3459));
  AOI32xp33_ASAP7_75t_L     g03203(.A1(new_n1998), .A2(new_n2001), .A3(new_n597), .B1(new_n600), .B2(\b[23] ), .Y(new_n3460));
  OAI221xp5_ASAP7_75t_L     g03204(.A1(new_n721), .A2(new_n1857), .B1(new_n1709), .B2(new_n1620), .C(new_n3460), .Y(new_n3461));
  XNOR2x2_ASAP7_75t_L       g03205(.A(\a[11] ), .B(new_n3461), .Y(new_n3462));
  NAND3xp33_ASAP7_75t_L     g03206(.A(new_n3352), .B(new_n3341), .C(new_n3333), .Y(new_n3463));
  INVx1_ASAP7_75t_L         g03207(.A(new_n3463), .Y(new_n3464));
  A2O1A1O1Ixp25_ASAP7_75t_L g03208(.A1(new_n3165), .A2(new_n3155), .B(new_n3354), .C(new_n3357), .D(new_n3464), .Y(new_n3465));
  OAI21xp33_ASAP7_75t_L     g03209(.A1(new_n3315), .A2(new_n3317), .B(new_n3320), .Y(new_n3466));
  NAND2xp33_ASAP7_75t_L     g03210(.A(\b[12] ), .B(new_n1548), .Y(new_n3467));
  NAND2xp33_ASAP7_75t_L     g03211(.A(\b[13] ), .B(new_n1410), .Y(new_n3468));
  AOI32xp33_ASAP7_75t_L     g03212(.A1(new_n877), .A2(new_n874), .A3(new_n1404), .B1(\b[14] ), .B2(new_n1406), .Y(new_n3469));
  NAND4xp25_ASAP7_75t_L     g03213(.A(new_n3469), .B(\a[20] ), .C(new_n3467), .D(new_n3468), .Y(new_n3470));
  NAND2xp33_ASAP7_75t_L     g03214(.A(new_n3468), .B(new_n3469), .Y(new_n3471));
  A2O1A1Ixp33_ASAP7_75t_L   g03215(.A1(\b[12] ), .A2(new_n1548), .B(new_n3471), .C(new_n1401), .Y(new_n3472));
  AND2x2_ASAP7_75t_L        g03216(.A(new_n3470), .B(new_n3472), .Y(new_n3473));
  NAND3xp33_ASAP7_75t_L     g03217(.A(new_n3281), .B(new_n3287), .C(new_n3298), .Y(new_n3474));
  INVx1_ASAP7_75t_L         g03218(.A(new_n3474), .Y(new_n3475));
  O2A1O1Ixp33_ASAP7_75t_L   g03219(.A1(new_n3303), .A2(new_n3304), .B(new_n3306), .C(new_n3475), .Y(new_n3476));
  AOI21xp33_ASAP7_75t_L     g03220(.A1(new_n3229), .A2(new_n3280), .B(new_n3285), .Y(new_n3477));
  NOR2xp33_ASAP7_75t_L      g03221(.A(new_n382), .B(new_n2387), .Y(new_n3478));
  NAND2xp33_ASAP7_75t_L     g03222(.A(\b[7] ), .B(new_n2232), .Y(new_n3479));
  OAI221xp5_ASAP7_75t_L     g03223(.A1(new_n2234), .A2(new_n503), .B1(new_n2233), .B2(new_n509), .C(new_n3479), .Y(new_n3480));
  OR3x1_ASAP7_75t_L         g03224(.A(new_n3480), .B(new_n2223), .C(new_n3478), .Y(new_n3481));
  A2O1A1Ixp33_ASAP7_75t_L   g03225(.A1(\b[6] ), .A2(new_n2386), .B(new_n3480), .C(new_n2223), .Y(new_n3482));
  OAI21xp33_ASAP7_75t_L     g03226(.A1(new_n3242), .A2(new_n3244), .B(new_n3268), .Y(new_n3483));
  NAND2xp33_ASAP7_75t_L     g03227(.A(\b[3] ), .B(new_n2931), .Y(new_n3484));
  NAND2xp33_ASAP7_75t_L     g03228(.A(\b[4] ), .B(new_n2706), .Y(new_n3485));
  AOI32xp33_ASAP7_75t_L     g03229(.A1(new_n358), .A2(new_n356), .A3(new_n2700), .B1(\b[5] ), .B2(new_n2702), .Y(new_n3486));
  NAND3xp33_ASAP7_75t_L     g03230(.A(new_n3486), .B(new_n3485), .C(new_n3484), .Y(new_n3487));
  NOR2xp33_ASAP7_75t_L      g03231(.A(new_n2697), .B(new_n3487), .Y(new_n3488));
  AOI31xp33_ASAP7_75t_L     g03232(.A1(new_n3486), .A2(new_n3485), .A3(new_n3484), .B(\a[29] ), .Y(new_n3489));
  A2O1A1O1Ixp25_ASAP7_75t_L g03233(.A1(new_n3246), .A2(new_n3065), .B(new_n258), .C(new_n3257), .D(new_n3251), .Y(new_n3490));
  NOR3xp33_ASAP7_75t_L      g03234(.A(new_n3253), .B(new_n3247), .C(new_n3259), .Y(new_n3491));
  INVx1_ASAP7_75t_L         g03235(.A(new_n3491), .Y(new_n3492));
  NOR2xp33_ASAP7_75t_L      g03236(.A(new_n258), .B(new_n3492), .Y(new_n3493));
  NAND2xp33_ASAP7_75t_L     g03237(.A(\b[1] ), .B(new_n3260), .Y(new_n3494));
  OAI221xp5_ASAP7_75t_L     g03238(.A1(new_n3261), .A2(new_n283), .B1(new_n278), .B2(new_n3262), .C(new_n3494), .Y(new_n3495));
  OR3x1_ASAP7_75t_L         g03239(.A(new_n3490), .B(new_n3493), .C(new_n3495), .Y(new_n3496));
  A2O1A1Ixp33_ASAP7_75t_L   g03240(.A1(\b[0] ), .A2(new_n3491), .B(new_n3495), .C(new_n3490), .Y(new_n3497));
  AOI211xp5_ASAP7_75t_L     g03241(.A1(new_n3496), .A2(new_n3497), .B(new_n3489), .C(new_n3488), .Y(new_n3498));
  INVx1_ASAP7_75t_L         g03242(.A(new_n3498), .Y(new_n3499));
  OAI211xp5_ASAP7_75t_L     g03243(.A1(new_n3489), .A2(new_n3488), .B(new_n3496), .C(new_n3497), .Y(new_n3500));
  NAND4xp25_ASAP7_75t_L     g03244(.A(new_n3270), .B(new_n3499), .C(new_n3500), .D(new_n3483), .Y(new_n3501));
  A2O1A1Ixp33_ASAP7_75t_L   g03245(.A1(new_n3273), .A2(new_n3274), .B(new_n3272), .C(new_n3483), .Y(new_n3502));
  INVx1_ASAP7_75t_L         g03246(.A(new_n3500), .Y(new_n3503));
  OAI21xp33_ASAP7_75t_L     g03247(.A1(new_n3498), .A2(new_n3503), .B(new_n3502), .Y(new_n3504));
  AOI22xp33_ASAP7_75t_L     g03248(.A1(new_n3481), .A2(new_n3482), .B1(new_n3501), .B2(new_n3504), .Y(new_n3505));
  NAND4xp25_ASAP7_75t_L     g03249(.A(new_n3504), .B(new_n3481), .C(new_n3501), .D(new_n3482), .Y(new_n3506));
  INVx1_ASAP7_75t_L         g03250(.A(new_n3506), .Y(new_n3507));
  OAI21xp33_ASAP7_75t_L     g03251(.A1(new_n3505), .A2(new_n3507), .B(new_n3477), .Y(new_n3508));
  A2O1A1Ixp33_ASAP7_75t_L   g03252(.A1(new_n3284), .A2(new_n3228), .B(new_n3286), .C(new_n3276), .Y(new_n3509));
  INVx1_ASAP7_75t_L         g03253(.A(new_n3505), .Y(new_n3510));
  NAND3xp33_ASAP7_75t_L     g03254(.A(new_n3509), .B(new_n3510), .C(new_n3506), .Y(new_n3511));
  NAND2xp33_ASAP7_75t_L     g03255(.A(\b[9] ), .B(new_n1910), .Y(new_n3512));
  NAND2xp33_ASAP7_75t_L     g03256(.A(\b[10] ), .B(new_n1770), .Y(new_n3513));
  AOI32xp33_ASAP7_75t_L     g03257(.A1(new_n700), .A2(new_n698), .A3(new_n1764), .B1(\b[11] ), .B2(new_n1766), .Y(new_n3514));
  NAND4xp25_ASAP7_75t_L     g03258(.A(new_n3514), .B(\a[23] ), .C(new_n3512), .D(new_n3513), .Y(new_n3515));
  AOI31xp33_ASAP7_75t_L     g03259(.A1(new_n3514), .A2(new_n3513), .A3(new_n3512), .B(\a[23] ), .Y(new_n3516));
  INVx1_ASAP7_75t_L         g03260(.A(new_n3516), .Y(new_n3517));
  NAND2xp33_ASAP7_75t_L     g03261(.A(new_n3515), .B(new_n3517), .Y(new_n3518));
  AO21x2_ASAP7_75t_L        g03262(.A1(new_n3508), .A2(new_n3511), .B(new_n3518), .Y(new_n3519));
  NAND3xp33_ASAP7_75t_L     g03263(.A(new_n3518), .B(new_n3511), .C(new_n3508), .Y(new_n3520));
  NAND3xp33_ASAP7_75t_L     g03264(.A(new_n3476), .B(new_n3519), .C(new_n3520), .Y(new_n3521));
  A2O1A1Ixp33_ASAP7_75t_L   g03265(.A1(new_n3299), .A2(new_n3295), .B(new_n3301), .C(new_n3474), .Y(new_n3522));
  AOI21xp33_ASAP7_75t_L     g03266(.A1(new_n3511), .A2(new_n3508), .B(new_n3518), .Y(new_n3523));
  INVx1_ASAP7_75t_L         g03267(.A(new_n3520), .Y(new_n3524));
  OAI21xp33_ASAP7_75t_L     g03268(.A1(new_n3523), .A2(new_n3524), .B(new_n3522), .Y(new_n3525));
  NAND3xp33_ASAP7_75t_L     g03269(.A(new_n3473), .B(new_n3521), .C(new_n3525), .Y(new_n3526));
  NAND2xp33_ASAP7_75t_L     g03270(.A(new_n3470), .B(new_n3472), .Y(new_n3527));
  NOR3xp33_ASAP7_75t_L      g03271(.A(new_n3524), .B(new_n3523), .C(new_n3522), .Y(new_n3528));
  AOI21xp33_ASAP7_75t_L     g03272(.A1(new_n3520), .A2(new_n3519), .B(new_n3476), .Y(new_n3529));
  OAI21xp33_ASAP7_75t_L     g03273(.A1(new_n3529), .A2(new_n3528), .B(new_n3527), .Y(new_n3530));
  NAND3xp33_ASAP7_75t_L     g03274(.A(new_n3466), .B(new_n3526), .C(new_n3530), .Y(new_n3531));
  A2O1A1O1Ixp25_ASAP7_75t_L g03275(.A1(new_n3105), .A2(new_n3051), .B(new_n3115), .C(new_n3319), .D(new_n3316), .Y(new_n3532));
  NOR3xp33_ASAP7_75t_L      g03276(.A(new_n3528), .B(new_n3529), .C(new_n3527), .Y(new_n3533));
  AOI21xp33_ASAP7_75t_L     g03277(.A1(new_n3525), .A2(new_n3521), .B(new_n3473), .Y(new_n3534));
  OAI21xp33_ASAP7_75t_L     g03278(.A1(new_n3533), .A2(new_n3534), .B(new_n3532), .Y(new_n3535));
  NAND2xp33_ASAP7_75t_L     g03279(.A(\b[15] ), .B(new_n1194), .Y(new_n3536));
  NAND2xp33_ASAP7_75t_L     g03280(.A(\b[16] ), .B(new_n1103), .Y(new_n3537));
  AOI32xp33_ASAP7_75t_L     g03281(.A1(new_n1250), .A2(new_n1247), .A3(new_n1110), .B1(new_n1113), .B2(\b[17] ), .Y(new_n3538));
  NAND4xp25_ASAP7_75t_L     g03282(.A(new_n3538), .B(\a[17] ), .C(new_n3536), .D(new_n3537), .Y(new_n3539));
  NAND2xp33_ASAP7_75t_L     g03283(.A(new_n3537), .B(new_n3538), .Y(new_n3540));
  A2O1A1Ixp33_ASAP7_75t_L   g03284(.A1(\b[15] ), .A2(new_n1194), .B(new_n3540), .C(new_n1107), .Y(new_n3541));
  NAND4xp25_ASAP7_75t_L     g03285(.A(new_n3531), .B(new_n3541), .C(new_n3535), .D(new_n3539), .Y(new_n3542));
  NOR3xp33_ASAP7_75t_L      g03286(.A(new_n3532), .B(new_n3533), .C(new_n3534), .Y(new_n3543));
  AOI21xp33_ASAP7_75t_L     g03287(.A1(new_n3530), .A2(new_n3526), .B(new_n3466), .Y(new_n3544));
  NAND2xp33_ASAP7_75t_L     g03288(.A(new_n3539), .B(new_n3541), .Y(new_n3545));
  OAI21xp33_ASAP7_75t_L     g03289(.A1(new_n3544), .A2(new_n3543), .B(new_n3545), .Y(new_n3546));
  AND2x2_ASAP7_75t_L        g03290(.A(new_n3542), .B(new_n3546), .Y(new_n3547));
  NAND3xp33_ASAP7_75t_L     g03291(.A(new_n3335), .B(new_n3336), .C(new_n3328), .Y(new_n3548));
  INVx1_ASAP7_75t_L         g03292(.A(new_n3548), .Y(new_n3549));
  O2A1O1Ixp33_ASAP7_75t_L   g03293(.A1(new_n3329), .A2(new_n3330), .B(new_n3340), .C(new_n3549), .Y(new_n3550));
  NAND2xp33_ASAP7_75t_L     g03294(.A(new_n3550), .B(new_n3547), .Y(new_n3551));
  NAND2xp33_ASAP7_75t_L     g03295(.A(new_n3542), .B(new_n3546), .Y(new_n3552));
  A2O1A1Ixp33_ASAP7_75t_L   g03296(.A1(new_n3339), .A2(new_n3340), .B(new_n3549), .C(new_n3552), .Y(new_n3553));
  NOR2xp33_ASAP7_75t_L      g03297(.A(new_n1356), .B(new_n909), .Y(new_n3554));
  INVx1_ASAP7_75t_L         g03298(.A(new_n3554), .Y(new_n3555));
  NAND2xp33_ASAP7_75t_L     g03299(.A(\b[19] ), .B(new_n817), .Y(new_n3556));
  AOI22xp33_ASAP7_75t_L     g03300(.A1(new_n826), .A2(\b[20] ), .B1(new_n823), .B2(new_n1600), .Y(new_n3557));
  AND4x1_ASAP7_75t_L        g03301(.A(new_n3557), .B(new_n3556), .C(new_n3555), .D(\a[14] ), .Y(new_n3558));
  AOI31xp33_ASAP7_75t_L     g03302(.A1(new_n3557), .A2(new_n3556), .A3(new_n3555), .B(\a[14] ), .Y(new_n3559));
  OR2x4_ASAP7_75t_L         g03303(.A(new_n3559), .B(new_n3558), .Y(new_n3560));
  AOI21xp33_ASAP7_75t_L     g03304(.A1(new_n3553), .A2(new_n3551), .B(new_n3560), .Y(new_n3561));
  A2O1A1Ixp33_ASAP7_75t_L   g03305(.A1(new_n3145), .A2(new_n3332), .B(new_n3331), .C(new_n3548), .Y(new_n3562));
  NOR2xp33_ASAP7_75t_L      g03306(.A(new_n3552), .B(new_n3562), .Y(new_n3563));
  NOR2xp33_ASAP7_75t_L      g03307(.A(new_n3550), .B(new_n3547), .Y(new_n3564));
  NOR2xp33_ASAP7_75t_L      g03308(.A(new_n3559), .B(new_n3558), .Y(new_n3565));
  NOR3xp33_ASAP7_75t_L      g03309(.A(new_n3563), .B(new_n3564), .C(new_n3565), .Y(new_n3566));
  NOR2xp33_ASAP7_75t_L      g03310(.A(new_n3561), .B(new_n3566), .Y(new_n3567));
  NAND2xp33_ASAP7_75t_L     g03311(.A(new_n3567), .B(new_n3465), .Y(new_n3568));
  OAI21xp33_ASAP7_75t_L     g03312(.A1(new_n3564), .A2(new_n3563), .B(new_n3565), .Y(new_n3569));
  NAND3xp33_ASAP7_75t_L     g03313(.A(new_n3560), .B(new_n3553), .C(new_n3551), .Y(new_n3570));
  NAND2xp33_ASAP7_75t_L     g03314(.A(new_n3569), .B(new_n3570), .Y(new_n3571));
  A2O1A1Ixp33_ASAP7_75t_L   g03315(.A1(new_n3366), .A2(new_n3357), .B(new_n3464), .C(new_n3571), .Y(new_n3572));
  NAND3xp33_ASAP7_75t_L     g03316(.A(new_n3572), .B(new_n3568), .C(new_n3462), .Y(new_n3573));
  INVx1_ASAP7_75t_L         g03317(.A(new_n3462), .Y(new_n3574));
  A2O1A1Ixp33_ASAP7_75t_L   g03318(.A1(new_n3353), .A2(new_n3349), .B(new_n3355), .C(new_n3463), .Y(new_n3575));
  NOR2xp33_ASAP7_75t_L      g03319(.A(new_n3571), .B(new_n3575), .Y(new_n3576));
  NOR2xp33_ASAP7_75t_L      g03320(.A(new_n3567), .B(new_n3465), .Y(new_n3577));
  OAI21xp33_ASAP7_75t_L     g03321(.A1(new_n3576), .A2(new_n3577), .B(new_n3574), .Y(new_n3578));
  NAND2xp33_ASAP7_75t_L     g03322(.A(new_n3573), .B(new_n3578), .Y(new_n3579));
  XNOR2x2_ASAP7_75t_L       g03323(.A(new_n3459), .B(new_n3579), .Y(new_n3580));
  OAI22xp33_ASAP7_75t_L     g03324(.A1(new_n2487), .A2(new_n482), .B1(new_n2477), .B2(new_n667), .Y(new_n3581));
  AOI221xp5_ASAP7_75t_L     g03325(.A1(\b[24] ), .A2(new_n480), .B1(\b[25] ), .B2(new_n441), .C(new_n3581), .Y(new_n3582));
  XNOR2x2_ASAP7_75t_L       g03326(.A(new_n445), .B(new_n3582), .Y(new_n3583));
  INVx1_ASAP7_75t_L         g03327(.A(new_n3583), .Y(new_n3584));
  NOR2xp33_ASAP7_75t_L      g03328(.A(new_n3584), .B(new_n3580), .Y(new_n3585));
  NOR3xp33_ASAP7_75t_L      g03329(.A(new_n3577), .B(new_n3576), .C(new_n3574), .Y(new_n3586));
  AOI21xp33_ASAP7_75t_L     g03330(.A1(new_n3572), .A2(new_n3568), .B(new_n3462), .Y(new_n3587));
  NOR3xp33_ASAP7_75t_L      g03331(.A(new_n3459), .B(new_n3586), .C(new_n3587), .Y(new_n3588));
  NAND2xp33_ASAP7_75t_L     g03332(.A(new_n3370), .B(new_n3364), .Y(new_n3589));
  AOI211xp5_ASAP7_75t_L     g03333(.A1(new_n3362), .A2(new_n3363), .B(new_n3368), .C(new_n3367), .Y(new_n3590));
  AOI221xp5_ASAP7_75t_L     g03334(.A1(new_n3589), .A2(new_n3376), .B1(new_n3573), .B2(new_n3578), .C(new_n3590), .Y(new_n3591));
  OAI21xp33_ASAP7_75t_L     g03335(.A1(new_n3591), .A2(new_n3588), .B(new_n3584), .Y(new_n3592));
  INVx1_ASAP7_75t_L         g03336(.A(new_n3592), .Y(new_n3593));
  MAJIxp5_ASAP7_75t_L       g03337(.A(new_n3393), .B(new_n3387), .C(new_n3378), .Y(new_n3594));
  NOR3xp33_ASAP7_75t_L      g03338(.A(new_n3593), .B(new_n3585), .C(new_n3594), .Y(new_n3595));
  NOR2xp33_ASAP7_75t_L      g03339(.A(new_n3591), .B(new_n3588), .Y(new_n3596));
  NAND2xp33_ASAP7_75t_L     g03340(.A(new_n3583), .B(new_n3596), .Y(new_n3597));
  INVx1_ASAP7_75t_L         g03341(.A(new_n3594), .Y(new_n3598));
  AOI21xp33_ASAP7_75t_L     g03342(.A1(new_n3592), .A2(new_n3597), .B(new_n3598), .Y(new_n3599));
  OAI22xp33_ASAP7_75t_L     g03343(.A1(new_n2881), .A2(new_n367), .B1(new_n2871), .B2(new_n368), .Y(new_n3600));
  AOI221xp5_ASAP7_75t_L     g03344(.A1(\b[27] ), .A2(new_n366), .B1(\b[28] ), .B2(new_n334), .C(new_n3600), .Y(new_n3601));
  XNOR2x2_ASAP7_75t_L       g03345(.A(new_n339), .B(new_n3601), .Y(new_n3602));
  OAI21xp33_ASAP7_75t_L     g03346(.A1(new_n3599), .A2(new_n3595), .B(new_n3602), .Y(new_n3603));
  NAND3xp33_ASAP7_75t_L     g03347(.A(new_n3598), .B(new_n3592), .C(new_n3597), .Y(new_n3604));
  OAI21xp33_ASAP7_75t_L     g03348(.A1(new_n3585), .A2(new_n3593), .B(new_n3594), .Y(new_n3605));
  INVx1_ASAP7_75t_L         g03349(.A(new_n3602), .Y(new_n3606));
  NAND3xp33_ASAP7_75t_L     g03350(.A(new_n3605), .B(new_n3604), .C(new_n3606), .Y(new_n3607));
  NAND3xp33_ASAP7_75t_L     g03351(.A(new_n3457), .B(new_n3603), .C(new_n3607), .Y(new_n3608));
  O2A1O1Ixp33_ASAP7_75t_L   g03352(.A1(new_n3407), .A2(new_n3197), .B(new_n3208), .C(new_n3406), .Y(new_n3609));
  AOI21xp33_ASAP7_75t_L     g03353(.A1(new_n3605), .A2(new_n3604), .B(new_n3606), .Y(new_n3610));
  INVx1_ASAP7_75t_L         g03354(.A(new_n3607), .Y(new_n3611));
  OAI22xp33_ASAP7_75t_L     g03355(.A1(new_n3609), .A2(new_n3456), .B1(new_n3611), .B2(new_n3610), .Y(new_n3612));
  AOI21xp33_ASAP7_75t_L     g03356(.A1(new_n3612), .A2(new_n3608), .B(new_n3455), .Y(new_n3613));
  INVx1_ASAP7_75t_L         g03357(.A(new_n3613), .Y(new_n3614));
  NAND3xp33_ASAP7_75t_L     g03358(.A(new_n3612), .B(new_n3608), .C(new_n3455), .Y(new_n3615));
  NAND2xp33_ASAP7_75t_L     g03359(.A(new_n3615), .B(new_n3614), .Y(new_n3616));
  XNOR2x2_ASAP7_75t_L       g03360(.A(new_n3616), .B(new_n3439), .Y(\f[32] ));
  NOR2xp33_ASAP7_75t_L      g03361(.A(new_n3431), .B(new_n3437), .Y(new_n3618));
  A2O1A1O1Ixp25_ASAP7_75t_L g03362(.A1(new_n3434), .A2(new_n3435), .B(new_n3618), .C(new_n3615), .D(new_n3613), .Y(new_n3619));
  INVx1_ASAP7_75t_L         g03363(.A(new_n3590), .Y(new_n3620));
  A2O1A1Ixp33_ASAP7_75t_L   g03364(.A1(new_n3377), .A2(new_n3620), .B(new_n3586), .C(new_n3578), .Y(new_n3621));
  NOR2xp33_ASAP7_75t_L      g03365(.A(new_n1857), .B(new_n1620), .Y(new_n3622));
  INVx1_ASAP7_75t_L         g03366(.A(new_n3622), .Y(new_n3623));
  NOR2xp33_ASAP7_75t_L      g03367(.A(new_n1995), .B(new_n721), .Y(new_n3624));
  INVx1_ASAP7_75t_L         g03368(.A(new_n3624), .Y(new_n3625));
  AOI22xp33_ASAP7_75t_L     g03369(.A1(new_n600), .A2(\b[24] ), .B1(new_n597), .B2(new_n2027), .Y(new_n3626));
  NAND4xp25_ASAP7_75t_L     g03370(.A(new_n3626), .B(\a[11] ), .C(new_n3623), .D(new_n3625), .Y(new_n3627));
  AOI31xp33_ASAP7_75t_L     g03371(.A1(new_n3626), .A2(new_n3625), .A3(new_n3623), .B(\a[11] ), .Y(new_n3628));
  INVx1_ASAP7_75t_L         g03372(.A(new_n3628), .Y(new_n3629));
  NAND2xp33_ASAP7_75t_L     g03373(.A(new_n3627), .B(new_n3629), .Y(new_n3630));
  AOI211xp5_ASAP7_75t_L     g03374(.A1(new_n3539), .A2(new_n3541), .B(new_n3544), .C(new_n3543), .Y(new_n3631));
  A2O1A1O1Ixp25_ASAP7_75t_L g03375(.A1(new_n3340), .A2(new_n3339), .B(new_n3549), .C(new_n3552), .D(new_n3631), .Y(new_n3632));
  NAND2xp33_ASAP7_75t_L     g03376(.A(\b[16] ), .B(new_n1194), .Y(new_n3633));
  NAND2xp33_ASAP7_75t_L     g03377(.A(\b[17] ), .B(new_n1103), .Y(new_n3634));
  AOI22xp33_ASAP7_75t_L     g03378(.A1(new_n1113), .A2(\b[18] ), .B1(new_n1110), .B2(new_n1363), .Y(new_n3635));
  NAND4xp25_ASAP7_75t_L     g03379(.A(new_n3635), .B(\a[17] ), .C(new_n3633), .D(new_n3634), .Y(new_n3636));
  OAI221xp5_ASAP7_75t_L     g03380(.A1(new_n1198), .A2(new_n1356), .B1(new_n1197), .B2(new_n3138), .C(new_n3634), .Y(new_n3637));
  A2O1A1Ixp33_ASAP7_75t_L   g03381(.A1(\b[16] ), .A2(new_n1194), .B(new_n3637), .C(new_n1107), .Y(new_n3638));
  NAND2xp33_ASAP7_75t_L     g03382(.A(new_n3636), .B(new_n3638), .Y(new_n3639));
  OAI21xp33_ASAP7_75t_L     g03383(.A1(new_n3533), .A2(new_n3532), .B(new_n3530), .Y(new_n3640));
  NAND2xp33_ASAP7_75t_L     g03384(.A(new_n3273), .B(new_n3274), .Y(new_n3641));
  INVx1_ASAP7_75t_L         g03385(.A(new_n3483), .Y(new_n3642));
  O2A1O1Ixp33_ASAP7_75t_L   g03386(.A1(new_n3084), .A2(new_n3237), .B(new_n3641), .C(new_n3642), .Y(new_n3643));
  INVx1_ASAP7_75t_L         g03387(.A(new_n3066), .Y(new_n3644));
  NAND2xp33_ASAP7_75t_L     g03388(.A(\b[0] ), .B(new_n3260), .Y(new_n3645));
  NAND4xp25_ASAP7_75t_L     g03389(.A(new_n3257), .B(\a[32] ), .C(new_n3644), .D(new_n3645), .Y(new_n3646));
  INVx1_ASAP7_75t_L         g03390(.A(\a[33] ), .Y(new_n3647));
  NAND2xp33_ASAP7_75t_L     g03391(.A(\a[32] ), .B(new_n3647), .Y(new_n3648));
  NAND2xp33_ASAP7_75t_L     g03392(.A(\a[33] ), .B(new_n3251), .Y(new_n3649));
  AND2x2_ASAP7_75t_L        g03393(.A(new_n3648), .B(new_n3649), .Y(new_n3650));
  NOR2xp33_ASAP7_75t_L      g03394(.A(new_n258), .B(new_n3650), .Y(new_n3651));
  OAI31xp33_ASAP7_75t_L     g03395(.A1(new_n3646), .A2(new_n3495), .A3(new_n3493), .B(new_n3651), .Y(new_n3652));
  OR4x2_ASAP7_75t_L         g03396(.A(new_n3651), .B(new_n3646), .C(new_n3495), .D(new_n3493), .Y(new_n3653));
  NOR2xp33_ASAP7_75t_L      g03397(.A(new_n278), .B(new_n3248), .Y(new_n3654));
  AOI221xp5_ASAP7_75t_L     g03398(.A1(new_n3256), .A2(\b[3] ), .B1(new_n3254), .B2(new_n1000), .C(new_n3654), .Y(new_n3655));
  OAI211xp5_ASAP7_75t_L     g03399(.A1(new_n276), .A2(new_n3492), .B(new_n3655), .C(\a[32] ), .Y(new_n3656));
  NAND2xp33_ASAP7_75t_L     g03400(.A(\b[3] ), .B(new_n3256), .Y(new_n3657));
  OAI221xp5_ASAP7_75t_L     g03401(.A1(new_n278), .A2(new_n3248), .B1(new_n3261), .B2(new_n303), .C(new_n3657), .Y(new_n3658));
  A2O1A1Ixp33_ASAP7_75t_L   g03402(.A1(\b[1] ), .A2(new_n3491), .B(new_n3658), .C(new_n3251), .Y(new_n3659));
  AO22x1_ASAP7_75t_L        g03403(.A1(new_n3659), .A2(new_n3656), .B1(new_n3652), .B2(new_n3653), .Y(new_n3660));
  NAND4xp25_ASAP7_75t_L     g03404(.A(new_n3653), .B(new_n3652), .C(new_n3656), .D(new_n3659), .Y(new_n3661));
  NAND2xp33_ASAP7_75t_L     g03405(.A(\b[4] ), .B(new_n2931), .Y(new_n3662));
  NAND2xp33_ASAP7_75t_L     g03406(.A(\b[5] ), .B(new_n2706), .Y(new_n3663));
  AOI22xp33_ASAP7_75t_L     g03407(.A1(new_n2702), .A2(\b[6] ), .B1(new_n2700), .B2(new_n389), .Y(new_n3664));
  NAND4xp25_ASAP7_75t_L     g03408(.A(new_n3664), .B(\a[29] ), .C(new_n3662), .D(new_n3663), .Y(new_n3665));
  NAND2xp33_ASAP7_75t_L     g03409(.A(\b[6] ), .B(new_n2702), .Y(new_n3666));
  OAI211xp5_ASAP7_75t_L     g03410(.A1(new_n2707), .A2(new_n540), .B(new_n3663), .C(new_n3666), .Y(new_n3667));
  A2O1A1Ixp33_ASAP7_75t_L   g03411(.A1(\b[4] ), .A2(new_n2931), .B(new_n3667), .C(new_n2697), .Y(new_n3668));
  NAND4xp25_ASAP7_75t_L     g03412(.A(new_n3660), .B(new_n3668), .C(new_n3665), .D(new_n3661), .Y(new_n3669));
  AOI22xp33_ASAP7_75t_L     g03413(.A1(new_n3656), .A2(new_n3659), .B1(new_n3652), .B2(new_n3653), .Y(new_n3670));
  AND4x1_ASAP7_75t_L        g03414(.A(new_n3653), .B(new_n3652), .C(new_n3659), .D(new_n3656), .Y(new_n3671));
  AOI211xp5_ASAP7_75t_L     g03415(.A1(\b[4] ), .A2(new_n2931), .B(new_n2697), .C(new_n3667), .Y(new_n3672));
  AOI31xp33_ASAP7_75t_L     g03416(.A1(new_n3664), .A2(new_n3663), .A3(new_n3662), .B(\a[29] ), .Y(new_n3673));
  OAI22xp33_ASAP7_75t_L     g03417(.A1(new_n3672), .A2(new_n3673), .B1(new_n3670), .B2(new_n3671), .Y(new_n3674));
  NAND2xp33_ASAP7_75t_L     g03418(.A(new_n3669), .B(new_n3674), .Y(new_n3675));
  O2A1O1Ixp33_ASAP7_75t_L   g03419(.A1(new_n3643), .A2(new_n3498), .B(new_n3500), .C(new_n3675), .Y(new_n3676));
  NOR4xp25_ASAP7_75t_L      g03420(.A(new_n3672), .B(new_n3673), .C(new_n3671), .D(new_n3670), .Y(new_n3677));
  AOI22xp33_ASAP7_75t_L     g03421(.A1(new_n3668), .A2(new_n3665), .B1(new_n3660), .B2(new_n3661), .Y(new_n3678));
  NOR2xp33_ASAP7_75t_L      g03422(.A(new_n3678), .B(new_n3677), .Y(new_n3679));
  A2O1A1Ixp33_ASAP7_75t_L   g03423(.A1(new_n3270), .A2(new_n3483), .B(new_n3498), .C(new_n3500), .Y(new_n3680));
  NOR2xp33_ASAP7_75t_L      g03424(.A(new_n3680), .B(new_n3679), .Y(new_n3681));
  NOR2xp33_ASAP7_75t_L      g03425(.A(new_n421), .B(new_n2387), .Y(new_n3682));
  INVx1_ASAP7_75t_L         g03426(.A(new_n3682), .Y(new_n3683));
  NAND2xp33_ASAP7_75t_L     g03427(.A(\b[8] ), .B(new_n2232), .Y(new_n3684));
  AOI22xp33_ASAP7_75t_L     g03428(.A1(new_n2228), .A2(\b[9] ), .B1(new_n2226), .B2(new_n566), .Y(new_n3685));
  NAND4xp25_ASAP7_75t_L     g03429(.A(new_n3685), .B(\a[26] ), .C(new_n3683), .D(new_n3684), .Y(new_n3686));
  OAI221xp5_ASAP7_75t_L     g03430(.A1(new_n2234), .A2(new_n559), .B1(new_n2233), .B2(new_n978), .C(new_n3684), .Y(new_n3687));
  A2O1A1Ixp33_ASAP7_75t_L   g03431(.A1(\b[7] ), .A2(new_n2386), .B(new_n3687), .C(new_n2223), .Y(new_n3688));
  NAND2xp33_ASAP7_75t_L     g03432(.A(new_n3686), .B(new_n3688), .Y(new_n3689));
  OAI21xp33_ASAP7_75t_L     g03433(.A1(new_n3676), .A2(new_n3681), .B(new_n3689), .Y(new_n3690));
  NAND2xp33_ASAP7_75t_L     g03434(.A(new_n3680), .B(new_n3679), .Y(new_n3691));
  AND2x2_ASAP7_75t_L        g03435(.A(new_n3074), .B(new_n3071), .Y(new_n3692));
  A2O1A1Ixp33_ASAP7_75t_L   g03436(.A1(new_n3068), .A2(new_n3067), .B(new_n3692), .C(new_n3236), .Y(new_n3693));
  A2O1A1O1Ixp25_ASAP7_75t_L g03437(.A1(new_n3641), .A2(new_n3693), .B(new_n3642), .C(new_n3499), .D(new_n3503), .Y(new_n3694));
  NAND2xp33_ASAP7_75t_L     g03438(.A(new_n3694), .B(new_n3675), .Y(new_n3695));
  NAND4xp25_ASAP7_75t_L     g03439(.A(new_n3691), .B(new_n3695), .C(new_n3688), .D(new_n3686), .Y(new_n3696));
  AOI221xp5_ASAP7_75t_L     g03440(.A1(new_n3506), .A2(new_n3509), .B1(new_n3696), .B2(new_n3690), .C(new_n3505), .Y(new_n3697));
  A2O1A1O1Ixp25_ASAP7_75t_L g03441(.A1(new_n3280), .A2(new_n3229), .B(new_n3285), .C(new_n3506), .D(new_n3505), .Y(new_n3698));
  AOI22xp33_ASAP7_75t_L     g03442(.A1(new_n3686), .A2(new_n3688), .B1(new_n3695), .B2(new_n3691), .Y(new_n3699));
  AND4x1_ASAP7_75t_L        g03443(.A(new_n3691), .B(new_n3688), .C(new_n3695), .D(new_n3686), .Y(new_n3700));
  NOR3xp33_ASAP7_75t_L      g03444(.A(new_n3698), .B(new_n3700), .C(new_n3699), .Y(new_n3701));
  NOR2xp33_ASAP7_75t_L      g03445(.A(new_n631), .B(new_n1911), .Y(new_n3702));
  NAND2xp33_ASAP7_75t_L     g03446(.A(\b[12] ), .B(new_n1766), .Y(new_n3703));
  OAI221xp5_ASAP7_75t_L     g03447(.A1(new_n695), .A2(new_n1758), .B1(new_n1771), .B2(new_n775), .C(new_n3703), .Y(new_n3704));
  OR3x1_ASAP7_75t_L         g03448(.A(new_n3704), .B(new_n1761), .C(new_n3702), .Y(new_n3705));
  A2O1A1Ixp33_ASAP7_75t_L   g03449(.A1(\b[10] ), .A2(new_n1910), .B(new_n3704), .C(new_n1761), .Y(new_n3706));
  OA211x2_ASAP7_75t_L       g03450(.A1(new_n3701), .A2(new_n3697), .B(new_n3706), .C(new_n3705), .Y(new_n3707));
  AOI211xp5_ASAP7_75t_L     g03451(.A1(new_n3705), .A2(new_n3706), .B(new_n3701), .C(new_n3697), .Y(new_n3708));
  NAND2xp33_ASAP7_75t_L     g03452(.A(new_n3295), .B(new_n3299), .Y(new_n3709));
  A2O1A1Ixp33_ASAP7_75t_L   g03453(.A1(new_n3709), .A2(new_n3306), .B(new_n3475), .C(new_n3519), .Y(new_n3710));
  AOI211xp5_ASAP7_75t_L     g03454(.A1(new_n3710), .A2(new_n3520), .B(new_n3707), .C(new_n3708), .Y(new_n3711));
  OAI211xp5_ASAP7_75t_L     g03455(.A1(new_n3701), .A2(new_n3697), .B(new_n3705), .C(new_n3706), .Y(new_n3712));
  NOR2xp33_ASAP7_75t_L      g03456(.A(new_n3701), .B(new_n3697), .Y(new_n3713));
  NAND2xp33_ASAP7_75t_L     g03457(.A(new_n3706), .B(new_n3705), .Y(new_n3714));
  NAND2xp33_ASAP7_75t_L     g03458(.A(new_n3714), .B(new_n3713), .Y(new_n3715));
  A2O1A1Ixp33_ASAP7_75t_L   g03459(.A1(new_n3307), .A2(new_n3474), .B(new_n3523), .C(new_n3520), .Y(new_n3716));
  AOI21xp33_ASAP7_75t_L     g03460(.A1(new_n3715), .A2(new_n3712), .B(new_n3716), .Y(new_n3717));
  NAND2xp33_ASAP7_75t_L     g03461(.A(\b[13] ), .B(new_n1548), .Y(new_n3718));
  NAND2xp33_ASAP7_75t_L     g03462(.A(\b[14] ), .B(new_n1410), .Y(new_n3719));
  AOI22xp33_ASAP7_75t_L     g03463(.A1(new_n1406), .A2(\b[15] ), .B1(new_n1404), .B2(new_n959), .Y(new_n3720));
  NAND4xp25_ASAP7_75t_L     g03464(.A(new_n3720), .B(\a[20] ), .C(new_n3718), .D(new_n3719), .Y(new_n3721));
  OAI221xp5_ASAP7_75t_L     g03465(.A1(new_n1412), .A2(new_n952), .B1(new_n1411), .B2(new_n2573), .C(new_n3719), .Y(new_n3722));
  A2O1A1Ixp33_ASAP7_75t_L   g03466(.A1(\b[13] ), .A2(new_n1548), .B(new_n3722), .C(new_n1401), .Y(new_n3723));
  NAND2xp33_ASAP7_75t_L     g03467(.A(new_n3721), .B(new_n3723), .Y(new_n3724));
  NOR3xp33_ASAP7_75t_L      g03468(.A(new_n3711), .B(new_n3717), .C(new_n3724), .Y(new_n3725));
  NAND3xp33_ASAP7_75t_L     g03469(.A(new_n3716), .B(new_n3715), .C(new_n3712), .Y(new_n3726));
  OAI211xp5_ASAP7_75t_L     g03470(.A1(new_n3708), .A2(new_n3707), .B(new_n3520), .C(new_n3710), .Y(new_n3727));
  INVx1_ASAP7_75t_L         g03471(.A(new_n3724), .Y(new_n3728));
  AOI21xp33_ASAP7_75t_L     g03472(.A1(new_n3727), .A2(new_n3726), .B(new_n3728), .Y(new_n3729));
  OAI21xp33_ASAP7_75t_L     g03473(.A1(new_n3725), .A2(new_n3729), .B(new_n3640), .Y(new_n3730));
  A2O1A1O1Ixp25_ASAP7_75t_L g03474(.A1(new_n3319), .A2(new_n3334), .B(new_n3316), .C(new_n3526), .D(new_n3534), .Y(new_n3731));
  NAND3xp33_ASAP7_75t_L     g03475(.A(new_n3728), .B(new_n3727), .C(new_n3726), .Y(new_n3732));
  OAI21xp33_ASAP7_75t_L     g03476(.A1(new_n3717), .A2(new_n3711), .B(new_n3724), .Y(new_n3733));
  NAND3xp33_ASAP7_75t_L     g03477(.A(new_n3731), .B(new_n3732), .C(new_n3733), .Y(new_n3734));
  NAND3xp33_ASAP7_75t_L     g03478(.A(new_n3734), .B(new_n3730), .C(new_n3639), .Y(new_n3735));
  AO21x2_ASAP7_75t_L        g03479(.A1(new_n3730), .A2(new_n3734), .B(new_n3639), .Y(new_n3736));
  NAND2xp33_ASAP7_75t_L     g03480(.A(new_n3735), .B(new_n3736), .Y(new_n3737));
  NAND2xp33_ASAP7_75t_L     g03481(.A(new_n3737), .B(new_n3632), .Y(new_n3738));
  AND3x1_ASAP7_75t_L        g03482(.A(new_n3734), .B(new_n3730), .C(new_n3639), .Y(new_n3739));
  AOI21xp33_ASAP7_75t_L     g03483(.A1(new_n3734), .A2(new_n3730), .B(new_n3639), .Y(new_n3740));
  NOR2xp33_ASAP7_75t_L      g03484(.A(new_n3740), .B(new_n3739), .Y(new_n3741));
  A2O1A1Ixp33_ASAP7_75t_L   g03485(.A1(new_n3562), .A2(new_n3552), .B(new_n3631), .C(new_n3741), .Y(new_n3742));
  NOR2xp33_ASAP7_75t_L      g03486(.A(new_n1493), .B(new_n909), .Y(new_n3743));
  INVx1_ASAP7_75t_L         g03487(.A(new_n3743), .Y(new_n3744));
  NOR2xp33_ASAP7_75t_L      g03488(.A(new_n1594), .B(new_n994), .Y(new_n3745));
  INVx1_ASAP7_75t_L         g03489(.A(new_n3745), .Y(new_n3746));
  AOI22xp33_ASAP7_75t_L     g03490(.A1(new_n826), .A2(\b[21] ), .B1(new_n823), .B2(new_n1715), .Y(new_n3747));
  NAND4xp25_ASAP7_75t_L     g03491(.A(new_n3747), .B(\a[14] ), .C(new_n3744), .D(new_n3746), .Y(new_n3748));
  INVx1_ASAP7_75t_L         g03492(.A(new_n3748), .Y(new_n3749));
  AOI31xp33_ASAP7_75t_L     g03493(.A1(new_n3747), .A2(new_n3746), .A3(new_n3744), .B(\a[14] ), .Y(new_n3750));
  NOR2xp33_ASAP7_75t_L      g03494(.A(new_n3750), .B(new_n3749), .Y(new_n3751));
  NAND3xp33_ASAP7_75t_L     g03495(.A(new_n3742), .B(new_n3751), .C(new_n3738), .Y(new_n3752));
  AOI221xp5_ASAP7_75t_L     g03496(.A1(new_n3736), .A2(new_n3735), .B1(new_n3552), .B2(new_n3562), .C(new_n3631), .Y(new_n3753));
  NOR2xp33_ASAP7_75t_L      g03497(.A(new_n3737), .B(new_n3632), .Y(new_n3754));
  INVx1_ASAP7_75t_L         g03498(.A(new_n3750), .Y(new_n3755));
  NAND2xp33_ASAP7_75t_L     g03499(.A(new_n3748), .B(new_n3755), .Y(new_n3756));
  OAI21xp33_ASAP7_75t_L     g03500(.A1(new_n3753), .A2(new_n3754), .B(new_n3756), .Y(new_n3757));
  NAND2xp33_ASAP7_75t_L     g03501(.A(new_n3757), .B(new_n3752), .Y(new_n3758));
  A2O1A1O1Ixp25_ASAP7_75t_L g03502(.A1(new_n3353), .A2(new_n3349), .B(new_n3355), .C(new_n3463), .D(new_n3561), .Y(new_n3759));
  OAI21xp33_ASAP7_75t_L     g03503(.A1(new_n3759), .A2(new_n3566), .B(new_n3758), .Y(new_n3760));
  A2O1A1O1Ixp25_ASAP7_75t_L g03504(.A1(new_n3357), .A2(new_n3366), .B(new_n3464), .C(new_n3569), .D(new_n3566), .Y(new_n3761));
  NAND3xp33_ASAP7_75t_L     g03505(.A(new_n3761), .B(new_n3757), .C(new_n3752), .Y(new_n3762));
  AOI21xp33_ASAP7_75t_L     g03506(.A1(new_n3760), .A2(new_n3762), .B(new_n3630), .Y(new_n3763));
  INVx1_ASAP7_75t_L         g03507(.A(new_n3627), .Y(new_n3764));
  NOR2xp33_ASAP7_75t_L      g03508(.A(new_n3628), .B(new_n3764), .Y(new_n3765));
  AOI21xp33_ASAP7_75t_L     g03509(.A1(new_n3757), .A2(new_n3752), .B(new_n3761), .Y(new_n3766));
  A2O1A1Ixp33_ASAP7_75t_L   g03510(.A1(new_n3366), .A2(new_n3357), .B(new_n3464), .C(new_n3569), .Y(new_n3767));
  AND4x1_ASAP7_75t_L        g03511(.A(new_n3767), .B(new_n3757), .C(new_n3752), .D(new_n3570), .Y(new_n3768));
  NOR3xp33_ASAP7_75t_L      g03512(.A(new_n3768), .B(new_n3766), .C(new_n3765), .Y(new_n3769));
  NOR2xp33_ASAP7_75t_L      g03513(.A(new_n3769), .B(new_n3763), .Y(new_n3770));
  NAND2xp33_ASAP7_75t_L     g03514(.A(new_n3621), .B(new_n3770), .Y(new_n3771));
  A2O1A1O1Ixp25_ASAP7_75t_L g03515(.A1(new_n3376), .A2(new_n3589), .B(new_n3590), .C(new_n3573), .D(new_n3587), .Y(new_n3772));
  OAI21xp33_ASAP7_75t_L     g03516(.A1(new_n3766), .A2(new_n3768), .B(new_n3765), .Y(new_n3773));
  NAND3xp33_ASAP7_75t_L     g03517(.A(new_n3760), .B(new_n3630), .C(new_n3762), .Y(new_n3774));
  NAND2xp33_ASAP7_75t_L     g03518(.A(new_n3773), .B(new_n3774), .Y(new_n3775));
  NAND2xp33_ASAP7_75t_L     g03519(.A(new_n3772), .B(new_n3775), .Y(new_n3776));
  NAND2xp33_ASAP7_75t_L     g03520(.A(\b[25] ), .B(new_n480), .Y(new_n3777));
  NAND2xp33_ASAP7_75t_L     g03521(.A(\b[26] ), .B(new_n441), .Y(new_n3778));
  AOI22xp33_ASAP7_75t_L     g03522(.A1(new_n451), .A2(\b[27] ), .B1(new_n448), .B2(new_n2657), .Y(new_n3779));
  AND4x1_ASAP7_75t_L        g03523(.A(new_n3779), .B(new_n3778), .C(new_n3777), .D(\a[8] ), .Y(new_n3780));
  AOI31xp33_ASAP7_75t_L     g03524(.A1(new_n3779), .A2(new_n3778), .A3(new_n3777), .B(\a[8] ), .Y(new_n3781));
  NOR2xp33_ASAP7_75t_L      g03525(.A(new_n3781), .B(new_n3780), .Y(new_n3782));
  NAND3xp33_ASAP7_75t_L     g03526(.A(new_n3771), .B(new_n3776), .C(new_n3782), .Y(new_n3783));
  AO21x2_ASAP7_75t_L        g03527(.A1(new_n3776), .A2(new_n3771), .B(new_n3782), .Y(new_n3784));
  MAJIxp5_ASAP7_75t_L       g03528(.A(new_n3594), .B(new_n3584), .C(new_n3596), .Y(new_n3785));
  NAND3xp33_ASAP7_75t_L     g03529(.A(new_n3785), .B(new_n3784), .C(new_n3783), .Y(new_n3786));
  AOI21xp33_ASAP7_75t_L     g03530(.A1(new_n3784), .A2(new_n3783), .B(new_n3785), .Y(new_n3787));
  INVx1_ASAP7_75t_L         g03531(.A(new_n3787), .Y(new_n3788));
  NAND2xp33_ASAP7_75t_L     g03532(.A(new_n342), .B(new_n3219), .Y(new_n3789));
  OAI221xp5_ASAP7_75t_L     g03533(.A1(new_n368), .A2(new_n3212), .B1(new_n2871), .B2(new_n406), .C(new_n3789), .Y(new_n3790));
  AOI21xp33_ASAP7_75t_L     g03534(.A1(new_n366), .A2(\b[28] ), .B(new_n3790), .Y(new_n3791));
  NAND2xp33_ASAP7_75t_L     g03535(.A(\a[5] ), .B(new_n3791), .Y(new_n3792));
  A2O1A1Ixp33_ASAP7_75t_L   g03536(.A1(\b[28] ), .A2(new_n366), .B(new_n3790), .C(new_n339), .Y(new_n3793));
  AND2x2_ASAP7_75t_L        g03537(.A(new_n3793), .B(new_n3792), .Y(new_n3794));
  NAND3xp33_ASAP7_75t_L     g03538(.A(new_n3794), .B(new_n3788), .C(new_n3786), .Y(new_n3795));
  INVx1_ASAP7_75t_L         g03539(.A(new_n3786), .Y(new_n3796));
  NAND2xp33_ASAP7_75t_L     g03540(.A(new_n3793), .B(new_n3792), .Y(new_n3797));
  OAI21xp33_ASAP7_75t_L     g03541(.A1(new_n3787), .A2(new_n3796), .B(new_n3797), .Y(new_n3798));
  NAND2xp33_ASAP7_75t_L     g03542(.A(new_n3798), .B(new_n3795), .Y(new_n3799));
  O2A1O1Ixp33_ASAP7_75t_L   g03543(.A1(new_n3457), .A2(new_n3610), .B(new_n3607), .C(new_n3799), .Y(new_n3800));
  INVx1_ASAP7_75t_L         g03544(.A(new_n3456), .Y(new_n3801));
  A2O1A1Ixp33_ASAP7_75t_L   g03545(.A1(new_n3415), .A2(new_n3801), .B(new_n3610), .C(new_n3607), .Y(new_n3802));
  AOI21xp33_ASAP7_75t_L     g03546(.A1(new_n3798), .A2(new_n3795), .B(new_n3802), .Y(new_n3803));
  O2A1O1Ixp33_ASAP7_75t_L   g03547(.A1(new_n3213), .A2(new_n3216), .B(new_n3421), .C(new_n3420), .Y(new_n3804));
  INVx1_ASAP7_75t_L         g03548(.A(new_n3444), .Y(new_n3805));
  NOR2xp33_ASAP7_75t_L      g03549(.A(\b[32] ), .B(\b[33] ), .Y(new_n3806));
  INVx1_ASAP7_75t_L         g03550(.A(\b[33] ), .Y(new_n3807));
  NOR2xp33_ASAP7_75t_L      g03551(.A(new_n3443), .B(new_n3807), .Y(new_n3808));
  NOR2xp33_ASAP7_75t_L      g03552(.A(new_n3806), .B(new_n3808), .Y(new_n3809));
  INVx1_ASAP7_75t_L         g03553(.A(new_n3809), .Y(new_n3810));
  O2A1O1Ixp33_ASAP7_75t_L   g03554(.A1(new_n3446), .A2(new_n3804), .B(new_n3805), .C(new_n3810), .Y(new_n3811));
  NOR3xp33_ASAP7_75t_L      g03555(.A(new_n3447), .B(new_n3809), .C(new_n3444), .Y(new_n3812));
  NOR2xp33_ASAP7_75t_L      g03556(.A(new_n3811), .B(new_n3812), .Y(new_n3813));
  AOI22xp33_ASAP7_75t_L     g03557(.A1(new_n272), .A2(\b[33] ), .B1(new_n269), .B2(new_n3813), .Y(new_n3814));
  OAI221xp5_ASAP7_75t_L     g03558(.A1(new_n261), .A2(new_n3443), .B1(new_n3419), .B2(new_n277), .C(new_n3814), .Y(new_n3815));
  XNOR2x2_ASAP7_75t_L       g03559(.A(new_n265), .B(new_n3815), .Y(new_n3816));
  OAI21xp33_ASAP7_75t_L     g03560(.A1(new_n3803), .A2(new_n3800), .B(new_n3816), .Y(new_n3817));
  INVx1_ASAP7_75t_L         g03561(.A(new_n3817), .Y(new_n3818));
  NOR3xp33_ASAP7_75t_L      g03562(.A(new_n3800), .B(new_n3803), .C(new_n3816), .Y(new_n3819));
  NOR3xp33_ASAP7_75t_L      g03563(.A(new_n3818), .B(new_n3819), .C(new_n3619), .Y(new_n3820));
  INVx1_ASAP7_75t_L         g03564(.A(new_n3619), .Y(new_n3821));
  NOR2xp33_ASAP7_75t_L      g03565(.A(new_n3819), .B(new_n3818), .Y(new_n3822));
  NOR2xp33_ASAP7_75t_L      g03566(.A(new_n3821), .B(new_n3822), .Y(new_n3823));
  NOR2xp33_ASAP7_75t_L      g03567(.A(new_n3820), .B(new_n3823), .Y(\f[33] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03568(.A1(new_n3448), .A2(new_n3445), .B(new_n3444), .C(new_n3809), .Y(new_n3825));
  NOR2xp33_ASAP7_75t_L      g03569(.A(\b[33] ), .B(\b[34] ), .Y(new_n3826));
  INVx1_ASAP7_75t_L         g03570(.A(\b[34] ), .Y(new_n3827));
  NOR2xp33_ASAP7_75t_L      g03571(.A(new_n3807), .B(new_n3827), .Y(new_n3828));
  NOR2xp33_ASAP7_75t_L      g03572(.A(new_n3826), .B(new_n3828), .Y(new_n3829));
  INVx1_ASAP7_75t_L         g03573(.A(new_n3829), .Y(new_n3830));
  O2A1O1Ixp33_ASAP7_75t_L   g03574(.A1(new_n3443), .A2(new_n3807), .B(new_n3825), .C(new_n3830), .Y(new_n3831));
  NOR3xp33_ASAP7_75t_L      g03575(.A(new_n3811), .B(new_n3829), .C(new_n3808), .Y(new_n3832));
  NOR2xp33_ASAP7_75t_L      g03576(.A(new_n3832), .B(new_n3831), .Y(new_n3833));
  AOI22xp33_ASAP7_75t_L     g03577(.A1(new_n272), .A2(\b[34] ), .B1(new_n269), .B2(new_n3833), .Y(new_n3834));
  OAI221xp5_ASAP7_75t_L     g03578(.A1(new_n261), .A2(new_n3807), .B1(new_n3443), .B2(new_n277), .C(new_n3834), .Y(new_n3835));
  XNOR2x2_ASAP7_75t_L       g03579(.A(\a[2] ), .B(new_n3835), .Y(new_n3836));
  O2A1O1Ixp33_ASAP7_75t_L   g03580(.A1(new_n3406), .A2(new_n3409), .B(new_n3801), .C(new_n3610), .Y(new_n3837));
  NOR3xp33_ASAP7_75t_L      g03581(.A(new_n3794), .B(new_n3787), .C(new_n3796), .Y(new_n3838));
  O2A1O1Ixp33_ASAP7_75t_L   g03582(.A1(new_n3611), .A2(new_n3837), .B(new_n3799), .C(new_n3838), .Y(new_n3839));
  AOI22xp33_ASAP7_75t_L     g03583(.A1(new_n451), .A2(\b[28] ), .B1(new_n448), .B2(new_n2858), .Y(new_n3840));
  OAI221xp5_ASAP7_75t_L     g03584(.A1(new_n529), .A2(new_n2650), .B1(new_n2477), .B2(new_n481), .C(new_n3840), .Y(new_n3841));
  XNOR2x2_ASAP7_75t_L       g03585(.A(\a[8] ), .B(new_n3841), .Y(new_n3842));
  OAI21xp33_ASAP7_75t_L     g03586(.A1(new_n3763), .A2(new_n3772), .B(new_n3774), .Y(new_n3843));
  NAND3xp33_ASAP7_75t_L     g03587(.A(new_n3726), .B(new_n3727), .C(new_n3724), .Y(new_n3844));
  NAND2xp33_ASAP7_75t_L     g03588(.A(\b[14] ), .B(new_n1548), .Y(new_n3845));
  NAND2xp33_ASAP7_75t_L     g03589(.A(\b[15] ), .B(new_n1410), .Y(new_n3846));
  AOI22xp33_ASAP7_75t_L     g03590(.A1(new_n1406), .A2(\b[16] ), .B1(new_n1404), .B2(new_n1058), .Y(new_n3847));
  AND4x1_ASAP7_75t_L        g03591(.A(new_n3847), .B(new_n3846), .C(new_n3845), .D(\a[20] ), .Y(new_n3848));
  AOI31xp33_ASAP7_75t_L     g03592(.A1(new_n3847), .A2(new_n3846), .A3(new_n3845), .B(\a[20] ), .Y(new_n3849));
  OR2x4_ASAP7_75t_L         g03593(.A(new_n3849), .B(new_n3848), .Y(new_n3850));
  A2O1A1O1Ixp25_ASAP7_75t_L g03594(.A1(new_n3519), .A2(new_n3522), .B(new_n3524), .C(new_n3712), .D(new_n3708), .Y(new_n3851));
  AOI211xp5_ASAP7_75t_L     g03595(.A1(new_n3668), .A2(new_n3665), .B(new_n3670), .C(new_n3671), .Y(new_n3852));
  INVx1_ASAP7_75t_L         g03596(.A(new_n3852), .Y(new_n3853));
  A2O1A1Ixp33_ASAP7_75t_L   g03597(.A1(new_n3674), .A2(new_n3669), .B(new_n3694), .C(new_n3853), .Y(new_n3854));
  NAND2xp33_ASAP7_75t_L     g03598(.A(\b[5] ), .B(new_n2931), .Y(new_n3855));
  NAND2xp33_ASAP7_75t_L     g03599(.A(\b[6] ), .B(new_n2706), .Y(new_n3856));
  AOI32xp33_ASAP7_75t_L     g03600(.A1(new_n424), .A2(new_n426), .A3(new_n2700), .B1(new_n2702), .B2(\b[7] ), .Y(new_n3857));
  NAND4xp25_ASAP7_75t_L     g03601(.A(new_n3857), .B(\a[29] ), .C(new_n3855), .D(new_n3856), .Y(new_n3858));
  NAND2xp33_ASAP7_75t_L     g03602(.A(new_n3856), .B(new_n3857), .Y(new_n3859));
  A2O1A1Ixp33_ASAP7_75t_L   g03603(.A1(\b[5] ), .A2(new_n2931), .B(new_n3859), .C(new_n2697), .Y(new_n3860));
  NOR3xp33_ASAP7_75t_L      g03604(.A(new_n3646), .B(new_n3493), .C(new_n3495), .Y(new_n3861));
  NAND2xp33_ASAP7_75t_L     g03605(.A(new_n3659), .B(new_n3656), .Y(new_n3862));
  MAJIxp5_ASAP7_75t_L       g03606(.A(new_n3862), .B(new_n3651), .C(new_n3861), .Y(new_n3863));
  NAND2xp33_ASAP7_75t_L     g03607(.A(\b[2] ), .B(new_n3491), .Y(new_n3864));
  INVx1_ASAP7_75t_L         g03608(.A(new_n3864), .Y(new_n3865));
  NOR2xp33_ASAP7_75t_L      g03609(.A(new_n299), .B(new_n3248), .Y(new_n3866));
  OAI32xp33_ASAP7_75t_L     g03610(.A1(new_n325), .A2(new_n327), .A3(new_n3261), .B1(new_n323), .B2(new_n3262), .Y(new_n3867));
  NOR4xp25_ASAP7_75t_L      g03611(.A(new_n3865), .B(new_n3867), .C(new_n3251), .D(new_n3866), .Y(new_n3868));
  NOR2xp33_ASAP7_75t_L      g03612(.A(new_n3866), .B(new_n3867), .Y(new_n3869));
  AOI21xp33_ASAP7_75t_L     g03613(.A1(new_n3869), .A2(new_n3864), .B(\a[32] ), .Y(new_n3870));
  NAND2xp33_ASAP7_75t_L     g03614(.A(\a[35] ), .B(new_n3651), .Y(new_n3871));
  NAND2xp33_ASAP7_75t_L     g03615(.A(new_n3649), .B(new_n3648), .Y(new_n3872));
  XNOR2x2_ASAP7_75t_L       g03616(.A(\a[34] ), .B(\a[33] ), .Y(new_n3873));
  NOR2xp33_ASAP7_75t_L      g03617(.A(new_n3873), .B(new_n3872), .Y(new_n3874));
  NAND2xp33_ASAP7_75t_L     g03618(.A(\b[0] ), .B(new_n3874), .Y(new_n3875));
  INVx1_ASAP7_75t_L         g03619(.A(\a[34] ), .Y(new_n3876));
  NAND2xp33_ASAP7_75t_L     g03620(.A(\a[35] ), .B(new_n3876), .Y(new_n3877));
  INVx1_ASAP7_75t_L         g03621(.A(\a[35] ), .Y(new_n3878));
  NAND2xp33_ASAP7_75t_L     g03622(.A(\a[34] ), .B(new_n3878), .Y(new_n3879));
  AND2x2_ASAP7_75t_L        g03623(.A(new_n3877), .B(new_n3879), .Y(new_n3880));
  NOR2xp33_ASAP7_75t_L      g03624(.A(new_n3650), .B(new_n3880), .Y(new_n3881));
  NAND2xp33_ASAP7_75t_L     g03625(.A(new_n271), .B(new_n3881), .Y(new_n3882));
  NAND2xp33_ASAP7_75t_L     g03626(.A(new_n3879), .B(new_n3877), .Y(new_n3883));
  NOR2xp33_ASAP7_75t_L      g03627(.A(new_n3883), .B(new_n3650), .Y(new_n3884));
  NAND2xp33_ASAP7_75t_L     g03628(.A(\b[1] ), .B(new_n3884), .Y(new_n3885));
  NAND3xp33_ASAP7_75t_L     g03629(.A(new_n3882), .B(new_n3885), .C(new_n3875), .Y(new_n3886));
  XNOR2x2_ASAP7_75t_L       g03630(.A(new_n3871), .B(new_n3886), .Y(new_n3887));
  NOR3xp33_ASAP7_75t_L      g03631(.A(new_n3887), .B(new_n3870), .C(new_n3868), .Y(new_n3888));
  OA21x2_ASAP7_75t_L        g03632(.A1(new_n3868), .A2(new_n3870), .B(new_n3887), .Y(new_n3889));
  NOR3xp33_ASAP7_75t_L      g03633(.A(new_n3863), .B(new_n3888), .C(new_n3889), .Y(new_n3890));
  NAND2xp33_ASAP7_75t_L     g03634(.A(new_n3651), .B(new_n3861), .Y(new_n3891));
  INVx1_ASAP7_75t_L         g03635(.A(new_n3891), .Y(new_n3892));
  NAND3xp33_ASAP7_75t_L     g03636(.A(new_n3886), .B(new_n3651), .C(\a[35] ), .Y(new_n3893));
  AND3x1_ASAP7_75t_L        g03637(.A(new_n3882), .B(new_n3885), .C(new_n3875), .Y(new_n3894));
  NAND2xp33_ASAP7_75t_L     g03638(.A(new_n3871), .B(new_n3894), .Y(new_n3895));
  AO211x2_ASAP7_75t_L       g03639(.A1(new_n3895), .A2(new_n3893), .B(new_n3868), .C(new_n3870), .Y(new_n3896));
  OAI21xp33_ASAP7_75t_L     g03640(.A1(new_n3870), .A2(new_n3868), .B(new_n3887), .Y(new_n3897));
  AOI211xp5_ASAP7_75t_L     g03641(.A1(new_n3896), .A2(new_n3897), .B(new_n3892), .C(new_n3670), .Y(new_n3898));
  OAI211xp5_ASAP7_75t_L     g03642(.A1(new_n3898), .A2(new_n3890), .B(new_n3860), .C(new_n3858), .Y(new_n3899));
  INVx1_ASAP7_75t_L         g03643(.A(new_n3858), .Y(new_n3900));
  INVx1_ASAP7_75t_L         g03644(.A(new_n3860), .Y(new_n3901));
  AND2x2_ASAP7_75t_L        g03645(.A(new_n3659), .B(new_n3656), .Y(new_n3902));
  A2O1A1Ixp33_ASAP7_75t_L   g03646(.A1(new_n3653), .A2(new_n3652), .B(new_n3902), .C(new_n3891), .Y(new_n3903));
  NAND3xp33_ASAP7_75t_L     g03647(.A(new_n3903), .B(new_n3896), .C(new_n3897), .Y(new_n3904));
  OAI21xp33_ASAP7_75t_L     g03648(.A1(new_n3888), .A2(new_n3889), .B(new_n3863), .Y(new_n3905));
  OAI211xp5_ASAP7_75t_L     g03649(.A1(new_n3900), .A2(new_n3901), .B(new_n3904), .C(new_n3905), .Y(new_n3906));
  NAND3xp33_ASAP7_75t_L     g03650(.A(new_n3854), .B(new_n3899), .C(new_n3906), .Y(new_n3907));
  A2O1A1O1Ixp25_ASAP7_75t_L g03651(.A1(new_n3273), .A2(new_n3274), .B(new_n3272), .C(new_n3483), .D(new_n3498), .Y(new_n3908));
  O2A1O1Ixp33_ASAP7_75t_L   g03652(.A1(new_n3503), .A2(new_n3908), .B(new_n3675), .C(new_n3852), .Y(new_n3909));
  AOI211xp5_ASAP7_75t_L     g03653(.A1(new_n3904), .A2(new_n3905), .B(new_n3901), .C(new_n3900), .Y(new_n3910));
  AOI211xp5_ASAP7_75t_L     g03654(.A1(new_n3860), .A2(new_n3858), .B(new_n3898), .C(new_n3890), .Y(new_n3911));
  OAI21xp33_ASAP7_75t_L     g03655(.A1(new_n3910), .A2(new_n3911), .B(new_n3909), .Y(new_n3912));
  NAND2xp33_ASAP7_75t_L     g03656(.A(\b[9] ), .B(new_n2232), .Y(new_n3913));
  NAND2xp33_ASAP7_75t_L     g03657(.A(\b[10] ), .B(new_n2228), .Y(new_n3914));
  OAI311xp33_ASAP7_75t_L    g03658(.A1(new_n639), .A2(new_n851), .A3(new_n2233), .B1(new_n3914), .C1(new_n3913), .Y(new_n3915));
  AOI21xp33_ASAP7_75t_L     g03659(.A1(new_n2386), .A2(\b[8] ), .B(new_n3915), .Y(new_n3916));
  NAND2xp33_ASAP7_75t_L     g03660(.A(\a[26] ), .B(new_n3916), .Y(new_n3917));
  A2O1A1Ixp33_ASAP7_75t_L   g03661(.A1(\b[8] ), .A2(new_n2386), .B(new_n3915), .C(new_n2223), .Y(new_n3918));
  AND2x2_ASAP7_75t_L        g03662(.A(new_n3918), .B(new_n3917), .Y(new_n3919));
  NAND3xp33_ASAP7_75t_L     g03663(.A(new_n3919), .B(new_n3912), .C(new_n3907), .Y(new_n3920));
  OAI22xp33_ASAP7_75t_L     g03664(.A1(new_n3908), .A2(new_n3503), .B1(new_n3677), .B2(new_n3678), .Y(new_n3921));
  AOI211xp5_ASAP7_75t_L     g03665(.A1(new_n3921), .A2(new_n3853), .B(new_n3911), .C(new_n3910), .Y(new_n3922));
  AOI21xp33_ASAP7_75t_L     g03666(.A1(new_n3906), .A2(new_n3899), .B(new_n3854), .Y(new_n3923));
  NAND2xp33_ASAP7_75t_L     g03667(.A(new_n3918), .B(new_n3917), .Y(new_n3924));
  OAI21xp33_ASAP7_75t_L     g03668(.A1(new_n3922), .A2(new_n3923), .B(new_n3924), .Y(new_n3925));
  A2O1A1O1Ixp25_ASAP7_75t_L g03669(.A1(new_n3506), .A2(new_n3509), .B(new_n3505), .C(new_n3696), .D(new_n3699), .Y(new_n3926));
  NAND3xp33_ASAP7_75t_L     g03670(.A(new_n3926), .B(new_n3925), .C(new_n3920), .Y(new_n3927));
  NOR3xp33_ASAP7_75t_L      g03671(.A(new_n3923), .B(new_n3922), .C(new_n3924), .Y(new_n3928));
  AOI21xp33_ASAP7_75t_L     g03672(.A1(new_n3912), .A2(new_n3907), .B(new_n3919), .Y(new_n3929));
  OAI21xp33_ASAP7_75t_L     g03673(.A1(new_n3700), .A2(new_n3698), .B(new_n3690), .Y(new_n3930));
  OAI21xp33_ASAP7_75t_L     g03674(.A1(new_n3928), .A2(new_n3929), .B(new_n3930), .Y(new_n3931));
  NAND2xp33_ASAP7_75t_L     g03675(.A(\b[12] ), .B(new_n1770), .Y(new_n3932));
  NAND2xp33_ASAP7_75t_L     g03676(.A(\b[13] ), .B(new_n1766), .Y(new_n3933));
  OAI311xp33_ASAP7_75t_L    g03677(.A1(new_n799), .A2(new_n797), .A3(new_n1771), .B1(new_n3933), .C1(new_n3932), .Y(new_n3934));
  AOI21xp33_ASAP7_75t_L     g03678(.A1(new_n1910), .A2(\b[11] ), .B(new_n3934), .Y(new_n3935));
  NAND2xp33_ASAP7_75t_L     g03679(.A(\a[23] ), .B(new_n3935), .Y(new_n3936));
  A2O1A1Ixp33_ASAP7_75t_L   g03680(.A1(\b[11] ), .A2(new_n1910), .B(new_n3934), .C(new_n1761), .Y(new_n3937));
  NAND2xp33_ASAP7_75t_L     g03681(.A(new_n3937), .B(new_n3936), .Y(new_n3938));
  AO21x2_ASAP7_75t_L        g03682(.A1(new_n3931), .A2(new_n3927), .B(new_n3938), .Y(new_n3939));
  NAND3xp33_ASAP7_75t_L     g03683(.A(new_n3927), .B(new_n3938), .C(new_n3931), .Y(new_n3940));
  AND3x1_ASAP7_75t_L        g03684(.A(new_n3851), .B(new_n3940), .C(new_n3939), .Y(new_n3941));
  AOI21xp33_ASAP7_75t_L     g03685(.A1(new_n3940), .A2(new_n3939), .B(new_n3851), .Y(new_n3942));
  OAI21xp33_ASAP7_75t_L     g03686(.A1(new_n3942), .A2(new_n3941), .B(new_n3850), .Y(new_n3943));
  NOR2xp33_ASAP7_75t_L      g03687(.A(new_n3849), .B(new_n3848), .Y(new_n3944));
  NAND3xp33_ASAP7_75t_L     g03688(.A(new_n3851), .B(new_n3939), .C(new_n3940), .Y(new_n3945));
  A2O1A1Ixp33_ASAP7_75t_L   g03689(.A1(new_n3710), .A2(new_n3520), .B(new_n3707), .C(new_n3715), .Y(new_n3946));
  AOI21xp33_ASAP7_75t_L     g03690(.A1(new_n3927), .A2(new_n3931), .B(new_n3938), .Y(new_n3947));
  INVx1_ASAP7_75t_L         g03691(.A(new_n3940), .Y(new_n3948));
  OAI21xp33_ASAP7_75t_L     g03692(.A1(new_n3947), .A2(new_n3948), .B(new_n3946), .Y(new_n3949));
  NAND3xp33_ASAP7_75t_L     g03693(.A(new_n3949), .B(new_n3945), .C(new_n3944), .Y(new_n3950));
  NAND2xp33_ASAP7_75t_L     g03694(.A(new_n3950), .B(new_n3943), .Y(new_n3951));
  NAND3xp33_ASAP7_75t_L     g03695(.A(new_n3951), .B(new_n3844), .C(new_n3730), .Y(new_n3952));
  NAND2xp33_ASAP7_75t_L     g03696(.A(new_n3727), .B(new_n3726), .Y(new_n3953));
  MAJIxp5_ASAP7_75t_L       g03697(.A(new_n3731), .B(new_n3728), .C(new_n3953), .Y(new_n3954));
  NAND3xp33_ASAP7_75t_L     g03698(.A(new_n3954), .B(new_n3943), .C(new_n3950), .Y(new_n3955));
  NOR2xp33_ASAP7_75t_L      g03699(.A(new_n1244), .B(new_n1195), .Y(new_n3956));
  NOR2xp33_ASAP7_75t_L      g03700(.A(new_n1356), .B(new_n1298), .Y(new_n3957));
  INVx1_ASAP7_75t_L         g03701(.A(new_n3957), .Y(new_n3958));
  OAI221xp5_ASAP7_75t_L     g03702(.A1(new_n1198), .A2(new_n1493), .B1(new_n1197), .B2(new_n2793), .C(new_n3958), .Y(new_n3959));
  NOR3xp33_ASAP7_75t_L      g03703(.A(new_n3959), .B(new_n3956), .C(new_n1107), .Y(new_n3960));
  INVx1_ASAP7_75t_L         g03704(.A(new_n3956), .Y(new_n3961));
  AOI22xp33_ASAP7_75t_L     g03705(.A1(new_n1113), .A2(\b[19] ), .B1(new_n1110), .B2(new_n1499), .Y(new_n3962));
  AOI31xp33_ASAP7_75t_L     g03706(.A1(new_n3962), .A2(new_n3958), .A3(new_n3961), .B(\a[17] ), .Y(new_n3963));
  NOR2xp33_ASAP7_75t_L      g03707(.A(new_n3963), .B(new_n3960), .Y(new_n3964));
  NAND3xp33_ASAP7_75t_L     g03708(.A(new_n3952), .B(new_n3955), .C(new_n3964), .Y(new_n3965));
  AOI21xp33_ASAP7_75t_L     g03709(.A1(new_n3950), .A2(new_n3943), .B(new_n3954), .Y(new_n3966));
  O2A1O1Ixp33_ASAP7_75t_L   g03710(.A1(new_n3953), .A2(new_n3728), .B(new_n3730), .C(new_n3951), .Y(new_n3967));
  NAND4xp25_ASAP7_75t_L     g03711(.A(new_n3962), .B(\a[17] ), .C(new_n3961), .D(new_n3958), .Y(new_n3968));
  A2O1A1Ixp33_ASAP7_75t_L   g03712(.A1(\b[17] ), .A2(new_n1194), .B(new_n3959), .C(new_n1107), .Y(new_n3969));
  NAND2xp33_ASAP7_75t_L     g03713(.A(new_n3968), .B(new_n3969), .Y(new_n3970));
  OAI21xp33_ASAP7_75t_L     g03714(.A1(new_n3966), .A2(new_n3967), .B(new_n3970), .Y(new_n3971));
  NAND2xp33_ASAP7_75t_L     g03715(.A(new_n3965), .B(new_n3971), .Y(new_n3972));
  OAI21xp33_ASAP7_75t_L     g03716(.A1(new_n3737), .A2(new_n3632), .B(new_n3735), .Y(new_n3973));
  NOR2xp33_ASAP7_75t_L      g03717(.A(new_n3972), .B(new_n3973), .Y(new_n3974));
  NOR3xp33_ASAP7_75t_L      g03718(.A(new_n3967), .B(new_n3966), .C(new_n3970), .Y(new_n3975));
  AOI21xp33_ASAP7_75t_L     g03719(.A1(new_n3952), .A2(new_n3955), .B(new_n3964), .Y(new_n3976));
  NOR2xp33_ASAP7_75t_L      g03720(.A(new_n3976), .B(new_n3975), .Y(new_n3977));
  A2O1A1O1Ixp25_ASAP7_75t_L g03721(.A1(new_n3552), .A2(new_n3562), .B(new_n3631), .C(new_n3736), .D(new_n3739), .Y(new_n3978));
  NOR2xp33_ASAP7_75t_L      g03722(.A(new_n3978), .B(new_n3977), .Y(new_n3979));
  NAND2xp33_ASAP7_75t_L     g03723(.A(\b[20] ), .B(new_n908), .Y(new_n3980));
  NAND2xp33_ASAP7_75t_L     g03724(.A(\b[21] ), .B(new_n817), .Y(new_n3981));
  AOI32xp33_ASAP7_75t_L     g03725(.A1(new_n1862), .A2(new_n1860), .A3(new_n823), .B1(new_n826), .B2(\b[22] ), .Y(new_n3982));
  NAND4xp25_ASAP7_75t_L     g03726(.A(new_n3982), .B(\a[14] ), .C(new_n3980), .D(new_n3981), .Y(new_n3983));
  NAND2xp33_ASAP7_75t_L     g03727(.A(new_n3981), .B(new_n3982), .Y(new_n3984));
  A2O1A1Ixp33_ASAP7_75t_L   g03728(.A1(\b[20] ), .A2(new_n908), .B(new_n3984), .C(new_n813), .Y(new_n3985));
  NAND2xp33_ASAP7_75t_L     g03729(.A(new_n3983), .B(new_n3985), .Y(new_n3986));
  NOR3xp33_ASAP7_75t_L      g03730(.A(new_n3974), .B(new_n3979), .C(new_n3986), .Y(new_n3987));
  NAND2xp33_ASAP7_75t_L     g03731(.A(new_n3978), .B(new_n3977), .Y(new_n3988));
  NAND2xp33_ASAP7_75t_L     g03732(.A(new_n3972), .B(new_n3973), .Y(new_n3989));
  AND2x2_ASAP7_75t_L        g03733(.A(new_n3983), .B(new_n3985), .Y(new_n3990));
  AOI21xp33_ASAP7_75t_L     g03734(.A1(new_n3989), .A2(new_n3988), .B(new_n3990), .Y(new_n3991));
  NOR2xp33_ASAP7_75t_L      g03735(.A(new_n3991), .B(new_n3987), .Y(new_n3992));
  NAND2xp33_ASAP7_75t_L     g03736(.A(new_n3738), .B(new_n3742), .Y(new_n3993));
  NOR2xp33_ASAP7_75t_L      g03737(.A(new_n3751), .B(new_n3993), .Y(new_n3994));
  O2A1O1Ixp33_ASAP7_75t_L   g03738(.A1(new_n3566), .A2(new_n3759), .B(new_n3758), .C(new_n3994), .Y(new_n3995));
  NAND2xp33_ASAP7_75t_L     g03739(.A(new_n3992), .B(new_n3995), .Y(new_n3996));
  INVx1_ASAP7_75t_L         g03740(.A(new_n3761), .Y(new_n3997));
  NAND3xp33_ASAP7_75t_L     g03741(.A(new_n3989), .B(new_n3988), .C(new_n3990), .Y(new_n3998));
  OAI21xp33_ASAP7_75t_L     g03742(.A1(new_n3979), .A2(new_n3974), .B(new_n3986), .Y(new_n3999));
  NAND2xp33_ASAP7_75t_L     g03743(.A(new_n3998), .B(new_n3999), .Y(new_n4000));
  A2O1A1Ixp33_ASAP7_75t_L   g03744(.A1(new_n3758), .A2(new_n3997), .B(new_n3994), .C(new_n4000), .Y(new_n4001));
  NAND2xp33_ASAP7_75t_L     g03745(.A(\b[24] ), .B(new_n590), .Y(new_n4002));
  OAI221xp5_ASAP7_75t_L     g03746(.A1(new_n676), .A2(new_n2180), .B1(new_n675), .B2(new_n2187), .C(new_n4002), .Y(new_n4003));
  AOI21xp33_ASAP7_75t_L     g03747(.A1(new_n674), .A2(\b[23] ), .B(new_n4003), .Y(new_n4004));
  NAND2xp33_ASAP7_75t_L     g03748(.A(\a[11] ), .B(new_n4004), .Y(new_n4005));
  A2O1A1Ixp33_ASAP7_75t_L   g03749(.A1(\b[23] ), .A2(new_n674), .B(new_n4003), .C(new_n594), .Y(new_n4006));
  NAND2xp33_ASAP7_75t_L     g03750(.A(new_n4006), .B(new_n4005), .Y(new_n4007));
  NAND3xp33_ASAP7_75t_L     g03751(.A(new_n3996), .B(new_n4001), .C(new_n4007), .Y(new_n4008));
  MAJIxp5_ASAP7_75t_L       g03752(.A(new_n3761), .B(new_n3993), .C(new_n3751), .Y(new_n4009));
  NOR2xp33_ASAP7_75t_L      g03753(.A(new_n4009), .B(new_n4000), .Y(new_n4010));
  O2A1O1Ixp33_ASAP7_75t_L   g03754(.A1(new_n3993), .A2(new_n3751), .B(new_n3760), .C(new_n3992), .Y(new_n4011));
  AND2x2_ASAP7_75t_L        g03755(.A(new_n4006), .B(new_n4005), .Y(new_n4012));
  OAI21xp33_ASAP7_75t_L     g03756(.A1(new_n4010), .A2(new_n4011), .B(new_n4012), .Y(new_n4013));
  NAND2xp33_ASAP7_75t_L     g03757(.A(new_n4008), .B(new_n4013), .Y(new_n4014));
  XNOR2x2_ASAP7_75t_L       g03758(.A(new_n3843), .B(new_n4014), .Y(new_n4015));
  NAND2xp33_ASAP7_75t_L     g03759(.A(new_n3842), .B(new_n4015), .Y(new_n4016));
  NAND3xp33_ASAP7_75t_L     g03760(.A(new_n4014), .B(new_n3771), .C(new_n3774), .Y(new_n4017));
  NOR3xp33_ASAP7_75t_L      g03761(.A(new_n4011), .B(new_n4012), .C(new_n4010), .Y(new_n4018));
  AOI21xp33_ASAP7_75t_L     g03762(.A1(new_n3996), .A2(new_n4001), .B(new_n4007), .Y(new_n4019));
  NOR2xp33_ASAP7_75t_L      g03763(.A(new_n4019), .B(new_n4018), .Y(new_n4020));
  A2O1A1Ixp33_ASAP7_75t_L   g03764(.A1(new_n3773), .A2(new_n3621), .B(new_n3769), .C(new_n4020), .Y(new_n4021));
  AO21x2_ASAP7_75t_L        g03765(.A1(new_n4017), .A2(new_n4021), .B(new_n3842), .Y(new_n4022));
  NAND2xp33_ASAP7_75t_L     g03766(.A(new_n3776), .B(new_n3771), .Y(new_n4023));
  MAJIxp5_ASAP7_75t_L       g03767(.A(new_n3785), .B(new_n4023), .C(new_n3782), .Y(new_n4024));
  INVx1_ASAP7_75t_L         g03768(.A(new_n4024), .Y(new_n4025));
  NAND3xp33_ASAP7_75t_L     g03769(.A(new_n4025), .B(new_n4022), .C(new_n4016), .Y(new_n4026));
  AND3x1_ASAP7_75t_L        g03770(.A(new_n4021), .B(new_n4017), .C(new_n3842), .Y(new_n4027));
  NOR2xp33_ASAP7_75t_L      g03771(.A(new_n3842), .B(new_n4015), .Y(new_n4028));
  OAI21xp33_ASAP7_75t_L     g03772(.A1(new_n4027), .A2(new_n4028), .B(new_n4024), .Y(new_n4029));
  NAND2xp33_ASAP7_75t_L     g03773(.A(new_n3422), .B(new_n3425), .Y(new_n4030));
  NAND2xp33_ASAP7_75t_L     g03774(.A(\b[31] ), .B(new_n345), .Y(new_n4031));
  OAI221xp5_ASAP7_75t_L     g03775(.A1(new_n3212), .A2(new_n406), .B1(new_n367), .B2(new_n4030), .C(new_n4031), .Y(new_n4032));
  AOI21xp33_ASAP7_75t_L     g03776(.A1(new_n366), .A2(\b[29] ), .B(new_n4032), .Y(new_n4033));
  NAND2xp33_ASAP7_75t_L     g03777(.A(\a[5] ), .B(new_n4033), .Y(new_n4034));
  A2O1A1Ixp33_ASAP7_75t_L   g03778(.A1(\b[29] ), .A2(new_n366), .B(new_n4032), .C(new_n339), .Y(new_n4035));
  NAND2xp33_ASAP7_75t_L     g03779(.A(new_n4035), .B(new_n4034), .Y(new_n4036));
  AO21x2_ASAP7_75t_L        g03780(.A1(new_n4029), .A2(new_n4026), .B(new_n4036), .Y(new_n4037));
  NAND3xp33_ASAP7_75t_L     g03781(.A(new_n4026), .B(new_n4036), .C(new_n4029), .Y(new_n4038));
  NAND3xp33_ASAP7_75t_L     g03782(.A(new_n3839), .B(new_n4037), .C(new_n4038), .Y(new_n4039));
  NAND2xp33_ASAP7_75t_L     g03783(.A(new_n4038), .B(new_n4037), .Y(new_n4040));
  A2O1A1Ixp33_ASAP7_75t_L   g03784(.A1(new_n3802), .A2(new_n3799), .B(new_n3838), .C(new_n4040), .Y(new_n4041));
  AOI21xp33_ASAP7_75t_L     g03785(.A1(new_n4041), .A2(new_n4039), .B(new_n3836), .Y(new_n4042));
  INVx1_ASAP7_75t_L         g03786(.A(new_n4042), .Y(new_n4043));
  NAND3xp33_ASAP7_75t_L     g03787(.A(new_n4041), .B(new_n4039), .C(new_n3836), .Y(new_n4044));
  NAND2xp33_ASAP7_75t_L     g03788(.A(new_n4044), .B(new_n4043), .Y(new_n4045));
  O2A1O1Ixp33_ASAP7_75t_L   g03789(.A1(new_n3619), .A2(new_n3819), .B(new_n3817), .C(new_n4045), .Y(new_n4046));
  OAI21xp33_ASAP7_75t_L     g03790(.A1(new_n3819), .A2(new_n3619), .B(new_n3817), .Y(new_n4047));
  AOI21xp33_ASAP7_75t_L     g03791(.A1(new_n4043), .A2(new_n4044), .B(new_n4047), .Y(new_n4048));
  NOR2xp33_ASAP7_75t_L      g03792(.A(new_n4048), .B(new_n4046), .Y(\f[34] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03793(.A1(new_n3615), .A2(new_n3439), .B(new_n3613), .C(new_n3822), .Y(new_n4050));
  NOR2xp33_ASAP7_75t_L      g03794(.A(new_n3807), .B(new_n277), .Y(new_n4051));
  NOR2xp33_ASAP7_75t_L      g03795(.A(\b[34] ), .B(\b[35] ), .Y(new_n4052));
  INVx1_ASAP7_75t_L         g03796(.A(\b[35] ), .Y(new_n4053));
  NOR2xp33_ASAP7_75t_L      g03797(.A(new_n3827), .B(new_n4053), .Y(new_n4054));
  NOR2xp33_ASAP7_75t_L      g03798(.A(new_n4052), .B(new_n4054), .Y(new_n4055));
  A2O1A1Ixp33_ASAP7_75t_L   g03799(.A1(\b[34] ), .A2(\b[33] ), .B(new_n3831), .C(new_n4055), .Y(new_n4056));
  O2A1O1Ixp33_ASAP7_75t_L   g03800(.A1(new_n3808), .A2(new_n3811), .B(new_n3829), .C(new_n3828), .Y(new_n4057));
  INVx1_ASAP7_75t_L         g03801(.A(new_n4055), .Y(new_n4058));
  NAND2xp33_ASAP7_75t_L     g03802(.A(new_n4058), .B(new_n4057), .Y(new_n4059));
  NAND2xp33_ASAP7_75t_L     g03803(.A(new_n4059), .B(new_n4056), .Y(new_n4060));
  NAND2xp33_ASAP7_75t_L     g03804(.A(\b[35] ), .B(new_n272), .Y(new_n4061));
  OAI221xp5_ASAP7_75t_L     g03805(.A1(new_n3827), .A2(new_n261), .B1(new_n292), .B2(new_n4060), .C(new_n4061), .Y(new_n4062));
  OR3x1_ASAP7_75t_L         g03806(.A(new_n4062), .B(new_n265), .C(new_n4051), .Y(new_n4063));
  A2O1A1Ixp33_ASAP7_75t_L   g03807(.A1(\b[33] ), .A2(new_n291), .B(new_n4062), .C(new_n265), .Y(new_n4064));
  AND2x2_ASAP7_75t_L        g03808(.A(new_n4064), .B(new_n4063), .Y(new_n4065));
  AOI32xp33_ASAP7_75t_L     g03809(.A1(new_n2483), .A2(new_n2486), .A3(new_n597), .B1(new_n600), .B2(\b[26] ), .Y(new_n4066));
  OAI221xp5_ASAP7_75t_L     g03810(.A1(new_n721), .A2(new_n2180), .B1(new_n2019), .B2(new_n1620), .C(new_n4066), .Y(new_n4067));
  XNOR2x2_ASAP7_75t_L       g03811(.A(\a[11] ), .B(new_n4067), .Y(new_n4068));
  INVx1_ASAP7_75t_L         g03812(.A(new_n4068), .Y(new_n4069));
  NOR3xp33_ASAP7_75t_L      g03813(.A(new_n3974), .B(new_n3979), .C(new_n3990), .Y(new_n4070));
  NOR2xp33_ASAP7_75t_L      g03814(.A(new_n1709), .B(new_n909), .Y(new_n4071));
  INVx1_ASAP7_75t_L         g03815(.A(new_n4071), .Y(new_n4072));
  NAND2xp33_ASAP7_75t_L     g03816(.A(\b[22] ), .B(new_n817), .Y(new_n4073));
  AOI22xp33_ASAP7_75t_L     g03817(.A1(new_n826), .A2(\b[23] ), .B1(new_n823), .B2(new_n2002), .Y(new_n4074));
  AND4x1_ASAP7_75t_L        g03818(.A(new_n4074), .B(new_n4073), .C(new_n4072), .D(\a[14] ), .Y(new_n4075));
  AOI31xp33_ASAP7_75t_L     g03819(.A1(new_n4074), .A2(new_n4073), .A3(new_n4072), .B(\a[14] ), .Y(new_n4076));
  OR2x4_ASAP7_75t_L         g03820(.A(new_n4076), .B(new_n4075), .Y(new_n4077));
  NOR3xp33_ASAP7_75t_L      g03821(.A(new_n3967), .B(new_n3966), .C(new_n3964), .Y(new_n4078));
  INVx1_ASAP7_75t_L         g03822(.A(new_n4078), .Y(new_n4079));
  A2O1A1Ixp33_ASAP7_75t_L   g03823(.A1(new_n3971), .A2(new_n3965), .B(new_n3978), .C(new_n4079), .Y(new_n4080));
  NAND2xp33_ASAP7_75t_L     g03824(.A(\b[12] ), .B(new_n1910), .Y(new_n4081));
  NAND2xp33_ASAP7_75t_L     g03825(.A(\b[13] ), .B(new_n1770), .Y(new_n4082));
  AOI32xp33_ASAP7_75t_L     g03826(.A1(new_n877), .A2(new_n874), .A3(new_n1764), .B1(\b[14] ), .B2(new_n1766), .Y(new_n4083));
  AND4x1_ASAP7_75t_L        g03827(.A(new_n4083), .B(new_n4082), .C(new_n4081), .D(\a[23] ), .Y(new_n4084));
  AOI31xp33_ASAP7_75t_L     g03828(.A1(new_n4083), .A2(new_n4082), .A3(new_n4081), .B(\a[23] ), .Y(new_n4085));
  NOR2xp33_ASAP7_75t_L      g03829(.A(new_n4085), .B(new_n4084), .Y(new_n4086));
  NOR2xp33_ASAP7_75t_L      g03830(.A(new_n3922), .B(new_n3923), .Y(new_n4087));
  MAJIxp5_ASAP7_75t_L       g03831(.A(new_n3930), .B(new_n3924), .C(new_n4087), .Y(new_n4088));
  NAND2xp33_ASAP7_75t_L     g03832(.A(\b[9] ), .B(new_n2386), .Y(new_n4089));
  NAND2xp33_ASAP7_75t_L     g03833(.A(\b[10] ), .B(new_n2232), .Y(new_n4090));
  AOI32xp33_ASAP7_75t_L     g03834(.A1(new_n700), .A2(new_n698), .A3(new_n2226), .B1(\b[11] ), .B2(new_n2228), .Y(new_n4091));
  NAND4xp25_ASAP7_75t_L     g03835(.A(new_n4091), .B(\a[26] ), .C(new_n4089), .D(new_n4090), .Y(new_n4092));
  AOI31xp33_ASAP7_75t_L     g03836(.A1(new_n4091), .A2(new_n4090), .A3(new_n4089), .B(\a[26] ), .Y(new_n4093));
  INVx1_ASAP7_75t_L         g03837(.A(new_n4093), .Y(new_n4094));
  NAND2xp33_ASAP7_75t_L     g03838(.A(new_n4092), .B(new_n4094), .Y(new_n4095));
  A2O1A1O1Ixp25_ASAP7_75t_L g03839(.A1(new_n3675), .A2(new_n3680), .B(new_n3852), .C(new_n3899), .D(new_n3911), .Y(new_n4096));
  NOR2xp33_ASAP7_75t_L      g03840(.A(new_n382), .B(new_n2932), .Y(new_n4097));
  NAND2xp33_ASAP7_75t_L     g03841(.A(\b[7] ), .B(new_n2706), .Y(new_n4098));
  OAI221xp5_ASAP7_75t_L     g03842(.A1(new_n2708), .A2(new_n503), .B1(new_n2707), .B2(new_n509), .C(new_n4098), .Y(new_n4099));
  NOR3xp33_ASAP7_75t_L      g03843(.A(new_n4099), .B(new_n4097), .C(new_n2697), .Y(new_n4100));
  INVx1_ASAP7_75t_L         g03844(.A(new_n4100), .Y(new_n4101));
  A2O1A1Ixp33_ASAP7_75t_L   g03845(.A1(\b[6] ), .A2(new_n2931), .B(new_n4099), .C(new_n2697), .Y(new_n4102));
  O2A1O1Ixp33_ASAP7_75t_L   g03846(.A1(new_n3892), .A2(new_n3670), .B(new_n3896), .C(new_n3889), .Y(new_n4103));
  NAND2xp33_ASAP7_75t_L     g03847(.A(\b[4] ), .B(new_n3260), .Y(new_n4104));
  OAI221xp5_ASAP7_75t_L     g03848(.A1(new_n3262), .A2(new_n353), .B1(new_n3261), .B2(new_n359), .C(new_n4104), .Y(new_n4105));
  AOI211xp5_ASAP7_75t_L     g03849(.A1(\b[3] ), .A2(new_n3491), .B(new_n3251), .C(new_n4105), .Y(new_n4106));
  INVx1_ASAP7_75t_L         g03850(.A(new_n4106), .Y(new_n4107));
  A2O1A1Ixp33_ASAP7_75t_L   g03851(.A1(\b[3] ), .A2(new_n3491), .B(new_n4105), .C(new_n3251), .Y(new_n4108));
  A2O1A1Ixp33_ASAP7_75t_L   g03852(.A1(\b[0] ), .A2(new_n3872), .B(new_n3886), .C(\a[35] ), .Y(new_n4109));
  INVx1_ASAP7_75t_L         g03853(.A(new_n3873), .Y(new_n4110));
  NOR3xp33_ASAP7_75t_L      g03854(.A(new_n3880), .B(new_n4110), .C(new_n3872), .Y(new_n4111));
  NAND2xp33_ASAP7_75t_L     g03855(.A(\b[0] ), .B(new_n4111), .Y(new_n4112));
  INVx1_ASAP7_75t_L         g03856(.A(new_n4112), .Y(new_n4113));
  NAND2xp33_ASAP7_75t_L     g03857(.A(new_n3883), .B(new_n3872), .Y(new_n4114));
  INVx1_ASAP7_75t_L         g03858(.A(new_n3884), .Y(new_n4115));
  NAND2xp33_ASAP7_75t_L     g03859(.A(\b[1] ), .B(new_n3874), .Y(new_n4116));
  OAI221xp5_ASAP7_75t_L     g03860(.A1(new_n4114), .A2(new_n283), .B1(new_n278), .B2(new_n4115), .C(new_n4116), .Y(new_n4117));
  NOR2xp33_ASAP7_75t_L      g03861(.A(new_n4113), .B(new_n4117), .Y(new_n4118));
  XNOR2x2_ASAP7_75t_L       g03862(.A(new_n4118), .B(new_n4109), .Y(new_n4119));
  NAND3xp33_ASAP7_75t_L     g03863(.A(new_n4119), .B(new_n4108), .C(new_n4107), .Y(new_n4120));
  INVx1_ASAP7_75t_L         g03864(.A(new_n4108), .Y(new_n4121));
  INVx1_ASAP7_75t_L         g03865(.A(new_n3651), .Y(new_n4122));
  A2O1A1Ixp33_ASAP7_75t_L   g03866(.A1(new_n4122), .A2(new_n3894), .B(new_n3878), .C(new_n4118), .Y(new_n4123));
  O2A1O1Ixp33_ASAP7_75t_L   g03867(.A1(new_n258), .A2(new_n3650), .B(new_n3894), .C(new_n3878), .Y(new_n4124));
  A2O1A1Ixp33_ASAP7_75t_L   g03868(.A1(\b[0] ), .A2(new_n4111), .B(new_n4117), .C(new_n4124), .Y(new_n4125));
  OAI211xp5_ASAP7_75t_L     g03869(.A1(new_n4106), .A2(new_n4121), .B(new_n4123), .C(new_n4125), .Y(new_n4126));
  NAND3xp33_ASAP7_75t_L     g03870(.A(new_n4103), .B(new_n4126), .C(new_n4120), .Y(new_n4127));
  A2O1A1Ixp33_ASAP7_75t_L   g03871(.A1(new_n3660), .A2(new_n3891), .B(new_n3888), .C(new_n3897), .Y(new_n4128));
  AOI211xp5_ASAP7_75t_L     g03872(.A1(new_n4125), .A2(new_n4123), .B(new_n4106), .C(new_n4121), .Y(new_n4129));
  AOI21xp33_ASAP7_75t_L     g03873(.A1(new_n4108), .A2(new_n4107), .B(new_n4119), .Y(new_n4130));
  OAI21xp33_ASAP7_75t_L     g03874(.A1(new_n4129), .A2(new_n4130), .B(new_n4128), .Y(new_n4131));
  AOI22xp33_ASAP7_75t_L     g03875(.A1(new_n4127), .A2(new_n4131), .B1(new_n4102), .B2(new_n4101), .Y(new_n4132));
  OA21x2_ASAP7_75t_L        g03876(.A1(new_n4097), .A2(new_n4099), .B(new_n2697), .Y(new_n4133));
  NOR3xp33_ASAP7_75t_L      g03877(.A(new_n4128), .B(new_n4129), .C(new_n4130), .Y(new_n4134));
  AOI21xp33_ASAP7_75t_L     g03878(.A1(new_n4126), .A2(new_n4120), .B(new_n4103), .Y(new_n4135));
  NOR4xp25_ASAP7_75t_L      g03879(.A(new_n4134), .B(new_n4100), .C(new_n4135), .D(new_n4133), .Y(new_n4136));
  NOR3xp33_ASAP7_75t_L      g03880(.A(new_n4096), .B(new_n4136), .C(new_n4132), .Y(new_n4137));
  A2O1A1Ixp33_ASAP7_75t_L   g03881(.A1(new_n3921), .A2(new_n3853), .B(new_n3910), .C(new_n3906), .Y(new_n4138));
  OAI22xp33_ASAP7_75t_L     g03882(.A1(new_n4134), .A2(new_n4135), .B1(new_n4100), .B2(new_n4133), .Y(new_n4139));
  NAND4xp25_ASAP7_75t_L     g03883(.A(new_n4101), .B(new_n4131), .C(new_n4127), .D(new_n4102), .Y(new_n4140));
  AOI21xp33_ASAP7_75t_L     g03884(.A1(new_n4140), .A2(new_n4139), .B(new_n4138), .Y(new_n4141));
  OAI21xp33_ASAP7_75t_L     g03885(.A1(new_n4137), .A2(new_n4141), .B(new_n4095), .Y(new_n4142));
  NAND3xp33_ASAP7_75t_L     g03886(.A(new_n4138), .B(new_n4139), .C(new_n4140), .Y(new_n4143));
  OAI21xp33_ASAP7_75t_L     g03887(.A1(new_n4132), .A2(new_n4136), .B(new_n4096), .Y(new_n4144));
  NAND4xp25_ASAP7_75t_L     g03888(.A(new_n4143), .B(new_n4092), .C(new_n4094), .D(new_n4144), .Y(new_n4145));
  AOI21xp33_ASAP7_75t_L     g03889(.A1(new_n4145), .A2(new_n4142), .B(new_n4088), .Y(new_n4146));
  NAND2xp33_ASAP7_75t_L     g03890(.A(new_n3907), .B(new_n3912), .Y(new_n4147));
  MAJIxp5_ASAP7_75t_L       g03891(.A(new_n3926), .B(new_n3919), .C(new_n4147), .Y(new_n4148));
  NAND2xp33_ASAP7_75t_L     g03892(.A(new_n4142), .B(new_n4145), .Y(new_n4149));
  NOR2xp33_ASAP7_75t_L      g03893(.A(new_n4148), .B(new_n4149), .Y(new_n4150));
  OAI21xp33_ASAP7_75t_L     g03894(.A1(new_n4146), .A2(new_n4150), .B(new_n4086), .Y(new_n4151));
  INVx1_ASAP7_75t_L         g03895(.A(new_n4086), .Y(new_n4152));
  NAND2xp33_ASAP7_75t_L     g03896(.A(new_n4148), .B(new_n4149), .Y(new_n4153));
  NAND3xp33_ASAP7_75t_L     g03897(.A(new_n4088), .B(new_n4142), .C(new_n4145), .Y(new_n4154));
  NAND3xp33_ASAP7_75t_L     g03898(.A(new_n4153), .B(new_n4154), .C(new_n4152), .Y(new_n4155));
  A2O1A1O1Ixp25_ASAP7_75t_L g03899(.A1(new_n3520), .A2(new_n3710), .B(new_n3707), .C(new_n3715), .D(new_n3947), .Y(new_n4156));
  OAI211xp5_ASAP7_75t_L     g03900(.A1(new_n3948), .A2(new_n4156), .B(new_n4151), .C(new_n4155), .Y(new_n4157));
  AOI21xp33_ASAP7_75t_L     g03901(.A1(new_n4153), .A2(new_n4154), .B(new_n4152), .Y(new_n4158));
  NOR3xp33_ASAP7_75t_L      g03902(.A(new_n4150), .B(new_n4146), .C(new_n4086), .Y(new_n4159));
  A2O1A1Ixp33_ASAP7_75t_L   g03903(.A1(new_n3716), .A2(new_n3712), .B(new_n3708), .C(new_n3939), .Y(new_n4160));
  OAI211xp5_ASAP7_75t_L     g03904(.A1(new_n4158), .A2(new_n4159), .B(new_n3940), .C(new_n4160), .Y(new_n4161));
  NOR2xp33_ASAP7_75t_L      g03905(.A(new_n952), .B(new_n1549), .Y(new_n4162));
  INVx1_ASAP7_75t_L         g03906(.A(new_n4162), .Y(new_n4163));
  NOR2xp33_ASAP7_75t_L      g03907(.A(new_n1051), .B(new_n1398), .Y(new_n4164));
  INVx1_ASAP7_75t_L         g03908(.A(new_n4164), .Y(new_n4165));
  AOI32xp33_ASAP7_75t_L     g03909(.A1(new_n1250), .A2(new_n1247), .A3(new_n1404), .B1(\b[17] ), .B2(new_n1406), .Y(new_n4166));
  AND4x1_ASAP7_75t_L        g03910(.A(new_n4166), .B(new_n4165), .C(new_n4163), .D(\a[20] ), .Y(new_n4167));
  AOI31xp33_ASAP7_75t_L     g03911(.A1(new_n4166), .A2(new_n4165), .A3(new_n4163), .B(\a[20] ), .Y(new_n4168));
  NOR2xp33_ASAP7_75t_L      g03912(.A(new_n4168), .B(new_n4167), .Y(new_n4169));
  NAND3xp33_ASAP7_75t_L     g03913(.A(new_n4161), .B(new_n4157), .C(new_n4169), .Y(new_n4170));
  AO21x2_ASAP7_75t_L        g03914(.A1(new_n4157), .A2(new_n4161), .B(new_n4169), .Y(new_n4171));
  NAND2xp33_ASAP7_75t_L     g03915(.A(new_n4170), .B(new_n4171), .Y(new_n4172));
  INVx1_ASAP7_75t_L         g03916(.A(new_n3950), .Y(new_n4173));
  A2O1A1Ixp33_ASAP7_75t_L   g03917(.A1(new_n3730), .A2(new_n3844), .B(new_n4173), .C(new_n3943), .Y(new_n4174));
  NOR2xp33_ASAP7_75t_L      g03918(.A(new_n4172), .B(new_n4174), .Y(new_n4175));
  AOI21xp33_ASAP7_75t_L     g03919(.A1(new_n3949), .A2(new_n3945), .B(new_n3944), .Y(new_n4176));
  AOI21xp33_ASAP7_75t_L     g03920(.A1(new_n3954), .A2(new_n3950), .B(new_n4176), .Y(new_n4177));
  AOI21xp33_ASAP7_75t_L     g03921(.A1(new_n4171), .A2(new_n4170), .B(new_n4177), .Y(new_n4178));
  NOR2xp33_ASAP7_75t_L      g03922(.A(new_n1356), .B(new_n1195), .Y(new_n4179));
  NAND2xp33_ASAP7_75t_L     g03923(.A(\b[19] ), .B(new_n1103), .Y(new_n4180));
  NAND2xp33_ASAP7_75t_L     g03924(.A(\b[20] ), .B(new_n1113), .Y(new_n4181));
  OAI311xp33_ASAP7_75t_L    g03925(.A1(new_n1599), .A2(new_n1598), .A3(new_n1197), .B1(new_n4181), .C1(new_n4180), .Y(new_n4182));
  OR3x1_ASAP7_75t_L         g03926(.A(new_n4182), .B(new_n1107), .C(new_n4179), .Y(new_n4183));
  A2O1A1Ixp33_ASAP7_75t_L   g03927(.A1(\b[18] ), .A2(new_n1194), .B(new_n4182), .C(new_n1107), .Y(new_n4184));
  AND2x2_ASAP7_75t_L        g03928(.A(new_n4184), .B(new_n4183), .Y(new_n4185));
  OAI21xp33_ASAP7_75t_L     g03929(.A1(new_n4175), .A2(new_n4178), .B(new_n4185), .Y(new_n4186));
  NAND3xp33_ASAP7_75t_L     g03930(.A(new_n4177), .B(new_n4171), .C(new_n4170), .Y(new_n4187));
  A2O1A1Ixp33_ASAP7_75t_L   g03931(.A1(new_n3950), .A2(new_n3954), .B(new_n4176), .C(new_n4172), .Y(new_n4188));
  NAND2xp33_ASAP7_75t_L     g03932(.A(new_n4184), .B(new_n4183), .Y(new_n4189));
  NAND3xp33_ASAP7_75t_L     g03933(.A(new_n4187), .B(new_n4188), .C(new_n4189), .Y(new_n4190));
  NAND2xp33_ASAP7_75t_L     g03934(.A(new_n4190), .B(new_n4186), .Y(new_n4191));
  NOR2xp33_ASAP7_75t_L      g03935(.A(new_n4191), .B(new_n4080), .Y(new_n4192));
  AOI21xp33_ASAP7_75t_L     g03936(.A1(new_n4187), .A2(new_n4188), .B(new_n4189), .Y(new_n4193));
  NOR3xp33_ASAP7_75t_L      g03937(.A(new_n4178), .B(new_n4175), .C(new_n4185), .Y(new_n4194));
  NOR2xp33_ASAP7_75t_L      g03938(.A(new_n4193), .B(new_n4194), .Y(new_n4195));
  O2A1O1Ixp33_ASAP7_75t_L   g03939(.A1(new_n3977), .A2(new_n3978), .B(new_n4079), .C(new_n4195), .Y(new_n4196));
  NOR3xp33_ASAP7_75t_L      g03940(.A(new_n4077), .B(new_n4196), .C(new_n4192), .Y(new_n4197));
  NOR2xp33_ASAP7_75t_L      g03941(.A(new_n4076), .B(new_n4075), .Y(new_n4198));
  O2A1O1Ixp33_ASAP7_75t_L   g03942(.A1(new_n3975), .A2(new_n3976), .B(new_n3973), .C(new_n4078), .Y(new_n4199));
  NAND2xp33_ASAP7_75t_L     g03943(.A(new_n4195), .B(new_n4199), .Y(new_n4200));
  A2O1A1Ixp33_ASAP7_75t_L   g03944(.A1(new_n3973), .A2(new_n3972), .B(new_n4078), .C(new_n4191), .Y(new_n4201));
  AOI21xp33_ASAP7_75t_L     g03945(.A1(new_n4200), .A2(new_n4201), .B(new_n4198), .Y(new_n4202));
  NOR2xp33_ASAP7_75t_L      g03946(.A(new_n4202), .B(new_n4197), .Y(new_n4203));
  A2O1A1Ixp33_ASAP7_75t_L   g03947(.A1(new_n4009), .A2(new_n4000), .B(new_n4070), .C(new_n4203), .Y(new_n4204));
  NAND3xp33_ASAP7_75t_L     g03948(.A(new_n4200), .B(new_n4198), .C(new_n4201), .Y(new_n4205));
  OAI21xp33_ASAP7_75t_L     g03949(.A1(new_n4192), .A2(new_n4196), .B(new_n4077), .Y(new_n4206));
  AOI221xp5_ASAP7_75t_L     g03950(.A1(new_n4000), .A2(new_n4009), .B1(new_n4205), .B2(new_n4206), .C(new_n4070), .Y(new_n4207));
  INVx1_ASAP7_75t_L         g03951(.A(new_n4207), .Y(new_n4208));
  AOI21xp33_ASAP7_75t_L     g03952(.A1(new_n4204), .A2(new_n4208), .B(new_n4069), .Y(new_n4209));
  NOR2xp33_ASAP7_75t_L      g03953(.A(new_n3979), .B(new_n3974), .Y(new_n4210));
  MAJIxp5_ASAP7_75t_L       g03954(.A(new_n4009), .B(new_n4210), .C(new_n3986), .Y(new_n4211));
  NAND2xp33_ASAP7_75t_L     g03955(.A(new_n4205), .B(new_n4206), .Y(new_n4212));
  NOR2xp33_ASAP7_75t_L      g03956(.A(new_n4211), .B(new_n4212), .Y(new_n4213));
  NOR3xp33_ASAP7_75t_L      g03957(.A(new_n4213), .B(new_n4207), .C(new_n4068), .Y(new_n4214));
  A2O1A1O1Ixp25_ASAP7_75t_L g03958(.A1(new_n3621), .A2(new_n3770), .B(new_n3769), .C(new_n4013), .D(new_n4018), .Y(new_n4215));
  NOR3xp33_ASAP7_75t_L      g03959(.A(new_n4215), .B(new_n4209), .C(new_n4214), .Y(new_n4216));
  OAI21xp33_ASAP7_75t_L     g03960(.A1(new_n4207), .A2(new_n4213), .B(new_n4068), .Y(new_n4217));
  NAND3xp33_ASAP7_75t_L     g03961(.A(new_n4204), .B(new_n4208), .C(new_n4069), .Y(new_n4218));
  AOI221xp5_ASAP7_75t_L     g03962(.A1(new_n4020), .A2(new_n3843), .B1(new_n4217), .B2(new_n4218), .C(new_n4018), .Y(new_n4219));
  NAND2xp33_ASAP7_75t_L     g03963(.A(\b[29] ), .B(new_n451), .Y(new_n4220));
  OAI221xp5_ASAP7_75t_L     g03964(.A1(new_n2852), .A2(new_n529), .B1(new_n482), .B2(new_n2881), .C(new_n4220), .Y(new_n4221));
  AOI21xp33_ASAP7_75t_L     g03965(.A1(new_n480), .A2(\b[27] ), .B(new_n4221), .Y(new_n4222));
  NAND2xp33_ASAP7_75t_L     g03966(.A(\a[8] ), .B(new_n4222), .Y(new_n4223));
  A2O1A1Ixp33_ASAP7_75t_L   g03967(.A1(\b[27] ), .A2(new_n480), .B(new_n4221), .C(new_n445), .Y(new_n4224));
  NAND2xp33_ASAP7_75t_L     g03968(.A(new_n4224), .B(new_n4223), .Y(new_n4225));
  OR3x1_ASAP7_75t_L         g03969(.A(new_n4219), .B(new_n4216), .C(new_n4225), .Y(new_n4226));
  OAI21xp33_ASAP7_75t_L     g03970(.A1(new_n4216), .A2(new_n4219), .B(new_n4225), .Y(new_n4227));
  INVx1_ASAP7_75t_L         g03971(.A(new_n3842), .Y(new_n4228));
  MAJIxp5_ASAP7_75t_L       g03972(.A(new_n4024), .B(new_n4228), .C(new_n4015), .Y(new_n4229));
  NAND3xp33_ASAP7_75t_L     g03973(.A(new_n4229), .B(new_n4227), .C(new_n4226), .Y(new_n4230));
  AOI21xp33_ASAP7_75t_L     g03974(.A1(new_n4227), .A2(new_n4226), .B(new_n4229), .Y(new_n4231));
  INVx1_ASAP7_75t_L         g03975(.A(new_n4231), .Y(new_n4232));
  NAND2xp33_ASAP7_75t_L     g03976(.A(new_n342), .B(new_n3450), .Y(new_n4233));
  OAI221xp5_ASAP7_75t_L     g03977(.A1(new_n368), .A2(new_n3443), .B1(new_n3419), .B2(new_n406), .C(new_n4233), .Y(new_n4234));
  AOI21xp33_ASAP7_75t_L     g03978(.A1(new_n366), .A2(\b[30] ), .B(new_n4234), .Y(new_n4235));
  NAND2xp33_ASAP7_75t_L     g03979(.A(\a[5] ), .B(new_n4235), .Y(new_n4236));
  A2O1A1Ixp33_ASAP7_75t_L   g03980(.A1(\b[30] ), .A2(new_n366), .B(new_n4234), .C(new_n339), .Y(new_n4237));
  NAND2xp33_ASAP7_75t_L     g03981(.A(new_n4237), .B(new_n4236), .Y(new_n4238));
  AOI21xp33_ASAP7_75t_L     g03982(.A1(new_n4232), .A2(new_n4230), .B(new_n4238), .Y(new_n4239));
  INVx1_ASAP7_75t_L         g03983(.A(new_n4230), .Y(new_n4240));
  INVx1_ASAP7_75t_L         g03984(.A(new_n4238), .Y(new_n4241));
  NOR3xp33_ASAP7_75t_L      g03985(.A(new_n4241), .B(new_n4240), .C(new_n4231), .Y(new_n4242));
  A2O1A1Ixp33_ASAP7_75t_L   g03986(.A1(new_n3802), .A2(new_n3799), .B(new_n3838), .C(new_n4037), .Y(new_n4243));
  AOI211xp5_ASAP7_75t_L     g03987(.A1(new_n4243), .A2(new_n4038), .B(new_n4239), .C(new_n4242), .Y(new_n4244));
  OAI21xp33_ASAP7_75t_L     g03988(.A1(new_n4231), .A2(new_n4240), .B(new_n4241), .Y(new_n4245));
  NAND3xp33_ASAP7_75t_L     g03989(.A(new_n4232), .B(new_n4238), .C(new_n4230), .Y(new_n4246));
  INVx1_ASAP7_75t_L         g03990(.A(new_n3838), .Y(new_n4247));
  NOR3xp33_ASAP7_75t_L      g03991(.A(new_n3796), .B(new_n3787), .C(new_n3797), .Y(new_n4248));
  AOI21xp33_ASAP7_75t_L     g03992(.A1(new_n3788), .A2(new_n3786), .B(new_n3794), .Y(new_n4249));
  OAI22xp33_ASAP7_75t_L     g03993(.A1(new_n3837), .A2(new_n3611), .B1(new_n4248), .B2(new_n4249), .Y(new_n4250));
  AOI21xp33_ASAP7_75t_L     g03994(.A1(new_n4026), .A2(new_n4029), .B(new_n4036), .Y(new_n4251));
  A2O1A1Ixp33_ASAP7_75t_L   g03995(.A1(new_n4250), .A2(new_n4247), .B(new_n4251), .C(new_n4038), .Y(new_n4252));
  AOI21xp33_ASAP7_75t_L     g03996(.A1(new_n4246), .A2(new_n4245), .B(new_n4252), .Y(new_n4253));
  NOR3xp33_ASAP7_75t_L      g03997(.A(new_n4244), .B(new_n4253), .C(new_n4065), .Y(new_n4254));
  INVx1_ASAP7_75t_L         g03998(.A(new_n4254), .Y(new_n4255));
  OAI21xp33_ASAP7_75t_L     g03999(.A1(new_n4253), .A2(new_n4244), .B(new_n4065), .Y(new_n4256));
  NAND2xp33_ASAP7_75t_L     g04000(.A(new_n4256), .B(new_n4255), .Y(new_n4257));
  A2O1A1O1Ixp25_ASAP7_75t_L g04001(.A1(new_n4050), .A2(new_n3817), .B(new_n4045), .C(new_n4043), .D(new_n4257), .Y(new_n4258));
  O2A1O1Ixp33_ASAP7_75t_L   g04002(.A1(new_n3818), .A2(new_n3820), .B(new_n4044), .C(new_n4042), .Y(new_n4259));
  INVx1_ASAP7_75t_L         g04003(.A(new_n4259), .Y(new_n4260));
  AOI21xp33_ASAP7_75t_L     g04004(.A1(new_n4256), .A2(new_n4255), .B(new_n4260), .Y(new_n4261));
  NOR2xp33_ASAP7_75t_L      g04005(.A(new_n4258), .B(new_n4261), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g04006(.A(new_n3807), .B(new_n368), .Y(new_n4263));
  AOI221xp5_ASAP7_75t_L     g04007(.A1(new_n334), .A2(\b[32] ), .B1(new_n342), .B2(new_n3813), .C(new_n4263), .Y(new_n4264));
  OA211x2_ASAP7_75t_L       g04008(.A1(new_n365), .A2(new_n3419), .B(new_n4264), .C(\a[5] ), .Y(new_n4265));
  O2A1O1Ixp33_ASAP7_75t_L   g04009(.A1(new_n3419), .A2(new_n365), .B(new_n4264), .C(\a[5] ), .Y(new_n4266));
  NOR2xp33_ASAP7_75t_L      g04010(.A(new_n4266), .B(new_n4265), .Y(new_n4267));
  NOR2xp33_ASAP7_75t_L      g04011(.A(new_n4216), .B(new_n4219), .Y(new_n4268));
  NAND2xp33_ASAP7_75t_L     g04012(.A(new_n4225), .B(new_n4268), .Y(new_n4269));
  A2O1A1Ixp33_ASAP7_75t_L   g04013(.A1(new_n4227), .A2(new_n4226), .B(new_n4229), .C(new_n4269), .Y(new_n4270));
  NOR2xp33_ASAP7_75t_L      g04014(.A(new_n2852), .B(new_n481), .Y(new_n4271));
  INVx1_ASAP7_75t_L         g04015(.A(new_n4271), .Y(new_n4272));
  NAND2xp33_ASAP7_75t_L     g04016(.A(\b[29] ), .B(new_n441), .Y(new_n4273));
  AOI22xp33_ASAP7_75t_L     g04017(.A1(new_n451), .A2(\b[30] ), .B1(new_n448), .B2(new_n3219), .Y(new_n4274));
  NAND4xp25_ASAP7_75t_L     g04018(.A(new_n4274), .B(\a[8] ), .C(new_n4272), .D(new_n4273), .Y(new_n4275));
  NAND2xp33_ASAP7_75t_L     g04019(.A(new_n4273), .B(new_n4274), .Y(new_n4276));
  A2O1A1Ixp33_ASAP7_75t_L   g04020(.A1(\b[28] ), .A2(new_n480), .B(new_n4276), .C(new_n445), .Y(new_n4277));
  NAND2xp33_ASAP7_75t_L     g04021(.A(new_n4275), .B(new_n4277), .Y(new_n4278));
  OAI21xp33_ASAP7_75t_L     g04022(.A1(new_n4209), .A2(new_n4215), .B(new_n4218), .Y(new_n4279));
  INVx1_ASAP7_75t_L         g04023(.A(new_n4070), .Y(new_n4280));
  A2O1A1Ixp33_ASAP7_75t_L   g04024(.A1(new_n3999), .A2(new_n3998), .B(new_n3995), .C(new_n4280), .Y(new_n4281));
  NAND2xp33_ASAP7_75t_L     g04025(.A(\b[23] ), .B(new_n817), .Y(new_n4282));
  NAND2xp33_ASAP7_75t_L     g04026(.A(\b[24] ), .B(new_n826), .Y(new_n4283));
  OAI311xp33_ASAP7_75t_L    g04027(.A1(new_n2026), .A2(new_n2023), .A3(new_n911), .B1(new_n4283), .C1(new_n4282), .Y(new_n4284));
  AOI21xp33_ASAP7_75t_L     g04028(.A1(new_n908), .A2(\b[22] ), .B(new_n4284), .Y(new_n4285));
  NAND2xp33_ASAP7_75t_L     g04029(.A(\a[14] ), .B(new_n4285), .Y(new_n4286));
  A2O1A1Ixp33_ASAP7_75t_L   g04030(.A1(\b[22] ), .A2(new_n908), .B(new_n4284), .C(new_n813), .Y(new_n4287));
  NAND2xp33_ASAP7_75t_L     g04031(.A(new_n4287), .B(new_n4286), .Y(new_n4288));
  OAI211xp5_ASAP7_75t_L     g04032(.A1(new_n4167), .A2(new_n4168), .B(new_n4161), .C(new_n4157), .Y(new_n4289));
  INVx1_ASAP7_75t_L         g04033(.A(new_n4289), .Y(new_n4290));
  NOR2xp33_ASAP7_75t_L      g04034(.A(new_n1356), .B(new_n1412), .Y(new_n4291));
  AOI221xp5_ASAP7_75t_L     g04035(.A1(new_n1410), .A2(\b[17] ), .B1(new_n1404), .B2(new_n1363), .C(new_n4291), .Y(new_n4292));
  OAI211xp5_ASAP7_75t_L     g04036(.A1(new_n1051), .A2(new_n1549), .B(new_n4292), .C(\a[20] ), .Y(new_n4293));
  INVx1_ASAP7_75t_L         g04037(.A(new_n4291), .Y(new_n4294));
  OAI221xp5_ASAP7_75t_L     g04038(.A1(new_n1244), .A2(new_n1398), .B1(new_n1411), .B2(new_n3138), .C(new_n4294), .Y(new_n4295));
  A2O1A1Ixp33_ASAP7_75t_L   g04039(.A1(\b[16] ), .A2(new_n1548), .B(new_n4295), .C(new_n1401), .Y(new_n4296));
  NAND2xp33_ASAP7_75t_L     g04040(.A(new_n4296), .B(new_n4293), .Y(new_n4297));
  A2O1A1Ixp33_ASAP7_75t_L   g04041(.A1(new_n4160), .A2(new_n3940), .B(new_n4158), .C(new_n4155), .Y(new_n4298));
  OAI21xp33_ASAP7_75t_L     g04042(.A1(new_n4136), .A2(new_n4096), .B(new_n4139), .Y(new_n4299));
  NAND5xp2_ASAP7_75t_L      g04043(.A(new_n3885), .B(new_n3882), .C(new_n3875), .D(new_n4122), .E(\a[35] ), .Y(new_n4300));
  INVx1_ASAP7_75t_L         g04044(.A(\a[36] ), .Y(new_n4301));
  NAND2xp33_ASAP7_75t_L     g04045(.A(\a[35] ), .B(new_n4301), .Y(new_n4302));
  NAND2xp33_ASAP7_75t_L     g04046(.A(\a[36] ), .B(new_n3878), .Y(new_n4303));
  AND2x2_ASAP7_75t_L        g04047(.A(new_n4302), .B(new_n4303), .Y(new_n4304));
  NOR2xp33_ASAP7_75t_L      g04048(.A(new_n258), .B(new_n4304), .Y(new_n4305));
  OAI31xp33_ASAP7_75t_L     g04049(.A1(new_n4300), .A2(new_n4117), .A3(new_n4113), .B(new_n4305), .Y(new_n4306));
  AND4x1_ASAP7_75t_L        g04050(.A(new_n3885), .B(new_n3882), .C(new_n3875), .D(\a[35] ), .Y(new_n4307));
  NOR2xp33_ASAP7_75t_L      g04051(.A(new_n4114), .B(new_n283), .Y(new_n4308));
  AOI221xp5_ASAP7_75t_L     g04052(.A1(\b[2] ), .A2(new_n3884), .B1(new_n3874), .B2(\b[1] ), .C(new_n4308), .Y(new_n4309));
  INVx1_ASAP7_75t_L         g04053(.A(new_n4305), .Y(new_n4310));
  NAND5xp2_ASAP7_75t_L      g04054(.A(new_n4307), .B(new_n4309), .C(new_n4112), .D(new_n4310), .E(new_n4122), .Y(new_n4311));
  NAND2xp33_ASAP7_75t_L     g04055(.A(new_n4110), .B(new_n3650), .Y(new_n4312));
  NAND2xp33_ASAP7_75t_L     g04056(.A(\b[3] ), .B(new_n3884), .Y(new_n4313));
  OAI221xp5_ASAP7_75t_L     g04057(.A1(new_n278), .A2(new_n4312), .B1(new_n4114), .B2(new_n303), .C(new_n4313), .Y(new_n4314));
  AO211x2_ASAP7_75t_L       g04058(.A1(\b[1] ), .A2(new_n4111), .B(new_n3878), .C(new_n4314), .Y(new_n4315));
  A2O1A1Ixp33_ASAP7_75t_L   g04059(.A1(\b[1] ), .A2(new_n4111), .B(new_n4314), .C(new_n3878), .Y(new_n4316));
  AO22x1_ASAP7_75t_L        g04060(.A1(new_n4316), .A2(new_n4315), .B1(new_n4306), .B2(new_n4311), .Y(new_n4317));
  NAND4xp25_ASAP7_75t_L     g04061(.A(new_n4311), .B(new_n4306), .C(new_n4315), .D(new_n4316), .Y(new_n4318));
  NAND2xp33_ASAP7_75t_L     g04062(.A(\b[4] ), .B(new_n3491), .Y(new_n4319));
  NAND2xp33_ASAP7_75t_L     g04063(.A(\b[5] ), .B(new_n3260), .Y(new_n4320));
  AOI22xp33_ASAP7_75t_L     g04064(.A1(new_n3256), .A2(\b[6] ), .B1(new_n3254), .B2(new_n389), .Y(new_n4321));
  NAND4xp25_ASAP7_75t_L     g04065(.A(new_n4321), .B(\a[32] ), .C(new_n4319), .D(new_n4320), .Y(new_n4322));
  NAND2xp33_ASAP7_75t_L     g04066(.A(\b[6] ), .B(new_n3256), .Y(new_n4323));
  OAI211xp5_ASAP7_75t_L     g04067(.A1(new_n3261), .A2(new_n540), .B(new_n4320), .C(new_n4323), .Y(new_n4324));
  A2O1A1Ixp33_ASAP7_75t_L   g04068(.A1(\b[4] ), .A2(new_n3491), .B(new_n4324), .C(new_n3251), .Y(new_n4325));
  NAND4xp25_ASAP7_75t_L     g04069(.A(new_n4325), .B(new_n4317), .C(new_n4318), .D(new_n4322), .Y(new_n4326));
  AOI22xp33_ASAP7_75t_L     g04070(.A1(new_n4315), .A2(new_n4316), .B1(new_n4306), .B2(new_n4311), .Y(new_n4327));
  AND4x1_ASAP7_75t_L        g04071(.A(new_n4311), .B(new_n4306), .C(new_n4315), .D(new_n4316), .Y(new_n4328));
  AOI211xp5_ASAP7_75t_L     g04072(.A1(\b[4] ), .A2(new_n3491), .B(new_n3251), .C(new_n4324), .Y(new_n4329));
  AOI31xp33_ASAP7_75t_L     g04073(.A1(new_n4321), .A2(new_n4320), .A3(new_n4319), .B(\a[32] ), .Y(new_n4330));
  OAI22xp33_ASAP7_75t_L     g04074(.A1(new_n4329), .A2(new_n4330), .B1(new_n4327), .B2(new_n4328), .Y(new_n4331));
  OAI21xp33_ASAP7_75t_L     g04075(.A1(new_n4129), .A2(new_n4103), .B(new_n4126), .Y(new_n4332));
  NAND3xp33_ASAP7_75t_L     g04076(.A(new_n4332), .B(new_n4331), .C(new_n4326), .Y(new_n4333));
  NAND2xp33_ASAP7_75t_L     g04077(.A(new_n4326), .B(new_n4331), .Y(new_n4334));
  A2O1A1O1Ixp25_ASAP7_75t_L g04078(.A1(new_n3896), .A2(new_n3903), .B(new_n3889), .C(new_n4120), .D(new_n4130), .Y(new_n4335));
  NAND2xp33_ASAP7_75t_L     g04079(.A(new_n4335), .B(new_n4334), .Y(new_n4336));
  NOR2xp33_ASAP7_75t_L      g04080(.A(new_n421), .B(new_n2932), .Y(new_n4337));
  NAND2xp33_ASAP7_75t_L     g04081(.A(\b[8] ), .B(new_n2706), .Y(new_n4338));
  OAI221xp5_ASAP7_75t_L     g04082(.A1(new_n2708), .A2(new_n559), .B1(new_n2707), .B2(new_n978), .C(new_n4338), .Y(new_n4339));
  OR3x1_ASAP7_75t_L         g04083(.A(new_n4339), .B(new_n2697), .C(new_n4337), .Y(new_n4340));
  A2O1A1Ixp33_ASAP7_75t_L   g04084(.A1(\b[7] ), .A2(new_n2931), .B(new_n4339), .C(new_n2697), .Y(new_n4341));
  AO22x1_ASAP7_75t_L        g04085(.A1(new_n4341), .A2(new_n4340), .B1(new_n4336), .B2(new_n4333), .Y(new_n4342));
  NAND4xp25_ASAP7_75t_L     g04086(.A(new_n4333), .B(new_n4336), .C(new_n4341), .D(new_n4340), .Y(new_n4343));
  AOI21xp33_ASAP7_75t_L     g04087(.A1(new_n4343), .A2(new_n4342), .B(new_n4299), .Y(new_n4344));
  A2O1A1O1Ixp25_ASAP7_75t_L g04088(.A1(new_n3899), .A2(new_n3854), .B(new_n3911), .C(new_n4140), .D(new_n4132), .Y(new_n4345));
  AOI22xp33_ASAP7_75t_L     g04089(.A1(new_n4341), .A2(new_n4340), .B1(new_n4336), .B2(new_n4333), .Y(new_n4346));
  AND4x1_ASAP7_75t_L        g04090(.A(new_n4333), .B(new_n4341), .C(new_n4336), .D(new_n4340), .Y(new_n4347));
  NOR3xp33_ASAP7_75t_L      g04091(.A(new_n4345), .B(new_n4346), .C(new_n4347), .Y(new_n4348));
  NOR2xp33_ASAP7_75t_L      g04092(.A(new_n631), .B(new_n2387), .Y(new_n4349));
  INVx1_ASAP7_75t_L         g04093(.A(new_n4349), .Y(new_n4350));
  NOR2xp33_ASAP7_75t_L      g04094(.A(new_n695), .B(new_n2220), .Y(new_n4351));
  INVx1_ASAP7_75t_L         g04095(.A(new_n4351), .Y(new_n4352));
  AOI22xp33_ASAP7_75t_L     g04096(.A1(new_n2228), .A2(\b[12] ), .B1(new_n2226), .B2(new_n970), .Y(new_n4353));
  NAND4xp25_ASAP7_75t_L     g04097(.A(new_n4353), .B(\a[26] ), .C(new_n4350), .D(new_n4352), .Y(new_n4354));
  OAI221xp5_ASAP7_75t_L     g04098(.A1(new_n2234), .A2(new_n763), .B1(new_n2233), .B2(new_n775), .C(new_n4352), .Y(new_n4355));
  A2O1A1Ixp33_ASAP7_75t_L   g04099(.A1(\b[10] ), .A2(new_n2386), .B(new_n4355), .C(new_n2223), .Y(new_n4356));
  OAI211xp5_ASAP7_75t_L     g04100(.A1(new_n4344), .A2(new_n4348), .B(new_n4354), .C(new_n4356), .Y(new_n4357));
  OAI21xp33_ASAP7_75t_L     g04101(.A1(new_n4346), .A2(new_n4347), .B(new_n4345), .Y(new_n4358));
  NAND3xp33_ASAP7_75t_L     g04102(.A(new_n4299), .B(new_n4342), .C(new_n4343), .Y(new_n4359));
  INVx1_ASAP7_75t_L         g04103(.A(new_n4354), .Y(new_n4360));
  AOI31xp33_ASAP7_75t_L     g04104(.A1(new_n4353), .A2(new_n4352), .A3(new_n4350), .B(\a[26] ), .Y(new_n4361));
  OAI211xp5_ASAP7_75t_L     g04105(.A1(new_n4361), .A2(new_n4360), .B(new_n4359), .C(new_n4358), .Y(new_n4362));
  NAND2xp33_ASAP7_75t_L     g04106(.A(new_n4362), .B(new_n4357), .Y(new_n4363));
  NOR2xp33_ASAP7_75t_L      g04107(.A(new_n4137), .B(new_n4141), .Y(new_n4364));
  MAJIxp5_ASAP7_75t_L       g04108(.A(new_n4148), .B(new_n4095), .C(new_n4364), .Y(new_n4365));
  NOR2xp33_ASAP7_75t_L      g04109(.A(new_n4365), .B(new_n4363), .Y(new_n4366));
  AOI211xp5_ASAP7_75t_L     g04110(.A1(new_n4359), .A2(new_n4358), .B(new_n4360), .C(new_n4361), .Y(new_n4367));
  AOI211xp5_ASAP7_75t_L     g04111(.A1(new_n4356), .A2(new_n4354), .B(new_n4344), .C(new_n4348), .Y(new_n4368));
  NOR2xp33_ASAP7_75t_L      g04112(.A(new_n4368), .B(new_n4367), .Y(new_n4369));
  NAND2xp33_ASAP7_75t_L     g04113(.A(new_n4095), .B(new_n4364), .Y(new_n4370));
  A2O1A1Ixp33_ASAP7_75t_L   g04114(.A1(new_n4142), .A2(new_n4145), .B(new_n4088), .C(new_n4370), .Y(new_n4371));
  NOR2xp33_ASAP7_75t_L      g04115(.A(new_n4371), .B(new_n4369), .Y(new_n4372));
  NAND2xp33_ASAP7_75t_L     g04116(.A(\b[13] ), .B(new_n1910), .Y(new_n4373));
  NAND2xp33_ASAP7_75t_L     g04117(.A(\b[14] ), .B(new_n1770), .Y(new_n4374));
  AOI22xp33_ASAP7_75t_L     g04118(.A1(new_n1766), .A2(\b[15] ), .B1(new_n1764), .B2(new_n959), .Y(new_n4375));
  NAND4xp25_ASAP7_75t_L     g04119(.A(new_n4375), .B(\a[23] ), .C(new_n4373), .D(new_n4374), .Y(new_n4376));
  OAI221xp5_ASAP7_75t_L     g04120(.A1(new_n1772), .A2(new_n952), .B1(new_n1771), .B2(new_n2573), .C(new_n4374), .Y(new_n4377));
  A2O1A1Ixp33_ASAP7_75t_L   g04121(.A1(\b[13] ), .A2(new_n1910), .B(new_n4377), .C(new_n1761), .Y(new_n4378));
  NAND2xp33_ASAP7_75t_L     g04122(.A(new_n4376), .B(new_n4378), .Y(new_n4379));
  NOR3xp33_ASAP7_75t_L      g04123(.A(new_n4372), .B(new_n4366), .C(new_n4379), .Y(new_n4380));
  NAND2xp33_ASAP7_75t_L     g04124(.A(new_n4371), .B(new_n4369), .Y(new_n4381));
  NAND2xp33_ASAP7_75t_L     g04125(.A(new_n4365), .B(new_n4363), .Y(new_n4382));
  AND2x2_ASAP7_75t_L        g04126(.A(new_n4376), .B(new_n4378), .Y(new_n4383));
  AOI21xp33_ASAP7_75t_L     g04127(.A1(new_n4381), .A2(new_n4382), .B(new_n4383), .Y(new_n4384));
  OAI21xp33_ASAP7_75t_L     g04128(.A1(new_n4384), .A2(new_n4380), .B(new_n4298), .Y(new_n4385));
  A2O1A1O1Ixp25_ASAP7_75t_L g04129(.A1(new_n3939), .A2(new_n3946), .B(new_n3948), .C(new_n4151), .D(new_n4159), .Y(new_n4386));
  NAND3xp33_ASAP7_75t_L     g04130(.A(new_n4381), .B(new_n4383), .C(new_n4382), .Y(new_n4387));
  OAI21xp33_ASAP7_75t_L     g04131(.A1(new_n4366), .A2(new_n4372), .B(new_n4379), .Y(new_n4388));
  NAND3xp33_ASAP7_75t_L     g04132(.A(new_n4386), .B(new_n4387), .C(new_n4388), .Y(new_n4389));
  NAND3xp33_ASAP7_75t_L     g04133(.A(new_n4297), .B(new_n4389), .C(new_n4385), .Y(new_n4390));
  AND2x2_ASAP7_75t_L        g04134(.A(new_n4296), .B(new_n4293), .Y(new_n4391));
  AOI21xp33_ASAP7_75t_L     g04135(.A1(new_n4388), .A2(new_n4387), .B(new_n4386), .Y(new_n4392));
  NOR3xp33_ASAP7_75t_L      g04136(.A(new_n4298), .B(new_n4380), .C(new_n4384), .Y(new_n4393));
  OAI21xp33_ASAP7_75t_L     g04137(.A1(new_n4392), .A2(new_n4393), .B(new_n4391), .Y(new_n4394));
  AOI221xp5_ASAP7_75t_L     g04138(.A1(new_n4394), .A2(new_n4390), .B1(new_n4172), .B2(new_n4174), .C(new_n4290), .Y(new_n4395));
  NAND2xp33_ASAP7_75t_L     g04139(.A(new_n4390), .B(new_n4394), .Y(new_n4396));
  A2O1A1O1Ixp25_ASAP7_75t_L g04140(.A1(new_n4171), .A2(new_n4170), .B(new_n4177), .C(new_n4289), .D(new_n4396), .Y(new_n4397));
  NOR2xp33_ASAP7_75t_L      g04141(.A(new_n1493), .B(new_n1195), .Y(new_n4398));
  INVx1_ASAP7_75t_L         g04142(.A(new_n4398), .Y(new_n4399));
  NOR2xp33_ASAP7_75t_L      g04143(.A(new_n1594), .B(new_n1298), .Y(new_n4400));
  INVx1_ASAP7_75t_L         g04144(.A(new_n4400), .Y(new_n4401));
  AOI22xp33_ASAP7_75t_L     g04145(.A1(new_n1113), .A2(\b[21] ), .B1(new_n1110), .B2(new_n1715), .Y(new_n4402));
  NAND4xp25_ASAP7_75t_L     g04146(.A(new_n4402), .B(\a[17] ), .C(new_n4399), .D(new_n4401), .Y(new_n4403));
  AOI31xp33_ASAP7_75t_L     g04147(.A1(new_n4402), .A2(new_n4401), .A3(new_n4399), .B(\a[17] ), .Y(new_n4404));
  INVx1_ASAP7_75t_L         g04148(.A(new_n4404), .Y(new_n4405));
  NAND2xp33_ASAP7_75t_L     g04149(.A(new_n4403), .B(new_n4405), .Y(new_n4406));
  NOR3xp33_ASAP7_75t_L      g04150(.A(new_n4397), .B(new_n4406), .C(new_n4395), .Y(new_n4407));
  INVx1_ASAP7_75t_L         g04151(.A(new_n4395), .Y(new_n4408));
  A2O1A1Ixp33_ASAP7_75t_L   g04152(.A1(new_n4171), .A2(new_n4170), .B(new_n4177), .C(new_n4289), .Y(new_n4409));
  NAND3xp33_ASAP7_75t_L     g04153(.A(new_n4409), .B(new_n4390), .C(new_n4394), .Y(new_n4410));
  AND2x2_ASAP7_75t_L        g04154(.A(new_n4403), .B(new_n4405), .Y(new_n4411));
  AOI21xp33_ASAP7_75t_L     g04155(.A1(new_n4408), .A2(new_n4410), .B(new_n4411), .Y(new_n4412));
  A2O1A1O1Ixp25_ASAP7_75t_L g04156(.A1(new_n3971), .A2(new_n3965), .B(new_n3978), .C(new_n4079), .D(new_n4193), .Y(new_n4413));
  OAI22xp33_ASAP7_75t_L     g04157(.A1(new_n4413), .A2(new_n4194), .B1(new_n4407), .B2(new_n4412), .Y(new_n4414));
  NAND3xp33_ASAP7_75t_L     g04158(.A(new_n4411), .B(new_n4408), .C(new_n4410), .Y(new_n4415));
  OAI21xp33_ASAP7_75t_L     g04159(.A1(new_n4395), .A2(new_n4397), .B(new_n4406), .Y(new_n4416));
  A2O1A1O1Ixp25_ASAP7_75t_L g04160(.A1(new_n3972), .A2(new_n3973), .B(new_n4078), .C(new_n4186), .D(new_n4194), .Y(new_n4417));
  NAND3xp33_ASAP7_75t_L     g04161(.A(new_n4417), .B(new_n4416), .C(new_n4415), .Y(new_n4418));
  AOI21xp33_ASAP7_75t_L     g04162(.A1(new_n4418), .A2(new_n4414), .B(new_n4288), .Y(new_n4419));
  AND2x2_ASAP7_75t_L        g04163(.A(new_n4287), .B(new_n4286), .Y(new_n4420));
  AOI21xp33_ASAP7_75t_L     g04164(.A1(new_n4416), .A2(new_n4415), .B(new_n4417), .Y(new_n4421));
  NOR4xp25_ASAP7_75t_L      g04165(.A(new_n4413), .B(new_n4412), .C(new_n4407), .D(new_n4194), .Y(new_n4422));
  NOR3xp33_ASAP7_75t_L      g04166(.A(new_n4421), .B(new_n4422), .C(new_n4420), .Y(new_n4423));
  NOR2xp33_ASAP7_75t_L      g04167(.A(new_n4419), .B(new_n4423), .Y(new_n4424));
  A2O1A1Ixp33_ASAP7_75t_L   g04168(.A1(new_n4203), .A2(new_n4281), .B(new_n4202), .C(new_n4424), .Y(new_n4425));
  A2O1A1O1Ixp25_ASAP7_75t_L g04169(.A1(new_n4009), .A2(new_n4000), .B(new_n4070), .C(new_n4205), .D(new_n4202), .Y(new_n4426));
  OAI21xp33_ASAP7_75t_L     g04170(.A1(new_n4422), .A2(new_n4421), .B(new_n4420), .Y(new_n4427));
  NAND3xp33_ASAP7_75t_L     g04171(.A(new_n4418), .B(new_n4414), .C(new_n4288), .Y(new_n4428));
  NAND2xp33_ASAP7_75t_L     g04172(.A(new_n4428), .B(new_n4427), .Y(new_n4429));
  NAND2xp33_ASAP7_75t_L     g04173(.A(new_n4426), .B(new_n4429), .Y(new_n4430));
  NAND2xp33_ASAP7_75t_L     g04174(.A(\b[25] ), .B(new_n674), .Y(new_n4431));
  NAND2xp33_ASAP7_75t_L     g04175(.A(\b[26] ), .B(new_n590), .Y(new_n4432));
  AOI22xp33_ASAP7_75t_L     g04176(.A1(new_n600), .A2(\b[27] ), .B1(new_n597), .B2(new_n2657), .Y(new_n4433));
  AND4x1_ASAP7_75t_L        g04177(.A(new_n4433), .B(new_n4432), .C(new_n4431), .D(\a[11] ), .Y(new_n4434));
  AOI31xp33_ASAP7_75t_L     g04178(.A1(new_n4433), .A2(new_n4432), .A3(new_n4431), .B(\a[11] ), .Y(new_n4435));
  NOR2xp33_ASAP7_75t_L      g04179(.A(new_n4435), .B(new_n4434), .Y(new_n4436));
  NAND3xp33_ASAP7_75t_L     g04180(.A(new_n4425), .B(new_n4430), .C(new_n4436), .Y(new_n4437));
  NOR2xp33_ASAP7_75t_L      g04181(.A(new_n4426), .B(new_n4429), .Y(new_n4438));
  AOI221xp5_ASAP7_75t_L     g04182(.A1(new_n4428), .A2(new_n4427), .B1(new_n4205), .B2(new_n4281), .C(new_n4202), .Y(new_n4439));
  INVx1_ASAP7_75t_L         g04183(.A(new_n4436), .Y(new_n4440));
  OAI21xp33_ASAP7_75t_L     g04184(.A1(new_n4438), .A2(new_n4439), .B(new_n4440), .Y(new_n4441));
  NAND2xp33_ASAP7_75t_L     g04185(.A(new_n4441), .B(new_n4437), .Y(new_n4442));
  NAND2xp33_ASAP7_75t_L     g04186(.A(new_n4279), .B(new_n4442), .Y(new_n4443));
  A2O1A1O1Ixp25_ASAP7_75t_L g04187(.A1(new_n4013), .A2(new_n3843), .B(new_n4018), .C(new_n4217), .D(new_n4214), .Y(new_n4444));
  NAND3xp33_ASAP7_75t_L     g04188(.A(new_n4444), .B(new_n4437), .C(new_n4441), .Y(new_n4445));
  AOI21xp33_ASAP7_75t_L     g04189(.A1(new_n4443), .A2(new_n4445), .B(new_n4278), .Y(new_n4446));
  AND2x2_ASAP7_75t_L        g04190(.A(new_n4275), .B(new_n4277), .Y(new_n4447));
  AOI21xp33_ASAP7_75t_L     g04191(.A1(new_n4441), .A2(new_n4437), .B(new_n4444), .Y(new_n4448));
  NOR2xp33_ASAP7_75t_L      g04192(.A(new_n4279), .B(new_n4442), .Y(new_n4449));
  NOR3xp33_ASAP7_75t_L      g04193(.A(new_n4449), .B(new_n4448), .C(new_n4447), .Y(new_n4450));
  NOR2xp33_ASAP7_75t_L      g04194(.A(new_n4446), .B(new_n4450), .Y(new_n4451));
  AND2x2_ASAP7_75t_L        g04195(.A(new_n4451), .B(new_n4270), .Y(new_n4452));
  NOR2xp33_ASAP7_75t_L      g04196(.A(new_n4451), .B(new_n4270), .Y(new_n4453));
  NOR3xp33_ASAP7_75t_L      g04197(.A(new_n4452), .B(new_n4267), .C(new_n4453), .Y(new_n4454));
  INVx1_ASAP7_75t_L         g04198(.A(new_n4454), .Y(new_n4455));
  OAI21xp33_ASAP7_75t_L     g04199(.A1(new_n4453), .A2(new_n4452), .B(new_n4267), .Y(new_n4456));
  A2O1A1Ixp33_ASAP7_75t_L   g04200(.A1(new_n4243), .A2(new_n4038), .B(new_n4239), .C(new_n4246), .Y(new_n4457));
  NAND3xp33_ASAP7_75t_L     g04201(.A(new_n4457), .B(new_n4455), .C(new_n4456), .Y(new_n4458));
  OA21x2_ASAP7_75t_L        g04202(.A1(new_n4453), .A2(new_n4452), .B(new_n4267), .Y(new_n4459));
  A2O1A1Ixp33_ASAP7_75t_L   g04203(.A1(new_n4232), .A2(new_n4230), .B(new_n4238), .C(new_n4252), .Y(new_n4460));
  OAI211xp5_ASAP7_75t_L     g04204(.A1(new_n4454), .A2(new_n4459), .B(new_n4460), .C(new_n4246), .Y(new_n4461));
  NAND2xp33_ASAP7_75t_L     g04205(.A(new_n4458), .B(new_n4461), .Y(new_n4462));
  INVx1_ASAP7_75t_L         g04206(.A(new_n4054), .Y(new_n4463));
  NOR2xp33_ASAP7_75t_L      g04207(.A(\b[35] ), .B(\b[36] ), .Y(new_n4464));
  INVx1_ASAP7_75t_L         g04208(.A(\b[36] ), .Y(new_n4465));
  NOR2xp33_ASAP7_75t_L      g04209(.A(new_n4053), .B(new_n4465), .Y(new_n4466));
  NOR2xp33_ASAP7_75t_L      g04210(.A(new_n4464), .B(new_n4466), .Y(new_n4467));
  INVx1_ASAP7_75t_L         g04211(.A(new_n4467), .Y(new_n4468));
  O2A1O1Ixp33_ASAP7_75t_L   g04212(.A1(new_n4058), .A2(new_n4057), .B(new_n4463), .C(new_n4468), .Y(new_n4469));
  A2O1A1Ixp33_ASAP7_75t_L   g04213(.A1(\b[33] ), .A2(\b[32] ), .B(new_n3811), .C(new_n3829), .Y(new_n4470));
  O2A1O1Ixp33_ASAP7_75t_L   g04214(.A1(new_n3807), .A2(new_n3827), .B(new_n4470), .C(new_n4058), .Y(new_n4471));
  NOR3xp33_ASAP7_75t_L      g04215(.A(new_n4471), .B(new_n4467), .C(new_n4054), .Y(new_n4472));
  NOR2xp33_ASAP7_75t_L      g04216(.A(new_n4469), .B(new_n4472), .Y(new_n4473));
  NOR2xp33_ASAP7_75t_L      g04217(.A(new_n4465), .B(new_n632), .Y(new_n4474));
  AOI221xp5_ASAP7_75t_L     g04218(.A1(new_n380), .A2(\b[35] ), .B1(new_n269), .B2(new_n4473), .C(new_n4474), .Y(new_n4475));
  OA211x2_ASAP7_75t_L       g04219(.A1(new_n277), .A2(new_n3827), .B(new_n4475), .C(\a[2] ), .Y(new_n4476));
  O2A1O1Ixp33_ASAP7_75t_L   g04220(.A1(new_n3827), .A2(new_n277), .B(new_n4475), .C(\a[2] ), .Y(new_n4477));
  NOR2xp33_ASAP7_75t_L      g04221(.A(new_n4477), .B(new_n4476), .Y(new_n4478));
  XOR2x2_ASAP7_75t_L        g04222(.A(new_n4478), .B(new_n4462), .Y(new_n4479));
  A2O1A1O1Ixp25_ASAP7_75t_L g04223(.A1(new_n4044), .A2(new_n4047), .B(new_n4042), .C(new_n4256), .D(new_n4254), .Y(new_n4480));
  XNOR2x2_ASAP7_75t_L       g04224(.A(new_n4480), .B(new_n4479), .Y(\f[36] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04225(.A1(new_n4256), .A2(new_n4260), .B(new_n4254), .C(new_n4479), .Y(new_n4482));
  AOI21xp33_ASAP7_75t_L     g04226(.A1(new_n4270), .A2(new_n4451), .B(new_n4450), .Y(new_n4483));
  AOI22xp33_ASAP7_75t_L     g04227(.A1(new_n451), .A2(\b[31] ), .B1(new_n448), .B2(new_n3426), .Y(new_n4484));
  OAI221xp5_ASAP7_75t_L     g04228(.A1(new_n529), .A2(new_n3212), .B1(new_n2871), .B2(new_n481), .C(new_n4484), .Y(new_n4485));
  XNOR2x2_ASAP7_75t_L       g04229(.A(new_n445), .B(new_n4485), .Y(new_n4486));
  NOR3xp33_ASAP7_75t_L      g04230(.A(new_n4439), .B(new_n4438), .C(new_n4436), .Y(new_n4487));
  INVx1_ASAP7_75t_L         g04231(.A(new_n4487), .Y(new_n4488));
  A2O1A1Ixp33_ASAP7_75t_L   g04232(.A1(new_n4437), .A2(new_n4441), .B(new_n4444), .C(new_n4488), .Y(new_n4489));
  NOR2xp33_ASAP7_75t_L      g04233(.A(new_n2852), .B(new_n676), .Y(new_n4490));
  AOI221xp5_ASAP7_75t_L     g04234(.A1(new_n590), .A2(\b[27] ), .B1(new_n597), .B2(new_n2858), .C(new_n4490), .Y(new_n4491));
  OA211x2_ASAP7_75t_L       g04235(.A1(new_n1620), .A2(new_n2477), .B(new_n4491), .C(\a[11] ), .Y(new_n4492));
  O2A1O1Ixp33_ASAP7_75t_L   g04236(.A1(new_n2477), .A2(new_n1620), .B(new_n4491), .C(\a[11] ), .Y(new_n4493));
  NOR2xp33_ASAP7_75t_L      g04237(.A(new_n4493), .B(new_n4492), .Y(new_n4494));
  A2O1A1O1Ixp25_ASAP7_75t_L g04238(.A1(new_n4205), .A2(new_n4281), .B(new_n4202), .C(new_n4427), .D(new_n4423), .Y(new_n4495));
  NOR2xp33_ASAP7_75t_L      g04239(.A(new_n695), .B(new_n2387), .Y(new_n4496));
  NAND2xp33_ASAP7_75t_L     g04240(.A(\b[12] ), .B(new_n2232), .Y(new_n4497));
  NAND2xp33_ASAP7_75t_L     g04241(.A(\b[13] ), .B(new_n2228), .Y(new_n4498));
  OAI311xp33_ASAP7_75t_L    g04242(.A1(new_n799), .A2(new_n797), .A3(new_n2233), .B1(new_n4498), .C1(new_n4497), .Y(new_n4499));
  OR3x1_ASAP7_75t_L         g04243(.A(new_n4499), .B(new_n2223), .C(new_n4496), .Y(new_n4500));
  A2O1A1Ixp33_ASAP7_75t_L   g04244(.A1(\b[11] ), .A2(new_n2386), .B(new_n4499), .C(new_n2223), .Y(new_n4501));
  NAND2xp33_ASAP7_75t_L     g04245(.A(new_n4501), .B(new_n4500), .Y(new_n4502));
  OAI21xp33_ASAP7_75t_L     g04246(.A1(new_n4347), .A2(new_n4345), .B(new_n4342), .Y(new_n4503));
  NAND2xp33_ASAP7_75t_L     g04247(.A(\b[9] ), .B(new_n2706), .Y(new_n4504));
  NAND2xp33_ASAP7_75t_L     g04248(.A(\b[10] ), .B(new_n2702), .Y(new_n4505));
  OAI311xp33_ASAP7_75t_L    g04249(.A1(new_n639), .A2(new_n851), .A3(new_n2707), .B1(new_n4505), .C1(new_n4504), .Y(new_n4506));
  AOI211xp5_ASAP7_75t_L     g04250(.A1(\b[8] ), .A2(new_n2931), .B(new_n2697), .C(new_n4506), .Y(new_n4507));
  NOR2xp33_ASAP7_75t_L      g04251(.A(new_n503), .B(new_n2932), .Y(new_n4508));
  OA21x2_ASAP7_75t_L        g04252(.A1(new_n4508), .A2(new_n4506), .B(new_n2697), .Y(new_n4509));
  NOR2xp33_ASAP7_75t_L      g04253(.A(new_n4507), .B(new_n4509), .Y(new_n4510));
  AOI211xp5_ASAP7_75t_L     g04254(.A1(new_n4325), .A2(new_n4322), .B(new_n4327), .C(new_n4328), .Y(new_n4511));
  INVx1_ASAP7_75t_L         g04255(.A(new_n4511), .Y(new_n4512));
  NOR4xp25_ASAP7_75t_L      g04256(.A(new_n4329), .B(new_n4330), .C(new_n4327), .D(new_n4328), .Y(new_n4513));
  AOI22xp33_ASAP7_75t_L     g04257(.A1(new_n4317), .A2(new_n4318), .B1(new_n4322), .B2(new_n4325), .Y(new_n4514));
  O2A1O1Ixp33_ASAP7_75t_L   g04258(.A1(new_n3888), .A2(new_n3863), .B(new_n3897), .C(new_n4129), .Y(new_n4515));
  OAI22xp33_ASAP7_75t_L     g04259(.A1(new_n4515), .A2(new_n4130), .B1(new_n4513), .B2(new_n4514), .Y(new_n4516));
  NAND2xp33_ASAP7_75t_L     g04260(.A(\b[5] ), .B(new_n3491), .Y(new_n4517));
  NAND2xp33_ASAP7_75t_L     g04261(.A(\b[6] ), .B(new_n3260), .Y(new_n4518));
  AOI32xp33_ASAP7_75t_L     g04262(.A1(new_n424), .A2(new_n426), .A3(new_n3254), .B1(new_n3256), .B2(\b[7] ), .Y(new_n4519));
  NAND3xp33_ASAP7_75t_L     g04263(.A(new_n4519), .B(new_n4518), .C(new_n4517), .Y(new_n4520));
  NOR2xp33_ASAP7_75t_L      g04264(.A(new_n3251), .B(new_n4520), .Y(new_n4521));
  NAND2xp33_ASAP7_75t_L     g04265(.A(new_n3251), .B(new_n4520), .Y(new_n4522));
  INVx1_ASAP7_75t_L         g04266(.A(new_n4522), .Y(new_n4523));
  NOR3xp33_ASAP7_75t_L      g04267(.A(new_n4300), .B(new_n4113), .C(new_n4117), .Y(new_n4524));
  NAND2xp33_ASAP7_75t_L     g04268(.A(\b[2] ), .B(new_n4111), .Y(new_n4525));
  INVx1_ASAP7_75t_L         g04269(.A(new_n4525), .Y(new_n4526));
  NOR2xp33_ASAP7_75t_L      g04270(.A(new_n299), .B(new_n4312), .Y(new_n4527));
  OAI32xp33_ASAP7_75t_L     g04271(.A1(new_n325), .A2(new_n327), .A3(new_n4114), .B1(new_n4115), .B2(new_n323), .Y(new_n4528));
  NOR4xp25_ASAP7_75t_L      g04272(.A(new_n4528), .B(new_n3878), .C(new_n4526), .D(new_n4527), .Y(new_n4529));
  INVx1_ASAP7_75t_L         g04273(.A(new_n4527), .Y(new_n4530));
  AOI22xp33_ASAP7_75t_L     g04274(.A1(new_n3884), .A2(\b[4] ), .B1(new_n3881), .B2(new_n328), .Y(new_n4531));
  AOI31xp33_ASAP7_75t_L     g04275(.A1(new_n4531), .A2(new_n4530), .A3(new_n4525), .B(\a[35] ), .Y(new_n4532));
  NAND2xp33_ASAP7_75t_L     g04276(.A(\a[38] ), .B(new_n4305), .Y(new_n4533));
  XNOR2x2_ASAP7_75t_L       g04277(.A(\a[37] ), .B(\a[36] ), .Y(new_n4534));
  INVx1_ASAP7_75t_L         g04278(.A(new_n4534), .Y(new_n4535));
  NAND2xp33_ASAP7_75t_L     g04279(.A(new_n4535), .B(new_n4304), .Y(new_n4536));
  INVx1_ASAP7_75t_L         g04280(.A(\a[37] ), .Y(new_n4537));
  NAND2xp33_ASAP7_75t_L     g04281(.A(\a[38] ), .B(new_n4537), .Y(new_n4538));
  INVx1_ASAP7_75t_L         g04282(.A(\a[38] ), .Y(new_n4539));
  NAND2xp33_ASAP7_75t_L     g04283(.A(\a[37] ), .B(new_n4539), .Y(new_n4540));
  AND2x2_ASAP7_75t_L        g04284(.A(new_n4538), .B(new_n4540), .Y(new_n4541));
  NOR2xp33_ASAP7_75t_L      g04285(.A(new_n4304), .B(new_n4541), .Y(new_n4542));
  NAND2xp33_ASAP7_75t_L     g04286(.A(new_n4540), .B(new_n4538), .Y(new_n4543));
  NOR2xp33_ASAP7_75t_L      g04287(.A(new_n4543), .B(new_n4304), .Y(new_n4544));
  AOI22xp33_ASAP7_75t_L     g04288(.A1(new_n4544), .A2(\b[1] ), .B1(new_n271), .B2(new_n4542), .Y(new_n4545));
  O2A1O1Ixp33_ASAP7_75t_L   g04289(.A1(new_n4536), .A2(new_n258), .B(new_n4545), .C(new_n4533), .Y(new_n4546));
  NAND2xp33_ASAP7_75t_L     g04290(.A(new_n4303), .B(new_n4302), .Y(new_n4547));
  NOR2xp33_ASAP7_75t_L      g04291(.A(new_n4534), .B(new_n4547), .Y(new_n4548));
  NAND2xp33_ASAP7_75t_L     g04292(.A(new_n4543), .B(new_n4547), .Y(new_n4549));
  NAND2xp33_ASAP7_75t_L     g04293(.A(new_n4547), .B(new_n4541), .Y(new_n4550));
  OAI22xp33_ASAP7_75t_L     g04294(.A1(new_n4550), .A2(new_n276), .B1(new_n270), .B2(new_n4549), .Y(new_n4551));
  A2O1A1O1Ixp25_ASAP7_75t_L g04295(.A1(new_n4547), .A2(\a[38] ), .B(new_n4548), .C(\b[0] ), .D(new_n4551), .Y(new_n4552));
  NOR2xp33_ASAP7_75t_L      g04296(.A(new_n4552), .B(new_n4546), .Y(new_n4553));
  NOR3xp33_ASAP7_75t_L      g04297(.A(new_n4532), .B(new_n4553), .C(new_n4529), .Y(new_n4554));
  NAND4xp25_ASAP7_75t_L     g04298(.A(new_n4531), .B(\a[35] ), .C(new_n4525), .D(new_n4530), .Y(new_n4555));
  OAI31xp33_ASAP7_75t_L     g04299(.A1(new_n4528), .A2(new_n4527), .A3(new_n4526), .B(new_n3878), .Y(new_n4556));
  OR2x4_ASAP7_75t_L         g04300(.A(new_n4552), .B(new_n4546), .Y(new_n4557));
  AOI21xp33_ASAP7_75t_L     g04301(.A1(new_n4556), .A2(new_n4555), .B(new_n4557), .Y(new_n4558));
  NOR2xp33_ASAP7_75t_L      g04302(.A(new_n4554), .B(new_n4558), .Y(new_n4559));
  A2O1A1Ixp33_ASAP7_75t_L   g04303(.A1(new_n4524), .A2(new_n4305), .B(new_n4327), .C(new_n4559), .Y(new_n4560));
  NAND2xp33_ASAP7_75t_L     g04304(.A(new_n4305), .B(new_n4524), .Y(new_n4561));
  OAI211xp5_ASAP7_75t_L     g04305(.A1(new_n4554), .A2(new_n4558), .B(new_n4317), .C(new_n4561), .Y(new_n4562));
  AOI211xp5_ASAP7_75t_L     g04306(.A1(new_n4560), .A2(new_n4562), .B(new_n4523), .C(new_n4521), .Y(new_n4563));
  INVx1_ASAP7_75t_L         g04307(.A(new_n4521), .Y(new_n4564));
  AOI211xp5_ASAP7_75t_L     g04308(.A1(new_n4317), .A2(new_n4561), .B(new_n4554), .C(new_n4558), .Y(new_n4565));
  NAND3xp33_ASAP7_75t_L     g04309(.A(new_n4557), .B(new_n4556), .C(new_n4555), .Y(new_n4566));
  OAI21xp33_ASAP7_75t_L     g04310(.A1(new_n4529), .A2(new_n4532), .B(new_n4553), .Y(new_n4567));
  AOI221xp5_ASAP7_75t_L     g04311(.A1(new_n4305), .A2(new_n4524), .B1(new_n4567), .B2(new_n4566), .C(new_n4327), .Y(new_n4568));
  AOI211xp5_ASAP7_75t_L     g04312(.A1(new_n4564), .A2(new_n4522), .B(new_n4565), .C(new_n4568), .Y(new_n4569));
  AOI211xp5_ASAP7_75t_L     g04313(.A1(new_n4516), .A2(new_n4512), .B(new_n4569), .C(new_n4563), .Y(new_n4570));
  OAI211xp5_ASAP7_75t_L     g04314(.A1(new_n4568), .A2(new_n4565), .B(new_n4522), .C(new_n4564), .Y(new_n4571));
  OAI211xp5_ASAP7_75t_L     g04315(.A1(new_n4523), .A2(new_n4521), .B(new_n4560), .C(new_n4562), .Y(new_n4572));
  AOI221xp5_ASAP7_75t_L     g04316(.A1(new_n4334), .A2(new_n4332), .B1(new_n4571), .B2(new_n4572), .C(new_n4511), .Y(new_n4573));
  OAI21xp33_ASAP7_75t_L     g04317(.A1(new_n4573), .A2(new_n4570), .B(new_n4510), .Y(new_n4574));
  INVx1_ASAP7_75t_L         g04318(.A(new_n4510), .Y(new_n4575));
  A2O1A1Ixp33_ASAP7_75t_L   g04319(.A1(new_n4331), .A2(new_n4326), .B(new_n4335), .C(new_n4512), .Y(new_n4576));
  NAND3xp33_ASAP7_75t_L     g04320(.A(new_n4576), .B(new_n4571), .C(new_n4572), .Y(new_n4577));
  O2A1O1Ixp33_ASAP7_75t_L   g04321(.A1(new_n4130), .A2(new_n4515), .B(new_n4334), .C(new_n4511), .Y(new_n4578));
  OAI21xp33_ASAP7_75t_L     g04322(.A1(new_n4563), .A2(new_n4569), .B(new_n4578), .Y(new_n4579));
  NAND3xp33_ASAP7_75t_L     g04323(.A(new_n4575), .B(new_n4579), .C(new_n4577), .Y(new_n4580));
  NAND3xp33_ASAP7_75t_L     g04324(.A(new_n4503), .B(new_n4574), .C(new_n4580), .Y(new_n4581));
  A2O1A1O1Ixp25_ASAP7_75t_L g04325(.A1(new_n4138), .A2(new_n4140), .B(new_n4132), .C(new_n4343), .D(new_n4346), .Y(new_n4582));
  AOI21xp33_ASAP7_75t_L     g04326(.A1(new_n4579), .A2(new_n4577), .B(new_n4575), .Y(new_n4583));
  NOR3xp33_ASAP7_75t_L      g04327(.A(new_n4570), .B(new_n4510), .C(new_n4573), .Y(new_n4584));
  OAI21xp33_ASAP7_75t_L     g04328(.A1(new_n4584), .A2(new_n4583), .B(new_n4582), .Y(new_n4585));
  AOI21xp33_ASAP7_75t_L     g04329(.A1(new_n4581), .A2(new_n4585), .B(new_n4502), .Y(new_n4586));
  AND2x2_ASAP7_75t_L        g04330(.A(new_n4501), .B(new_n4500), .Y(new_n4587));
  NOR3xp33_ASAP7_75t_L      g04331(.A(new_n4582), .B(new_n4583), .C(new_n4584), .Y(new_n4588));
  AOI21xp33_ASAP7_75t_L     g04332(.A1(new_n4580), .A2(new_n4574), .B(new_n4503), .Y(new_n4589));
  NOR3xp33_ASAP7_75t_L      g04333(.A(new_n4589), .B(new_n4588), .C(new_n4587), .Y(new_n4590));
  NOR2xp33_ASAP7_75t_L      g04334(.A(new_n4590), .B(new_n4586), .Y(new_n4591));
  A2O1A1Ixp33_ASAP7_75t_L   g04335(.A1(new_n4371), .A2(new_n4357), .B(new_n4368), .C(new_n4591), .Y(new_n4592));
  INVx1_ASAP7_75t_L         g04336(.A(new_n4095), .Y(new_n4593));
  NAND2xp33_ASAP7_75t_L     g04337(.A(new_n4144), .B(new_n4143), .Y(new_n4594));
  NOR2xp33_ASAP7_75t_L      g04338(.A(new_n4593), .B(new_n4594), .Y(new_n4595));
  A2O1A1O1Ixp25_ASAP7_75t_L g04339(.A1(new_n4148), .A2(new_n4149), .B(new_n4595), .C(new_n4357), .D(new_n4368), .Y(new_n4596));
  OAI21xp33_ASAP7_75t_L     g04340(.A1(new_n4588), .A2(new_n4589), .B(new_n4587), .Y(new_n4597));
  NAND3xp33_ASAP7_75t_L     g04341(.A(new_n4581), .B(new_n4502), .C(new_n4585), .Y(new_n4598));
  NAND2xp33_ASAP7_75t_L     g04342(.A(new_n4598), .B(new_n4597), .Y(new_n4599));
  NAND2xp33_ASAP7_75t_L     g04343(.A(new_n4596), .B(new_n4599), .Y(new_n4600));
  AOI22xp33_ASAP7_75t_L     g04344(.A1(new_n1766), .A2(\b[16] ), .B1(new_n1764), .B2(new_n1058), .Y(new_n4601));
  OAI221xp5_ASAP7_75t_L     g04345(.A1(new_n1758), .A2(new_n952), .B1(new_n871), .B2(new_n1911), .C(new_n4601), .Y(new_n4602));
  XNOR2x2_ASAP7_75t_L       g04346(.A(\a[23] ), .B(new_n4602), .Y(new_n4603));
  NAND3xp33_ASAP7_75t_L     g04347(.A(new_n4603), .B(new_n4592), .C(new_n4600), .Y(new_n4604));
  O2A1O1Ixp33_ASAP7_75t_L   g04348(.A1(new_n4367), .A2(new_n4365), .B(new_n4362), .C(new_n4599), .Y(new_n4605));
  OAI21xp33_ASAP7_75t_L     g04349(.A1(new_n4367), .A2(new_n4365), .B(new_n4362), .Y(new_n4606));
  NOR2xp33_ASAP7_75t_L      g04350(.A(new_n4591), .B(new_n4606), .Y(new_n4607));
  XNOR2x2_ASAP7_75t_L       g04351(.A(new_n1761), .B(new_n4602), .Y(new_n4608));
  OAI21xp33_ASAP7_75t_L     g04352(.A1(new_n4605), .A2(new_n4607), .B(new_n4608), .Y(new_n4609));
  XNOR2x2_ASAP7_75t_L       g04353(.A(new_n4371), .B(new_n4363), .Y(new_n4610));
  MAJIxp5_ASAP7_75t_L       g04354(.A(new_n4298), .B(new_n4379), .C(new_n4610), .Y(new_n4611));
  NAND3xp33_ASAP7_75t_L     g04355(.A(new_n4611), .B(new_n4609), .C(new_n4604), .Y(new_n4612));
  NOR3xp33_ASAP7_75t_L      g04356(.A(new_n4608), .B(new_n4607), .C(new_n4605), .Y(new_n4613));
  AOI21xp33_ASAP7_75t_L     g04357(.A1(new_n4592), .A2(new_n4600), .B(new_n4603), .Y(new_n4614));
  NAND3xp33_ASAP7_75t_L     g04358(.A(new_n4381), .B(new_n4382), .C(new_n4379), .Y(new_n4615));
  A2O1A1Ixp33_ASAP7_75t_L   g04359(.A1(new_n4388), .A2(new_n4387), .B(new_n4386), .C(new_n4615), .Y(new_n4616));
  OAI21xp33_ASAP7_75t_L     g04360(.A1(new_n4613), .A2(new_n4614), .B(new_n4616), .Y(new_n4617));
  NAND2xp33_ASAP7_75t_L     g04361(.A(\b[17] ), .B(new_n1548), .Y(new_n4618));
  NAND2xp33_ASAP7_75t_L     g04362(.A(\b[18] ), .B(new_n1410), .Y(new_n4619));
  AOI32xp33_ASAP7_75t_L     g04363(.A1(new_n2792), .A2(new_n1496), .A3(new_n1404), .B1(new_n1406), .B2(\b[19] ), .Y(new_n4620));
  NAND3xp33_ASAP7_75t_L     g04364(.A(new_n4620), .B(new_n4619), .C(new_n4618), .Y(new_n4621));
  XNOR2x2_ASAP7_75t_L       g04365(.A(\a[20] ), .B(new_n4621), .Y(new_n4622));
  NAND3xp33_ASAP7_75t_L     g04366(.A(new_n4612), .B(new_n4617), .C(new_n4622), .Y(new_n4623));
  NOR3xp33_ASAP7_75t_L      g04367(.A(new_n4616), .B(new_n4614), .C(new_n4613), .Y(new_n4624));
  AOI22xp33_ASAP7_75t_L     g04368(.A1(new_n4604), .A2(new_n4609), .B1(new_n4615), .B2(new_n4385), .Y(new_n4625));
  XNOR2x2_ASAP7_75t_L       g04369(.A(new_n1401), .B(new_n4621), .Y(new_n4626));
  OAI21xp33_ASAP7_75t_L     g04370(.A1(new_n4625), .A2(new_n4624), .B(new_n4626), .Y(new_n4627));
  NOR3xp33_ASAP7_75t_L      g04371(.A(new_n4391), .B(new_n4393), .C(new_n4392), .Y(new_n4628));
  A2O1A1O1Ixp25_ASAP7_75t_L g04372(.A1(new_n4172), .A2(new_n4174), .B(new_n4290), .C(new_n4394), .D(new_n4628), .Y(new_n4629));
  AND3x1_ASAP7_75t_L        g04373(.A(new_n4629), .B(new_n4627), .C(new_n4623), .Y(new_n4630));
  AOI21xp33_ASAP7_75t_L     g04374(.A1(new_n4627), .A2(new_n4623), .B(new_n4629), .Y(new_n4631));
  NAND2xp33_ASAP7_75t_L     g04375(.A(\b[20] ), .B(new_n1194), .Y(new_n4632));
  NAND2xp33_ASAP7_75t_L     g04376(.A(\b[21] ), .B(new_n1103), .Y(new_n4633));
  AOI32xp33_ASAP7_75t_L     g04377(.A1(new_n1862), .A2(new_n1860), .A3(new_n1110), .B1(new_n1113), .B2(\b[22] ), .Y(new_n4634));
  NAND4xp25_ASAP7_75t_L     g04378(.A(new_n4634), .B(\a[17] ), .C(new_n4632), .D(new_n4633), .Y(new_n4635));
  AOI31xp33_ASAP7_75t_L     g04379(.A1(new_n4634), .A2(new_n4633), .A3(new_n4632), .B(\a[17] ), .Y(new_n4636));
  INVx1_ASAP7_75t_L         g04380(.A(new_n4636), .Y(new_n4637));
  NAND2xp33_ASAP7_75t_L     g04381(.A(new_n4635), .B(new_n4637), .Y(new_n4638));
  NOR3xp33_ASAP7_75t_L      g04382(.A(new_n4630), .B(new_n4631), .C(new_n4638), .Y(new_n4639));
  NAND3xp33_ASAP7_75t_L     g04383(.A(new_n4629), .B(new_n4627), .C(new_n4623), .Y(new_n4640));
  NAND2xp33_ASAP7_75t_L     g04384(.A(new_n4623), .B(new_n4627), .Y(new_n4641));
  A2O1A1Ixp33_ASAP7_75t_L   g04385(.A1(new_n4394), .A2(new_n4409), .B(new_n4628), .C(new_n4641), .Y(new_n4642));
  AND2x2_ASAP7_75t_L        g04386(.A(new_n4635), .B(new_n4637), .Y(new_n4643));
  AOI21xp33_ASAP7_75t_L     g04387(.A1(new_n4642), .A2(new_n4640), .B(new_n4643), .Y(new_n4644));
  NOR2xp33_ASAP7_75t_L      g04388(.A(new_n4639), .B(new_n4644), .Y(new_n4645));
  NAND3xp33_ASAP7_75t_L     g04389(.A(new_n4408), .B(new_n4410), .C(new_n4406), .Y(new_n4646));
  NAND3xp33_ASAP7_75t_L     g04390(.A(new_n4645), .B(new_n4414), .C(new_n4646), .Y(new_n4647));
  NAND3xp33_ASAP7_75t_L     g04391(.A(new_n4642), .B(new_n4640), .C(new_n4643), .Y(new_n4648));
  OAI21xp33_ASAP7_75t_L     g04392(.A1(new_n4631), .A2(new_n4630), .B(new_n4638), .Y(new_n4649));
  NAND2xp33_ASAP7_75t_L     g04393(.A(new_n4648), .B(new_n4649), .Y(new_n4650));
  A2O1A1Ixp33_ASAP7_75t_L   g04394(.A1(new_n4416), .A2(new_n4415), .B(new_n4417), .C(new_n4646), .Y(new_n4651));
  NAND2xp33_ASAP7_75t_L     g04395(.A(new_n4651), .B(new_n4650), .Y(new_n4652));
  NOR2xp33_ASAP7_75t_L      g04396(.A(new_n1995), .B(new_n909), .Y(new_n4653));
  NAND2xp33_ASAP7_75t_L     g04397(.A(\b[24] ), .B(new_n817), .Y(new_n4654));
  OAI221xp5_ASAP7_75t_L     g04398(.A1(new_n912), .A2(new_n2180), .B1(new_n911), .B2(new_n2187), .C(new_n4654), .Y(new_n4655));
  OR3x1_ASAP7_75t_L         g04399(.A(new_n4655), .B(new_n813), .C(new_n4653), .Y(new_n4656));
  A2O1A1Ixp33_ASAP7_75t_L   g04400(.A1(\b[23] ), .A2(new_n908), .B(new_n4655), .C(new_n813), .Y(new_n4657));
  NAND2xp33_ASAP7_75t_L     g04401(.A(new_n4657), .B(new_n4656), .Y(new_n4658));
  AOI21xp33_ASAP7_75t_L     g04402(.A1(new_n4647), .A2(new_n4652), .B(new_n4658), .Y(new_n4659));
  NOR2xp33_ASAP7_75t_L      g04403(.A(new_n4651), .B(new_n4650), .Y(new_n4660));
  AOI22xp33_ASAP7_75t_L     g04404(.A1(new_n4648), .A2(new_n4649), .B1(new_n4646), .B2(new_n4414), .Y(new_n4661));
  AND2x2_ASAP7_75t_L        g04405(.A(new_n4657), .B(new_n4656), .Y(new_n4662));
  NOR3xp33_ASAP7_75t_L      g04406(.A(new_n4660), .B(new_n4662), .C(new_n4661), .Y(new_n4663));
  NOR2xp33_ASAP7_75t_L      g04407(.A(new_n4663), .B(new_n4659), .Y(new_n4664));
  NAND2xp33_ASAP7_75t_L     g04408(.A(new_n4495), .B(new_n4664), .Y(new_n4665));
  OAI21xp33_ASAP7_75t_L     g04409(.A1(new_n4197), .A2(new_n4211), .B(new_n4206), .Y(new_n4666));
  OAI21xp33_ASAP7_75t_L     g04410(.A1(new_n4661), .A2(new_n4660), .B(new_n4662), .Y(new_n4667));
  NAND3xp33_ASAP7_75t_L     g04411(.A(new_n4647), .B(new_n4652), .C(new_n4658), .Y(new_n4668));
  NAND2xp33_ASAP7_75t_L     g04412(.A(new_n4667), .B(new_n4668), .Y(new_n4669));
  A2O1A1Ixp33_ASAP7_75t_L   g04413(.A1(new_n4427), .A2(new_n4666), .B(new_n4423), .C(new_n4669), .Y(new_n4670));
  NAND3xp33_ASAP7_75t_L     g04414(.A(new_n4670), .B(new_n4665), .C(new_n4494), .Y(new_n4671));
  OR2x4_ASAP7_75t_L         g04415(.A(new_n4493), .B(new_n4492), .Y(new_n4672));
  OAI21xp33_ASAP7_75t_L     g04416(.A1(new_n4419), .A2(new_n4426), .B(new_n4428), .Y(new_n4673));
  NOR2xp33_ASAP7_75t_L      g04417(.A(new_n4673), .B(new_n4669), .Y(new_n4674));
  O2A1O1Ixp33_ASAP7_75t_L   g04418(.A1(new_n4426), .A2(new_n4419), .B(new_n4428), .C(new_n4664), .Y(new_n4675));
  OAI21xp33_ASAP7_75t_L     g04419(.A1(new_n4674), .A2(new_n4675), .B(new_n4672), .Y(new_n4676));
  NAND3xp33_ASAP7_75t_L     g04420(.A(new_n4489), .B(new_n4671), .C(new_n4676), .Y(new_n4677));
  NOR2xp33_ASAP7_75t_L      g04421(.A(new_n4438), .B(new_n4439), .Y(new_n4678));
  MAJIxp5_ASAP7_75t_L       g04422(.A(new_n4279), .B(new_n4678), .C(new_n4440), .Y(new_n4679));
  NOR3xp33_ASAP7_75t_L      g04423(.A(new_n4672), .B(new_n4674), .C(new_n4675), .Y(new_n4680));
  AOI21xp33_ASAP7_75t_L     g04424(.A1(new_n4670), .A2(new_n4665), .B(new_n4494), .Y(new_n4681));
  OAI21xp33_ASAP7_75t_L     g04425(.A1(new_n4680), .A2(new_n4681), .B(new_n4679), .Y(new_n4682));
  AOI21xp33_ASAP7_75t_L     g04426(.A1(new_n4682), .A2(new_n4677), .B(new_n4486), .Y(new_n4683));
  AND3x1_ASAP7_75t_L        g04427(.A(new_n4682), .B(new_n4486), .C(new_n4677), .Y(new_n4684));
  NOR2xp33_ASAP7_75t_L      g04428(.A(new_n4683), .B(new_n4684), .Y(new_n4685));
  XNOR2x2_ASAP7_75t_L       g04429(.A(new_n4483), .B(new_n4685), .Y(new_n4686));
  NAND2xp33_ASAP7_75t_L     g04430(.A(new_n342), .B(new_n3833), .Y(new_n4687));
  OAI221xp5_ASAP7_75t_L     g04431(.A1(new_n368), .A2(new_n3827), .B1(new_n3807), .B2(new_n406), .C(new_n4687), .Y(new_n4688));
  AOI21xp33_ASAP7_75t_L     g04432(.A1(new_n366), .A2(\b[32] ), .B(new_n4688), .Y(new_n4689));
  NAND2xp33_ASAP7_75t_L     g04433(.A(\a[5] ), .B(new_n4689), .Y(new_n4690));
  A2O1A1Ixp33_ASAP7_75t_L   g04434(.A1(\b[32] ), .A2(new_n366), .B(new_n4688), .C(new_n339), .Y(new_n4691));
  NAND2xp33_ASAP7_75t_L     g04435(.A(new_n4691), .B(new_n4690), .Y(new_n4692));
  INVx1_ASAP7_75t_L         g04436(.A(new_n4692), .Y(new_n4693));
  NAND2xp33_ASAP7_75t_L     g04437(.A(new_n4693), .B(new_n4686), .Y(new_n4694));
  XOR2x2_ASAP7_75t_L        g04438(.A(new_n4483), .B(new_n4685), .Y(new_n4695));
  NAND2xp33_ASAP7_75t_L     g04439(.A(new_n4692), .B(new_n4695), .Y(new_n4696));
  A2O1A1O1Ixp25_ASAP7_75t_L g04440(.A1(new_n4245), .A2(new_n4252), .B(new_n4242), .C(new_n4456), .D(new_n4454), .Y(new_n4697));
  AND3x1_ASAP7_75t_L        g04441(.A(new_n4694), .B(new_n4696), .C(new_n4697), .Y(new_n4698));
  AOI21xp33_ASAP7_75t_L     g04442(.A1(new_n4694), .A2(new_n4696), .B(new_n4697), .Y(new_n4699));
  NOR2xp33_ASAP7_75t_L      g04443(.A(\b[36] ), .B(\b[37] ), .Y(new_n4700));
  INVx1_ASAP7_75t_L         g04444(.A(\b[37] ), .Y(new_n4701));
  NOR2xp33_ASAP7_75t_L      g04445(.A(new_n4465), .B(new_n4701), .Y(new_n4702));
  NOR2xp33_ASAP7_75t_L      g04446(.A(new_n4700), .B(new_n4702), .Y(new_n4703));
  A2O1A1Ixp33_ASAP7_75t_L   g04447(.A1(\b[36] ), .A2(\b[35] ), .B(new_n4469), .C(new_n4703), .Y(new_n4704));
  INVx1_ASAP7_75t_L         g04448(.A(new_n4704), .Y(new_n4705));
  INVx1_ASAP7_75t_L         g04449(.A(new_n4466), .Y(new_n4706));
  A2O1A1Ixp33_ASAP7_75t_L   g04450(.A1(new_n4056), .A2(new_n4463), .B(new_n4464), .C(new_n4706), .Y(new_n4707));
  NOR2xp33_ASAP7_75t_L      g04451(.A(new_n4703), .B(new_n4707), .Y(new_n4708));
  NOR2xp33_ASAP7_75t_L      g04452(.A(new_n4705), .B(new_n4708), .Y(new_n4709));
  NOR2xp33_ASAP7_75t_L      g04453(.A(new_n4701), .B(new_n632), .Y(new_n4710));
  AOI221xp5_ASAP7_75t_L     g04454(.A1(new_n380), .A2(\b[36] ), .B1(new_n269), .B2(new_n4709), .C(new_n4710), .Y(new_n4711));
  OA211x2_ASAP7_75t_L       g04455(.A1(new_n277), .A2(new_n4053), .B(new_n4711), .C(\a[2] ), .Y(new_n4712));
  O2A1O1Ixp33_ASAP7_75t_L   g04456(.A1(new_n4053), .A2(new_n277), .B(new_n4711), .C(\a[2] ), .Y(new_n4713));
  NOR2xp33_ASAP7_75t_L      g04457(.A(new_n4713), .B(new_n4712), .Y(new_n4714));
  OAI21xp33_ASAP7_75t_L     g04458(.A1(new_n4699), .A2(new_n4698), .B(new_n4714), .Y(new_n4715));
  NOR3xp33_ASAP7_75t_L      g04459(.A(new_n4698), .B(new_n4699), .C(new_n4714), .Y(new_n4716));
  INVx1_ASAP7_75t_L         g04460(.A(new_n4716), .Y(new_n4717));
  NAND2xp33_ASAP7_75t_L     g04461(.A(new_n4715), .B(new_n4717), .Y(new_n4718));
  O2A1O1Ixp33_ASAP7_75t_L   g04462(.A1(new_n4462), .A2(new_n4478), .B(new_n4482), .C(new_n4718), .Y(new_n4719));
  MAJIxp5_ASAP7_75t_L       g04463(.A(new_n4480), .B(new_n4478), .C(new_n4462), .Y(new_n4720));
  AOI21xp33_ASAP7_75t_L     g04464(.A1(new_n4717), .A2(new_n4715), .B(new_n4720), .Y(new_n4721));
  NOR2xp33_ASAP7_75t_L      g04465(.A(new_n4721), .B(new_n4719), .Y(\f[37] ));
  INVx1_ASAP7_75t_L         g04466(.A(new_n4720), .Y(new_n4723));
  MAJIxp5_ASAP7_75t_L       g04467(.A(new_n4697), .B(new_n4695), .C(new_n4693), .Y(new_n4724));
  NAND2xp33_ASAP7_75t_L     g04468(.A(\b[35] ), .B(new_n345), .Y(new_n4725));
  OAI221xp5_ASAP7_75t_L     g04469(.A1(new_n3827), .A2(new_n406), .B1(new_n367), .B2(new_n4060), .C(new_n4725), .Y(new_n4726));
  AOI21xp33_ASAP7_75t_L     g04470(.A1(new_n366), .A2(\b[33] ), .B(new_n4726), .Y(new_n4727));
  NAND2xp33_ASAP7_75t_L     g04471(.A(\a[5] ), .B(new_n4727), .Y(new_n4728));
  A2O1A1Ixp33_ASAP7_75t_L   g04472(.A1(\b[33] ), .A2(new_n366), .B(new_n4726), .C(new_n339), .Y(new_n4729));
  NAND2xp33_ASAP7_75t_L     g04473(.A(new_n4729), .B(new_n4728), .Y(new_n4730));
  INVx1_ASAP7_75t_L         g04474(.A(new_n4730), .Y(new_n4731));
  INVx1_ASAP7_75t_L         g04475(.A(new_n4684), .Y(new_n4732));
  NOR2xp33_ASAP7_75t_L      g04476(.A(new_n3212), .B(new_n481), .Y(new_n4733));
  INVx1_ASAP7_75t_L         g04477(.A(new_n4733), .Y(new_n4734));
  NAND2xp33_ASAP7_75t_L     g04478(.A(\b[31] ), .B(new_n441), .Y(new_n4735));
  AOI22xp33_ASAP7_75t_L     g04479(.A1(new_n451), .A2(\b[32] ), .B1(new_n448), .B2(new_n3450), .Y(new_n4736));
  NAND4xp25_ASAP7_75t_L     g04480(.A(new_n4736), .B(\a[8] ), .C(new_n4734), .D(new_n4735), .Y(new_n4737));
  NAND2xp33_ASAP7_75t_L     g04481(.A(new_n4735), .B(new_n4736), .Y(new_n4738));
  A2O1A1Ixp33_ASAP7_75t_L   g04482(.A1(\b[30] ), .A2(new_n480), .B(new_n4738), .C(new_n445), .Y(new_n4739));
  AND2x2_ASAP7_75t_L        g04483(.A(new_n4737), .B(new_n4739), .Y(new_n4740));
  NAND2xp33_ASAP7_75t_L     g04484(.A(\b[28] ), .B(new_n590), .Y(new_n4741));
  OAI221xp5_ASAP7_75t_L     g04485(.A1(new_n676), .A2(new_n2871), .B1(new_n675), .B2(new_n2881), .C(new_n4741), .Y(new_n4742));
  AOI21xp33_ASAP7_75t_L     g04486(.A1(new_n674), .A2(\b[27] ), .B(new_n4742), .Y(new_n4743));
  NAND2xp33_ASAP7_75t_L     g04487(.A(\a[11] ), .B(new_n4743), .Y(new_n4744));
  A2O1A1Ixp33_ASAP7_75t_L   g04488(.A1(\b[27] ), .A2(new_n674), .B(new_n4742), .C(new_n594), .Y(new_n4745));
  NAND2xp33_ASAP7_75t_L     g04489(.A(new_n4745), .B(new_n4744), .Y(new_n4746));
  AOI32xp33_ASAP7_75t_L     g04490(.A1(new_n2483), .A2(new_n2486), .A3(new_n823), .B1(new_n826), .B2(\b[26] ), .Y(new_n4747));
  OAI221xp5_ASAP7_75t_L     g04491(.A1(new_n994), .A2(new_n2180), .B1(new_n2019), .B2(new_n909), .C(new_n4747), .Y(new_n4748));
  XNOR2x2_ASAP7_75t_L       g04492(.A(\a[14] ), .B(new_n4748), .Y(new_n4749));
  NOR3xp33_ASAP7_75t_L      g04493(.A(new_n4630), .B(new_n4631), .C(new_n4643), .Y(new_n4750));
  INVx1_ASAP7_75t_L         g04494(.A(new_n4750), .Y(new_n4751));
  OAI21xp33_ASAP7_75t_L     g04495(.A1(new_n4586), .A2(new_n4596), .B(new_n4598), .Y(new_n4752));
  NAND2xp33_ASAP7_75t_L     g04496(.A(\b[12] ), .B(new_n2386), .Y(new_n4753));
  NAND2xp33_ASAP7_75t_L     g04497(.A(\b[13] ), .B(new_n2232), .Y(new_n4754));
  AOI32xp33_ASAP7_75t_L     g04498(.A1(new_n877), .A2(new_n874), .A3(new_n2226), .B1(\b[14] ), .B2(new_n2228), .Y(new_n4755));
  AND4x1_ASAP7_75t_L        g04499(.A(new_n4755), .B(new_n4754), .C(new_n4753), .D(\a[26] ), .Y(new_n4756));
  AOI31xp33_ASAP7_75t_L     g04500(.A1(new_n4755), .A2(new_n4754), .A3(new_n4753), .B(\a[26] ), .Y(new_n4757));
  NOR2xp33_ASAP7_75t_L      g04501(.A(new_n4757), .B(new_n4756), .Y(new_n4758));
  A2O1A1O1Ixp25_ASAP7_75t_L g04502(.A1(new_n4299), .A2(new_n4343), .B(new_n4346), .C(new_n4574), .D(new_n4584), .Y(new_n4759));
  NAND2xp33_ASAP7_75t_L     g04503(.A(\b[9] ), .B(new_n2931), .Y(new_n4760));
  NAND2xp33_ASAP7_75t_L     g04504(.A(\b[10] ), .B(new_n2706), .Y(new_n4761));
  AOI32xp33_ASAP7_75t_L     g04505(.A1(new_n700), .A2(new_n698), .A3(new_n2700), .B1(\b[11] ), .B2(new_n2702), .Y(new_n4762));
  AND4x1_ASAP7_75t_L        g04506(.A(new_n4762), .B(new_n4761), .C(new_n4760), .D(\a[29] ), .Y(new_n4763));
  AOI31xp33_ASAP7_75t_L     g04507(.A1(new_n4762), .A2(new_n4761), .A3(new_n4760), .B(\a[29] ), .Y(new_n4764));
  OR2x4_ASAP7_75t_L         g04508(.A(new_n4764), .B(new_n4763), .Y(new_n4765));
  A2O1A1O1Ixp25_ASAP7_75t_L g04509(.A1(new_n4334), .A2(new_n4332), .B(new_n4511), .C(new_n4571), .D(new_n4569), .Y(new_n4766));
  NOR2xp33_ASAP7_75t_L      g04510(.A(new_n382), .B(new_n3492), .Y(new_n4767));
  NAND2xp33_ASAP7_75t_L     g04511(.A(\b[7] ), .B(new_n3260), .Y(new_n4768));
  OAI221xp5_ASAP7_75t_L     g04512(.A1(new_n3262), .A2(new_n503), .B1(new_n3261), .B2(new_n509), .C(new_n4768), .Y(new_n4769));
  OR3x1_ASAP7_75t_L         g04513(.A(new_n4769), .B(new_n3251), .C(new_n4767), .Y(new_n4770));
  A2O1A1Ixp33_ASAP7_75t_L   g04514(.A1(\b[6] ), .A2(new_n3491), .B(new_n4769), .C(new_n3251), .Y(new_n4771));
  A2O1A1O1Ixp25_ASAP7_75t_L g04515(.A1(new_n4524), .A2(new_n4305), .B(new_n4327), .C(new_n4566), .D(new_n4558), .Y(new_n4772));
  NAND2xp33_ASAP7_75t_L     g04516(.A(\b[3] ), .B(new_n4111), .Y(new_n4773));
  NAND2xp33_ASAP7_75t_L     g04517(.A(\b[4] ), .B(new_n3874), .Y(new_n4774));
  AOI22xp33_ASAP7_75t_L     g04518(.A1(new_n3884), .A2(\b[5] ), .B1(new_n3881), .B2(new_n360), .Y(new_n4775));
  NAND4xp25_ASAP7_75t_L     g04519(.A(new_n4775), .B(\a[35] ), .C(new_n4773), .D(new_n4774), .Y(new_n4776));
  OAI221xp5_ASAP7_75t_L     g04520(.A1(new_n4115), .A2(new_n353), .B1(new_n4114), .B2(new_n359), .C(new_n4774), .Y(new_n4777));
  A2O1A1Ixp33_ASAP7_75t_L   g04521(.A1(\b[3] ), .A2(new_n4111), .B(new_n4777), .C(new_n3878), .Y(new_n4778));
  A2O1A1O1Ixp25_ASAP7_75t_L g04522(.A1(new_n4534), .A2(new_n4304), .B(new_n258), .C(new_n4545), .D(new_n4539), .Y(new_n4779));
  NOR3xp33_ASAP7_75t_L      g04523(.A(new_n4541), .B(new_n4535), .C(new_n4547), .Y(new_n4780));
  INVx1_ASAP7_75t_L         g04524(.A(new_n4780), .Y(new_n4781));
  NOR2xp33_ASAP7_75t_L      g04525(.A(new_n258), .B(new_n4781), .Y(new_n4782));
  NAND2xp33_ASAP7_75t_L     g04526(.A(\b[1] ), .B(new_n4548), .Y(new_n4783));
  OAI221xp5_ASAP7_75t_L     g04527(.A1(new_n4549), .A2(new_n283), .B1(new_n278), .B2(new_n4550), .C(new_n4783), .Y(new_n4784));
  OR3x1_ASAP7_75t_L         g04528(.A(new_n4779), .B(new_n4782), .C(new_n4784), .Y(new_n4785));
  A2O1A1Ixp33_ASAP7_75t_L   g04529(.A1(\b[0] ), .A2(new_n4780), .B(new_n4784), .C(new_n4779), .Y(new_n4786));
  NAND4xp25_ASAP7_75t_L     g04530(.A(new_n4776), .B(new_n4785), .C(new_n4778), .D(new_n4786), .Y(new_n4787));
  AO22x1_ASAP7_75t_L        g04531(.A1(new_n4786), .A2(new_n4785), .B1(new_n4778), .B2(new_n4776), .Y(new_n4788));
  AOI21xp33_ASAP7_75t_L     g04532(.A1(new_n4788), .A2(new_n4787), .B(new_n4772), .Y(new_n4789));
  A2O1A1Ixp33_ASAP7_75t_L   g04533(.A1(new_n4317), .A2(new_n4561), .B(new_n4554), .C(new_n4567), .Y(new_n4790));
  NAND2xp33_ASAP7_75t_L     g04534(.A(new_n4787), .B(new_n4788), .Y(new_n4791));
  NOR2xp33_ASAP7_75t_L      g04535(.A(new_n4790), .B(new_n4791), .Y(new_n4792));
  AOI211xp5_ASAP7_75t_L     g04536(.A1(new_n4770), .A2(new_n4771), .B(new_n4789), .C(new_n4792), .Y(new_n4793));
  NOR3xp33_ASAP7_75t_L      g04537(.A(new_n4769), .B(new_n4767), .C(new_n3251), .Y(new_n4794));
  OA21x2_ASAP7_75t_L        g04538(.A1(new_n4767), .A2(new_n4769), .B(new_n3251), .Y(new_n4795));
  NAND2xp33_ASAP7_75t_L     g04539(.A(new_n4790), .B(new_n4791), .Y(new_n4796));
  NAND3xp33_ASAP7_75t_L     g04540(.A(new_n4772), .B(new_n4787), .C(new_n4788), .Y(new_n4797));
  AOI211xp5_ASAP7_75t_L     g04541(.A1(new_n4796), .A2(new_n4797), .B(new_n4795), .C(new_n4794), .Y(new_n4798));
  NOR3xp33_ASAP7_75t_L      g04542(.A(new_n4766), .B(new_n4793), .C(new_n4798), .Y(new_n4799));
  OAI211xp5_ASAP7_75t_L     g04543(.A1(new_n4794), .A2(new_n4795), .B(new_n4796), .C(new_n4797), .Y(new_n4800));
  OAI211xp5_ASAP7_75t_L     g04544(.A1(new_n4789), .A2(new_n4792), .B(new_n4771), .C(new_n4770), .Y(new_n4801));
  AOI221xp5_ASAP7_75t_L     g04545(.A1(new_n4576), .A2(new_n4571), .B1(new_n4800), .B2(new_n4801), .C(new_n4569), .Y(new_n4802));
  OAI21xp33_ASAP7_75t_L     g04546(.A1(new_n4802), .A2(new_n4799), .B(new_n4765), .Y(new_n4803));
  NOR2xp33_ASAP7_75t_L      g04547(.A(new_n4764), .B(new_n4763), .Y(new_n4804));
  A2O1A1Ixp33_ASAP7_75t_L   g04548(.A1(new_n4516), .A2(new_n4512), .B(new_n4563), .C(new_n4572), .Y(new_n4805));
  NAND3xp33_ASAP7_75t_L     g04549(.A(new_n4805), .B(new_n4800), .C(new_n4801), .Y(new_n4806));
  OAI21xp33_ASAP7_75t_L     g04550(.A1(new_n4793), .A2(new_n4798), .B(new_n4766), .Y(new_n4807));
  NAND3xp33_ASAP7_75t_L     g04551(.A(new_n4806), .B(new_n4804), .C(new_n4807), .Y(new_n4808));
  AOI21xp33_ASAP7_75t_L     g04552(.A1(new_n4808), .A2(new_n4803), .B(new_n4759), .Y(new_n4809));
  OAI21xp33_ASAP7_75t_L     g04553(.A1(new_n4583), .A2(new_n4582), .B(new_n4580), .Y(new_n4810));
  NAND2xp33_ASAP7_75t_L     g04554(.A(new_n4803), .B(new_n4808), .Y(new_n4811));
  NOR2xp33_ASAP7_75t_L      g04555(.A(new_n4810), .B(new_n4811), .Y(new_n4812));
  OAI21xp33_ASAP7_75t_L     g04556(.A1(new_n4809), .A2(new_n4812), .B(new_n4758), .Y(new_n4813));
  AOI21xp33_ASAP7_75t_L     g04557(.A1(new_n4806), .A2(new_n4807), .B(new_n4804), .Y(new_n4814));
  NOR3xp33_ASAP7_75t_L      g04558(.A(new_n4765), .B(new_n4799), .C(new_n4802), .Y(new_n4815));
  OAI21xp33_ASAP7_75t_L     g04559(.A1(new_n4814), .A2(new_n4815), .B(new_n4810), .Y(new_n4816));
  NAND3xp33_ASAP7_75t_L     g04560(.A(new_n4759), .B(new_n4803), .C(new_n4808), .Y(new_n4817));
  OAI211xp5_ASAP7_75t_L     g04561(.A1(new_n4757), .A2(new_n4756), .B(new_n4816), .C(new_n4817), .Y(new_n4818));
  NAND3xp33_ASAP7_75t_L     g04562(.A(new_n4752), .B(new_n4813), .C(new_n4818), .Y(new_n4819));
  A2O1A1O1Ixp25_ASAP7_75t_L g04563(.A1(new_n4357), .A2(new_n4371), .B(new_n4368), .C(new_n4597), .D(new_n4590), .Y(new_n4820));
  AOI211xp5_ASAP7_75t_L     g04564(.A1(new_n4816), .A2(new_n4817), .B(new_n4757), .C(new_n4756), .Y(new_n4821));
  NOR3xp33_ASAP7_75t_L      g04565(.A(new_n4812), .B(new_n4809), .C(new_n4758), .Y(new_n4822));
  OAI21xp33_ASAP7_75t_L     g04566(.A1(new_n4821), .A2(new_n4822), .B(new_n4820), .Y(new_n4823));
  NAND2xp33_ASAP7_75t_L     g04567(.A(\b[15] ), .B(new_n1910), .Y(new_n4824));
  NAND2xp33_ASAP7_75t_L     g04568(.A(\b[16] ), .B(new_n1770), .Y(new_n4825));
  AOI32xp33_ASAP7_75t_L     g04569(.A1(new_n1250), .A2(new_n1247), .A3(new_n1764), .B1(\b[17] ), .B2(new_n1766), .Y(new_n4826));
  NAND4xp25_ASAP7_75t_L     g04570(.A(new_n4826), .B(\a[23] ), .C(new_n4824), .D(new_n4825), .Y(new_n4827));
  INVx1_ASAP7_75t_L         g04571(.A(new_n4827), .Y(new_n4828));
  AOI31xp33_ASAP7_75t_L     g04572(.A1(new_n4826), .A2(new_n4825), .A3(new_n4824), .B(\a[23] ), .Y(new_n4829));
  NOR2xp33_ASAP7_75t_L      g04573(.A(new_n4829), .B(new_n4828), .Y(new_n4830));
  NAND3xp33_ASAP7_75t_L     g04574(.A(new_n4819), .B(new_n4823), .C(new_n4830), .Y(new_n4831));
  NOR3xp33_ASAP7_75t_L      g04575(.A(new_n4820), .B(new_n4821), .C(new_n4822), .Y(new_n4832));
  AOI21xp33_ASAP7_75t_L     g04576(.A1(new_n4818), .A2(new_n4813), .B(new_n4752), .Y(new_n4833));
  INVx1_ASAP7_75t_L         g04577(.A(new_n4830), .Y(new_n4834));
  OAI21xp33_ASAP7_75t_L     g04578(.A1(new_n4832), .A2(new_n4833), .B(new_n4834), .Y(new_n4835));
  NOR2xp33_ASAP7_75t_L      g04579(.A(new_n4605), .B(new_n4607), .Y(new_n4836));
  MAJIxp5_ASAP7_75t_L       g04580(.A(new_n4616), .B(new_n4608), .C(new_n4836), .Y(new_n4837));
  NAND3xp33_ASAP7_75t_L     g04581(.A(new_n4837), .B(new_n4835), .C(new_n4831), .Y(new_n4838));
  NAND2xp33_ASAP7_75t_L     g04582(.A(new_n4831), .B(new_n4835), .Y(new_n4839));
  NAND2xp33_ASAP7_75t_L     g04583(.A(new_n4600), .B(new_n4592), .Y(new_n4840));
  MAJIxp5_ASAP7_75t_L       g04584(.A(new_n4611), .B(new_n4840), .C(new_n4603), .Y(new_n4841));
  NAND2xp33_ASAP7_75t_L     g04585(.A(new_n4839), .B(new_n4841), .Y(new_n4842));
  NOR2xp33_ASAP7_75t_L      g04586(.A(new_n1594), .B(new_n1412), .Y(new_n4843));
  AOI221xp5_ASAP7_75t_L     g04587(.A1(new_n1410), .A2(\b[19] ), .B1(new_n1404), .B2(new_n1600), .C(new_n4843), .Y(new_n4844));
  OAI211xp5_ASAP7_75t_L     g04588(.A1(new_n1356), .A2(new_n1549), .B(new_n4844), .C(\a[20] ), .Y(new_n4845));
  O2A1O1Ixp33_ASAP7_75t_L   g04589(.A1(new_n1356), .A2(new_n1549), .B(new_n4844), .C(\a[20] ), .Y(new_n4846));
  INVx1_ASAP7_75t_L         g04590(.A(new_n4846), .Y(new_n4847));
  AND4x1_ASAP7_75t_L        g04591(.A(new_n4842), .B(new_n4838), .C(new_n4847), .D(new_n4845), .Y(new_n4848));
  INVx1_ASAP7_75t_L         g04592(.A(new_n4845), .Y(new_n4849));
  NOR2xp33_ASAP7_75t_L      g04593(.A(new_n4846), .B(new_n4849), .Y(new_n4850));
  AOI21xp33_ASAP7_75t_L     g04594(.A1(new_n4838), .A2(new_n4842), .B(new_n4850), .Y(new_n4851));
  NAND3xp33_ASAP7_75t_L     g04595(.A(new_n4612), .B(new_n4617), .C(new_n4626), .Y(new_n4852));
  A2O1A1Ixp33_ASAP7_75t_L   g04596(.A1(new_n4627), .A2(new_n4623), .B(new_n4629), .C(new_n4852), .Y(new_n4853));
  NOR3xp33_ASAP7_75t_L      g04597(.A(new_n4853), .B(new_n4851), .C(new_n4848), .Y(new_n4854));
  OA21x2_ASAP7_75t_L        g04598(.A1(new_n4848), .A2(new_n4851), .B(new_n4853), .Y(new_n4855));
  NAND2xp33_ASAP7_75t_L     g04599(.A(\b[21] ), .B(new_n1194), .Y(new_n4856));
  NAND2xp33_ASAP7_75t_L     g04600(.A(\b[22] ), .B(new_n1103), .Y(new_n4857));
  AOI22xp33_ASAP7_75t_L     g04601(.A1(new_n1113), .A2(\b[23] ), .B1(new_n1110), .B2(new_n2002), .Y(new_n4858));
  NAND4xp25_ASAP7_75t_L     g04602(.A(new_n4858), .B(\a[17] ), .C(new_n4856), .D(new_n4857), .Y(new_n4859));
  NAND2xp33_ASAP7_75t_L     g04603(.A(new_n2001), .B(new_n1998), .Y(new_n4860));
  OAI221xp5_ASAP7_75t_L     g04604(.A1(new_n1198), .A2(new_n1995), .B1(new_n1197), .B2(new_n4860), .C(new_n4857), .Y(new_n4861));
  A2O1A1Ixp33_ASAP7_75t_L   g04605(.A1(\b[21] ), .A2(new_n1194), .B(new_n4861), .C(new_n1107), .Y(new_n4862));
  AND2x2_ASAP7_75t_L        g04606(.A(new_n4862), .B(new_n4859), .Y(new_n4863));
  OAI21xp33_ASAP7_75t_L     g04607(.A1(new_n4854), .A2(new_n4855), .B(new_n4863), .Y(new_n4864));
  NOR3xp33_ASAP7_75t_L      g04608(.A(new_n4855), .B(new_n4863), .C(new_n4854), .Y(new_n4865));
  INVx1_ASAP7_75t_L         g04609(.A(new_n4865), .Y(new_n4866));
  NAND4xp25_ASAP7_75t_L     g04610(.A(new_n4652), .B(new_n4866), .C(new_n4864), .D(new_n4751), .Y(new_n4867));
  XNOR2x2_ASAP7_75t_L       g04611(.A(new_n4837), .B(new_n4839), .Y(new_n4868));
  NAND2xp33_ASAP7_75t_L     g04612(.A(new_n4850), .B(new_n4868), .Y(new_n4869));
  NAND2xp33_ASAP7_75t_L     g04613(.A(new_n4842), .B(new_n4838), .Y(new_n4870));
  NAND2xp33_ASAP7_75t_L     g04614(.A(new_n4845), .B(new_n4847), .Y(new_n4871));
  NAND2xp33_ASAP7_75t_L     g04615(.A(new_n4871), .B(new_n4870), .Y(new_n4872));
  NAND4xp25_ASAP7_75t_L     g04616(.A(new_n4642), .B(new_n4852), .C(new_n4872), .D(new_n4869), .Y(new_n4873));
  OAI21xp33_ASAP7_75t_L     g04617(.A1(new_n4848), .A2(new_n4851), .B(new_n4853), .Y(new_n4874));
  NAND2xp33_ASAP7_75t_L     g04618(.A(new_n4862), .B(new_n4859), .Y(new_n4875));
  AOI21xp33_ASAP7_75t_L     g04619(.A1(new_n4873), .A2(new_n4874), .B(new_n4875), .Y(new_n4876));
  OAI22xp33_ASAP7_75t_L     g04620(.A1(new_n4661), .A2(new_n4750), .B1(new_n4865), .B2(new_n4876), .Y(new_n4877));
  NAND3xp33_ASAP7_75t_L     g04621(.A(new_n4867), .B(new_n4877), .C(new_n4749), .Y(new_n4878));
  INVx1_ASAP7_75t_L         g04622(.A(new_n4749), .Y(new_n4879));
  A2O1A1Ixp33_ASAP7_75t_L   g04623(.A1(new_n4646), .A2(new_n4414), .B(new_n4645), .C(new_n4751), .Y(new_n4880));
  NOR3xp33_ASAP7_75t_L      g04624(.A(new_n4880), .B(new_n4876), .C(new_n4865), .Y(new_n4881));
  NOR2xp33_ASAP7_75t_L      g04625(.A(new_n4876), .B(new_n4865), .Y(new_n4882));
  A2O1A1O1Ixp25_ASAP7_75t_L g04626(.A1(new_n4414), .A2(new_n4646), .B(new_n4645), .C(new_n4751), .D(new_n4882), .Y(new_n4883));
  OAI21xp33_ASAP7_75t_L     g04627(.A1(new_n4881), .A2(new_n4883), .B(new_n4879), .Y(new_n4884));
  O2A1O1Ixp33_ASAP7_75t_L   g04628(.A1(new_n4426), .A2(new_n4429), .B(new_n4428), .C(new_n4659), .Y(new_n4885));
  OAI211xp5_ASAP7_75t_L     g04629(.A1(new_n4663), .A2(new_n4885), .B(new_n4884), .C(new_n4878), .Y(new_n4886));
  NOR3xp33_ASAP7_75t_L      g04630(.A(new_n4883), .B(new_n4881), .C(new_n4879), .Y(new_n4887));
  AOI21xp33_ASAP7_75t_L     g04631(.A1(new_n4867), .A2(new_n4877), .B(new_n4749), .Y(new_n4888));
  A2O1A1O1Ixp25_ASAP7_75t_L g04632(.A1(new_n4427), .A2(new_n4666), .B(new_n4423), .C(new_n4667), .D(new_n4663), .Y(new_n4889));
  OAI21xp33_ASAP7_75t_L     g04633(.A1(new_n4887), .A2(new_n4888), .B(new_n4889), .Y(new_n4890));
  AO21x2_ASAP7_75t_L        g04634(.A1(new_n4886), .A2(new_n4890), .B(new_n4746), .Y(new_n4891));
  NAND3xp33_ASAP7_75t_L     g04635(.A(new_n4890), .B(new_n4886), .C(new_n4746), .Y(new_n4892));
  NAND2xp33_ASAP7_75t_L     g04636(.A(new_n4892), .B(new_n4891), .Y(new_n4893));
  O2A1O1Ixp33_ASAP7_75t_L   g04637(.A1(new_n4679), .A2(new_n4680), .B(new_n4676), .C(new_n4893), .Y(new_n4894));
  OAI21xp33_ASAP7_75t_L     g04638(.A1(new_n4680), .A2(new_n4679), .B(new_n4676), .Y(new_n4895));
  AOI21xp33_ASAP7_75t_L     g04639(.A1(new_n4892), .A2(new_n4891), .B(new_n4895), .Y(new_n4896));
  OAI21xp33_ASAP7_75t_L     g04640(.A1(new_n4894), .A2(new_n4896), .B(new_n4740), .Y(new_n4897));
  OR3x1_ASAP7_75t_L         g04641(.A(new_n4896), .B(new_n4894), .C(new_n4740), .Y(new_n4898));
  NAND2xp33_ASAP7_75t_L     g04642(.A(new_n4897), .B(new_n4898), .Y(new_n4899));
  O2A1O1Ixp33_ASAP7_75t_L   g04643(.A1(new_n4483), .A2(new_n4683), .B(new_n4732), .C(new_n4899), .Y(new_n4900));
  AO21x2_ASAP7_75t_L        g04644(.A1(new_n4677), .A2(new_n4682), .B(new_n4486), .Y(new_n4901));
  A2O1A1O1Ixp25_ASAP7_75t_L g04645(.A1(new_n4451), .A2(new_n4270), .B(new_n4450), .C(new_n4901), .D(new_n4684), .Y(new_n4902));
  INVx1_ASAP7_75t_L         g04646(.A(new_n4902), .Y(new_n4903));
  OA21x2_ASAP7_75t_L        g04647(.A1(new_n4894), .A2(new_n4896), .B(new_n4740), .Y(new_n4904));
  NOR3xp33_ASAP7_75t_L      g04648(.A(new_n4896), .B(new_n4894), .C(new_n4740), .Y(new_n4905));
  NOR2xp33_ASAP7_75t_L      g04649(.A(new_n4905), .B(new_n4904), .Y(new_n4906));
  NOR2xp33_ASAP7_75t_L      g04650(.A(new_n4903), .B(new_n4906), .Y(new_n4907));
  OAI21xp33_ASAP7_75t_L     g04651(.A1(new_n4907), .A2(new_n4900), .B(new_n4731), .Y(new_n4908));
  NAND2xp33_ASAP7_75t_L     g04652(.A(new_n4903), .B(new_n4906), .Y(new_n4909));
  NAND2xp33_ASAP7_75t_L     g04653(.A(new_n4902), .B(new_n4899), .Y(new_n4910));
  NAND3xp33_ASAP7_75t_L     g04654(.A(new_n4910), .B(new_n4730), .C(new_n4909), .Y(new_n4911));
  NAND2xp33_ASAP7_75t_L     g04655(.A(new_n4911), .B(new_n4908), .Y(new_n4912));
  XNOR2x2_ASAP7_75t_L       g04656(.A(new_n4724), .B(new_n4912), .Y(new_n4913));
  NOR2xp33_ASAP7_75t_L      g04657(.A(\b[37] ), .B(\b[38] ), .Y(new_n4914));
  INVx1_ASAP7_75t_L         g04658(.A(\b[38] ), .Y(new_n4915));
  NOR2xp33_ASAP7_75t_L      g04659(.A(new_n4701), .B(new_n4915), .Y(new_n4916));
  NOR2xp33_ASAP7_75t_L      g04660(.A(new_n4914), .B(new_n4916), .Y(new_n4917));
  A2O1A1Ixp33_ASAP7_75t_L   g04661(.A1(new_n4707), .A2(new_n4703), .B(new_n4702), .C(new_n4917), .Y(new_n4918));
  INVx1_ASAP7_75t_L         g04662(.A(new_n4918), .Y(new_n4919));
  O2A1O1Ixp33_ASAP7_75t_L   g04663(.A1(new_n4466), .A2(new_n4469), .B(new_n4703), .C(new_n4702), .Y(new_n4920));
  INVx1_ASAP7_75t_L         g04664(.A(new_n4920), .Y(new_n4921));
  NOR2xp33_ASAP7_75t_L      g04665(.A(new_n4917), .B(new_n4921), .Y(new_n4922));
  NOR2xp33_ASAP7_75t_L      g04666(.A(new_n4922), .B(new_n4919), .Y(new_n4923));
  AOI22xp33_ASAP7_75t_L     g04667(.A1(new_n272), .A2(\b[38] ), .B1(new_n269), .B2(new_n4923), .Y(new_n4924));
  OAI221xp5_ASAP7_75t_L     g04668(.A1(new_n261), .A2(new_n4701), .B1(new_n4465), .B2(new_n277), .C(new_n4924), .Y(new_n4925));
  XNOR2x2_ASAP7_75t_L       g04669(.A(new_n265), .B(new_n4925), .Y(new_n4926));
  XNOR2x2_ASAP7_75t_L       g04670(.A(new_n4926), .B(new_n4913), .Y(new_n4927));
  O2A1O1Ixp33_ASAP7_75t_L   g04671(.A1(new_n4723), .A2(new_n4718), .B(new_n4717), .C(new_n4927), .Y(new_n4928));
  INVx1_ASAP7_75t_L         g04672(.A(new_n4927), .Y(new_n4929));
  AO21x2_ASAP7_75t_L        g04673(.A1(new_n4715), .A2(new_n4720), .B(new_n4716), .Y(new_n4930));
  NOR2xp33_ASAP7_75t_L      g04674(.A(new_n4930), .B(new_n4929), .Y(new_n4931));
  NOR2xp33_ASAP7_75t_L      g04675(.A(new_n4928), .B(new_n4931), .Y(\f[38] ));
  NOR3xp33_ASAP7_75t_L      g04676(.A(new_n4900), .B(new_n4907), .C(new_n4731), .Y(new_n4933));
  AOI21xp33_ASAP7_75t_L     g04677(.A1(new_n4724), .A2(new_n4908), .B(new_n4933), .Y(new_n4934));
  NAND2xp33_ASAP7_75t_L     g04678(.A(\b[34] ), .B(new_n366), .Y(new_n4935));
  NAND2xp33_ASAP7_75t_L     g04679(.A(\b[35] ), .B(new_n334), .Y(new_n4936));
  AOI22xp33_ASAP7_75t_L     g04680(.A1(new_n345), .A2(\b[36] ), .B1(new_n342), .B2(new_n4473), .Y(new_n4937));
  AND4x1_ASAP7_75t_L        g04681(.A(new_n4937), .B(new_n4936), .C(new_n4935), .D(\a[5] ), .Y(new_n4938));
  AOI31xp33_ASAP7_75t_L     g04682(.A1(new_n4937), .A2(new_n4936), .A3(new_n4935), .B(\a[5] ), .Y(new_n4939));
  NOR2xp33_ASAP7_75t_L      g04683(.A(new_n4939), .B(new_n4938), .Y(new_n4940));
  OAI21xp33_ASAP7_75t_L     g04684(.A1(new_n4904), .A2(new_n4902), .B(new_n4898), .Y(new_n4941));
  A2O1A1O1Ixp25_ASAP7_75t_L g04685(.A1(new_n4279), .A2(new_n4442), .B(new_n4487), .C(new_n4671), .D(new_n4681), .Y(new_n4942));
  AOI21xp33_ASAP7_75t_L     g04686(.A1(new_n4890), .A2(new_n4886), .B(new_n4746), .Y(new_n4943));
  OAI21xp33_ASAP7_75t_L     g04687(.A1(new_n4943), .A2(new_n4942), .B(new_n4892), .Y(new_n4944));
  NOR2xp33_ASAP7_75t_L      g04688(.A(new_n2852), .B(new_n1620), .Y(new_n4945));
  INVx1_ASAP7_75t_L         g04689(.A(new_n4945), .Y(new_n4946));
  NOR2xp33_ASAP7_75t_L      g04690(.A(new_n2871), .B(new_n721), .Y(new_n4947));
  INVx1_ASAP7_75t_L         g04691(.A(new_n4947), .Y(new_n4948));
  AOI22xp33_ASAP7_75t_L     g04692(.A1(new_n600), .A2(\b[30] ), .B1(new_n597), .B2(new_n3219), .Y(new_n4949));
  AND4x1_ASAP7_75t_L        g04693(.A(new_n4949), .B(new_n4948), .C(new_n4946), .D(\a[11] ), .Y(new_n4950));
  AOI31xp33_ASAP7_75t_L     g04694(.A1(new_n4949), .A2(new_n4948), .A3(new_n4946), .B(\a[11] ), .Y(new_n4951));
  NOR2xp33_ASAP7_75t_L      g04695(.A(new_n4951), .B(new_n4950), .Y(new_n4952));
  INVx1_ASAP7_75t_L         g04696(.A(new_n4952), .Y(new_n4953));
  INVx1_ASAP7_75t_L         g04697(.A(new_n4889), .Y(new_n4954));
  NAND2xp33_ASAP7_75t_L     g04698(.A(new_n4823), .B(new_n4819), .Y(new_n4955));
  NOR2xp33_ASAP7_75t_L      g04699(.A(new_n4830), .B(new_n4955), .Y(new_n4956));
  NAND2xp33_ASAP7_75t_L     g04700(.A(\b[16] ), .B(new_n1910), .Y(new_n4957));
  NAND2xp33_ASAP7_75t_L     g04701(.A(\b[17] ), .B(new_n1770), .Y(new_n4958));
  AOI22xp33_ASAP7_75t_L     g04702(.A1(new_n1766), .A2(\b[18] ), .B1(new_n1764), .B2(new_n1363), .Y(new_n4959));
  NAND4xp25_ASAP7_75t_L     g04703(.A(new_n4959), .B(\a[23] ), .C(new_n4957), .D(new_n4958), .Y(new_n4960));
  OAI221xp5_ASAP7_75t_L     g04704(.A1(new_n1772), .A2(new_n1356), .B1(new_n1771), .B2(new_n3138), .C(new_n4958), .Y(new_n4961));
  A2O1A1Ixp33_ASAP7_75t_L   g04705(.A1(\b[16] ), .A2(new_n1910), .B(new_n4961), .C(new_n1761), .Y(new_n4962));
  NAND2xp33_ASAP7_75t_L     g04706(.A(new_n4960), .B(new_n4962), .Y(new_n4963));
  OAI21xp33_ASAP7_75t_L     g04707(.A1(new_n4821), .A2(new_n4820), .B(new_n4818), .Y(new_n4964));
  NAND2xp33_ASAP7_75t_L     g04708(.A(\b[0] ), .B(new_n4548), .Y(new_n4965));
  NAND4xp25_ASAP7_75t_L     g04709(.A(new_n4545), .B(\a[38] ), .C(new_n4310), .D(new_n4965), .Y(new_n4966));
  INVx1_ASAP7_75t_L         g04710(.A(\a[39] ), .Y(new_n4967));
  NAND2xp33_ASAP7_75t_L     g04711(.A(\a[38] ), .B(new_n4967), .Y(new_n4968));
  NAND2xp33_ASAP7_75t_L     g04712(.A(\a[39] ), .B(new_n4539), .Y(new_n4969));
  AND2x2_ASAP7_75t_L        g04713(.A(new_n4968), .B(new_n4969), .Y(new_n4970));
  NOR2xp33_ASAP7_75t_L      g04714(.A(new_n258), .B(new_n4970), .Y(new_n4971));
  OAI31xp33_ASAP7_75t_L     g04715(.A1(new_n4966), .A2(new_n4784), .A3(new_n4782), .B(new_n4971), .Y(new_n4972));
  OR4x2_ASAP7_75t_L         g04716(.A(new_n4971), .B(new_n4966), .C(new_n4784), .D(new_n4782), .Y(new_n4973));
  NOR2xp33_ASAP7_75t_L      g04717(.A(new_n278), .B(new_n4536), .Y(new_n4974));
  AOI221xp5_ASAP7_75t_L     g04718(.A1(new_n4544), .A2(\b[3] ), .B1(new_n4542), .B2(new_n1000), .C(new_n4974), .Y(new_n4975));
  OAI211xp5_ASAP7_75t_L     g04719(.A1(new_n276), .A2(new_n4781), .B(new_n4975), .C(\a[38] ), .Y(new_n4976));
  NAND2xp33_ASAP7_75t_L     g04720(.A(\b[3] ), .B(new_n4544), .Y(new_n4977));
  OAI221xp5_ASAP7_75t_L     g04721(.A1(new_n278), .A2(new_n4536), .B1(new_n4549), .B2(new_n303), .C(new_n4977), .Y(new_n4978));
  A2O1A1Ixp33_ASAP7_75t_L   g04722(.A1(\b[1] ), .A2(new_n4780), .B(new_n4978), .C(new_n4539), .Y(new_n4979));
  AOI22xp33_ASAP7_75t_L     g04723(.A1(new_n4976), .A2(new_n4979), .B1(new_n4972), .B2(new_n4973), .Y(new_n4980));
  OA31x2_ASAP7_75t_L        g04724(.A1(new_n4782), .A2(new_n4784), .A3(new_n4966), .B1(new_n4971), .Y(new_n4981));
  NOR4xp25_ASAP7_75t_L      g04725(.A(new_n4966), .B(new_n4971), .C(new_n4784), .D(new_n4782), .Y(new_n4982));
  AOI211xp5_ASAP7_75t_L     g04726(.A1(\b[1] ), .A2(new_n4780), .B(new_n4539), .C(new_n4978), .Y(new_n4983));
  O2A1O1Ixp33_ASAP7_75t_L   g04727(.A1(new_n276), .A2(new_n4781), .B(new_n4975), .C(\a[38] ), .Y(new_n4984));
  NOR4xp25_ASAP7_75t_L      g04728(.A(new_n4981), .B(new_n4984), .C(new_n4983), .D(new_n4982), .Y(new_n4985));
  INVx1_ASAP7_75t_L         g04729(.A(new_n4111), .Y(new_n4986));
  NOR2xp33_ASAP7_75t_L      g04730(.A(new_n323), .B(new_n4986), .Y(new_n4987));
  NAND2xp33_ASAP7_75t_L     g04731(.A(\b[5] ), .B(new_n3874), .Y(new_n4988));
  NAND2xp33_ASAP7_75t_L     g04732(.A(\b[6] ), .B(new_n3884), .Y(new_n4989));
  OAI311xp33_ASAP7_75t_L    g04733(.A1(new_n388), .A2(new_n386), .A3(new_n4114), .B1(new_n4989), .C1(new_n4988), .Y(new_n4990));
  NOR3xp33_ASAP7_75t_L      g04734(.A(new_n4990), .B(new_n4987), .C(new_n3878), .Y(new_n4991));
  A2O1A1Ixp33_ASAP7_75t_L   g04735(.A1(\b[4] ), .A2(new_n4111), .B(new_n4990), .C(new_n3878), .Y(new_n4992));
  INVx1_ASAP7_75t_L         g04736(.A(new_n4992), .Y(new_n4993));
  NOR4xp25_ASAP7_75t_L      g04737(.A(new_n4980), .B(new_n4985), .C(new_n4993), .D(new_n4991), .Y(new_n4994));
  OAI22xp33_ASAP7_75t_L     g04738(.A1(new_n4981), .A2(new_n4982), .B1(new_n4984), .B2(new_n4983), .Y(new_n4995));
  NAND4xp25_ASAP7_75t_L     g04739(.A(new_n4973), .B(new_n4972), .C(new_n4976), .D(new_n4979), .Y(new_n4996));
  INVx1_ASAP7_75t_L         g04740(.A(new_n4991), .Y(new_n4997));
  AOI22xp33_ASAP7_75t_L     g04741(.A1(new_n4997), .A2(new_n4992), .B1(new_n4996), .B2(new_n4995), .Y(new_n4998));
  NOR2xp33_ASAP7_75t_L      g04742(.A(new_n4998), .B(new_n4994), .Y(new_n4999));
  NAND2xp33_ASAP7_75t_L     g04743(.A(new_n4778), .B(new_n4776), .Y(new_n5000));
  NOR2xp33_ASAP7_75t_L      g04744(.A(new_n4549), .B(new_n283), .Y(new_n5001));
  AOI221xp5_ASAP7_75t_L     g04745(.A1(\b[2] ), .A2(new_n4544), .B1(new_n4548), .B2(\b[1] ), .C(new_n5001), .Y(new_n5002));
  OAI21xp33_ASAP7_75t_L     g04746(.A1(new_n258), .A2(new_n4781), .B(new_n5002), .Y(new_n5003));
  NOR2xp33_ASAP7_75t_L      g04747(.A(new_n4779), .B(new_n5003), .Y(new_n5004));
  INVx1_ASAP7_75t_L         g04748(.A(new_n4786), .Y(new_n5005));
  NOR2xp33_ASAP7_75t_L      g04749(.A(new_n5004), .B(new_n5005), .Y(new_n5006));
  MAJIxp5_ASAP7_75t_L       g04750(.A(new_n4790), .B(new_n5000), .C(new_n5006), .Y(new_n5007));
  NAND2xp33_ASAP7_75t_L     g04751(.A(new_n4999), .B(new_n5007), .Y(new_n5008));
  NAND4xp25_ASAP7_75t_L     g04752(.A(new_n4996), .B(new_n4995), .C(new_n4997), .D(new_n4992), .Y(new_n5009));
  OAI22xp33_ASAP7_75t_L     g04753(.A1(new_n4980), .A2(new_n4985), .B1(new_n4993), .B2(new_n4991), .Y(new_n5010));
  NAND2xp33_ASAP7_75t_L     g04754(.A(new_n5009), .B(new_n5010), .Y(new_n5011));
  A2O1A1Ixp33_ASAP7_75t_L   g04755(.A1(new_n5006), .A2(new_n5000), .B(new_n4789), .C(new_n5011), .Y(new_n5012));
  NOR2xp33_ASAP7_75t_L      g04756(.A(new_n421), .B(new_n3492), .Y(new_n5013));
  INVx1_ASAP7_75t_L         g04757(.A(new_n5013), .Y(new_n5014));
  NAND2xp33_ASAP7_75t_L     g04758(.A(\b[8] ), .B(new_n3260), .Y(new_n5015));
  AOI32xp33_ASAP7_75t_L     g04759(.A1(new_n765), .A2(new_n977), .A3(new_n3254), .B1(new_n3256), .B2(\b[9] ), .Y(new_n5016));
  NAND4xp25_ASAP7_75t_L     g04760(.A(new_n5016), .B(\a[32] ), .C(new_n5014), .D(new_n5015), .Y(new_n5017));
  AOI31xp33_ASAP7_75t_L     g04761(.A1(new_n5016), .A2(new_n5015), .A3(new_n5014), .B(\a[32] ), .Y(new_n5018));
  INVx1_ASAP7_75t_L         g04762(.A(new_n5018), .Y(new_n5019));
  NAND4xp25_ASAP7_75t_L     g04763(.A(new_n5008), .B(new_n5012), .C(new_n5019), .D(new_n5017), .Y(new_n5020));
  NAND2xp33_ASAP7_75t_L     g04764(.A(new_n5000), .B(new_n5006), .Y(new_n5021));
  A2O1A1Ixp33_ASAP7_75t_L   g04765(.A1(new_n4787), .A2(new_n4788), .B(new_n4772), .C(new_n5021), .Y(new_n5022));
  NOR2xp33_ASAP7_75t_L      g04766(.A(new_n5011), .B(new_n5022), .Y(new_n5023));
  NOR2xp33_ASAP7_75t_L      g04767(.A(new_n4999), .B(new_n5007), .Y(new_n5024));
  INVx1_ASAP7_75t_L         g04768(.A(new_n5017), .Y(new_n5025));
  OAI22xp33_ASAP7_75t_L     g04769(.A1(new_n5024), .A2(new_n5023), .B1(new_n5018), .B2(new_n5025), .Y(new_n5026));
  NAND2xp33_ASAP7_75t_L     g04770(.A(new_n5020), .B(new_n5026), .Y(new_n5027));
  OAI21xp33_ASAP7_75t_L     g04771(.A1(new_n4798), .A2(new_n4766), .B(new_n4800), .Y(new_n5028));
  NOR2xp33_ASAP7_75t_L      g04772(.A(new_n5028), .B(new_n5027), .Y(new_n5029));
  A2O1A1O1Ixp25_ASAP7_75t_L g04773(.A1(new_n4571), .A2(new_n4576), .B(new_n4569), .C(new_n4801), .D(new_n4793), .Y(new_n5030));
  AOI21xp33_ASAP7_75t_L     g04774(.A1(new_n5026), .A2(new_n5020), .B(new_n5030), .Y(new_n5031));
  NAND2xp33_ASAP7_75t_L     g04775(.A(\b[10] ), .B(new_n2931), .Y(new_n5032));
  NAND2xp33_ASAP7_75t_L     g04776(.A(\b[11] ), .B(new_n2706), .Y(new_n5033));
  AOI32xp33_ASAP7_75t_L     g04777(.A1(new_n771), .A2(new_n774), .A3(new_n2700), .B1(new_n2702), .B2(\b[12] ), .Y(new_n5034));
  AND4x1_ASAP7_75t_L        g04778(.A(new_n5034), .B(new_n5033), .C(new_n5032), .D(\a[29] ), .Y(new_n5035));
  AOI31xp33_ASAP7_75t_L     g04779(.A1(new_n5034), .A2(new_n5033), .A3(new_n5032), .B(\a[29] ), .Y(new_n5036));
  NOR2xp33_ASAP7_75t_L      g04780(.A(new_n5036), .B(new_n5035), .Y(new_n5037));
  OAI21xp33_ASAP7_75t_L     g04781(.A1(new_n5031), .A2(new_n5029), .B(new_n5037), .Y(new_n5038));
  NAND3xp33_ASAP7_75t_L     g04782(.A(new_n5030), .B(new_n5026), .C(new_n5020), .Y(new_n5039));
  NOR4xp25_ASAP7_75t_L      g04783(.A(new_n5024), .B(new_n5023), .C(new_n5018), .D(new_n5025), .Y(new_n5040));
  NOR2xp33_ASAP7_75t_L      g04784(.A(new_n5018), .B(new_n5025), .Y(new_n5041));
  AOI21xp33_ASAP7_75t_L     g04785(.A1(new_n5012), .A2(new_n5008), .B(new_n5041), .Y(new_n5042));
  OAI21xp33_ASAP7_75t_L     g04786(.A1(new_n5040), .A2(new_n5042), .B(new_n5028), .Y(new_n5043));
  OAI211xp5_ASAP7_75t_L     g04787(.A1(new_n5035), .A2(new_n5036), .B(new_n5043), .C(new_n5039), .Y(new_n5044));
  NAND3xp33_ASAP7_75t_L     g04788(.A(new_n4806), .B(new_n4765), .C(new_n4807), .Y(new_n5045));
  A2O1A1Ixp33_ASAP7_75t_L   g04789(.A1(new_n4803), .A2(new_n4808), .B(new_n4759), .C(new_n5045), .Y(new_n5046));
  NAND3xp33_ASAP7_75t_L     g04790(.A(new_n5046), .B(new_n5044), .C(new_n5038), .Y(new_n5047));
  NAND2xp33_ASAP7_75t_L     g04791(.A(new_n5044), .B(new_n5038), .Y(new_n5048));
  INVx1_ASAP7_75t_L         g04792(.A(new_n5045), .Y(new_n5049));
  O2A1O1Ixp33_ASAP7_75t_L   g04793(.A1(new_n4814), .A2(new_n4815), .B(new_n4810), .C(new_n5049), .Y(new_n5050));
  NAND2xp33_ASAP7_75t_L     g04794(.A(new_n5050), .B(new_n5048), .Y(new_n5051));
  NAND2xp33_ASAP7_75t_L     g04795(.A(\b[13] ), .B(new_n2386), .Y(new_n5052));
  NAND2xp33_ASAP7_75t_L     g04796(.A(\b[14] ), .B(new_n2232), .Y(new_n5053));
  AOI22xp33_ASAP7_75t_L     g04797(.A1(new_n2228), .A2(\b[15] ), .B1(new_n2226), .B2(new_n959), .Y(new_n5054));
  NAND4xp25_ASAP7_75t_L     g04798(.A(new_n5054), .B(\a[26] ), .C(new_n5052), .D(new_n5053), .Y(new_n5055));
  OAI221xp5_ASAP7_75t_L     g04799(.A1(new_n2234), .A2(new_n952), .B1(new_n2233), .B2(new_n2573), .C(new_n5053), .Y(new_n5056));
  A2O1A1Ixp33_ASAP7_75t_L   g04800(.A1(\b[13] ), .A2(new_n2386), .B(new_n5056), .C(new_n2223), .Y(new_n5057));
  AND2x2_ASAP7_75t_L        g04801(.A(new_n5055), .B(new_n5057), .Y(new_n5058));
  AND3x1_ASAP7_75t_L        g04802(.A(new_n5058), .B(new_n5051), .C(new_n5047), .Y(new_n5059));
  AOI21xp33_ASAP7_75t_L     g04803(.A1(new_n5051), .A2(new_n5047), .B(new_n5058), .Y(new_n5060));
  OAI21xp33_ASAP7_75t_L     g04804(.A1(new_n5059), .A2(new_n5060), .B(new_n4964), .Y(new_n5061));
  A2O1A1O1Ixp25_ASAP7_75t_L g04805(.A1(new_n4597), .A2(new_n4606), .B(new_n4590), .C(new_n4813), .D(new_n4822), .Y(new_n5062));
  NAND3xp33_ASAP7_75t_L     g04806(.A(new_n5058), .B(new_n5051), .C(new_n5047), .Y(new_n5063));
  AO21x2_ASAP7_75t_L        g04807(.A1(new_n5047), .A2(new_n5051), .B(new_n5058), .Y(new_n5064));
  NAND3xp33_ASAP7_75t_L     g04808(.A(new_n5062), .B(new_n5063), .C(new_n5064), .Y(new_n5065));
  NAND3xp33_ASAP7_75t_L     g04809(.A(new_n5065), .B(new_n5061), .C(new_n4963), .Y(new_n5066));
  AND2x2_ASAP7_75t_L        g04810(.A(new_n4960), .B(new_n4962), .Y(new_n5067));
  AOI21xp33_ASAP7_75t_L     g04811(.A1(new_n5064), .A2(new_n5063), .B(new_n5062), .Y(new_n5068));
  NOR3xp33_ASAP7_75t_L      g04812(.A(new_n4964), .B(new_n5059), .C(new_n5060), .Y(new_n5069));
  OAI21xp33_ASAP7_75t_L     g04813(.A1(new_n5068), .A2(new_n5069), .B(new_n5067), .Y(new_n5070));
  AO221x2_ASAP7_75t_L       g04814(.A1(new_n4841), .A2(new_n4839), .B1(new_n5066), .B2(new_n5070), .C(new_n4956), .Y(new_n5071));
  AOI21xp33_ASAP7_75t_L     g04815(.A1(new_n4835), .A2(new_n4831), .B(new_n4837), .Y(new_n5072));
  NOR3xp33_ASAP7_75t_L      g04816(.A(new_n5069), .B(new_n5067), .C(new_n5068), .Y(new_n5073));
  AOI21xp33_ASAP7_75t_L     g04817(.A1(new_n5065), .A2(new_n5061), .B(new_n4963), .Y(new_n5074));
  NOR2xp33_ASAP7_75t_L      g04818(.A(new_n5074), .B(new_n5073), .Y(new_n5075));
  OAI21xp33_ASAP7_75t_L     g04819(.A1(new_n4956), .A2(new_n5072), .B(new_n5075), .Y(new_n5076));
  NAND2xp33_ASAP7_75t_L     g04820(.A(\b[19] ), .B(new_n1548), .Y(new_n5077));
  NAND2xp33_ASAP7_75t_L     g04821(.A(\b[20] ), .B(new_n1410), .Y(new_n5078));
  AOI22xp33_ASAP7_75t_L     g04822(.A1(new_n1406), .A2(\b[21] ), .B1(new_n1404), .B2(new_n1715), .Y(new_n5079));
  AND4x1_ASAP7_75t_L        g04823(.A(new_n5079), .B(new_n5078), .C(new_n5077), .D(\a[20] ), .Y(new_n5080));
  AOI31xp33_ASAP7_75t_L     g04824(.A1(new_n5079), .A2(new_n5078), .A3(new_n5077), .B(\a[20] ), .Y(new_n5081));
  NOR2xp33_ASAP7_75t_L      g04825(.A(new_n5081), .B(new_n5080), .Y(new_n5082));
  NAND3xp33_ASAP7_75t_L     g04826(.A(new_n5076), .B(new_n5071), .C(new_n5082), .Y(new_n5083));
  AOI221xp5_ASAP7_75t_L     g04827(.A1(new_n4841), .A2(new_n4839), .B1(new_n5066), .B2(new_n5070), .C(new_n4956), .Y(new_n5084));
  INVx1_ASAP7_75t_L         g04828(.A(new_n4956), .Y(new_n5085));
  NAND2xp33_ASAP7_75t_L     g04829(.A(new_n5066), .B(new_n5070), .Y(new_n5086));
  AOI21xp33_ASAP7_75t_L     g04830(.A1(new_n4842), .A2(new_n5085), .B(new_n5086), .Y(new_n5087));
  INVx1_ASAP7_75t_L         g04831(.A(new_n5082), .Y(new_n5088));
  OAI21xp33_ASAP7_75t_L     g04832(.A1(new_n5084), .A2(new_n5087), .B(new_n5088), .Y(new_n5089));
  NAND2xp33_ASAP7_75t_L     g04833(.A(new_n5083), .B(new_n5089), .Y(new_n5090));
  NOR2xp33_ASAP7_75t_L      g04834(.A(new_n4850), .B(new_n4870), .Y(new_n5091));
  NOR3xp33_ASAP7_75t_L      g04835(.A(new_n4855), .B(new_n5090), .C(new_n5091), .Y(new_n5092));
  MAJIxp5_ASAP7_75t_L       g04836(.A(new_n4853), .B(new_n4868), .C(new_n4871), .Y(new_n5093));
  AOI21xp33_ASAP7_75t_L     g04837(.A1(new_n5089), .A2(new_n5083), .B(new_n5093), .Y(new_n5094));
  NAND2xp33_ASAP7_75t_L     g04838(.A(\b[22] ), .B(new_n1194), .Y(new_n5095));
  NAND2xp33_ASAP7_75t_L     g04839(.A(\b[23] ), .B(new_n1103), .Y(new_n5096));
  AOI22xp33_ASAP7_75t_L     g04840(.A1(new_n1113), .A2(\b[24] ), .B1(new_n1110), .B2(new_n2027), .Y(new_n5097));
  NAND4xp25_ASAP7_75t_L     g04841(.A(new_n5097), .B(\a[17] ), .C(new_n5095), .D(new_n5096), .Y(new_n5098));
  NAND2xp33_ASAP7_75t_L     g04842(.A(new_n5096), .B(new_n5097), .Y(new_n5099));
  A2O1A1Ixp33_ASAP7_75t_L   g04843(.A1(\b[22] ), .A2(new_n1194), .B(new_n5099), .C(new_n1107), .Y(new_n5100));
  AND2x2_ASAP7_75t_L        g04844(.A(new_n5098), .B(new_n5100), .Y(new_n5101));
  OAI21xp33_ASAP7_75t_L     g04845(.A1(new_n5094), .A2(new_n5092), .B(new_n5101), .Y(new_n5102));
  NAND3xp33_ASAP7_75t_L     g04846(.A(new_n5093), .B(new_n5089), .C(new_n5083), .Y(new_n5103));
  NAND2xp33_ASAP7_75t_L     g04847(.A(new_n4869), .B(new_n4872), .Y(new_n5104));
  A2O1A1Ixp33_ASAP7_75t_L   g04848(.A1(new_n5104), .A2(new_n4853), .B(new_n5091), .C(new_n5090), .Y(new_n5105));
  NAND2xp33_ASAP7_75t_L     g04849(.A(new_n5098), .B(new_n5100), .Y(new_n5106));
  NAND3xp33_ASAP7_75t_L     g04850(.A(new_n5105), .B(new_n5103), .C(new_n5106), .Y(new_n5107));
  A2O1A1O1Ixp25_ASAP7_75t_L g04851(.A1(new_n4414), .A2(new_n4646), .B(new_n4645), .C(new_n4751), .D(new_n4876), .Y(new_n5108));
  OAI211xp5_ASAP7_75t_L     g04852(.A1(new_n4865), .A2(new_n5108), .B(new_n5102), .C(new_n5107), .Y(new_n5109));
  AOI21xp33_ASAP7_75t_L     g04853(.A1(new_n5105), .A2(new_n5103), .B(new_n5106), .Y(new_n5110));
  NOR3xp33_ASAP7_75t_L      g04854(.A(new_n5092), .B(new_n5101), .C(new_n5094), .Y(new_n5111));
  A2O1A1O1Ixp25_ASAP7_75t_L g04855(.A1(new_n4651), .A2(new_n4650), .B(new_n4750), .C(new_n4864), .D(new_n4865), .Y(new_n5112));
  OAI21xp33_ASAP7_75t_L     g04856(.A1(new_n5110), .A2(new_n5111), .B(new_n5112), .Y(new_n5113));
  NAND2xp33_ASAP7_75t_L     g04857(.A(\b[25] ), .B(new_n908), .Y(new_n5114));
  NAND2xp33_ASAP7_75t_L     g04858(.A(\b[26] ), .B(new_n817), .Y(new_n5115));
  NOR2xp33_ASAP7_75t_L      g04859(.A(new_n2650), .B(new_n912), .Y(new_n5116));
  AOI21xp33_ASAP7_75t_L     g04860(.A1(new_n2657), .A2(new_n823), .B(new_n5116), .Y(new_n5117));
  NAND4xp25_ASAP7_75t_L     g04861(.A(new_n5117), .B(\a[14] ), .C(new_n5114), .D(new_n5115), .Y(new_n5118));
  NAND2xp33_ASAP7_75t_L     g04862(.A(new_n5115), .B(new_n5117), .Y(new_n5119));
  A2O1A1Ixp33_ASAP7_75t_L   g04863(.A1(\b[25] ), .A2(new_n908), .B(new_n5119), .C(new_n813), .Y(new_n5120));
  AND2x2_ASAP7_75t_L        g04864(.A(new_n5118), .B(new_n5120), .Y(new_n5121));
  NAND3xp33_ASAP7_75t_L     g04865(.A(new_n5109), .B(new_n5121), .C(new_n5113), .Y(new_n5122));
  NOR3xp33_ASAP7_75t_L      g04866(.A(new_n5112), .B(new_n5111), .C(new_n5110), .Y(new_n5123));
  AOI211xp5_ASAP7_75t_L     g04867(.A1(new_n5102), .A2(new_n5107), .B(new_n4865), .C(new_n5108), .Y(new_n5124));
  NAND2xp33_ASAP7_75t_L     g04868(.A(new_n5118), .B(new_n5120), .Y(new_n5125));
  OAI21xp33_ASAP7_75t_L     g04869(.A1(new_n5123), .A2(new_n5124), .B(new_n5125), .Y(new_n5126));
  NAND2xp33_ASAP7_75t_L     g04870(.A(new_n5126), .B(new_n5122), .Y(new_n5127));
  A2O1A1Ixp33_ASAP7_75t_L   g04871(.A1(new_n4954), .A2(new_n4878), .B(new_n4888), .C(new_n5127), .Y(new_n5128));
  A2O1A1O1Ixp25_ASAP7_75t_L g04872(.A1(new_n4667), .A2(new_n4673), .B(new_n4663), .C(new_n4878), .D(new_n4888), .Y(new_n5129));
  AND2x2_ASAP7_75t_L        g04873(.A(new_n5126), .B(new_n5122), .Y(new_n5130));
  NAND2xp33_ASAP7_75t_L     g04874(.A(new_n5129), .B(new_n5130), .Y(new_n5131));
  NAND3xp33_ASAP7_75t_L     g04875(.A(new_n5131), .B(new_n5128), .C(new_n4953), .Y(new_n5132));
  O2A1O1Ixp33_ASAP7_75t_L   g04876(.A1(new_n4887), .A2(new_n4889), .B(new_n4884), .C(new_n5130), .Y(new_n5133));
  A2O1A1Ixp33_ASAP7_75t_L   g04877(.A1(new_n4666), .A2(new_n4424), .B(new_n4423), .C(new_n4667), .Y(new_n5134));
  A2O1A1Ixp33_ASAP7_75t_L   g04878(.A1(new_n5134), .A2(new_n4668), .B(new_n4887), .C(new_n4884), .Y(new_n5135));
  NOR2xp33_ASAP7_75t_L      g04879(.A(new_n5127), .B(new_n5135), .Y(new_n5136));
  OAI21xp33_ASAP7_75t_L     g04880(.A1(new_n5136), .A2(new_n5133), .B(new_n4952), .Y(new_n5137));
  NAND3xp33_ASAP7_75t_L     g04881(.A(new_n4944), .B(new_n5132), .C(new_n5137), .Y(new_n5138));
  AND3x1_ASAP7_75t_L        g04882(.A(new_n4890), .B(new_n4746), .C(new_n4886), .Y(new_n5139));
  A2O1A1O1Ixp25_ASAP7_75t_L g04883(.A1(new_n4671), .A2(new_n4489), .B(new_n4681), .C(new_n4891), .D(new_n5139), .Y(new_n5140));
  NOR3xp33_ASAP7_75t_L      g04884(.A(new_n5133), .B(new_n5136), .C(new_n4952), .Y(new_n5141));
  AOI21xp33_ASAP7_75t_L     g04885(.A1(new_n5131), .A2(new_n5128), .B(new_n4953), .Y(new_n5142));
  OAI21xp33_ASAP7_75t_L     g04886(.A1(new_n5142), .A2(new_n5141), .B(new_n5140), .Y(new_n5143));
  NAND2xp33_ASAP7_75t_L     g04887(.A(\b[31] ), .B(new_n480), .Y(new_n5144));
  NAND2xp33_ASAP7_75t_L     g04888(.A(\b[32] ), .B(new_n441), .Y(new_n5145));
  AOI22xp33_ASAP7_75t_L     g04889(.A1(new_n451), .A2(\b[33] ), .B1(new_n448), .B2(new_n3813), .Y(new_n5146));
  NAND4xp25_ASAP7_75t_L     g04890(.A(new_n5146), .B(\a[8] ), .C(new_n5144), .D(new_n5145), .Y(new_n5147));
  NAND2xp33_ASAP7_75t_L     g04891(.A(new_n5145), .B(new_n5146), .Y(new_n5148));
  A2O1A1Ixp33_ASAP7_75t_L   g04892(.A1(\b[31] ), .A2(new_n480), .B(new_n5148), .C(new_n445), .Y(new_n5149));
  AND2x2_ASAP7_75t_L        g04893(.A(new_n5147), .B(new_n5149), .Y(new_n5150));
  NAND3xp33_ASAP7_75t_L     g04894(.A(new_n5138), .B(new_n5150), .C(new_n5143), .Y(new_n5151));
  NOR3xp33_ASAP7_75t_L      g04895(.A(new_n5140), .B(new_n5141), .C(new_n5142), .Y(new_n5152));
  AOI21xp33_ASAP7_75t_L     g04896(.A1(new_n5137), .A2(new_n5132), .B(new_n4944), .Y(new_n5153));
  NAND2xp33_ASAP7_75t_L     g04897(.A(new_n5147), .B(new_n5149), .Y(new_n5154));
  OAI21xp33_ASAP7_75t_L     g04898(.A1(new_n5152), .A2(new_n5153), .B(new_n5154), .Y(new_n5155));
  NAND2xp33_ASAP7_75t_L     g04899(.A(new_n5151), .B(new_n5155), .Y(new_n5156));
  AND2x2_ASAP7_75t_L        g04900(.A(new_n5156), .B(new_n4941), .Y(new_n5157));
  NOR2xp33_ASAP7_75t_L      g04901(.A(new_n5156), .B(new_n4941), .Y(new_n5158));
  OAI21xp33_ASAP7_75t_L     g04902(.A1(new_n5158), .A2(new_n5157), .B(new_n4940), .Y(new_n5159));
  NOR3xp33_ASAP7_75t_L      g04903(.A(new_n5157), .B(new_n5158), .C(new_n4940), .Y(new_n5160));
  INVx1_ASAP7_75t_L         g04904(.A(new_n5160), .Y(new_n5161));
  NAND2xp33_ASAP7_75t_L     g04905(.A(new_n5159), .B(new_n5161), .Y(new_n5162));
  XNOR2x2_ASAP7_75t_L       g04906(.A(new_n4934), .B(new_n5162), .Y(new_n5163));
  INVx1_ASAP7_75t_L         g04907(.A(new_n4916), .Y(new_n5164));
  NOR2xp33_ASAP7_75t_L      g04908(.A(\b[38] ), .B(\b[39] ), .Y(new_n5165));
  INVx1_ASAP7_75t_L         g04909(.A(\b[39] ), .Y(new_n5166));
  NOR2xp33_ASAP7_75t_L      g04910(.A(new_n4915), .B(new_n5166), .Y(new_n5167));
  NOR2xp33_ASAP7_75t_L      g04911(.A(new_n5165), .B(new_n5167), .Y(new_n5168));
  INVx1_ASAP7_75t_L         g04912(.A(new_n5168), .Y(new_n5169));
  O2A1O1Ixp33_ASAP7_75t_L   g04913(.A1(new_n4914), .A2(new_n4920), .B(new_n5164), .C(new_n5169), .Y(new_n5170));
  INVx1_ASAP7_75t_L         g04914(.A(new_n4702), .Y(new_n5171));
  A2O1A1Ixp33_ASAP7_75t_L   g04915(.A1(new_n4704), .A2(new_n5171), .B(new_n4914), .C(new_n5164), .Y(new_n5172));
  NOR2xp33_ASAP7_75t_L      g04916(.A(new_n5168), .B(new_n5172), .Y(new_n5173));
  NOR2xp33_ASAP7_75t_L      g04917(.A(new_n5170), .B(new_n5173), .Y(new_n5174));
  AOI22xp33_ASAP7_75t_L     g04918(.A1(new_n272), .A2(\b[39] ), .B1(new_n269), .B2(new_n5174), .Y(new_n5175));
  OAI221xp5_ASAP7_75t_L     g04919(.A1(new_n261), .A2(new_n4915), .B1(new_n4701), .B2(new_n277), .C(new_n5175), .Y(new_n5176));
  XNOR2x2_ASAP7_75t_L       g04920(.A(\a[2] ), .B(new_n5176), .Y(new_n5177));
  XOR2x2_ASAP7_75t_L        g04921(.A(new_n5177), .B(new_n5163), .Y(new_n5178));
  MAJIxp5_ASAP7_75t_L       g04922(.A(new_n4930), .B(new_n4913), .C(new_n4926), .Y(new_n5179));
  XNOR2x2_ASAP7_75t_L       g04923(.A(new_n5179), .B(new_n5178), .Y(\f[39] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04924(.A1(new_n4926), .A2(new_n4913), .B(new_n4928), .C(new_n5178), .Y(new_n5181));
  NOR2xp33_ASAP7_75t_L      g04925(.A(new_n4915), .B(new_n277), .Y(new_n5182));
  INVx1_ASAP7_75t_L         g04926(.A(new_n5182), .Y(new_n5183));
  NAND2xp33_ASAP7_75t_L     g04927(.A(\b[39] ), .B(new_n380), .Y(new_n5184));
  NOR2xp33_ASAP7_75t_L      g04928(.A(\b[39] ), .B(\b[40] ), .Y(new_n5185));
  INVx1_ASAP7_75t_L         g04929(.A(\b[40] ), .Y(new_n5186));
  NOR2xp33_ASAP7_75t_L      g04930(.A(new_n5166), .B(new_n5186), .Y(new_n5187));
  NOR2xp33_ASAP7_75t_L      g04931(.A(new_n5185), .B(new_n5187), .Y(new_n5188));
  A2O1A1Ixp33_ASAP7_75t_L   g04932(.A1(new_n5172), .A2(new_n5168), .B(new_n5167), .C(new_n5188), .Y(new_n5189));
  INVx1_ASAP7_75t_L         g04933(.A(new_n5189), .Y(new_n5190));
  INVx1_ASAP7_75t_L         g04934(.A(new_n5167), .Y(new_n5191));
  A2O1A1Ixp33_ASAP7_75t_L   g04935(.A1(new_n4918), .A2(new_n5164), .B(new_n5165), .C(new_n5191), .Y(new_n5192));
  NOR2xp33_ASAP7_75t_L      g04936(.A(new_n5188), .B(new_n5192), .Y(new_n5193));
  NOR2xp33_ASAP7_75t_L      g04937(.A(new_n5190), .B(new_n5193), .Y(new_n5194));
  AOI22xp33_ASAP7_75t_L     g04938(.A1(new_n272), .A2(\b[40] ), .B1(new_n269), .B2(new_n5194), .Y(new_n5195));
  AND4x1_ASAP7_75t_L        g04939(.A(new_n5195), .B(new_n5184), .C(new_n5183), .D(\a[2] ), .Y(new_n5196));
  AOI31xp33_ASAP7_75t_L     g04940(.A1(new_n5195), .A2(new_n5184), .A3(new_n5183), .B(\a[2] ), .Y(new_n5197));
  NOR2xp33_ASAP7_75t_L      g04941(.A(new_n5197), .B(new_n5196), .Y(new_n5198));
  A2O1A1O1Ixp25_ASAP7_75t_L g04942(.A1(new_n4908), .A2(new_n4724), .B(new_n4933), .C(new_n5159), .D(new_n5160), .Y(new_n5199));
  NOR3xp33_ASAP7_75t_L      g04943(.A(new_n5153), .B(new_n5152), .C(new_n5150), .Y(new_n5200));
  NAND2xp33_ASAP7_75t_L     g04944(.A(\b[32] ), .B(new_n480), .Y(new_n5201));
  NAND2xp33_ASAP7_75t_L     g04945(.A(\b[33] ), .B(new_n441), .Y(new_n5202));
  AOI22xp33_ASAP7_75t_L     g04946(.A1(new_n451), .A2(\b[34] ), .B1(new_n448), .B2(new_n3833), .Y(new_n5203));
  NAND4xp25_ASAP7_75t_L     g04947(.A(new_n5203), .B(\a[8] ), .C(new_n5201), .D(new_n5202), .Y(new_n5204));
  NAND2xp33_ASAP7_75t_L     g04948(.A(new_n5202), .B(new_n5203), .Y(new_n5205));
  A2O1A1Ixp33_ASAP7_75t_L   g04949(.A1(\b[32] ), .A2(new_n480), .B(new_n5205), .C(new_n445), .Y(new_n5206));
  NAND2xp33_ASAP7_75t_L     g04950(.A(new_n5204), .B(new_n5206), .Y(new_n5207));
  OAI21xp33_ASAP7_75t_L     g04951(.A1(new_n5142), .A2(new_n5140), .B(new_n5132), .Y(new_n5208));
  NAND3xp33_ASAP7_75t_L     g04952(.A(new_n5109), .B(new_n5113), .C(new_n5125), .Y(new_n5209));
  A2O1A1Ixp33_ASAP7_75t_L   g04953(.A1(new_n5122), .A2(new_n5126), .B(new_n5129), .C(new_n5209), .Y(new_n5210));
  NOR2xp33_ASAP7_75t_L      g04954(.A(new_n2477), .B(new_n909), .Y(new_n5211));
  NAND2xp33_ASAP7_75t_L     g04955(.A(new_n2855), .B(new_n2857), .Y(new_n5212));
  NAND2xp33_ASAP7_75t_L     g04956(.A(\b[27] ), .B(new_n817), .Y(new_n5213));
  OAI221xp5_ASAP7_75t_L     g04957(.A1(new_n912), .A2(new_n2852), .B1(new_n911), .B2(new_n5212), .C(new_n5213), .Y(new_n5214));
  OR3x1_ASAP7_75t_L         g04958(.A(new_n5214), .B(new_n813), .C(new_n5211), .Y(new_n5215));
  A2O1A1Ixp33_ASAP7_75t_L   g04959(.A1(\b[26] ), .A2(new_n908), .B(new_n5214), .C(new_n813), .Y(new_n5216));
  AND2x2_ASAP7_75t_L        g04960(.A(new_n5216), .B(new_n5215), .Y(new_n5217));
  AOI211xp5_ASAP7_75t_L     g04961(.A1(new_n5043), .A2(new_n5039), .B(new_n5035), .C(new_n5036), .Y(new_n5218));
  A2O1A1Ixp33_ASAP7_75t_L   g04962(.A1(new_n4816), .A2(new_n5045), .B(new_n5218), .C(new_n5044), .Y(new_n5219));
  NOR2xp33_ASAP7_75t_L      g04963(.A(new_n695), .B(new_n2932), .Y(new_n5220));
  INVx1_ASAP7_75t_L         g04964(.A(new_n5220), .Y(new_n5221));
  NAND2xp33_ASAP7_75t_L     g04965(.A(\b[12] ), .B(new_n2706), .Y(new_n5222));
  AOI22xp33_ASAP7_75t_L     g04966(.A1(new_n2702), .A2(\b[13] ), .B1(new_n2700), .B2(new_n800), .Y(new_n5223));
  AND4x1_ASAP7_75t_L        g04967(.A(new_n5223), .B(new_n5222), .C(new_n5221), .D(\a[29] ), .Y(new_n5224));
  AOI31xp33_ASAP7_75t_L     g04968(.A1(new_n5223), .A2(new_n5222), .A3(new_n5221), .B(\a[29] ), .Y(new_n5225));
  NOR2xp33_ASAP7_75t_L      g04969(.A(new_n5225), .B(new_n5224), .Y(new_n5226));
  OAI211xp5_ASAP7_75t_L     g04970(.A1(new_n5025), .A2(new_n5018), .B(new_n5008), .C(new_n5012), .Y(new_n5227));
  INVx1_ASAP7_75t_L         g04971(.A(new_n4971), .Y(new_n5228));
  NOR3xp33_ASAP7_75t_L      g04972(.A(new_n5003), .B(new_n5228), .C(new_n4966), .Y(new_n5229));
  NAND2xp33_ASAP7_75t_L     g04973(.A(\b[2] ), .B(new_n4780), .Y(new_n5230));
  INVx1_ASAP7_75t_L         g04974(.A(new_n5230), .Y(new_n5231));
  NOR2xp33_ASAP7_75t_L      g04975(.A(new_n299), .B(new_n4536), .Y(new_n5232));
  OAI32xp33_ASAP7_75t_L     g04976(.A1(new_n325), .A2(new_n327), .A3(new_n4549), .B1(new_n323), .B2(new_n4550), .Y(new_n5233));
  NOR4xp25_ASAP7_75t_L      g04977(.A(new_n5231), .B(new_n5233), .C(new_n4539), .D(new_n5232), .Y(new_n5234));
  INVx1_ASAP7_75t_L         g04978(.A(new_n5234), .Y(new_n5235));
  OAI31xp33_ASAP7_75t_L     g04979(.A1(new_n5231), .A2(new_n5233), .A3(new_n5232), .B(new_n4539), .Y(new_n5236));
  NAND2xp33_ASAP7_75t_L     g04980(.A(\a[41] ), .B(new_n4971), .Y(new_n5237));
  NAND2xp33_ASAP7_75t_L     g04981(.A(new_n4969), .B(new_n4968), .Y(new_n5238));
  XNOR2x2_ASAP7_75t_L       g04982(.A(\a[40] ), .B(\a[39] ), .Y(new_n5239));
  NOR2xp33_ASAP7_75t_L      g04983(.A(new_n5239), .B(new_n5238), .Y(new_n5240));
  INVx1_ASAP7_75t_L         g04984(.A(new_n5240), .Y(new_n5241));
  INVx1_ASAP7_75t_L         g04985(.A(\a[40] ), .Y(new_n5242));
  NAND2xp33_ASAP7_75t_L     g04986(.A(\a[41] ), .B(new_n5242), .Y(new_n5243));
  INVx1_ASAP7_75t_L         g04987(.A(\a[41] ), .Y(new_n5244));
  NAND2xp33_ASAP7_75t_L     g04988(.A(\a[40] ), .B(new_n5244), .Y(new_n5245));
  AND2x2_ASAP7_75t_L        g04989(.A(new_n5243), .B(new_n5245), .Y(new_n5246));
  NOR2xp33_ASAP7_75t_L      g04990(.A(new_n4970), .B(new_n5246), .Y(new_n5247));
  NAND2xp33_ASAP7_75t_L     g04991(.A(new_n5245), .B(new_n5243), .Y(new_n5248));
  NOR2xp33_ASAP7_75t_L      g04992(.A(new_n5248), .B(new_n4970), .Y(new_n5249));
  AOI22xp33_ASAP7_75t_L     g04993(.A1(new_n5249), .A2(\b[1] ), .B1(new_n271), .B2(new_n5247), .Y(new_n5250));
  O2A1O1Ixp33_ASAP7_75t_L   g04994(.A1(new_n5241), .A2(new_n258), .B(new_n5250), .C(new_n5237), .Y(new_n5251));
  NAND2xp33_ASAP7_75t_L     g04995(.A(new_n5248), .B(new_n5238), .Y(new_n5252));
  NAND2xp33_ASAP7_75t_L     g04996(.A(new_n5238), .B(new_n5246), .Y(new_n5253));
  OAI22xp33_ASAP7_75t_L     g04997(.A1(new_n5253), .A2(new_n276), .B1(new_n270), .B2(new_n5252), .Y(new_n5254));
  A2O1A1O1Ixp25_ASAP7_75t_L g04998(.A1(new_n5238), .A2(\a[41] ), .B(new_n5240), .C(\b[0] ), .D(new_n5254), .Y(new_n5255));
  OR2x4_ASAP7_75t_L         g04999(.A(new_n5255), .B(new_n5251), .Y(new_n5256));
  NAND3xp33_ASAP7_75t_L     g05000(.A(new_n5256), .B(new_n5235), .C(new_n5236), .Y(new_n5257));
  INVx1_ASAP7_75t_L         g05001(.A(new_n5236), .Y(new_n5258));
  NOR2xp33_ASAP7_75t_L      g05002(.A(new_n5255), .B(new_n5251), .Y(new_n5259));
  OAI21xp33_ASAP7_75t_L     g05003(.A1(new_n5234), .A2(new_n5258), .B(new_n5259), .Y(new_n5260));
  OAI211xp5_ASAP7_75t_L     g05004(.A1(new_n5229), .A2(new_n4980), .B(new_n5257), .C(new_n5260), .Y(new_n5261));
  INVx1_ASAP7_75t_L         g05005(.A(new_n5229), .Y(new_n5262));
  NOR3xp33_ASAP7_75t_L      g05006(.A(new_n5258), .B(new_n5259), .C(new_n5234), .Y(new_n5263));
  AOI21xp33_ASAP7_75t_L     g05007(.A1(new_n5236), .A2(new_n5235), .B(new_n5256), .Y(new_n5264));
  OAI211xp5_ASAP7_75t_L     g05008(.A1(new_n5264), .A2(new_n5263), .B(new_n5262), .C(new_n4995), .Y(new_n5265));
  NAND2xp33_ASAP7_75t_L     g05009(.A(\b[5] ), .B(new_n4111), .Y(new_n5266));
  NAND2xp33_ASAP7_75t_L     g05010(.A(\b[6] ), .B(new_n3874), .Y(new_n5267));
  AOI32xp33_ASAP7_75t_L     g05011(.A1(new_n424), .A2(new_n426), .A3(new_n3881), .B1(new_n3884), .B2(\b[7] ), .Y(new_n5268));
  NAND4xp25_ASAP7_75t_L     g05012(.A(new_n5268), .B(\a[35] ), .C(new_n5266), .D(new_n5267), .Y(new_n5269));
  AOI31xp33_ASAP7_75t_L     g05013(.A1(new_n5268), .A2(new_n5267), .A3(new_n5266), .B(\a[35] ), .Y(new_n5270));
  INVx1_ASAP7_75t_L         g05014(.A(new_n5270), .Y(new_n5271));
  NAND4xp25_ASAP7_75t_L     g05015(.A(new_n5261), .B(new_n5271), .C(new_n5269), .D(new_n5265), .Y(new_n5272));
  AOI211xp5_ASAP7_75t_L     g05016(.A1(new_n4995), .A2(new_n5262), .B(new_n5263), .C(new_n5264), .Y(new_n5273));
  AOI211xp5_ASAP7_75t_L     g05017(.A1(new_n5257), .A2(new_n5260), .B(new_n5229), .C(new_n4980), .Y(new_n5274));
  INVx1_ASAP7_75t_L         g05018(.A(new_n5269), .Y(new_n5275));
  OAI22xp33_ASAP7_75t_L     g05019(.A1(new_n5273), .A2(new_n5274), .B1(new_n5270), .B2(new_n5275), .Y(new_n5276));
  NAND2xp33_ASAP7_75t_L     g05020(.A(new_n5272), .B(new_n5276), .Y(new_n5277));
  AOI211xp5_ASAP7_75t_L     g05021(.A1(new_n4997), .A2(new_n4992), .B(new_n4985), .C(new_n4980), .Y(new_n5278));
  INVx1_ASAP7_75t_L         g05022(.A(new_n5278), .Y(new_n5279));
  A2O1A1Ixp33_ASAP7_75t_L   g05023(.A1(new_n5010), .A2(new_n5009), .B(new_n5007), .C(new_n5279), .Y(new_n5280));
  NOR2xp33_ASAP7_75t_L      g05024(.A(new_n5277), .B(new_n5280), .Y(new_n5281));
  O2A1O1Ixp33_ASAP7_75t_L   g05025(.A1(new_n4994), .A2(new_n4998), .B(new_n5022), .C(new_n5278), .Y(new_n5282));
  AOI21xp33_ASAP7_75t_L     g05026(.A1(new_n5276), .A2(new_n5272), .B(new_n5282), .Y(new_n5283));
  NAND2xp33_ASAP7_75t_L     g05027(.A(\b[9] ), .B(new_n3260), .Y(new_n5284));
  NAND2xp33_ASAP7_75t_L     g05028(.A(\b[10] ), .B(new_n3256), .Y(new_n5285));
  OAI311xp33_ASAP7_75t_L    g05029(.A1(new_n639), .A2(new_n851), .A3(new_n3261), .B1(new_n5285), .C1(new_n5284), .Y(new_n5286));
  AOI21xp33_ASAP7_75t_L     g05030(.A1(new_n3491), .A2(\b[8] ), .B(new_n5286), .Y(new_n5287));
  NAND2xp33_ASAP7_75t_L     g05031(.A(\a[32] ), .B(new_n5287), .Y(new_n5288));
  A2O1A1Ixp33_ASAP7_75t_L   g05032(.A1(\b[8] ), .A2(new_n3491), .B(new_n5286), .C(new_n3251), .Y(new_n5289));
  AND2x2_ASAP7_75t_L        g05033(.A(new_n5289), .B(new_n5288), .Y(new_n5290));
  OAI21xp33_ASAP7_75t_L     g05034(.A1(new_n5283), .A2(new_n5281), .B(new_n5290), .Y(new_n5291));
  NAND3xp33_ASAP7_75t_L     g05035(.A(new_n5282), .B(new_n5276), .C(new_n5272), .Y(new_n5292));
  A2O1A1Ixp33_ASAP7_75t_L   g05036(.A1(new_n5011), .A2(new_n5022), .B(new_n5278), .C(new_n5277), .Y(new_n5293));
  NAND2xp33_ASAP7_75t_L     g05037(.A(new_n5289), .B(new_n5288), .Y(new_n5294));
  NAND3xp33_ASAP7_75t_L     g05038(.A(new_n5292), .B(new_n5293), .C(new_n5294), .Y(new_n5295));
  NAND4xp25_ASAP7_75t_L     g05039(.A(new_n5043), .B(new_n5295), .C(new_n5291), .D(new_n5227), .Y(new_n5296));
  A2O1A1Ixp33_ASAP7_75t_L   g05040(.A1(new_n5026), .A2(new_n5020), .B(new_n5030), .C(new_n5227), .Y(new_n5297));
  AOI21xp33_ASAP7_75t_L     g05041(.A1(new_n5292), .A2(new_n5293), .B(new_n5294), .Y(new_n5298));
  NOR3xp33_ASAP7_75t_L      g05042(.A(new_n5290), .B(new_n5281), .C(new_n5283), .Y(new_n5299));
  OAI21xp33_ASAP7_75t_L     g05043(.A1(new_n5298), .A2(new_n5299), .B(new_n5297), .Y(new_n5300));
  NAND3xp33_ASAP7_75t_L     g05044(.A(new_n5296), .B(new_n5300), .C(new_n5226), .Y(new_n5301));
  INVx1_ASAP7_75t_L         g05045(.A(new_n5226), .Y(new_n5302));
  NOR3xp33_ASAP7_75t_L      g05046(.A(new_n5297), .B(new_n5298), .C(new_n5299), .Y(new_n5303));
  INVx1_ASAP7_75t_L         g05047(.A(new_n5227), .Y(new_n5304));
  O2A1O1Ixp33_ASAP7_75t_L   g05048(.A1(new_n5040), .A2(new_n5042), .B(new_n5028), .C(new_n5304), .Y(new_n5305));
  AOI21xp33_ASAP7_75t_L     g05049(.A1(new_n5295), .A2(new_n5291), .B(new_n5305), .Y(new_n5306));
  OAI21xp33_ASAP7_75t_L     g05050(.A1(new_n5306), .A2(new_n5303), .B(new_n5302), .Y(new_n5307));
  NAND3xp33_ASAP7_75t_L     g05051(.A(new_n5219), .B(new_n5301), .C(new_n5307), .Y(new_n5308));
  NOR3xp33_ASAP7_75t_L      g05052(.A(new_n5029), .B(new_n5031), .C(new_n5037), .Y(new_n5309));
  A2O1A1O1Ixp25_ASAP7_75t_L g05053(.A1(new_n4810), .A2(new_n4811), .B(new_n5049), .C(new_n5038), .D(new_n5309), .Y(new_n5310));
  NOR3xp33_ASAP7_75t_L      g05054(.A(new_n5302), .B(new_n5306), .C(new_n5303), .Y(new_n5311));
  AOI21xp33_ASAP7_75t_L     g05055(.A1(new_n5296), .A2(new_n5300), .B(new_n5226), .Y(new_n5312));
  OAI21xp33_ASAP7_75t_L     g05056(.A1(new_n5312), .A2(new_n5311), .B(new_n5310), .Y(new_n5313));
  NAND2xp33_ASAP7_75t_L     g05057(.A(\b[14] ), .B(new_n2386), .Y(new_n5314));
  NAND2xp33_ASAP7_75t_L     g05058(.A(\b[15] ), .B(new_n2232), .Y(new_n5315));
  AOI22xp33_ASAP7_75t_L     g05059(.A1(new_n2228), .A2(\b[16] ), .B1(new_n2226), .B2(new_n1058), .Y(new_n5316));
  AND4x1_ASAP7_75t_L        g05060(.A(new_n5316), .B(new_n5315), .C(new_n5314), .D(\a[26] ), .Y(new_n5317));
  AOI31xp33_ASAP7_75t_L     g05061(.A1(new_n5316), .A2(new_n5315), .A3(new_n5314), .B(\a[26] ), .Y(new_n5318));
  NOR2xp33_ASAP7_75t_L      g05062(.A(new_n5318), .B(new_n5317), .Y(new_n5319));
  NAND3xp33_ASAP7_75t_L     g05063(.A(new_n5308), .B(new_n5313), .C(new_n5319), .Y(new_n5320));
  NOR3xp33_ASAP7_75t_L      g05064(.A(new_n5310), .B(new_n5311), .C(new_n5312), .Y(new_n5321));
  AOI221xp5_ASAP7_75t_L     g05065(.A1(new_n5038), .A2(new_n5046), .B1(new_n5301), .B2(new_n5307), .C(new_n5309), .Y(new_n5322));
  OR2x4_ASAP7_75t_L         g05066(.A(new_n5318), .B(new_n5317), .Y(new_n5323));
  OAI21xp33_ASAP7_75t_L     g05067(.A1(new_n5321), .A2(new_n5322), .B(new_n5323), .Y(new_n5324));
  XNOR2x2_ASAP7_75t_L       g05068(.A(new_n5046), .B(new_n5048), .Y(new_n5325));
  INVx1_ASAP7_75t_L         g05069(.A(new_n5058), .Y(new_n5326));
  MAJIxp5_ASAP7_75t_L       g05070(.A(new_n4964), .B(new_n5325), .C(new_n5326), .Y(new_n5327));
  NAND3xp33_ASAP7_75t_L     g05071(.A(new_n5327), .B(new_n5324), .C(new_n5320), .Y(new_n5328));
  NAND2xp33_ASAP7_75t_L     g05072(.A(new_n5324), .B(new_n5320), .Y(new_n5329));
  A2O1A1Ixp33_ASAP7_75t_L   g05073(.A1(new_n5326), .A2(new_n5325), .B(new_n5068), .C(new_n5329), .Y(new_n5330));
  NOR2xp33_ASAP7_75t_L      g05074(.A(new_n1244), .B(new_n1911), .Y(new_n5331));
  NAND2xp33_ASAP7_75t_L     g05075(.A(\b[18] ), .B(new_n1770), .Y(new_n5332));
  OAI221xp5_ASAP7_75t_L     g05076(.A1(new_n1772), .A2(new_n1493), .B1(new_n1771), .B2(new_n2793), .C(new_n5332), .Y(new_n5333));
  OR3x1_ASAP7_75t_L         g05077(.A(new_n5333), .B(new_n1761), .C(new_n5331), .Y(new_n5334));
  A2O1A1Ixp33_ASAP7_75t_L   g05078(.A1(\b[17] ), .A2(new_n1910), .B(new_n5333), .C(new_n1761), .Y(new_n5335));
  AND2x2_ASAP7_75t_L        g05079(.A(new_n5335), .B(new_n5334), .Y(new_n5336));
  NAND3xp33_ASAP7_75t_L     g05080(.A(new_n5336), .B(new_n5330), .C(new_n5328), .Y(new_n5337));
  NAND2xp33_ASAP7_75t_L     g05081(.A(new_n5047), .B(new_n5051), .Y(new_n5338));
  MAJIxp5_ASAP7_75t_L       g05082(.A(new_n5062), .B(new_n5338), .C(new_n5058), .Y(new_n5339));
  NOR2xp33_ASAP7_75t_L      g05083(.A(new_n5339), .B(new_n5329), .Y(new_n5340));
  AOI21xp33_ASAP7_75t_L     g05084(.A1(new_n5324), .A2(new_n5320), .B(new_n5327), .Y(new_n5341));
  NAND2xp33_ASAP7_75t_L     g05085(.A(new_n5335), .B(new_n5334), .Y(new_n5342));
  OAI21xp33_ASAP7_75t_L     g05086(.A1(new_n5341), .A2(new_n5340), .B(new_n5342), .Y(new_n5343));
  A2O1A1O1Ixp25_ASAP7_75t_L g05087(.A1(new_n4839), .A2(new_n4841), .B(new_n4956), .C(new_n5070), .D(new_n5073), .Y(new_n5344));
  NAND3xp33_ASAP7_75t_L     g05088(.A(new_n5344), .B(new_n5337), .C(new_n5343), .Y(new_n5345));
  AO21x2_ASAP7_75t_L        g05089(.A1(new_n5337), .A2(new_n5343), .B(new_n5344), .Y(new_n5346));
  NAND2xp33_ASAP7_75t_L     g05090(.A(\b[20] ), .B(new_n1548), .Y(new_n5347));
  NAND2xp33_ASAP7_75t_L     g05091(.A(\b[21] ), .B(new_n1410), .Y(new_n5348));
  AOI32xp33_ASAP7_75t_L     g05092(.A1(new_n1862), .A2(new_n1860), .A3(new_n1404), .B1(new_n1406), .B2(\b[22] ), .Y(new_n5349));
  NAND4xp25_ASAP7_75t_L     g05093(.A(new_n5349), .B(\a[20] ), .C(new_n5347), .D(new_n5348), .Y(new_n5350));
  NAND2xp33_ASAP7_75t_L     g05094(.A(new_n5348), .B(new_n5349), .Y(new_n5351));
  A2O1A1Ixp33_ASAP7_75t_L   g05095(.A1(\b[20] ), .A2(new_n1548), .B(new_n5351), .C(new_n1401), .Y(new_n5352));
  AND2x2_ASAP7_75t_L        g05096(.A(new_n5350), .B(new_n5352), .Y(new_n5353));
  NAND3xp33_ASAP7_75t_L     g05097(.A(new_n5346), .B(new_n5353), .C(new_n5345), .Y(new_n5354));
  AND3x1_ASAP7_75t_L        g05098(.A(new_n5344), .B(new_n5343), .C(new_n5337), .Y(new_n5355));
  AOI21xp33_ASAP7_75t_L     g05099(.A1(new_n5337), .A2(new_n5343), .B(new_n5344), .Y(new_n5356));
  NAND2xp33_ASAP7_75t_L     g05100(.A(new_n5350), .B(new_n5352), .Y(new_n5357));
  OAI21xp33_ASAP7_75t_L     g05101(.A1(new_n5356), .A2(new_n5355), .B(new_n5357), .Y(new_n5358));
  NAND2xp33_ASAP7_75t_L     g05102(.A(new_n5354), .B(new_n5358), .Y(new_n5359));
  NAND3xp33_ASAP7_75t_L     g05103(.A(new_n5088), .B(new_n5076), .C(new_n5071), .Y(new_n5360));
  A2O1A1Ixp33_ASAP7_75t_L   g05104(.A1(new_n5089), .A2(new_n5083), .B(new_n5093), .C(new_n5360), .Y(new_n5361));
  NOR2xp33_ASAP7_75t_L      g05105(.A(new_n5359), .B(new_n5361), .Y(new_n5362));
  INVx1_ASAP7_75t_L         g05106(.A(new_n5090), .Y(new_n5363));
  NOR3xp33_ASAP7_75t_L      g05107(.A(new_n5355), .B(new_n5356), .C(new_n5357), .Y(new_n5364));
  AOI21xp33_ASAP7_75t_L     g05108(.A1(new_n5346), .A2(new_n5345), .B(new_n5353), .Y(new_n5365));
  NOR2xp33_ASAP7_75t_L      g05109(.A(new_n5365), .B(new_n5364), .Y(new_n5366));
  O2A1O1Ixp33_ASAP7_75t_L   g05110(.A1(new_n5093), .A2(new_n5363), .B(new_n5360), .C(new_n5366), .Y(new_n5367));
  NOR2xp33_ASAP7_75t_L      g05111(.A(new_n1995), .B(new_n1195), .Y(new_n5368));
  NAND2xp33_ASAP7_75t_L     g05112(.A(\b[24] ), .B(new_n1103), .Y(new_n5369));
  OAI221xp5_ASAP7_75t_L     g05113(.A1(new_n1198), .A2(new_n2180), .B1(new_n1197), .B2(new_n2187), .C(new_n5369), .Y(new_n5370));
  OR3x1_ASAP7_75t_L         g05114(.A(new_n5370), .B(new_n1107), .C(new_n5368), .Y(new_n5371));
  A2O1A1Ixp33_ASAP7_75t_L   g05115(.A1(\b[23] ), .A2(new_n1194), .B(new_n5370), .C(new_n1107), .Y(new_n5372));
  NAND2xp33_ASAP7_75t_L     g05116(.A(new_n5372), .B(new_n5371), .Y(new_n5373));
  NOR3xp33_ASAP7_75t_L      g05117(.A(new_n5367), .B(new_n5362), .C(new_n5373), .Y(new_n5374));
  NAND3xp33_ASAP7_75t_L     g05118(.A(new_n5105), .B(new_n5366), .C(new_n5360), .Y(new_n5375));
  NAND2xp33_ASAP7_75t_L     g05119(.A(new_n5359), .B(new_n5361), .Y(new_n5376));
  AND2x2_ASAP7_75t_L        g05120(.A(new_n5372), .B(new_n5371), .Y(new_n5377));
  AOI21xp33_ASAP7_75t_L     g05121(.A1(new_n5375), .A2(new_n5376), .B(new_n5377), .Y(new_n5378));
  A2O1A1Ixp33_ASAP7_75t_L   g05122(.A1(new_n4650), .A2(new_n4651), .B(new_n4750), .C(new_n4864), .Y(new_n5379));
  A2O1A1Ixp33_ASAP7_75t_L   g05123(.A1(new_n5379), .A2(new_n4866), .B(new_n5110), .C(new_n5107), .Y(new_n5380));
  OAI21xp33_ASAP7_75t_L     g05124(.A1(new_n5374), .A2(new_n5378), .B(new_n5380), .Y(new_n5381));
  NAND3xp33_ASAP7_75t_L     g05125(.A(new_n5375), .B(new_n5376), .C(new_n5377), .Y(new_n5382));
  OAI21xp33_ASAP7_75t_L     g05126(.A1(new_n5362), .A2(new_n5367), .B(new_n5373), .Y(new_n5383));
  A2O1A1O1Ixp25_ASAP7_75t_L g05127(.A1(new_n4864), .A2(new_n4880), .B(new_n4865), .C(new_n5102), .D(new_n5111), .Y(new_n5384));
  NAND3xp33_ASAP7_75t_L     g05128(.A(new_n5384), .B(new_n5383), .C(new_n5382), .Y(new_n5385));
  AOI21xp33_ASAP7_75t_L     g05129(.A1(new_n5385), .A2(new_n5381), .B(new_n5217), .Y(new_n5386));
  NAND2xp33_ASAP7_75t_L     g05130(.A(new_n5216), .B(new_n5215), .Y(new_n5387));
  AOI21xp33_ASAP7_75t_L     g05131(.A1(new_n5383), .A2(new_n5382), .B(new_n5384), .Y(new_n5388));
  NOR3xp33_ASAP7_75t_L      g05132(.A(new_n5380), .B(new_n5378), .C(new_n5374), .Y(new_n5389));
  NOR3xp33_ASAP7_75t_L      g05133(.A(new_n5388), .B(new_n5389), .C(new_n5387), .Y(new_n5390));
  NOR2xp33_ASAP7_75t_L      g05134(.A(new_n5390), .B(new_n5386), .Y(new_n5391));
  NAND2xp33_ASAP7_75t_L     g05135(.A(new_n5210), .B(new_n5391), .Y(new_n5392));
  OAI221xp5_ASAP7_75t_L     g05136(.A1(new_n5386), .A2(new_n5390), .B1(new_n5129), .B2(new_n5130), .C(new_n5209), .Y(new_n5393));
  NOR2xp33_ASAP7_75t_L      g05137(.A(new_n2871), .B(new_n1620), .Y(new_n5394));
  NOR2xp33_ASAP7_75t_L      g05138(.A(new_n3212), .B(new_n721), .Y(new_n5395));
  OAI22xp33_ASAP7_75t_L     g05139(.A1(new_n4030), .A2(new_n675), .B1(new_n3419), .B2(new_n676), .Y(new_n5396));
  NOR4xp25_ASAP7_75t_L      g05140(.A(new_n5396), .B(new_n594), .C(new_n5394), .D(new_n5395), .Y(new_n5397));
  NOR2xp33_ASAP7_75t_L      g05141(.A(new_n5395), .B(new_n5396), .Y(new_n5398));
  O2A1O1Ixp33_ASAP7_75t_L   g05142(.A1(new_n2871), .A2(new_n1620), .B(new_n5398), .C(\a[11] ), .Y(new_n5399));
  NOR2xp33_ASAP7_75t_L      g05143(.A(new_n5397), .B(new_n5399), .Y(new_n5400));
  NAND3xp33_ASAP7_75t_L     g05144(.A(new_n5392), .B(new_n5400), .C(new_n5393), .Y(new_n5401));
  OAI21xp33_ASAP7_75t_L     g05145(.A1(new_n5389), .A2(new_n5388), .B(new_n5387), .Y(new_n5402));
  NAND3xp33_ASAP7_75t_L     g05146(.A(new_n5385), .B(new_n5217), .C(new_n5381), .Y(new_n5403));
  NAND2xp33_ASAP7_75t_L     g05147(.A(new_n5403), .B(new_n5402), .Y(new_n5404));
  O2A1O1Ixp33_ASAP7_75t_L   g05148(.A1(new_n5129), .A2(new_n5130), .B(new_n5209), .C(new_n5404), .Y(new_n5405));
  INVx1_ASAP7_75t_L         g05149(.A(new_n5393), .Y(new_n5406));
  INVx1_ASAP7_75t_L         g05150(.A(new_n5400), .Y(new_n5407));
  OAI21xp33_ASAP7_75t_L     g05151(.A1(new_n5405), .A2(new_n5406), .B(new_n5407), .Y(new_n5408));
  NAND3xp33_ASAP7_75t_L     g05152(.A(new_n5208), .B(new_n5408), .C(new_n5401), .Y(new_n5409));
  A2O1A1O1Ixp25_ASAP7_75t_L g05153(.A1(new_n4891), .A2(new_n4895), .B(new_n5139), .C(new_n5137), .D(new_n5141), .Y(new_n5410));
  NOR3xp33_ASAP7_75t_L      g05154(.A(new_n5406), .B(new_n5407), .C(new_n5405), .Y(new_n5411));
  AOI21xp33_ASAP7_75t_L     g05155(.A1(new_n5392), .A2(new_n5393), .B(new_n5400), .Y(new_n5412));
  OAI21xp33_ASAP7_75t_L     g05156(.A1(new_n5411), .A2(new_n5412), .B(new_n5410), .Y(new_n5413));
  AO21x2_ASAP7_75t_L        g05157(.A1(new_n5409), .A2(new_n5413), .B(new_n5207), .Y(new_n5414));
  NAND3xp33_ASAP7_75t_L     g05158(.A(new_n5413), .B(new_n5409), .C(new_n5207), .Y(new_n5415));
  AND2x2_ASAP7_75t_L        g05159(.A(new_n5415), .B(new_n5414), .Y(new_n5416));
  A2O1A1Ixp33_ASAP7_75t_L   g05160(.A1(new_n5156), .A2(new_n4941), .B(new_n5200), .C(new_n5416), .Y(new_n5417));
  A2O1A1O1Ixp25_ASAP7_75t_L g05161(.A1(new_n4897), .A2(new_n4903), .B(new_n4905), .C(new_n5156), .D(new_n5200), .Y(new_n5418));
  NAND2xp33_ASAP7_75t_L     g05162(.A(new_n5415), .B(new_n5414), .Y(new_n5419));
  NAND2xp33_ASAP7_75t_L     g05163(.A(new_n5419), .B(new_n5418), .Y(new_n5420));
  NAND2xp33_ASAP7_75t_L     g05164(.A(\b[36] ), .B(new_n334), .Y(new_n5421));
  AOI22xp33_ASAP7_75t_L     g05165(.A1(new_n345), .A2(\b[37] ), .B1(new_n342), .B2(new_n4709), .Y(new_n5422));
  NAND2xp33_ASAP7_75t_L     g05166(.A(new_n5421), .B(new_n5422), .Y(new_n5423));
  AOI211xp5_ASAP7_75t_L     g05167(.A1(\b[35] ), .A2(new_n366), .B(new_n339), .C(new_n5423), .Y(new_n5424));
  AND2x2_ASAP7_75t_L        g05168(.A(new_n5421), .B(new_n5422), .Y(new_n5425));
  O2A1O1Ixp33_ASAP7_75t_L   g05169(.A1(new_n4053), .A2(new_n365), .B(new_n5425), .C(\a[5] ), .Y(new_n5426));
  NOR2xp33_ASAP7_75t_L      g05170(.A(new_n5424), .B(new_n5426), .Y(new_n5427));
  NAND3xp33_ASAP7_75t_L     g05171(.A(new_n5417), .B(new_n5427), .C(new_n5420), .Y(new_n5428));
  AO21x2_ASAP7_75t_L        g05172(.A1(new_n5420), .A2(new_n5417), .B(new_n5427), .Y(new_n5429));
  AOI21xp33_ASAP7_75t_L     g05173(.A1(new_n5429), .A2(new_n5428), .B(new_n5199), .Y(new_n5430));
  NAND3xp33_ASAP7_75t_L     g05174(.A(new_n5429), .B(new_n5199), .C(new_n5428), .Y(new_n5431));
  INVx1_ASAP7_75t_L         g05175(.A(new_n5431), .Y(new_n5432));
  NOR3xp33_ASAP7_75t_L      g05176(.A(new_n5432), .B(new_n5198), .C(new_n5430), .Y(new_n5433));
  INVx1_ASAP7_75t_L         g05177(.A(new_n5198), .Y(new_n5434));
  INVx1_ASAP7_75t_L         g05178(.A(new_n5430), .Y(new_n5435));
  AOI21xp33_ASAP7_75t_L     g05179(.A1(new_n5435), .A2(new_n5431), .B(new_n5434), .Y(new_n5436));
  NOR2xp33_ASAP7_75t_L      g05180(.A(new_n5433), .B(new_n5436), .Y(new_n5437));
  INVx1_ASAP7_75t_L         g05181(.A(new_n5437), .Y(new_n5438));
  O2A1O1Ixp33_ASAP7_75t_L   g05182(.A1(new_n5163), .A2(new_n5177), .B(new_n5181), .C(new_n5438), .Y(new_n5439));
  MAJIxp5_ASAP7_75t_L       g05183(.A(new_n5179), .B(new_n5163), .C(new_n5177), .Y(new_n5440));
  NOR2xp33_ASAP7_75t_L      g05184(.A(new_n5437), .B(new_n5440), .Y(new_n5441));
  NOR2xp33_ASAP7_75t_L      g05185(.A(new_n5441), .B(new_n5439), .Y(\f[40] ));
  NOR2xp33_ASAP7_75t_L      g05186(.A(new_n5433), .B(new_n5439), .Y(new_n5443));
  XNOR2x2_ASAP7_75t_L       g05187(.A(new_n5419), .B(new_n5418), .Y(new_n5444));
  MAJIxp5_ASAP7_75t_L       g05188(.A(new_n5199), .B(new_n5427), .C(new_n5444), .Y(new_n5445));
  NAND2xp33_ASAP7_75t_L     g05189(.A(\b[36] ), .B(new_n366), .Y(new_n5446));
  NAND2xp33_ASAP7_75t_L     g05190(.A(\b[37] ), .B(new_n334), .Y(new_n5447));
  AOI22xp33_ASAP7_75t_L     g05191(.A1(new_n345), .A2(\b[38] ), .B1(new_n342), .B2(new_n4923), .Y(new_n5448));
  NAND4xp25_ASAP7_75t_L     g05192(.A(new_n5448), .B(\a[5] ), .C(new_n5446), .D(new_n5447), .Y(new_n5449));
  NAND2xp33_ASAP7_75t_L     g05193(.A(new_n5447), .B(new_n5448), .Y(new_n5450));
  A2O1A1Ixp33_ASAP7_75t_L   g05194(.A1(\b[36] ), .A2(new_n366), .B(new_n5450), .C(new_n339), .Y(new_n5451));
  AND2x2_ASAP7_75t_L        g05195(.A(new_n5449), .B(new_n5451), .Y(new_n5452));
  AND3x1_ASAP7_75t_L        g05196(.A(new_n5413), .B(new_n5409), .C(new_n5207), .Y(new_n5453));
  A2O1A1O1Ixp25_ASAP7_75t_L g05197(.A1(new_n5156), .A2(new_n4941), .B(new_n5200), .C(new_n5414), .D(new_n5453), .Y(new_n5454));
  A2O1A1O1Ixp25_ASAP7_75t_L g05198(.A1(new_n5137), .A2(new_n4944), .B(new_n5141), .C(new_n5401), .D(new_n5412), .Y(new_n5455));
  NOR2xp33_ASAP7_75t_L      g05199(.A(new_n3212), .B(new_n1620), .Y(new_n5456));
  INVx1_ASAP7_75t_L         g05200(.A(new_n5456), .Y(new_n5457));
  NAND2xp33_ASAP7_75t_L     g05201(.A(\b[31] ), .B(new_n590), .Y(new_n5458));
  AOI22xp33_ASAP7_75t_L     g05202(.A1(new_n600), .A2(\b[32] ), .B1(new_n597), .B2(new_n3450), .Y(new_n5459));
  AND4x1_ASAP7_75t_L        g05203(.A(new_n5459), .B(new_n5458), .C(new_n5457), .D(\a[11] ), .Y(new_n5460));
  AOI31xp33_ASAP7_75t_L     g05204(.A1(new_n5459), .A2(new_n5458), .A3(new_n5457), .B(\a[11] ), .Y(new_n5461));
  NOR2xp33_ASAP7_75t_L      g05205(.A(new_n5461), .B(new_n5460), .Y(new_n5462));
  INVx1_ASAP7_75t_L         g05206(.A(new_n5462), .Y(new_n5463));
  INVx1_ASAP7_75t_L         g05207(.A(new_n5209), .Y(new_n5464));
  AOI21xp33_ASAP7_75t_L     g05208(.A1(new_n5135), .A2(new_n5127), .B(new_n5464), .Y(new_n5465));
  NOR3xp33_ASAP7_75t_L      g05209(.A(new_n5388), .B(new_n5389), .C(new_n5217), .Y(new_n5466));
  INVx1_ASAP7_75t_L         g05210(.A(new_n5466), .Y(new_n5467));
  OAI21xp33_ASAP7_75t_L     g05211(.A1(new_n5465), .A2(new_n5391), .B(new_n5467), .Y(new_n5468));
  NOR2xp33_ASAP7_75t_L      g05212(.A(new_n2650), .B(new_n909), .Y(new_n5469));
  INVx1_ASAP7_75t_L         g05213(.A(new_n5469), .Y(new_n5470));
  NAND2xp33_ASAP7_75t_L     g05214(.A(\b[28] ), .B(new_n817), .Y(new_n5471));
  AND2x2_ASAP7_75t_L        g05215(.A(new_n2880), .B(new_n2877), .Y(new_n5472));
  AOI22xp33_ASAP7_75t_L     g05216(.A1(new_n826), .A2(\b[29] ), .B1(new_n823), .B2(new_n5472), .Y(new_n5473));
  AND4x1_ASAP7_75t_L        g05217(.A(new_n5473), .B(new_n5471), .C(new_n5470), .D(\a[14] ), .Y(new_n5474));
  AOI31xp33_ASAP7_75t_L     g05218(.A1(new_n5473), .A2(new_n5471), .A3(new_n5470), .B(\a[14] ), .Y(new_n5475));
  NOR2xp33_ASAP7_75t_L      g05219(.A(new_n5475), .B(new_n5474), .Y(new_n5476));
  NOR2xp33_ASAP7_75t_L      g05220(.A(new_n5362), .B(new_n5367), .Y(new_n5477));
  MAJIxp5_ASAP7_75t_L       g05221(.A(new_n5380), .B(new_n5373), .C(new_n5477), .Y(new_n5478));
  AOI22xp33_ASAP7_75t_L     g05222(.A1(new_n1113), .A2(\b[26] ), .B1(new_n1110), .B2(new_n2888), .Y(new_n5479));
  OAI221xp5_ASAP7_75t_L     g05223(.A1(new_n1298), .A2(new_n2180), .B1(new_n2019), .B2(new_n1195), .C(new_n5479), .Y(new_n5480));
  XNOR2x2_ASAP7_75t_L       g05224(.A(new_n1107), .B(new_n5480), .Y(new_n5481));
  NOR3xp33_ASAP7_75t_L      g05225(.A(new_n5355), .B(new_n5353), .C(new_n5356), .Y(new_n5482));
  INVx1_ASAP7_75t_L         g05226(.A(new_n5482), .Y(new_n5483));
  A2O1A1Ixp33_ASAP7_75t_L   g05227(.A1(new_n5105), .A2(new_n5360), .B(new_n5366), .C(new_n5483), .Y(new_n5484));
  AND2x2_ASAP7_75t_L        g05228(.A(new_n5324), .B(new_n5320), .Y(new_n5485));
  NOR2xp33_ASAP7_75t_L      g05229(.A(new_n5321), .B(new_n5322), .Y(new_n5486));
  NAND2xp33_ASAP7_75t_L     g05230(.A(new_n5323), .B(new_n5486), .Y(new_n5487));
  NAND2xp33_ASAP7_75t_L     g05231(.A(\b[15] ), .B(new_n2386), .Y(new_n5488));
  NAND2xp33_ASAP7_75t_L     g05232(.A(\b[16] ), .B(new_n2232), .Y(new_n5489));
  AOI32xp33_ASAP7_75t_L     g05233(.A1(new_n1250), .A2(new_n1247), .A3(new_n2226), .B1(\b[17] ), .B2(new_n2228), .Y(new_n5490));
  NAND4xp25_ASAP7_75t_L     g05234(.A(new_n5490), .B(\a[26] ), .C(new_n5488), .D(new_n5489), .Y(new_n5491));
  INVx1_ASAP7_75t_L         g05235(.A(new_n5491), .Y(new_n5492));
  AOI31xp33_ASAP7_75t_L     g05236(.A1(new_n5490), .A2(new_n5489), .A3(new_n5488), .B(\a[26] ), .Y(new_n5493));
  NOR2xp33_ASAP7_75t_L      g05237(.A(new_n5493), .B(new_n5492), .Y(new_n5494));
  A2O1A1O1Ixp25_ASAP7_75t_L g05238(.A1(new_n5038), .A2(new_n5046), .B(new_n5309), .C(new_n5301), .D(new_n5312), .Y(new_n5495));
  NOR2xp33_ASAP7_75t_L      g05239(.A(new_n763), .B(new_n2932), .Y(new_n5496));
  INVx1_ASAP7_75t_L         g05240(.A(new_n5496), .Y(new_n5497));
  NAND2xp33_ASAP7_75t_L     g05241(.A(\b[13] ), .B(new_n2706), .Y(new_n5498));
  AOI32xp33_ASAP7_75t_L     g05242(.A1(new_n877), .A2(new_n874), .A3(new_n2700), .B1(\b[14] ), .B2(new_n2702), .Y(new_n5499));
  NAND4xp25_ASAP7_75t_L     g05243(.A(new_n5499), .B(\a[29] ), .C(new_n5497), .D(new_n5498), .Y(new_n5500));
  AOI31xp33_ASAP7_75t_L     g05244(.A1(new_n5499), .A2(new_n5498), .A3(new_n5497), .B(\a[29] ), .Y(new_n5501));
  INVx1_ASAP7_75t_L         g05245(.A(new_n5501), .Y(new_n5502));
  NAND2xp33_ASAP7_75t_L     g05246(.A(new_n5500), .B(new_n5502), .Y(new_n5503));
  OAI211xp5_ASAP7_75t_L     g05247(.A1(new_n5275), .A2(new_n5270), .B(new_n5261), .C(new_n5265), .Y(new_n5504));
  A2O1A1Ixp33_ASAP7_75t_L   g05248(.A1(new_n5276), .A2(new_n5272), .B(new_n5282), .C(new_n5504), .Y(new_n5505));
  NOR2xp33_ASAP7_75t_L      g05249(.A(new_n382), .B(new_n4986), .Y(new_n5506));
  INVx1_ASAP7_75t_L         g05250(.A(new_n5506), .Y(new_n5507));
  NAND2xp33_ASAP7_75t_L     g05251(.A(\b[7] ), .B(new_n3874), .Y(new_n5508));
  AOI32xp33_ASAP7_75t_L     g05252(.A1(new_n508), .A2(new_n506), .A3(new_n3881), .B1(\b[8] ), .B2(new_n3884), .Y(new_n5509));
  NAND4xp25_ASAP7_75t_L     g05253(.A(new_n5509), .B(\a[35] ), .C(new_n5507), .D(new_n5508), .Y(new_n5510));
  AOI31xp33_ASAP7_75t_L     g05254(.A1(new_n5509), .A2(new_n5508), .A3(new_n5507), .B(\a[35] ), .Y(new_n5511));
  INVx1_ASAP7_75t_L         g05255(.A(new_n5511), .Y(new_n5512));
  A2O1A1Ixp33_ASAP7_75t_L   g05256(.A1(new_n4995), .A2(new_n5262), .B(new_n5263), .C(new_n5260), .Y(new_n5513));
  NAND2xp33_ASAP7_75t_L     g05257(.A(\b[3] ), .B(new_n4780), .Y(new_n5514));
  NAND2xp33_ASAP7_75t_L     g05258(.A(\b[4] ), .B(new_n4548), .Y(new_n5515));
  AOI32xp33_ASAP7_75t_L     g05259(.A1(new_n358), .A2(new_n356), .A3(new_n4542), .B1(\b[5] ), .B2(new_n4544), .Y(new_n5516));
  NAND4xp25_ASAP7_75t_L     g05260(.A(new_n5516), .B(\a[38] ), .C(new_n5514), .D(new_n5515), .Y(new_n5517));
  AOI31xp33_ASAP7_75t_L     g05261(.A1(new_n5516), .A2(new_n5515), .A3(new_n5514), .B(\a[38] ), .Y(new_n5518));
  INVx1_ASAP7_75t_L         g05262(.A(new_n5518), .Y(new_n5519));
  A2O1A1O1Ixp25_ASAP7_75t_L g05263(.A1(new_n5239), .A2(new_n4970), .B(new_n258), .C(new_n5250), .D(new_n5244), .Y(new_n5520));
  NAND3xp33_ASAP7_75t_L     g05264(.A(new_n4970), .B(new_n5239), .C(new_n5248), .Y(new_n5521));
  NOR2xp33_ASAP7_75t_L      g05265(.A(new_n258), .B(new_n5521), .Y(new_n5522));
  NAND2xp33_ASAP7_75t_L     g05266(.A(\b[1] ), .B(new_n5240), .Y(new_n5523));
  OAI221xp5_ASAP7_75t_L     g05267(.A1(new_n5252), .A2(new_n283), .B1(new_n278), .B2(new_n5253), .C(new_n5523), .Y(new_n5524));
  OR3x1_ASAP7_75t_L         g05268(.A(new_n5520), .B(new_n5522), .C(new_n5524), .Y(new_n5525));
  INVx1_ASAP7_75t_L         g05269(.A(new_n5521), .Y(new_n5526));
  A2O1A1Ixp33_ASAP7_75t_L   g05270(.A1(\b[0] ), .A2(new_n5526), .B(new_n5524), .C(new_n5520), .Y(new_n5527));
  NAND4xp25_ASAP7_75t_L     g05271(.A(new_n5525), .B(new_n5517), .C(new_n5519), .D(new_n5527), .Y(new_n5528));
  AO22x1_ASAP7_75t_L        g05272(.A1(new_n5517), .A2(new_n5519), .B1(new_n5527), .B2(new_n5525), .Y(new_n5529));
  NAND2xp33_ASAP7_75t_L     g05273(.A(new_n5528), .B(new_n5529), .Y(new_n5530));
  NAND2xp33_ASAP7_75t_L     g05274(.A(new_n5513), .B(new_n5530), .Y(new_n5531));
  NAND2xp33_ASAP7_75t_L     g05275(.A(new_n4972), .B(new_n4973), .Y(new_n5532));
  NAND2xp33_ASAP7_75t_L     g05276(.A(new_n4979), .B(new_n4976), .Y(new_n5533));
  A2O1A1O1Ixp25_ASAP7_75t_L g05277(.A1(new_n5533), .A2(new_n5532), .B(new_n5229), .C(new_n5257), .D(new_n5264), .Y(new_n5534));
  NAND3xp33_ASAP7_75t_L     g05278(.A(new_n5534), .B(new_n5528), .C(new_n5529), .Y(new_n5535));
  AOI22xp33_ASAP7_75t_L     g05279(.A1(new_n5510), .A2(new_n5512), .B1(new_n5531), .B2(new_n5535), .Y(new_n5536));
  INVx1_ASAP7_75t_L         g05280(.A(new_n5510), .Y(new_n5537));
  AOI21xp33_ASAP7_75t_L     g05281(.A1(new_n5529), .A2(new_n5528), .B(new_n5534), .Y(new_n5538));
  NOR2xp33_ASAP7_75t_L      g05282(.A(new_n5513), .B(new_n5530), .Y(new_n5539));
  NOR4xp25_ASAP7_75t_L      g05283(.A(new_n5538), .B(new_n5539), .C(new_n5537), .D(new_n5511), .Y(new_n5540));
  NOR2xp33_ASAP7_75t_L      g05284(.A(new_n5536), .B(new_n5540), .Y(new_n5541));
  NAND2xp33_ASAP7_75t_L     g05285(.A(new_n5541), .B(new_n5505), .Y(new_n5542));
  INVx1_ASAP7_75t_L         g05286(.A(new_n5504), .Y(new_n5543));
  A2O1A1O1Ixp25_ASAP7_75t_L g05287(.A1(new_n5022), .A2(new_n5011), .B(new_n5278), .C(new_n5277), .D(new_n5543), .Y(new_n5544));
  OAI22xp33_ASAP7_75t_L     g05288(.A1(new_n5538), .A2(new_n5539), .B1(new_n5537), .B2(new_n5511), .Y(new_n5545));
  NAND4xp25_ASAP7_75t_L     g05289(.A(new_n5535), .B(new_n5510), .C(new_n5531), .D(new_n5512), .Y(new_n5546));
  NAND2xp33_ASAP7_75t_L     g05290(.A(new_n5546), .B(new_n5545), .Y(new_n5547));
  NAND2xp33_ASAP7_75t_L     g05291(.A(new_n5547), .B(new_n5544), .Y(new_n5548));
  NAND2xp33_ASAP7_75t_L     g05292(.A(\b[9] ), .B(new_n3491), .Y(new_n5549));
  NAND2xp33_ASAP7_75t_L     g05293(.A(\b[10] ), .B(new_n3260), .Y(new_n5550));
  AOI32xp33_ASAP7_75t_L     g05294(.A1(new_n700), .A2(new_n698), .A3(new_n3254), .B1(\b[11] ), .B2(new_n3256), .Y(new_n5551));
  AND4x1_ASAP7_75t_L        g05295(.A(new_n5551), .B(new_n5550), .C(new_n5549), .D(\a[32] ), .Y(new_n5552));
  AOI31xp33_ASAP7_75t_L     g05296(.A1(new_n5551), .A2(new_n5550), .A3(new_n5549), .B(\a[32] ), .Y(new_n5553));
  NOR2xp33_ASAP7_75t_L      g05297(.A(new_n5553), .B(new_n5552), .Y(new_n5554));
  NAND3xp33_ASAP7_75t_L     g05298(.A(new_n5548), .B(new_n5542), .C(new_n5554), .Y(new_n5555));
  A2O1A1O1Ixp25_ASAP7_75t_L g05299(.A1(new_n5276), .A2(new_n5272), .B(new_n5282), .C(new_n5504), .D(new_n5547), .Y(new_n5556));
  NOR2xp33_ASAP7_75t_L      g05300(.A(new_n5541), .B(new_n5505), .Y(new_n5557));
  INVx1_ASAP7_75t_L         g05301(.A(new_n5554), .Y(new_n5558));
  OAI21xp33_ASAP7_75t_L     g05302(.A1(new_n5557), .A2(new_n5556), .B(new_n5558), .Y(new_n5559));
  A2O1A1Ixp33_ASAP7_75t_L   g05303(.A1(new_n5043), .A2(new_n5227), .B(new_n5298), .C(new_n5295), .Y(new_n5560));
  NAND3xp33_ASAP7_75t_L     g05304(.A(new_n5560), .B(new_n5559), .C(new_n5555), .Y(new_n5561));
  NOR3xp33_ASAP7_75t_L      g05305(.A(new_n5556), .B(new_n5557), .C(new_n5558), .Y(new_n5562));
  AOI21xp33_ASAP7_75t_L     g05306(.A1(new_n5548), .A2(new_n5542), .B(new_n5554), .Y(new_n5563));
  A2O1A1O1Ixp25_ASAP7_75t_L g05307(.A1(new_n5028), .A2(new_n5027), .B(new_n5304), .C(new_n5291), .D(new_n5299), .Y(new_n5564));
  OAI21xp33_ASAP7_75t_L     g05308(.A1(new_n5562), .A2(new_n5563), .B(new_n5564), .Y(new_n5565));
  AOI21xp33_ASAP7_75t_L     g05309(.A1(new_n5561), .A2(new_n5565), .B(new_n5503), .Y(new_n5566));
  INVx1_ASAP7_75t_L         g05310(.A(new_n5500), .Y(new_n5567));
  NOR2xp33_ASAP7_75t_L      g05311(.A(new_n5501), .B(new_n5567), .Y(new_n5568));
  NOR3xp33_ASAP7_75t_L      g05312(.A(new_n5564), .B(new_n5563), .C(new_n5562), .Y(new_n5569));
  A2O1A1O1Ixp25_ASAP7_75t_L g05313(.A1(new_n5026), .A2(new_n5020), .B(new_n5030), .C(new_n5227), .D(new_n5298), .Y(new_n5570));
  AOI211xp5_ASAP7_75t_L     g05314(.A1(new_n5559), .A2(new_n5555), .B(new_n5299), .C(new_n5570), .Y(new_n5571));
  NOR3xp33_ASAP7_75t_L      g05315(.A(new_n5569), .B(new_n5571), .C(new_n5568), .Y(new_n5572));
  NOR3xp33_ASAP7_75t_L      g05316(.A(new_n5495), .B(new_n5566), .C(new_n5572), .Y(new_n5573));
  OAI21xp33_ASAP7_75t_L     g05317(.A1(new_n5311), .A2(new_n5310), .B(new_n5307), .Y(new_n5574));
  OAI21xp33_ASAP7_75t_L     g05318(.A1(new_n5571), .A2(new_n5569), .B(new_n5568), .Y(new_n5575));
  NAND3xp33_ASAP7_75t_L     g05319(.A(new_n5561), .B(new_n5503), .C(new_n5565), .Y(new_n5576));
  AOI21xp33_ASAP7_75t_L     g05320(.A1(new_n5576), .A2(new_n5575), .B(new_n5574), .Y(new_n5577));
  OAI21xp33_ASAP7_75t_L     g05321(.A1(new_n5573), .A2(new_n5577), .B(new_n5494), .Y(new_n5578));
  INVx1_ASAP7_75t_L         g05322(.A(new_n5493), .Y(new_n5579));
  NAND2xp33_ASAP7_75t_L     g05323(.A(new_n5491), .B(new_n5579), .Y(new_n5580));
  NAND3xp33_ASAP7_75t_L     g05324(.A(new_n5574), .B(new_n5575), .C(new_n5576), .Y(new_n5581));
  OAI21xp33_ASAP7_75t_L     g05325(.A1(new_n5572), .A2(new_n5566), .B(new_n5495), .Y(new_n5582));
  NAND3xp33_ASAP7_75t_L     g05326(.A(new_n5581), .B(new_n5580), .C(new_n5582), .Y(new_n5583));
  NAND2xp33_ASAP7_75t_L     g05327(.A(new_n5583), .B(new_n5578), .Y(new_n5584));
  O2A1O1Ixp33_ASAP7_75t_L   g05328(.A1(new_n5485), .A2(new_n5327), .B(new_n5487), .C(new_n5584), .Y(new_n5585));
  NAND2xp33_ASAP7_75t_L     g05329(.A(new_n5313), .B(new_n5308), .Y(new_n5586));
  MAJIxp5_ASAP7_75t_L       g05330(.A(new_n5327), .B(new_n5586), .C(new_n5319), .Y(new_n5587));
  AOI21xp33_ASAP7_75t_L     g05331(.A1(new_n5581), .A2(new_n5582), .B(new_n5580), .Y(new_n5588));
  NOR3xp33_ASAP7_75t_L      g05332(.A(new_n5577), .B(new_n5573), .C(new_n5494), .Y(new_n5589));
  NOR2xp33_ASAP7_75t_L      g05333(.A(new_n5589), .B(new_n5588), .Y(new_n5590));
  NOR2xp33_ASAP7_75t_L      g05334(.A(new_n5590), .B(new_n5587), .Y(new_n5591));
  NAND2xp33_ASAP7_75t_L     g05335(.A(\b[18] ), .B(new_n1910), .Y(new_n5592));
  NAND2xp33_ASAP7_75t_L     g05336(.A(\b[19] ), .B(new_n1770), .Y(new_n5593));
  AOI22xp33_ASAP7_75t_L     g05337(.A1(new_n1766), .A2(\b[20] ), .B1(new_n1764), .B2(new_n1600), .Y(new_n5594));
  NAND4xp25_ASAP7_75t_L     g05338(.A(new_n5594), .B(\a[23] ), .C(new_n5592), .D(new_n5593), .Y(new_n5595));
  OAI221xp5_ASAP7_75t_L     g05339(.A1(new_n1772), .A2(new_n1594), .B1(new_n1771), .B2(new_n3001), .C(new_n5593), .Y(new_n5596));
  A2O1A1Ixp33_ASAP7_75t_L   g05340(.A1(\b[18] ), .A2(new_n1910), .B(new_n5596), .C(new_n1761), .Y(new_n5597));
  NAND2xp33_ASAP7_75t_L     g05341(.A(new_n5595), .B(new_n5597), .Y(new_n5598));
  NOR3xp33_ASAP7_75t_L      g05342(.A(new_n5591), .B(new_n5585), .C(new_n5598), .Y(new_n5599));
  OA21x2_ASAP7_75t_L        g05343(.A1(new_n5585), .A2(new_n5591), .B(new_n5598), .Y(new_n5600));
  NAND2xp33_ASAP7_75t_L     g05344(.A(new_n5328), .B(new_n5330), .Y(new_n5601));
  MAJIxp5_ASAP7_75t_L       g05345(.A(new_n5344), .B(new_n5336), .C(new_n5601), .Y(new_n5602));
  NOR3xp33_ASAP7_75t_L      g05346(.A(new_n5602), .B(new_n5600), .C(new_n5599), .Y(new_n5603));
  OA21x2_ASAP7_75t_L        g05347(.A1(new_n5599), .A2(new_n5600), .B(new_n5602), .Y(new_n5604));
  NOR2xp33_ASAP7_75t_L      g05348(.A(new_n1709), .B(new_n1549), .Y(new_n5605));
  INVx1_ASAP7_75t_L         g05349(.A(new_n5605), .Y(new_n5606));
  NAND2xp33_ASAP7_75t_L     g05350(.A(\b[22] ), .B(new_n1410), .Y(new_n5607));
  AOI22xp33_ASAP7_75t_L     g05351(.A1(new_n1406), .A2(\b[23] ), .B1(new_n1404), .B2(new_n2002), .Y(new_n5608));
  AND4x1_ASAP7_75t_L        g05352(.A(new_n5608), .B(new_n5607), .C(new_n5606), .D(\a[20] ), .Y(new_n5609));
  AOI31xp33_ASAP7_75t_L     g05353(.A1(new_n5608), .A2(new_n5607), .A3(new_n5606), .B(\a[20] ), .Y(new_n5610));
  NOR2xp33_ASAP7_75t_L      g05354(.A(new_n5610), .B(new_n5609), .Y(new_n5611));
  OAI21xp33_ASAP7_75t_L     g05355(.A1(new_n5603), .A2(new_n5604), .B(new_n5611), .Y(new_n5612));
  OR3x1_ASAP7_75t_L         g05356(.A(new_n5602), .B(new_n5599), .C(new_n5600), .Y(new_n5613));
  OAI21xp33_ASAP7_75t_L     g05357(.A1(new_n5599), .A2(new_n5600), .B(new_n5602), .Y(new_n5614));
  OAI211xp5_ASAP7_75t_L     g05358(.A1(new_n5609), .A2(new_n5610), .B(new_n5613), .C(new_n5614), .Y(new_n5615));
  NAND2xp33_ASAP7_75t_L     g05359(.A(new_n5612), .B(new_n5615), .Y(new_n5616));
  NOR2xp33_ASAP7_75t_L      g05360(.A(new_n5616), .B(new_n5484), .Y(new_n5617));
  AOI22xp33_ASAP7_75t_L     g05361(.A1(new_n5612), .A2(new_n5615), .B1(new_n5483), .B2(new_n5376), .Y(new_n5618));
  NOR3xp33_ASAP7_75t_L      g05362(.A(new_n5617), .B(new_n5481), .C(new_n5618), .Y(new_n5619));
  XNOR2x2_ASAP7_75t_L       g05363(.A(\a[17] ), .B(new_n5480), .Y(new_n5620));
  NAND4xp25_ASAP7_75t_L     g05364(.A(new_n5376), .B(new_n5615), .C(new_n5612), .D(new_n5483), .Y(new_n5621));
  NAND2xp33_ASAP7_75t_L     g05365(.A(new_n5616), .B(new_n5484), .Y(new_n5622));
  AOI21xp33_ASAP7_75t_L     g05366(.A1(new_n5622), .A2(new_n5621), .B(new_n5620), .Y(new_n5623));
  NOR3xp33_ASAP7_75t_L      g05367(.A(new_n5478), .B(new_n5619), .C(new_n5623), .Y(new_n5624));
  NAND2xp33_ASAP7_75t_L     g05368(.A(new_n5376), .B(new_n5375), .Y(new_n5625));
  MAJIxp5_ASAP7_75t_L       g05369(.A(new_n5384), .B(new_n5625), .C(new_n5377), .Y(new_n5626));
  NAND3xp33_ASAP7_75t_L     g05370(.A(new_n5622), .B(new_n5620), .C(new_n5621), .Y(new_n5627));
  OAI21xp33_ASAP7_75t_L     g05371(.A1(new_n5618), .A2(new_n5617), .B(new_n5481), .Y(new_n5628));
  AOI21xp33_ASAP7_75t_L     g05372(.A1(new_n5628), .A2(new_n5627), .B(new_n5626), .Y(new_n5629));
  OAI21xp33_ASAP7_75t_L     g05373(.A1(new_n5624), .A2(new_n5629), .B(new_n5476), .Y(new_n5630));
  INVx1_ASAP7_75t_L         g05374(.A(new_n5476), .Y(new_n5631));
  NAND3xp33_ASAP7_75t_L     g05375(.A(new_n5626), .B(new_n5627), .C(new_n5628), .Y(new_n5632));
  OAI21xp33_ASAP7_75t_L     g05376(.A1(new_n5619), .A2(new_n5623), .B(new_n5478), .Y(new_n5633));
  NAND3xp33_ASAP7_75t_L     g05377(.A(new_n5632), .B(new_n5631), .C(new_n5633), .Y(new_n5634));
  NAND3xp33_ASAP7_75t_L     g05378(.A(new_n5468), .B(new_n5630), .C(new_n5634), .Y(new_n5635));
  NOR2xp33_ASAP7_75t_L      g05379(.A(new_n5389), .B(new_n5388), .Y(new_n5636));
  MAJIxp5_ASAP7_75t_L       g05380(.A(new_n5210), .B(new_n5387), .C(new_n5636), .Y(new_n5637));
  AOI21xp33_ASAP7_75t_L     g05381(.A1(new_n5632), .A2(new_n5633), .B(new_n5631), .Y(new_n5638));
  NOR3xp33_ASAP7_75t_L      g05382(.A(new_n5629), .B(new_n5624), .C(new_n5476), .Y(new_n5639));
  OAI21xp33_ASAP7_75t_L     g05383(.A1(new_n5638), .A2(new_n5639), .B(new_n5637), .Y(new_n5640));
  AOI21xp33_ASAP7_75t_L     g05384(.A1(new_n5635), .A2(new_n5640), .B(new_n5463), .Y(new_n5641));
  NOR3xp33_ASAP7_75t_L      g05385(.A(new_n5637), .B(new_n5638), .C(new_n5639), .Y(new_n5642));
  AOI221xp5_ASAP7_75t_L     g05386(.A1(new_n5210), .A2(new_n5404), .B1(new_n5634), .B2(new_n5630), .C(new_n5466), .Y(new_n5643));
  NOR3xp33_ASAP7_75t_L      g05387(.A(new_n5642), .B(new_n5462), .C(new_n5643), .Y(new_n5644));
  OR3x1_ASAP7_75t_L         g05388(.A(new_n5455), .B(new_n5641), .C(new_n5644), .Y(new_n5645));
  OAI21xp33_ASAP7_75t_L     g05389(.A1(new_n5644), .A2(new_n5641), .B(new_n5455), .Y(new_n5646));
  NAND2xp33_ASAP7_75t_L     g05390(.A(\b[33] ), .B(new_n480), .Y(new_n5647));
  NAND2xp33_ASAP7_75t_L     g05391(.A(\b[34] ), .B(new_n441), .Y(new_n5648));
  AND2x2_ASAP7_75t_L        g05392(.A(new_n4059), .B(new_n4056), .Y(new_n5649));
  AOI22xp33_ASAP7_75t_L     g05393(.A1(new_n451), .A2(\b[35] ), .B1(new_n448), .B2(new_n5649), .Y(new_n5650));
  NAND3xp33_ASAP7_75t_L     g05394(.A(new_n5650), .B(new_n5648), .C(new_n5647), .Y(new_n5651));
  XNOR2x2_ASAP7_75t_L       g05395(.A(\a[8] ), .B(new_n5651), .Y(new_n5652));
  NAND3xp33_ASAP7_75t_L     g05396(.A(new_n5645), .B(new_n5652), .C(new_n5646), .Y(new_n5653));
  AO21x2_ASAP7_75t_L        g05397(.A1(new_n5646), .A2(new_n5645), .B(new_n5652), .Y(new_n5654));
  AOI21xp33_ASAP7_75t_L     g05398(.A1(new_n5653), .A2(new_n5654), .B(new_n5454), .Y(new_n5655));
  INVx1_ASAP7_75t_L         g05399(.A(new_n5454), .Y(new_n5656));
  NAND2xp33_ASAP7_75t_L     g05400(.A(new_n5653), .B(new_n5654), .Y(new_n5657));
  NOR2xp33_ASAP7_75t_L      g05401(.A(new_n5657), .B(new_n5656), .Y(new_n5658));
  NOR3xp33_ASAP7_75t_L      g05402(.A(new_n5658), .B(new_n5452), .C(new_n5655), .Y(new_n5659));
  INVx1_ASAP7_75t_L         g05403(.A(new_n5659), .Y(new_n5660));
  OAI21xp33_ASAP7_75t_L     g05404(.A1(new_n5655), .A2(new_n5658), .B(new_n5452), .Y(new_n5661));
  AOI21xp33_ASAP7_75t_L     g05405(.A1(new_n5660), .A2(new_n5661), .B(new_n5445), .Y(new_n5662));
  AND3x1_ASAP7_75t_L        g05406(.A(new_n5660), .B(new_n5661), .C(new_n5445), .Y(new_n5663));
  A2O1A1O1Ixp25_ASAP7_75t_L g05407(.A1(new_n5168), .A2(new_n5172), .B(new_n5167), .C(new_n5188), .D(new_n5187), .Y(new_n5664));
  NOR2xp33_ASAP7_75t_L      g05408(.A(\b[40] ), .B(\b[41] ), .Y(new_n5665));
  INVx1_ASAP7_75t_L         g05409(.A(\b[41] ), .Y(new_n5666));
  NOR2xp33_ASAP7_75t_L      g05410(.A(new_n5186), .B(new_n5666), .Y(new_n5667));
  NOR2xp33_ASAP7_75t_L      g05411(.A(new_n5665), .B(new_n5667), .Y(new_n5668));
  XNOR2x2_ASAP7_75t_L       g05412(.A(new_n5668), .B(new_n5664), .Y(new_n5669));
  AOI22xp33_ASAP7_75t_L     g05413(.A1(new_n272), .A2(\b[41] ), .B1(new_n269), .B2(new_n5669), .Y(new_n5670));
  OAI221xp5_ASAP7_75t_L     g05414(.A1(new_n261), .A2(new_n5186), .B1(new_n5166), .B2(new_n277), .C(new_n5670), .Y(new_n5671));
  XNOR2x2_ASAP7_75t_L       g05415(.A(\a[2] ), .B(new_n5671), .Y(new_n5672));
  OAI21xp33_ASAP7_75t_L     g05416(.A1(new_n5662), .A2(new_n5663), .B(new_n5672), .Y(new_n5673));
  NOR3xp33_ASAP7_75t_L      g05417(.A(new_n5663), .B(new_n5672), .C(new_n5662), .Y(new_n5674));
  INVx1_ASAP7_75t_L         g05418(.A(new_n5674), .Y(new_n5675));
  NAND2xp33_ASAP7_75t_L     g05419(.A(new_n5673), .B(new_n5675), .Y(new_n5676));
  XOR2x2_ASAP7_75t_L        g05420(.A(new_n5676), .B(new_n5443), .Y(\f[41] ));
  INVx1_ASAP7_75t_L         g05421(.A(new_n5664), .Y(new_n5678));
  NOR2xp33_ASAP7_75t_L      g05422(.A(\b[41] ), .B(\b[42] ), .Y(new_n5679));
  INVx1_ASAP7_75t_L         g05423(.A(\b[42] ), .Y(new_n5680));
  NOR2xp33_ASAP7_75t_L      g05424(.A(new_n5666), .B(new_n5680), .Y(new_n5681));
  NOR2xp33_ASAP7_75t_L      g05425(.A(new_n5679), .B(new_n5681), .Y(new_n5682));
  A2O1A1Ixp33_ASAP7_75t_L   g05426(.A1(new_n5678), .A2(new_n5668), .B(new_n5667), .C(new_n5682), .Y(new_n5683));
  INVx1_ASAP7_75t_L         g05427(.A(new_n5667), .Y(new_n5684));
  A2O1A1Ixp33_ASAP7_75t_L   g05428(.A1(new_n5192), .A2(new_n5188), .B(new_n5187), .C(new_n5668), .Y(new_n5685));
  OAI211xp5_ASAP7_75t_L     g05429(.A1(new_n5679), .A2(new_n5681), .B(new_n5685), .C(new_n5684), .Y(new_n5686));
  NAND2xp33_ASAP7_75t_L     g05430(.A(new_n5683), .B(new_n5686), .Y(new_n5687));
  INVx1_ASAP7_75t_L         g05431(.A(new_n5687), .Y(new_n5688));
  AOI22xp33_ASAP7_75t_L     g05432(.A1(new_n272), .A2(\b[42] ), .B1(new_n269), .B2(new_n5688), .Y(new_n5689));
  OAI221xp5_ASAP7_75t_L     g05433(.A1(new_n261), .A2(new_n5666), .B1(new_n5186), .B2(new_n277), .C(new_n5689), .Y(new_n5690));
  XNOR2x2_ASAP7_75t_L       g05434(.A(\a[2] ), .B(new_n5690), .Y(new_n5691));
  NAND2xp33_ASAP7_75t_L     g05435(.A(\b[38] ), .B(new_n334), .Y(new_n5692));
  AOI22xp33_ASAP7_75t_L     g05436(.A1(new_n345), .A2(\b[39] ), .B1(new_n342), .B2(new_n5174), .Y(new_n5693));
  NAND2xp33_ASAP7_75t_L     g05437(.A(new_n5692), .B(new_n5693), .Y(new_n5694));
  AOI211xp5_ASAP7_75t_L     g05438(.A1(\b[37] ), .A2(new_n366), .B(new_n339), .C(new_n5694), .Y(new_n5695));
  INVx1_ASAP7_75t_L         g05439(.A(new_n5695), .Y(new_n5696));
  A2O1A1Ixp33_ASAP7_75t_L   g05440(.A1(\b[37] ), .A2(new_n366), .B(new_n5694), .C(new_n339), .Y(new_n5697));
  NAND2xp33_ASAP7_75t_L     g05441(.A(new_n5697), .B(new_n5696), .Y(new_n5698));
  NAND2xp33_ASAP7_75t_L     g05442(.A(new_n5646), .B(new_n5645), .Y(new_n5699));
  MAJIxp5_ASAP7_75t_L       g05443(.A(new_n5454), .B(new_n5652), .C(new_n5699), .Y(new_n5700));
  NAND2xp33_ASAP7_75t_L     g05444(.A(\b[34] ), .B(new_n480), .Y(new_n5701));
  NAND2xp33_ASAP7_75t_L     g05445(.A(\b[35] ), .B(new_n441), .Y(new_n5702));
  AOI22xp33_ASAP7_75t_L     g05446(.A1(new_n451), .A2(\b[36] ), .B1(new_n448), .B2(new_n4473), .Y(new_n5703));
  AND4x1_ASAP7_75t_L        g05447(.A(new_n5703), .B(new_n5702), .C(new_n5701), .D(\a[8] ), .Y(new_n5704));
  AOI31xp33_ASAP7_75t_L     g05448(.A1(new_n5703), .A2(new_n5702), .A3(new_n5701), .B(\a[8] ), .Y(new_n5705));
  NOR2xp33_ASAP7_75t_L      g05449(.A(new_n5705), .B(new_n5704), .Y(new_n5706));
  OAI21xp33_ASAP7_75t_L     g05450(.A1(new_n5643), .A2(new_n5642), .B(new_n5462), .Y(new_n5707));
  A2O1A1O1Ixp25_ASAP7_75t_L g05451(.A1(new_n5401), .A2(new_n5208), .B(new_n5412), .C(new_n5707), .D(new_n5644), .Y(new_n5708));
  A2O1A1O1Ixp25_ASAP7_75t_L g05452(.A1(new_n5210), .A2(new_n5404), .B(new_n5466), .C(new_n5630), .D(new_n5639), .Y(new_n5709));
  NOR2xp33_ASAP7_75t_L      g05453(.A(new_n2852), .B(new_n909), .Y(new_n5710));
  INVx1_ASAP7_75t_L         g05454(.A(new_n5710), .Y(new_n5711));
  NAND2xp33_ASAP7_75t_L     g05455(.A(\b[29] ), .B(new_n817), .Y(new_n5712));
  AOI22xp33_ASAP7_75t_L     g05456(.A1(new_n826), .A2(\b[30] ), .B1(new_n823), .B2(new_n3219), .Y(new_n5713));
  AND4x1_ASAP7_75t_L        g05457(.A(new_n5713), .B(new_n5712), .C(new_n5711), .D(\a[14] ), .Y(new_n5714));
  AOI31xp33_ASAP7_75t_L     g05458(.A1(new_n5713), .A2(new_n5712), .A3(new_n5711), .B(\a[14] ), .Y(new_n5715));
  NOR2xp33_ASAP7_75t_L      g05459(.A(new_n5715), .B(new_n5714), .Y(new_n5716));
  NAND2xp33_ASAP7_75t_L     g05460(.A(new_n5382), .B(new_n5383), .Y(new_n5717));
  NOR2xp33_ASAP7_75t_L      g05461(.A(new_n5377), .B(new_n5625), .Y(new_n5718));
  A2O1A1O1Ixp25_ASAP7_75t_L g05462(.A1(new_n5380), .A2(new_n5717), .B(new_n5718), .C(new_n5627), .D(new_n5623), .Y(new_n5719));
  OAI21xp33_ASAP7_75t_L     g05463(.A1(new_n5566), .A2(new_n5495), .B(new_n5576), .Y(new_n5720));
  NAND2xp33_ASAP7_75t_L     g05464(.A(\b[13] ), .B(new_n2931), .Y(new_n5721));
  NAND2xp33_ASAP7_75t_L     g05465(.A(\b[14] ), .B(new_n2706), .Y(new_n5722));
  AOI22xp33_ASAP7_75t_L     g05466(.A1(new_n2702), .A2(\b[15] ), .B1(new_n2700), .B2(new_n959), .Y(new_n5723));
  NAND4xp25_ASAP7_75t_L     g05467(.A(new_n5723), .B(\a[29] ), .C(new_n5721), .D(new_n5722), .Y(new_n5724));
  OAI221xp5_ASAP7_75t_L     g05468(.A1(new_n2708), .A2(new_n952), .B1(new_n2707), .B2(new_n2573), .C(new_n5722), .Y(new_n5725));
  A2O1A1Ixp33_ASAP7_75t_L   g05469(.A1(\b[13] ), .A2(new_n2931), .B(new_n5725), .C(new_n2697), .Y(new_n5726));
  AND2x2_ASAP7_75t_L        g05470(.A(new_n5724), .B(new_n5726), .Y(new_n5727));
  A2O1A1O1Ixp25_ASAP7_75t_L g05471(.A1(new_n5291), .A2(new_n5297), .B(new_n5299), .C(new_n5555), .D(new_n5563), .Y(new_n5728));
  NOR2xp33_ASAP7_75t_L      g05472(.A(new_n631), .B(new_n3492), .Y(new_n5729));
  NAND2xp33_ASAP7_75t_L     g05473(.A(\b[11] ), .B(new_n3260), .Y(new_n5730));
  OAI221xp5_ASAP7_75t_L     g05474(.A1(new_n3262), .A2(new_n763), .B1(new_n3261), .B2(new_n775), .C(new_n5730), .Y(new_n5731));
  OR3x1_ASAP7_75t_L         g05475(.A(new_n5731), .B(new_n3251), .C(new_n5729), .Y(new_n5732));
  A2O1A1Ixp33_ASAP7_75t_L   g05476(.A1(\b[10] ), .A2(new_n3491), .B(new_n5731), .C(new_n3251), .Y(new_n5733));
  NAND2xp33_ASAP7_75t_L     g05477(.A(new_n5733), .B(new_n5732), .Y(new_n5734));
  AOI211xp5_ASAP7_75t_L     g05478(.A1(new_n5512), .A2(new_n5510), .B(new_n5539), .C(new_n5538), .Y(new_n5735));
  A2O1A1O1Ixp25_ASAP7_75t_L g05479(.A1(new_n5280), .A2(new_n5277), .B(new_n5543), .C(new_n5547), .D(new_n5735), .Y(new_n5736));
  NAND2xp33_ASAP7_75t_L     g05480(.A(\b[0] ), .B(new_n5240), .Y(new_n5737));
  NAND2xp33_ASAP7_75t_L     g05481(.A(new_n271), .B(new_n5247), .Y(new_n5738));
  NAND2xp33_ASAP7_75t_L     g05482(.A(\b[1] ), .B(new_n5249), .Y(new_n5739));
  NAND5xp2_ASAP7_75t_L      g05483(.A(new_n5739), .B(new_n5738), .C(new_n5737), .D(new_n5228), .E(\a[41] ), .Y(new_n5740));
  INVx1_ASAP7_75t_L         g05484(.A(\a[42] ), .Y(new_n5741));
  NAND2xp33_ASAP7_75t_L     g05485(.A(\a[41] ), .B(new_n5741), .Y(new_n5742));
  NAND2xp33_ASAP7_75t_L     g05486(.A(\a[42] ), .B(new_n5244), .Y(new_n5743));
  AND2x2_ASAP7_75t_L        g05487(.A(new_n5742), .B(new_n5743), .Y(new_n5744));
  NOR2xp33_ASAP7_75t_L      g05488(.A(new_n258), .B(new_n5744), .Y(new_n5745));
  OAI31xp33_ASAP7_75t_L     g05489(.A1(new_n5740), .A2(new_n5524), .A3(new_n5522), .B(new_n5745), .Y(new_n5746));
  OR4x2_ASAP7_75t_L         g05490(.A(new_n5745), .B(new_n5740), .C(new_n5524), .D(new_n5522), .Y(new_n5747));
  NOR2xp33_ASAP7_75t_L      g05491(.A(new_n276), .B(new_n5521), .Y(new_n5748));
  NAND2xp33_ASAP7_75t_L     g05492(.A(\b[3] ), .B(new_n5249), .Y(new_n5749));
  OAI221xp5_ASAP7_75t_L     g05493(.A1(new_n278), .A2(new_n5241), .B1(new_n5252), .B2(new_n303), .C(new_n5749), .Y(new_n5750));
  OR3x1_ASAP7_75t_L         g05494(.A(new_n5750), .B(new_n5244), .C(new_n5748), .Y(new_n5751));
  A2O1A1Ixp33_ASAP7_75t_L   g05495(.A1(\b[1] ), .A2(new_n5526), .B(new_n5750), .C(new_n5244), .Y(new_n5752));
  AO22x1_ASAP7_75t_L        g05496(.A1(new_n5752), .A2(new_n5751), .B1(new_n5746), .B2(new_n5747), .Y(new_n5753));
  NAND4xp25_ASAP7_75t_L     g05497(.A(new_n5747), .B(new_n5746), .C(new_n5751), .D(new_n5752), .Y(new_n5754));
  NAND2xp33_ASAP7_75t_L     g05498(.A(\b[4] ), .B(new_n4780), .Y(new_n5755));
  NAND2xp33_ASAP7_75t_L     g05499(.A(\b[5] ), .B(new_n4548), .Y(new_n5756));
  AOI22xp33_ASAP7_75t_L     g05500(.A1(new_n4544), .A2(\b[6] ), .B1(new_n4542), .B2(new_n389), .Y(new_n5757));
  NAND4xp25_ASAP7_75t_L     g05501(.A(new_n5757), .B(\a[38] ), .C(new_n5755), .D(new_n5756), .Y(new_n5758));
  OAI221xp5_ASAP7_75t_L     g05502(.A1(new_n4550), .A2(new_n382), .B1(new_n4549), .B2(new_n540), .C(new_n5756), .Y(new_n5759));
  A2O1A1Ixp33_ASAP7_75t_L   g05503(.A1(\b[4] ), .A2(new_n4780), .B(new_n5759), .C(new_n4539), .Y(new_n5760));
  NAND4xp25_ASAP7_75t_L     g05504(.A(new_n5760), .B(new_n5753), .C(new_n5754), .D(new_n5758), .Y(new_n5761));
  AOI22xp33_ASAP7_75t_L     g05505(.A1(new_n5751), .A2(new_n5752), .B1(new_n5746), .B2(new_n5747), .Y(new_n5762));
  AND4x1_ASAP7_75t_L        g05506(.A(new_n5747), .B(new_n5746), .C(new_n5752), .D(new_n5751), .Y(new_n5763));
  AOI211xp5_ASAP7_75t_L     g05507(.A1(\b[4] ), .A2(new_n4780), .B(new_n4539), .C(new_n5759), .Y(new_n5764));
  AOI31xp33_ASAP7_75t_L     g05508(.A1(new_n5757), .A2(new_n5756), .A3(new_n5755), .B(\a[38] ), .Y(new_n5765));
  OAI22xp33_ASAP7_75t_L     g05509(.A1(new_n5764), .A2(new_n5765), .B1(new_n5762), .B2(new_n5763), .Y(new_n5766));
  NAND2xp33_ASAP7_75t_L     g05510(.A(new_n5761), .B(new_n5766), .Y(new_n5767));
  NAND2xp33_ASAP7_75t_L     g05511(.A(new_n5517), .B(new_n5519), .Y(new_n5768));
  INVx1_ASAP7_75t_L         g05512(.A(new_n5524), .Y(new_n5769));
  OAI21xp33_ASAP7_75t_L     g05513(.A1(new_n258), .A2(new_n5521), .B(new_n5769), .Y(new_n5770));
  NOR2xp33_ASAP7_75t_L      g05514(.A(new_n5520), .B(new_n5770), .Y(new_n5771));
  INVx1_ASAP7_75t_L         g05515(.A(new_n5527), .Y(new_n5772));
  NOR2xp33_ASAP7_75t_L      g05516(.A(new_n5772), .B(new_n5771), .Y(new_n5773));
  NAND2xp33_ASAP7_75t_L     g05517(.A(new_n5768), .B(new_n5773), .Y(new_n5774));
  A2O1A1Ixp33_ASAP7_75t_L   g05518(.A1(new_n5528), .A2(new_n5529), .B(new_n5534), .C(new_n5774), .Y(new_n5775));
  NOR2xp33_ASAP7_75t_L      g05519(.A(new_n5767), .B(new_n5775), .Y(new_n5776));
  MAJIxp5_ASAP7_75t_L       g05520(.A(new_n5513), .B(new_n5768), .C(new_n5773), .Y(new_n5777));
  AOI21xp33_ASAP7_75t_L     g05521(.A1(new_n5766), .A2(new_n5761), .B(new_n5777), .Y(new_n5778));
  NOR2xp33_ASAP7_75t_L      g05522(.A(new_n421), .B(new_n4986), .Y(new_n5779));
  INVx1_ASAP7_75t_L         g05523(.A(new_n5779), .Y(new_n5780));
  NAND2xp33_ASAP7_75t_L     g05524(.A(\b[8] ), .B(new_n3874), .Y(new_n5781));
  AOI22xp33_ASAP7_75t_L     g05525(.A1(new_n3884), .A2(\b[9] ), .B1(new_n3881), .B2(new_n566), .Y(new_n5782));
  NAND4xp25_ASAP7_75t_L     g05526(.A(new_n5782), .B(\a[35] ), .C(new_n5780), .D(new_n5781), .Y(new_n5783));
  OAI221xp5_ASAP7_75t_L     g05527(.A1(new_n4115), .A2(new_n559), .B1(new_n4114), .B2(new_n978), .C(new_n5781), .Y(new_n5784));
  A2O1A1Ixp33_ASAP7_75t_L   g05528(.A1(\b[7] ), .A2(new_n4111), .B(new_n5784), .C(new_n3878), .Y(new_n5785));
  OAI211xp5_ASAP7_75t_L     g05529(.A1(new_n5778), .A2(new_n5776), .B(new_n5783), .C(new_n5785), .Y(new_n5786));
  NAND3xp33_ASAP7_75t_L     g05530(.A(new_n5777), .B(new_n5766), .C(new_n5761), .Y(new_n5787));
  NAND2xp33_ASAP7_75t_L     g05531(.A(new_n5767), .B(new_n5775), .Y(new_n5788));
  NOR3xp33_ASAP7_75t_L      g05532(.A(new_n5784), .B(new_n5779), .C(new_n3878), .Y(new_n5789));
  AOI31xp33_ASAP7_75t_L     g05533(.A1(new_n5782), .A2(new_n5781), .A3(new_n5780), .B(\a[35] ), .Y(new_n5790));
  OAI211xp5_ASAP7_75t_L     g05534(.A1(new_n5790), .A2(new_n5789), .B(new_n5788), .C(new_n5787), .Y(new_n5791));
  NAND2xp33_ASAP7_75t_L     g05535(.A(new_n5791), .B(new_n5786), .Y(new_n5792));
  NOR2xp33_ASAP7_75t_L      g05536(.A(new_n5736), .B(new_n5792), .Y(new_n5793));
  AOI221xp5_ASAP7_75t_L     g05537(.A1(new_n5505), .A2(new_n5547), .B1(new_n5791), .B2(new_n5786), .C(new_n5735), .Y(new_n5794));
  OAI21xp33_ASAP7_75t_L     g05538(.A1(new_n5794), .A2(new_n5793), .B(new_n5734), .Y(new_n5795));
  INVx1_ASAP7_75t_L         g05539(.A(new_n5735), .Y(new_n5796));
  A2O1A1Ixp33_ASAP7_75t_L   g05540(.A1(new_n5293), .A2(new_n5504), .B(new_n5541), .C(new_n5796), .Y(new_n5797));
  AOI211xp5_ASAP7_75t_L     g05541(.A1(new_n5788), .A2(new_n5787), .B(new_n5789), .C(new_n5790), .Y(new_n5798));
  AOI211xp5_ASAP7_75t_L     g05542(.A1(new_n5783), .A2(new_n5785), .B(new_n5778), .C(new_n5776), .Y(new_n5799));
  NOR2xp33_ASAP7_75t_L      g05543(.A(new_n5799), .B(new_n5798), .Y(new_n5800));
  NAND2xp33_ASAP7_75t_L     g05544(.A(new_n5797), .B(new_n5800), .Y(new_n5801));
  NAND2xp33_ASAP7_75t_L     g05545(.A(new_n5736), .B(new_n5792), .Y(new_n5802));
  NAND4xp25_ASAP7_75t_L     g05546(.A(new_n5801), .B(new_n5802), .C(new_n5732), .D(new_n5733), .Y(new_n5803));
  AO21x2_ASAP7_75t_L        g05547(.A1(new_n5803), .A2(new_n5795), .B(new_n5728), .Y(new_n5804));
  NAND3xp33_ASAP7_75t_L     g05548(.A(new_n5728), .B(new_n5795), .C(new_n5803), .Y(new_n5805));
  NAND3xp33_ASAP7_75t_L     g05549(.A(new_n5727), .B(new_n5804), .C(new_n5805), .Y(new_n5806));
  NAND2xp33_ASAP7_75t_L     g05550(.A(new_n5724), .B(new_n5726), .Y(new_n5807));
  AOI21xp33_ASAP7_75t_L     g05551(.A1(new_n5795), .A2(new_n5803), .B(new_n5728), .Y(new_n5808));
  AND3x1_ASAP7_75t_L        g05552(.A(new_n5728), .B(new_n5795), .C(new_n5803), .Y(new_n5809));
  OAI21xp33_ASAP7_75t_L     g05553(.A1(new_n5808), .A2(new_n5809), .B(new_n5807), .Y(new_n5810));
  NAND3xp33_ASAP7_75t_L     g05554(.A(new_n5720), .B(new_n5810), .C(new_n5806), .Y(new_n5811));
  A2O1A1O1Ixp25_ASAP7_75t_L g05555(.A1(new_n5301), .A2(new_n5219), .B(new_n5312), .C(new_n5575), .D(new_n5572), .Y(new_n5812));
  NOR3xp33_ASAP7_75t_L      g05556(.A(new_n5809), .B(new_n5808), .C(new_n5807), .Y(new_n5813));
  AOI21xp33_ASAP7_75t_L     g05557(.A1(new_n5804), .A2(new_n5805), .B(new_n5727), .Y(new_n5814));
  OAI21xp33_ASAP7_75t_L     g05558(.A1(new_n5813), .A2(new_n5814), .B(new_n5812), .Y(new_n5815));
  NAND2xp33_ASAP7_75t_L     g05559(.A(\b[16] ), .B(new_n2386), .Y(new_n5816));
  NAND2xp33_ASAP7_75t_L     g05560(.A(\b[17] ), .B(new_n2232), .Y(new_n5817));
  AOI22xp33_ASAP7_75t_L     g05561(.A1(new_n2228), .A2(\b[18] ), .B1(new_n2226), .B2(new_n1363), .Y(new_n5818));
  NAND4xp25_ASAP7_75t_L     g05562(.A(new_n5818), .B(\a[26] ), .C(new_n5816), .D(new_n5817), .Y(new_n5819));
  OAI221xp5_ASAP7_75t_L     g05563(.A1(new_n2234), .A2(new_n1356), .B1(new_n2233), .B2(new_n3138), .C(new_n5817), .Y(new_n5820));
  A2O1A1Ixp33_ASAP7_75t_L   g05564(.A1(\b[16] ), .A2(new_n2386), .B(new_n5820), .C(new_n2223), .Y(new_n5821));
  AND2x2_ASAP7_75t_L        g05565(.A(new_n5819), .B(new_n5821), .Y(new_n5822));
  AOI21xp33_ASAP7_75t_L     g05566(.A1(new_n5811), .A2(new_n5815), .B(new_n5822), .Y(new_n5823));
  NOR3xp33_ASAP7_75t_L      g05567(.A(new_n5812), .B(new_n5813), .C(new_n5814), .Y(new_n5824));
  AOI21xp33_ASAP7_75t_L     g05568(.A1(new_n5810), .A2(new_n5806), .B(new_n5720), .Y(new_n5825));
  NAND2xp33_ASAP7_75t_L     g05569(.A(new_n5819), .B(new_n5821), .Y(new_n5826));
  NOR3xp33_ASAP7_75t_L      g05570(.A(new_n5824), .B(new_n5825), .C(new_n5826), .Y(new_n5827));
  NOR2xp33_ASAP7_75t_L      g05571(.A(new_n5823), .B(new_n5827), .Y(new_n5828));
  A2O1A1Ixp33_ASAP7_75t_L   g05572(.A1(new_n5590), .A2(new_n5587), .B(new_n5589), .C(new_n5828), .Y(new_n5829));
  NOR2xp33_ASAP7_75t_L      g05573(.A(new_n5319), .B(new_n5586), .Y(new_n5830));
  A2O1A1O1Ixp25_ASAP7_75t_L g05574(.A1(new_n5339), .A2(new_n5329), .B(new_n5830), .C(new_n5578), .D(new_n5589), .Y(new_n5831));
  OAI21xp33_ASAP7_75t_L     g05575(.A1(new_n5825), .A2(new_n5824), .B(new_n5826), .Y(new_n5832));
  NAND3xp33_ASAP7_75t_L     g05576(.A(new_n5822), .B(new_n5811), .C(new_n5815), .Y(new_n5833));
  NAND2xp33_ASAP7_75t_L     g05577(.A(new_n5833), .B(new_n5832), .Y(new_n5834));
  NAND2xp33_ASAP7_75t_L     g05578(.A(new_n5831), .B(new_n5834), .Y(new_n5835));
  NOR2xp33_ASAP7_75t_L      g05579(.A(new_n1493), .B(new_n1911), .Y(new_n5836));
  INVx1_ASAP7_75t_L         g05580(.A(new_n5836), .Y(new_n5837));
  NAND2xp33_ASAP7_75t_L     g05581(.A(\b[20] ), .B(new_n1770), .Y(new_n5838));
  AOI22xp33_ASAP7_75t_L     g05582(.A1(new_n1766), .A2(\b[21] ), .B1(new_n1764), .B2(new_n1715), .Y(new_n5839));
  AND4x1_ASAP7_75t_L        g05583(.A(new_n5839), .B(new_n5838), .C(new_n5837), .D(\a[23] ), .Y(new_n5840));
  AOI31xp33_ASAP7_75t_L     g05584(.A1(new_n5839), .A2(new_n5838), .A3(new_n5837), .B(\a[23] ), .Y(new_n5841));
  NOR2xp33_ASAP7_75t_L      g05585(.A(new_n5841), .B(new_n5840), .Y(new_n5842));
  NAND3xp33_ASAP7_75t_L     g05586(.A(new_n5829), .B(new_n5835), .C(new_n5842), .Y(new_n5843));
  NOR2xp33_ASAP7_75t_L      g05587(.A(new_n5831), .B(new_n5834), .Y(new_n5844));
  AOI221xp5_ASAP7_75t_L     g05588(.A1(new_n5833), .A2(new_n5832), .B1(new_n5590), .B2(new_n5587), .C(new_n5589), .Y(new_n5845));
  INVx1_ASAP7_75t_L         g05589(.A(new_n5842), .Y(new_n5846));
  OAI21xp33_ASAP7_75t_L     g05590(.A1(new_n5845), .A2(new_n5844), .B(new_n5846), .Y(new_n5847));
  AND2x2_ASAP7_75t_L        g05591(.A(new_n5847), .B(new_n5843), .Y(new_n5848));
  AOI211xp5_ASAP7_75t_L     g05592(.A1(new_n5597), .A2(new_n5595), .B(new_n5585), .C(new_n5591), .Y(new_n5849));
  O2A1O1Ixp33_ASAP7_75t_L   g05593(.A1(new_n5599), .A2(new_n5600), .B(new_n5602), .C(new_n5849), .Y(new_n5850));
  NAND2xp33_ASAP7_75t_L     g05594(.A(new_n5850), .B(new_n5848), .Y(new_n5851));
  OR3x1_ASAP7_75t_L         g05595(.A(new_n5591), .B(new_n5585), .C(new_n5598), .Y(new_n5852));
  OAI21xp33_ASAP7_75t_L     g05596(.A1(new_n5585), .A2(new_n5591), .B(new_n5598), .Y(new_n5853));
  NAND2xp33_ASAP7_75t_L     g05597(.A(new_n5853), .B(new_n5852), .Y(new_n5854));
  NAND2xp33_ASAP7_75t_L     g05598(.A(new_n5847), .B(new_n5843), .Y(new_n5855));
  A2O1A1Ixp33_ASAP7_75t_L   g05599(.A1(new_n5854), .A2(new_n5602), .B(new_n5849), .C(new_n5855), .Y(new_n5856));
  NAND2xp33_ASAP7_75t_L     g05600(.A(\b[22] ), .B(new_n1548), .Y(new_n5857));
  NAND2xp33_ASAP7_75t_L     g05601(.A(\b[23] ), .B(new_n1410), .Y(new_n5858));
  AOI22xp33_ASAP7_75t_L     g05602(.A1(new_n1406), .A2(\b[24] ), .B1(new_n1404), .B2(new_n2027), .Y(new_n5859));
  NAND4xp25_ASAP7_75t_L     g05603(.A(new_n5859), .B(\a[20] ), .C(new_n5857), .D(new_n5858), .Y(new_n5860));
  NAND2xp33_ASAP7_75t_L     g05604(.A(new_n5858), .B(new_n5859), .Y(new_n5861));
  A2O1A1Ixp33_ASAP7_75t_L   g05605(.A1(\b[22] ), .A2(new_n1548), .B(new_n5861), .C(new_n1401), .Y(new_n5862));
  NAND2xp33_ASAP7_75t_L     g05606(.A(new_n5860), .B(new_n5862), .Y(new_n5863));
  AOI21xp33_ASAP7_75t_L     g05607(.A1(new_n5851), .A2(new_n5856), .B(new_n5863), .Y(new_n5864));
  NOR3xp33_ASAP7_75t_L      g05608(.A(new_n5604), .B(new_n5855), .C(new_n5849), .Y(new_n5865));
  NOR2xp33_ASAP7_75t_L      g05609(.A(new_n5850), .B(new_n5848), .Y(new_n5866));
  AND2x2_ASAP7_75t_L        g05610(.A(new_n5860), .B(new_n5862), .Y(new_n5867));
  NOR3xp33_ASAP7_75t_L      g05611(.A(new_n5866), .B(new_n5867), .C(new_n5865), .Y(new_n5868));
  A2O1A1Ixp33_ASAP7_75t_L   g05612(.A1(new_n5361), .A2(new_n5359), .B(new_n5482), .C(new_n5612), .Y(new_n5869));
  AO211x2_ASAP7_75t_L       g05613(.A1(new_n5869), .A2(new_n5615), .B(new_n5864), .C(new_n5868), .Y(new_n5870));
  OAI211xp5_ASAP7_75t_L     g05614(.A1(new_n5864), .A2(new_n5868), .B(new_n5615), .C(new_n5869), .Y(new_n5871));
  NAND2xp33_ASAP7_75t_L     g05615(.A(\b[25] ), .B(new_n1194), .Y(new_n5872));
  NAND2xp33_ASAP7_75t_L     g05616(.A(\b[26] ), .B(new_n1103), .Y(new_n5873));
  AOI22xp33_ASAP7_75t_L     g05617(.A1(new_n1113), .A2(\b[27] ), .B1(new_n1110), .B2(new_n2657), .Y(new_n5874));
  AND4x1_ASAP7_75t_L        g05618(.A(new_n5874), .B(new_n5873), .C(new_n5872), .D(\a[17] ), .Y(new_n5875));
  AOI31xp33_ASAP7_75t_L     g05619(.A1(new_n5874), .A2(new_n5873), .A3(new_n5872), .B(\a[17] ), .Y(new_n5876));
  NOR2xp33_ASAP7_75t_L      g05620(.A(new_n5876), .B(new_n5875), .Y(new_n5877));
  NAND3xp33_ASAP7_75t_L     g05621(.A(new_n5870), .B(new_n5877), .C(new_n5871), .Y(new_n5878));
  AOI211xp5_ASAP7_75t_L     g05622(.A1(new_n5869), .A2(new_n5615), .B(new_n5864), .C(new_n5868), .Y(new_n5879));
  INVx1_ASAP7_75t_L         g05623(.A(new_n5615), .Y(new_n5880));
  OAI21xp33_ASAP7_75t_L     g05624(.A1(new_n5865), .A2(new_n5866), .B(new_n5867), .Y(new_n5881));
  NAND3xp33_ASAP7_75t_L     g05625(.A(new_n5851), .B(new_n5856), .C(new_n5863), .Y(new_n5882));
  AOI221xp5_ASAP7_75t_L     g05626(.A1(new_n5881), .A2(new_n5882), .B1(new_n5484), .B2(new_n5612), .C(new_n5880), .Y(new_n5883));
  INVx1_ASAP7_75t_L         g05627(.A(new_n5877), .Y(new_n5884));
  OAI21xp33_ASAP7_75t_L     g05628(.A1(new_n5879), .A2(new_n5883), .B(new_n5884), .Y(new_n5885));
  AOI21xp33_ASAP7_75t_L     g05629(.A1(new_n5885), .A2(new_n5878), .B(new_n5719), .Y(new_n5886));
  NAND2xp33_ASAP7_75t_L     g05630(.A(new_n5373), .B(new_n5477), .Y(new_n5887));
  A2O1A1Ixp33_ASAP7_75t_L   g05631(.A1(new_n5381), .A2(new_n5887), .B(new_n5619), .C(new_n5628), .Y(new_n5888));
  NAND2xp33_ASAP7_75t_L     g05632(.A(new_n5885), .B(new_n5878), .Y(new_n5889));
  NOR2xp33_ASAP7_75t_L      g05633(.A(new_n5888), .B(new_n5889), .Y(new_n5890));
  NOR3xp33_ASAP7_75t_L      g05634(.A(new_n5890), .B(new_n5886), .C(new_n5716), .Y(new_n5891));
  INVx1_ASAP7_75t_L         g05635(.A(new_n5716), .Y(new_n5892));
  A2O1A1Ixp33_ASAP7_75t_L   g05636(.A1(new_n5627), .A2(new_n5626), .B(new_n5623), .C(new_n5889), .Y(new_n5893));
  NAND3xp33_ASAP7_75t_L     g05637(.A(new_n5719), .B(new_n5878), .C(new_n5885), .Y(new_n5894));
  AOI21xp33_ASAP7_75t_L     g05638(.A1(new_n5893), .A2(new_n5894), .B(new_n5892), .Y(new_n5895));
  NOR3xp33_ASAP7_75t_L      g05639(.A(new_n5709), .B(new_n5891), .C(new_n5895), .Y(new_n5896));
  NAND3xp33_ASAP7_75t_L     g05640(.A(new_n5893), .B(new_n5892), .C(new_n5894), .Y(new_n5897));
  OAI21xp33_ASAP7_75t_L     g05641(.A1(new_n5886), .A2(new_n5890), .B(new_n5716), .Y(new_n5898));
  AOI221xp5_ASAP7_75t_L     g05642(.A1(new_n5468), .A2(new_n5630), .B1(new_n5897), .B2(new_n5898), .C(new_n5639), .Y(new_n5899));
  NAND2xp33_ASAP7_75t_L     g05643(.A(\b[32] ), .B(new_n590), .Y(new_n5900));
  AOI22xp33_ASAP7_75t_L     g05644(.A1(new_n600), .A2(\b[33] ), .B1(new_n597), .B2(new_n3813), .Y(new_n5901));
  NAND2xp33_ASAP7_75t_L     g05645(.A(new_n5900), .B(new_n5901), .Y(new_n5902));
  INVx1_ASAP7_75t_L         g05646(.A(new_n5902), .Y(new_n5903));
  OAI211xp5_ASAP7_75t_L     g05647(.A1(new_n3419), .A2(new_n1620), .B(new_n5903), .C(\a[11] ), .Y(new_n5904));
  A2O1A1Ixp33_ASAP7_75t_L   g05648(.A1(\b[31] ), .A2(new_n674), .B(new_n5902), .C(new_n594), .Y(new_n5905));
  NAND2xp33_ASAP7_75t_L     g05649(.A(new_n5905), .B(new_n5904), .Y(new_n5906));
  NOR3xp33_ASAP7_75t_L      g05650(.A(new_n5906), .B(new_n5899), .C(new_n5896), .Y(new_n5907));
  INVx1_ASAP7_75t_L         g05651(.A(new_n5907), .Y(new_n5908));
  OAI21xp33_ASAP7_75t_L     g05652(.A1(new_n5638), .A2(new_n5637), .B(new_n5634), .Y(new_n5909));
  NAND3xp33_ASAP7_75t_L     g05653(.A(new_n5909), .B(new_n5897), .C(new_n5898), .Y(new_n5910));
  OAI21xp33_ASAP7_75t_L     g05654(.A1(new_n5895), .A2(new_n5891), .B(new_n5709), .Y(new_n5911));
  NAND2xp33_ASAP7_75t_L     g05655(.A(new_n5911), .B(new_n5910), .Y(new_n5912));
  NAND2xp33_ASAP7_75t_L     g05656(.A(new_n5906), .B(new_n5912), .Y(new_n5913));
  AOI21xp33_ASAP7_75t_L     g05657(.A1(new_n5913), .A2(new_n5908), .B(new_n5708), .Y(new_n5914));
  NAND3xp33_ASAP7_75t_L     g05658(.A(new_n5635), .B(new_n5463), .C(new_n5640), .Y(new_n5915));
  OAI21xp33_ASAP7_75t_L     g05659(.A1(new_n5641), .A2(new_n5455), .B(new_n5915), .Y(new_n5916));
  NOR2xp33_ASAP7_75t_L      g05660(.A(new_n5896), .B(new_n5899), .Y(new_n5917));
  INVx1_ASAP7_75t_L         g05661(.A(new_n5906), .Y(new_n5918));
  NOR2xp33_ASAP7_75t_L      g05662(.A(new_n5918), .B(new_n5917), .Y(new_n5919));
  NOR3xp33_ASAP7_75t_L      g05663(.A(new_n5919), .B(new_n5907), .C(new_n5916), .Y(new_n5920));
  OAI21xp33_ASAP7_75t_L     g05664(.A1(new_n5920), .A2(new_n5914), .B(new_n5706), .Y(new_n5921));
  NOR3xp33_ASAP7_75t_L      g05665(.A(new_n5914), .B(new_n5920), .C(new_n5706), .Y(new_n5922));
  INVx1_ASAP7_75t_L         g05666(.A(new_n5922), .Y(new_n5923));
  AND3x1_ASAP7_75t_L        g05667(.A(new_n5923), .B(new_n5921), .C(new_n5700), .Y(new_n5924));
  INVx1_ASAP7_75t_L         g05668(.A(new_n5706), .Y(new_n5925));
  OAI21xp33_ASAP7_75t_L     g05669(.A1(new_n5907), .A2(new_n5919), .B(new_n5916), .Y(new_n5926));
  NAND3xp33_ASAP7_75t_L     g05670(.A(new_n5913), .B(new_n5908), .C(new_n5708), .Y(new_n5927));
  AOI21xp33_ASAP7_75t_L     g05671(.A1(new_n5927), .A2(new_n5926), .B(new_n5925), .Y(new_n5928));
  NOR2xp33_ASAP7_75t_L      g05672(.A(new_n5928), .B(new_n5922), .Y(new_n5929));
  NOR2xp33_ASAP7_75t_L      g05673(.A(new_n5700), .B(new_n5929), .Y(new_n5930));
  OAI21xp33_ASAP7_75t_L     g05674(.A1(new_n5930), .A2(new_n5924), .B(new_n5698), .Y(new_n5931));
  AND2x2_ASAP7_75t_L        g05675(.A(new_n5697), .B(new_n5696), .Y(new_n5932));
  NAND2xp33_ASAP7_75t_L     g05676(.A(new_n5700), .B(new_n5929), .Y(new_n5933));
  AO21x2_ASAP7_75t_L        g05677(.A1(new_n5921), .A2(new_n5923), .B(new_n5700), .Y(new_n5934));
  NAND3xp33_ASAP7_75t_L     g05678(.A(new_n5934), .B(new_n5932), .C(new_n5933), .Y(new_n5935));
  NAND2xp33_ASAP7_75t_L     g05679(.A(new_n5935), .B(new_n5931), .Y(new_n5936));
  A2O1A1Ixp33_ASAP7_75t_L   g05680(.A1(new_n5661), .A2(new_n5445), .B(new_n5659), .C(new_n5936), .Y(new_n5937));
  NOR2xp33_ASAP7_75t_L      g05681(.A(new_n5427), .B(new_n5444), .Y(new_n5938));
  O2A1O1Ixp33_ASAP7_75t_L   g05682(.A1(new_n5938), .A2(new_n5430), .B(new_n5661), .C(new_n5659), .Y(new_n5939));
  NAND3xp33_ASAP7_75t_L     g05683(.A(new_n5939), .B(new_n5931), .C(new_n5935), .Y(new_n5940));
  NAND2xp33_ASAP7_75t_L     g05684(.A(new_n5937), .B(new_n5940), .Y(new_n5941));
  XNOR2x2_ASAP7_75t_L       g05685(.A(new_n5691), .B(new_n5941), .Y(new_n5942));
  O2A1O1Ixp33_ASAP7_75t_L   g05686(.A1(new_n5676), .A2(new_n5443), .B(new_n5675), .C(new_n5942), .Y(new_n5943));
  A2O1A1O1Ixp25_ASAP7_75t_L g05687(.A1(new_n5437), .A2(new_n5440), .B(new_n5433), .C(new_n5673), .D(new_n5674), .Y(new_n5944));
  AND2x2_ASAP7_75t_L        g05688(.A(new_n5944), .B(new_n5942), .Y(new_n5945));
  NOR2xp33_ASAP7_75t_L      g05689(.A(new_n5945), .B(new_n5943), .Y(\f[42] ));
  NOR3xp33_ASAP7_75t_L      g05690(.A(new_n5930), .B(new_n5924), .C(new_n5932), .Y(new_n5947));
  INVx1_ASAP7_75t_L         g05691(.A(new_n5947), .Y(new_n5948));
  A2O1A1Ixp33_ASAP7_75t_L   g05692(.A1(new_n5931), .A2(new_n5935), .B(new_n5939), .C(new_n5948), .Y(new_n5949));
  NOR2xp33_ASAP7_75t_L      g05693(.A(new_n4915), .B(new_n365), .Y(new_n5950));
  INVx1_ASAP7_75t_L         g05694(.A(new_n5950), .Y(new_n5951));
  NOR2xp33_ASAP7_75t_L      g05695(.A(new_n5166), .B(new_n406), .Y(new_n5952));
  INVx1_ASAP7_75t_L         g05696(.A(new_n5952), .Y(new_n5953));
  AOI22xp33_ASAP7_75t_L     g05697(.A1(new_n345), .A2(\b[40] ), .B1(new_n342), .B2(new_n5194), .Y(new_n5954));
  AND4x1_ASAP7_75t_L        g05698(.A(new_n5954), .B(new_n5953), .C(new_n5951), .D(\a[5] ), .Y(new_n5955));
  AOI31xp33_ASAP7_75t_L     g05699(.A1(new_n5954), .A2(new_n5953), .A3(new_n5951), .B(\a[5] ), .Y(new_n5956));
  NOR2xp33_ASAP7_75t_L      g05700(.A(new_n5956), .B(new_n5955), .Y(new_n5957));
  NOR2xp33_ASAP7_75t_L      g05701(.A(new_n5652), .B(new_n5699), .Y(new_n5958));
  A2O1A1O1Ixp25_ASAP7_75t_L g05702(.A1(new_n5657), .A2(new_n5656), .B(new_n5958), .C(new_n5921), .D(new_n5922), .Y(new_n5959));
  OAI21xp33_ASAP7_75t_L     g05703(.A1(new_n5895), .A2(new_n5709), .B(new_n5897), .Y(new_n5960));
  NAND2xp33_ASAP7_75t_L     g05704(.A(new_n5871), .B(new_n5870), .Y(new_n5961));
  MAJIxp5_ASAP7_75t_L       g05705(.A(new_n5719), .B(new_n5961), .C(new_n5877), .Y(new_n5962));
  NAND2xp33_ASAP7_75t_L     g05706(.A(\b[26] ), .B(new_n1194), .Y(new_n5963));
  NOR2xp33_ASAP7_75t_L      g05707(.A(new_n2852), .B(new_n1198), .Y(new_n5964));
  AOI221xp5_ASAP7_75t_L     g05708(.A1(new_n1103), .A2(\b[27] ), .B1(new_n1110), .B2(new_n2858), .C(new_n5964), .Y(new_n5965));
  AND3x1_ASAP7_75t_L        g05709(.A(new_n5965), .B(new_n5963), .C(\a[17] ), .Y(new_n5966));
  O2A1O1Ixp33_ASAP7_75t_L   g05710(.A1(new_n2477), .A2(new_n1195), .B(new_n5965), .C(\a[17] ), .Y(new_n5967));
  NOR2xp33_ASAP7_75t_L      g05711(.A(new_n5967), .B(new_n5966), .Y(new_n5968));
  INVx1_ASAP7_75t_L         g05712(.A(new_n5968), .Y(new_n5969));
  NAND3xp33_ASAP7_75t_L     g05713(.A(new_n5734), .B(new_n5801), .C(new_n5802), .Y(new_n5970));
  A2O1A1Ixp33_ASAP7_75t_L   g05714(.A1(new_n5803), .A2(new_n5795), .B(new_n5728), .C(new_n5970), .Y(new_n5971));
  NOR2xp33_ASAP7_75t_L      g05715(.A(new_n695), .B(new_n3492), .Y(new_n5972));
  INVx1_ASAP7_75t_L         g05716(.A(new_n5972), .Y(new_n5973));
  NAND2xp33_ASAP7_75t_L     g05717(.A(\b[12] ), .B(new_n3260), .Y(new_n5974));
  AOI22xp33_ASAP7_75t_L     g05718(.A1(new_n3256), .A2(\b[13] ), .B1(new_n3254), .B2(new_n800), .Y(new_n5975));
  NAND4xp25_ASAP7_75t_L     g05719(.A(new_n5975), .B(\a[32] ), .C(new_n5973), .D(new_n5974), .Y(new_n5976));
  AOI31xp33_ASAP7_75t_L     g05720(.A1(new_n5975), .A2(new_n5974), .A3(new_n5973), .B(\a[32] ), .Y(new_n5977));
  INVx1_ASAP7_75t_L         g05721(.A(new_n5977), .Y(new_n5978));
  AND2x2_ASAP7_75t_L        g05722(.A(new_n5976), .B(new_n5978), .Y(new_n5979));
  A2O1A1O1Ixp25_ASAP7_75t_L g05723(.A1(new_n5547), .A2(new_n5505), .B(new_n5735), .C(new_n5786), .D(new_n5799), .Y(new_n5980));
  INVx1_ASAP7_75t_L         g05724(.A(new_n5745), .Y(new_n5981));
  NOR3xp33_ASAP7_75t_L      g05725(.A(new_n5770), .B(new_n5981), .C(new_n5740), .Y(new_n5982));
  NOR2xp33_ASAP7_75t_L      g05726(.A(new_n278), .B(new_n5521), .Y(new_n5983));
  NOR2xp33_ASAP7_75t_L      g05727(.A(new_n299), .B(new_n5241), .Y(new_n5984));
  OAI32xp33_ASAP7_75t_L     g05728(.A1(new_n325), .A2(new_n327), .A3(new_n5252), .B1(new_n323), .B2(new_n5253), .Y(new_n5985));
  NOR4xp25_ASAP7_75t_L      g05729(.A(new_n5985), .B(new_n5244), .C(new_n5983), .D(new_n5984), .Y(new_n5986));
  INVx1_ASAP7_75t_L         g05730(.A(new_n5986), .Y(new_n5987));
  OAI31xp33_ASAP7_75t_L     g05731(.A1(new_n5985), .A2(new_n5984), .A3(new_n5983), .B(new_n5244), .Y(new_n5988));
  NAND2xp33_ASAP7_75t_L     g05732(.A(\a[44] ), .B(new_n5745), .Y(new_n5989));
  NAND2xp33_ASAP7_75t_L     g05733(.A(new_n5743), .B(new_n5742), .Y(new_n5990));
  XNOR2x2_ASAP7_75t_L       g05734(.A(\a[43] ), .B(\a[42] ), .Y(new_n5991));
  NOR2xp33_ASAP7_75t_L      g05735(.A(new_n5991), .B(new_n5990), .Y(new_n5992));
  NAND2xp33_ASAP7_75t_L     g05736(.A(\b[0] ), .B(new_n5992), .Y(new_n5993));
  INVx1_ASAP7_75t_L         g05737(.A(\a[43] ), .Y(new_n5994));
  NAND2xp33_ASAP7_75t_L     g05738(.A(\a[44] ), .B(new_n5994), .Y(new_n5995));
  INVx1_ASAP7_75t_L         g05739(.A(\a[44] ), .Y(new_n5996));
  NAND2xp33_ASAP7_75t_L     g05740(.A(\a[43] ), .B(new_n5996), .Y(new_n5997));
  AND2x2_ASAP7_75t_L        g05741(.A(new_n5995), .B(new_n5997), .Y(new_n5998));
  NOR2xp33_ASAP7_75t_L      g05742(.A(new_n5744), .B(new_n5998), .Y(new_n5999));
  NAND2xp33_ASAP7_75t_L     g05743(.A(new_n271), .B(new_n5999), .Y(new_n6000));
  NAND2xp33_ASAP7_75t_L     g05744(.A(new_n5997), .B(new_n5995), .Y(new_n6001));
  NOR2xp33_ASAP7_75t_L      g05745(.A(new_n6001), .B(new_n5744), .Y(new_n6002));
  NAND2xp33_ASAP7_75t_L     g05746(.A(\b[1] ), .B(new_n6002), .Y(new_n6003));
  NAND3xp33_ASAP7_75t_L     g05747(.A(new_n6000), .B(new_n6003), .C(new_n5993), .Y(new_n6004));
  XOR2x2_ASAP7_75t_L        g05748(.A(new_n5989), .B(new_n6004), .Y(new_n6005));
  NAND3xp33_ASAP7_75t_L     g05749(.A(new_n6005), .B(new_n5988), .C(new_n5987), .Y(new_n6006));
  INVx1_ASAP7_75t_L         g05750(.A(new_n5988), .Y(new_n6007));
  XNOR2x2_ASAP7_75t_L       g05751(.A(new_n5989), .B(new_n6004), .Y(new_n6008));
  OAI21xp33_ASAP7_75t_L     g05752(.A1(new_n5986), .A2(new_n6007), .B(new_n6008), .Y(new_n6009));
  OAI211xp5_ASAP7_75t_L     g05753(.A1(new_n5982), .A2(new_n5762), .B(new_n6006), .C(new_n6009), .Y(new_n6010));
  INVx1_ASAP7_75t_L         g05754(.A(new_n5982), .Y(new_n6011));
  NOR3xp33_ASAP7_75t_L      g05755(.A(new_n6008), .B(new_n6007), .C(new_n5986), .Y(new_n6012));
  AOI21xp33_ASAP7_75t_L     g05756(.A1(new_n5988), .A2(new_n5987), .B(new_n6005), .Y(new_n6013));
  OAI211xp5_ASAP7_75t_L     g05757(.A1(new_n6012), .A2(new_n6013), .B(new_n5753), .C(new_n6011), .Y(new_n6014));
  NAND2xp33_ASAP7_75t_L     g05758(.A(\b[5] ), .B(new_n4780), .Y(new_n6015));
  NAND2xp33_ASAP7_75t_L     g05759(.A(\b[6] ), .B(new_n4548), .Y(new_n6016));
  AOI32xp33_ASAP7_75t_L     g05760(.A1(new_n424), .A2(new_n426), .A3(new_n4542), .B1(new_n4544), .B2(\b[7] ), .Y(new_n6017));
  NAND4xp25_ASAP7_75t_L     g05761(.A(new_n6017), .B(\a[38] ), .C(new_n6015), .D(new_n6016), .Y(new_n6018));
  INVx1_ASAP7_75t_L         g05762(.A(new_n6018), .Y(new_n6019));
  AOI31xp33_ASAP7_75t_L     g05763(.A1(new_n6017), .A2(new_n6016), .A3(new_n6015), .B(\a[38] ), .Y(new_n6020));
  NOR2xp33_ASAP7_75t_L      g05764(.A(new_n6020), .B(new_n6019), .Y(new_n6021));
  NAND3xp33_ASAP7_75t_L     g05765(.A(new_n6021), .B(new_n6014), .C(new_n6010), .Y(new_n6022));
  AO21x2_ASAP7_75t_L        g05766(.A1(new_n6010), .A2(new_n6014), .B(new_n6021), .Y(new_n6023));
  NAND2xp33_ASAP7_75t_L     g05767(.A(new_n6022), .B(new_n6023), .Y(new_n6024));
  AOI211xp5_ASAP7_75t_L     g05768(.A1(new_n5760), .A2(new_n5758), .B(new_n5762), .C(new_n5763), .Y(new_n6025));
  INVx1_ASAP7_75t_L         g05769(.A(new_n6025), .Y(new_n6026));
  A2O1A1Ixp33_ASAP7_75t_L   g05770(.A1(new_n5766), .A2(new_n5761), .B(new_n5777), .C(new_n6026), .Y(new_n6027));
  NOR2xp33_ASAP7_75t_L      g05771(.A(new_n6027), .B(new_n6024), .Y(new_n6028));
  AOI21xp33_ASAP7_75t_L     g05772(.A1(new_n5775), .A2(new_n5767), .B(new_n6025), .Y(new_n6029));
  AOI21xp33_ASAP7_75t_L     g05773(.A1(new_n6023), .A2(new_n6022), .B(new_n6029), .Y(new_n6030));
  NOR2xp33_ASAP7_75t_L      g05774(.A(new_n503), .B(new_n4986), .Y(new_n6031));
  INVx1_ASAP7_75t_L         g05775(.A(new_n6031), .Y(new_n6032));
  NAND2xp33_ASAP7_75t_L     g05776(.A(\b[9] ), .B(new_n3874), .Y(new_n6033));
  AOI22xp33_ASAP7_75t_L     g05777(.A1(new_n3884), .A2(\b[10] ), .B1(new_n3881), .B2(new_n852), .Y(new_n6034));
  AND4x1_ASAP7_75t_L        g05778(.A(new_n6034), .B(new_n6033), .C(new_n6032), .D(\a[35] ), .Y(new_n6035));
  AOI31xp33_ASAP7_75t_L     g05779(.A1(new_n6034), .A2(new_n6033), .A3(new_n6032), .B(\a[35] ), .Y(new_n6036));
  NOR2xp33_ASAP7_75t_L      g05780(.A(new_n6036), .B(new_n6035), .Y(new_n6037));
  OAI21xp33_ASAP7_75t_L     g05781(.A1(new_n6030), .A2(new_n6028), .B(new_n6037), .Y(new_n6038));
  NAND3xp33_ASAP7_75t_L     g05782(.A(new_n6029), .B(new_n6023), .C(new_n6022), .Y(new_n6039));
  A2O1A1Ixp33_ASAP7_75t_L   g05783(.A1(new_n5767), .A2(new_n5775), .B(new_n6025), .C(new_n6024), .Y(new_n6040));
  OAI211xp5_ASAP7_75t_L     g05784(.A1(new_n6035), .A2(new_n6036), .B(new_n6040), .C(new_n6039), .Y(new_n6041));
  NAND3xp33_ASAP7_75t_L     g05785(.A(new_n5980), .B(new_n6041), .C(new_n6038), .Y(new_n6042));
  AOI21xp33_ASAP7_75t_L     g05786(.A1(new_n6041), .A2(new_n6038), .B(new_n5980), .Y(new_n6043));
  INVx1_ASAP7_75t_L         g05787(.A(new_n6043), .Y(new_n6044));
  NAND3xp33_ASAP7_75t_L     g05788(.A(new_n5979), .B(new_n6044), .C(new_n6042), .Y(new_n6045));
  NAND2xp33_ASAP7_75t_L     g05789(.A(new_n5976), .B(new_n5978), .Y(new_n6046));
  INVx1_ASAP7_75t_L         g05790(.A(new_n6042), .Y(new_n6047));
  OAI21xp33_ASAP7_75t_L     g05791(.A1(new_n6043), .A2(new_n6047), .B(new_n6046), .Y(new_n6048));
  NAND3xp33_ASAP7_75t_L     g05792(.A(new_n5971), .B(new_n6045), .C(new_n6048), .Y(new_n6049));
  A2O1A1Ixp33_ASAP7_75t_L   g05793(.A1(new_n5027), .A2(new_n5028), .B(new_n5304), .C(new_n5291), .Y(new_n6050));
  A2O1A1Ixp33_ASAP7_75t_L   g05794(.A1(new_n6050), .A2(new_n5295), .B(new_n5562), .C(new_n5559), .Y(new_n6051));
  NOR2xp33_ASAP7_75t_L      g05795(.A(new_n5794), .B(new_n5793), .Y(new_n6052));
  MAJIxp5_ASAP7_75t_L       g05796(.A(new_n6051), .B(new_n5734), .C(new_n6052), .Y(new_n6053));
  NOR3xp33_ASAP7_75t_L      g05797(.A(new_n6047), .B(new_n6043), .C(new_n6046), .Y(new_n6054));
  AOI21xp33_ASAP7_75t_L     g05798(.A1(new_n6044), .A2(new_n6042), .B(new_n5979), .Y(new_n6055));
  OAI21xp33_ASAP7_75t_L     g05799(.A1(new_n6055), .A2(new_n6054), .B(new_n6053), .Y(new_n6056));
  NOR2xp33_ASAP7_75t_L      g05800(.A(new_n871), .B(new_n2932), .Y(new_n6057));
  INVx1_ASAP7_75t_L         g05801(.A(new_n6057), .Y(new_n6058));
  AOI22xp33_ASAP7_75t_L     g05802(.A1(new_n2702), .A2(\b[16] ), .B1(new_n2700), .B2(new_n1058), .Y(new_n6059));
  OAI211xp5_ASAP7_75t_L     g05803(.A1(new_n952), .A2(new_n2694), .B(new_n6059), .C(new_n6058), .Y(new_n6060));
  XNOR2x2_ASAP7_75t_L       g05804(.A(\a[29] ), .B(new_n6060), .Y(new_n6061));
  NAND3xp33_ASAP7_75t_L     g05805(.A(new_n6061), .B(new_n6056), .C(new_n6049), .Y(new_n6062));
  NOR3xp33_ASAP7_75t_L      g05806(.A(new_n6053), .B(new_n6054), .C(new_n6055), .Y(new_n6063));
  AOI21xp33_ASAP7_75t_L     g05807(.A1(new_n6045), .A2(new_n6048), .B(new_n5971), .Y(new_n6064));
  XNOR2x2_ASAP7_75t_L       g05808(.A(new_n2697), .B(new_n6060), .Y(new_n6065));
  OAI21xp33_ASAP7_75t_L     g05809(.A1(new_n6064), .A2(new_n6063), .B(new_n6065), .Y(new_n6066));
  NOR2xp33_ASAP7_75t_L      g05810(.A(new_n5808), .B(new_n5809), .Y(new_n6067));
  MAJIxp5_ASAP7_75t_L       g05811(.A(new_n5720), .B(new_n5807), .C(new_n6067), .Y(new_n6068));
  NAND3xp33_ASAP7_75t_L     g05812(.A(new_n6068), .B(new_n6066), .C(new_n6062), .Y(new_n6069));
  NOR3xp33_ASAP7_75t_L      g05813(.A(new_n6065), .B(new_n6063), .C(new_n6064), .Y(new_n6070));
  AOI21xp33_ASAP7_75t_L     g05814(.A1(new_n6056), .A2(new_n6049), .B(new_n6061), .Y(new_n6071));
  NAND2xp33_ASAP7_75t_L     g05815(.A(new_n5805), .B(new_n5804), .Y(new_n6072));
  MAJIxp5_ASAP7_75t_L       g05816(.A(new_n5812), .B(new_n5727), .C(new_n6072), .Y(new_n6073));
  OAI21xp33_ASAP7_75t_L     g05817(.A1(new_n6070), .A2(new_n6071), .B(new_n6073), .Y(new_n6074));
  NOR2xp33_ASAP7_75t_L      g05818(.A(new_n1244), .B(new_n2387), .Y(new_n6075));
  INVx1_ASAP7_75t_L         g05819(.A(new_n6075), .Y(new_n6076));
  AOI32xp33_ASAP7_75t_L     g05820(.A1(new_n2792), .A2(new_n1496), .A3(new_n2226), .B1(\b[19] ), .B2(new_n2228), .Y(new_n6077));
  OAI311xp33_ASAP7_75t_L    g05821(.A1(new_n1356), .A2(new_n2218), .A3(new_n2231), .B1(new_n6076), .C1(new_n6077), .Y(new_n6078));
  XNOR2x2_ASAP7_75t_L       g05822(.A(\a[26] ), .B(new_n6078), .Y(new_n6079));
  NAND3xp33_ASAP7_75t_L     g05823(.A(new_n6069), .B(new_n6079), .C(new_n6074), .Y(new_n6080));
  NAND2xp33_ASAP7_75t_L     g05824(.A(new_n5807), .B(new_n6067), .Y(new_n6081));
  OAI21xp33_ASAP7_75t_L     g05825(.A1(new_n5813), .A2(new_n5814), .B(new_n5720), .Y(new_n6082));
  AND4x1_ASAP7_75t_L        g05826(.A(new_n6082), .B(new_n6081), .C(new_n6066), .D(new_n6062), .Y(new_n6083));
  AOI21xp33_ASAP7_75t_L     g05827(.A1(new_n6066), .A2(new_n6062), .B(new_n6068), .Y(new_n6084));
  XNOR2x2_ASAP7_75t_L       g05828(.A(new_n2223), .B(new_n6078), .Y(new_n6085));
  OAI21xp33_ASAP7_75t_L     g05829(.A1(new_n6084), .A2(new_n6083), .B(new_n6085), .Y(new_n6086));
  NAND2xp33_ASAP7_75t_L     g05830(.A(new_n6080), .B(new_n6086), .Y(new_n6087));
  OAI21xp33_ASAP7_75t_L     g05831(.A1(new_n5827), .A2(new_n5831), .B(new_n5832), .Y(new_n6088));
  NOR2xp33_ASAP7_75t_L      g05832(.A(new_n6088), .B(new_n6087), .Y(new_n6089));
  A2O1A1O1Ixp25_ASAP7_75t_L g05833(.A1(new_n5590), .A2(new_n5587), .B(new_n5589), .C(new_n5833), .D(new_n5823), .Y(new_n6090));
  AOI21xp33_ASAP7_75t_L     g05834(.A1(new_n6086), .A2(new_n6080), .B(new_n6090), .Y(new_n6091));
  NAND2xp33_ASAP7_75t_L     g05835(.A(\b[20] ), .B(new_n1910), .Y(new_n6092));
  NAND2xp33_ASAP7_75t_L     g05836(.A(\b[21] ), .B(new_n1770), .Y(new_n6093));
  AOI32xp33_ASAP7_75t_L     g05837(.A1(new_n1862), .A2(new_n1860), .A3(new_n1764), .B1(new_n1766), .B2(\b[22] ), .Y(new_n6094));
  NAND4xp25_ASAP7_75t_L     g05838(.A(new_n6094), .B(\a[23] ), .C(new_n6092), .D(new_n6093), .Y(new_n6095));
  NAND2xp33_ASAP7_75t_L     g05839(.A(new_n6093), .B(new_n6094), .Y(new_n6096));
  A2O1A1Ixp33_ASAP7_75t_L   g05840(.A1(\b[20] ), .A2(new_n1910), .B(new_n6096), .C(new_n1761), .Y(new_n6097));
  NAND2xp33_ASAP7_75t_L     g05841(.A(new_n6095), .B(new_n6097), .Y(new_n6098));
  NOR3xp33_ASAP7_75t_L      g05842(.A(new_n6089), .B(new_n6091), .C(new_n6098), .Y(new_n6099));
  NAND3xp33_ASAP7_75t_L     g05843(.A(new_n6090), .B(new_n6086), .C(new_n6080), .Y(new_n6100));
  NOR3xp33_ASAP7_75t_L      g05844(.A(new_n6083), .B(new_n6085), .C(new_n6084), .Y(new_n6101));
  AOI21xp33_ASAP7_75t_L     g05845(.A1(new_n6069), .A2(new_n6074), .B(new_n6079), .Y(new_n6102));
  OAI21xp33_ASAP7_75t_L     g05846(.A1(new_n6101), .A2(new_n6102), .B(new_n6088), .Y(new_n6103));
  AND2x2_ASAP7_75t_L        g05847(.A(new_n6095), .B(new_n6097), .Y(new_n6104));
  AOI21xp33_ASAP7_75t_L     g05848(.A1(new_n6100), .A2(new_n6103), .B(new_n6104), .Y(new_n6105));
  NOR2xp33_ASAP7_75t_L      g05849(.A(new_n6105), .B(new_n6099), .Y(new_n6106));
  NAND2xp33_ASAP7_75t_L     g05850(.A(new_n5835), .B(new_n5829), .Y(new_n6107));
  NOR2xp33_ASAP7_75t_L      g05851(.A(new_n5842), .B(new_n6107), .Y(new_n6108));
  INVx1_ASAP7_75t_L         g05852(.A(new_n6108), .Y(new_n6109));
  NAND3xp33_ASAP7_75t_L     g05853(.A(new_n5856), .B(new_n6106), .C(new_n6109), .Y(new_n6110));
  NAND3xp33_ASAP7_75t_L     g05854(.A(new_n6104), .B(new_n6100), .C(new_n6103), .Y(new_n6111));
  OAI21xp33_ASAP7_75t_L     g05855(.A1(new_n6091), .A2(new_n6089), .B(new_n6098), .Y(new_n6112));
  NAND2xp33_ASAP7_75t_L     g05856(.A(new_n6111), .B(new_n6112), .Y(new_n6113));
  MAJIxp5_ASAP7_75t_L       g05857(.A(new_n5850), .B(new_n6107), .C(new_n5842), .Y(new_n6114));
  NAND2xp33_ASAP7_75t_L     g05858(.A(new_n6113), .B(new_n6114), .Y(new_n6115));
  NOR2xp33_ASAP7_75t_L      g05859(.A(new_n1995), .B(new_n1549), .Y(new_n6116));
  NAND2xp33_ASAP7_75t_L     g05860(.A(\b[24] ), .B(new_n1410), .Y(new_n6117));
  OAI221xp5_ASAP7_75t_L     g05861(.A1(new_n1412), .A2(new_n2180), .B1(new_n1411), .B2(new_n2187), .C(new_n6117), .Y(new_n6118));
  OR3x1_ASAP7_75t_L         g05862(.A(new_n6118), .B(new_n1401), .C(new_n6116), .Y(new_n6119));
  A2O1A1Ixp33_ASAP7_75t_L   g05863(.A1(\b[23] ), .A2(new_n1548), .B(new_n6118), .C(new_n1401), .Y(new_n6120));
  AND2x2_ASAP7_75t_L        g05864(.A(new_n6120), .B(new_n6119), .Y(new_n6121));
  NAND3xp33_ASAP7_75t_L     g05865(.A(new_n6110), .B(new_n6115), .C(new_n6121), .Y(new_n6122));
  NOR2xp33_ASAP7_75t_L      g05866(.A(new_n6113), .B(new_n6114), .Y(new_n6123));
  O2A1O1Ixp33_ASAP7_75t_L   g05867(.A1(new_n5850), .A2(new_n5848), .B(new_n6109), .C(new_n6106), .Y(new_n6124));
  NAND2xp33_ASAP7_75t_L     g05868(.A(new_n6120), .B(new_n6119), .Y(new_n6125));
  OAI21xp33_ASAP7_75t_L     g05869(.A1(new_n6123), .A2(new_n6124), .B(new_n6125), .Y(new_n6126));
  A2O1A1O1Ixp25_ASAP7_75t_L g05870(.A1(new_n5612), .A2(new_n5484), .B(new_n5880), .C(new_n5881), .D(new_n5868), .Y(new_n6127));
  AOI21xp33_ASAP7_75t_L     g05871(.A1(new_n6126), .A2(new_n6122), .B(new_n6127), .Y(new_n6128));
  NAND2xp33_ASAP7_75t_L     g05872(.A(new_n6122), .B(new_n6126), .Y(new_n6129));
  A2O1A1Ixp33_ASAP7_75t_L   g05873(.A1(new_n5869), .A2(new_n5615), .B(new_n5864), .C(new_n5882), .Y(new_n6130));
  NOR2xp33_ASAP7_75t_L      g05874(.A(new_n6130), .B(new_n6129), .Y(new_n6131));
  OAI21xp33_ASAP7_75t_L     g05875(.A1(new_n6128), .A2(new_n6131), .B(new_n5969), .Y(new_n6132));
  NAND2xp33_ASAP7_75t_L     g05876(.A(new_n6130), .B(new_n6129), .Y(new_n6133));
  NAND3xp33_ASAP7_75t_L     g05877(.A(new_n6127), .B(new_n6126), .C(new_n6122), .Y(new_n6134));
  NAND3xp33_ASAP7_75t_L     g05878(.A(new_n6134), .B(new_n6133), .C(new_n5968), .Y(new_n6135));
  NAND3xp33_ASAP7_75t_L     g05879(.A(new_n5962), .B(new_n6132), .C(new_n6135), .Y(new_n6136));
  NOR2xp33_ASAP7_75t_L      g05880(.A(new_n5879), .B(new_n5883), .Y(new_n6137));
  MAJIxp5_ASAP7_75t_L       g05881(.A(new_n5888), .B(new_n6137), .C(new_n5884), .Y(new_n6138));
  NAND2xp33_ASAP7_75t_L     g05882(.A(new_n6135), .B(new_n6132), .Y(new_n6139));
  NAND2xp33_ASAP7_75t_L     g05883(.A(new_n6138), .B(new_n6139), .Y(new_n6140));
  NOR2xp33_ASAP7_75t_L      g05884(.A(new_n2871), .B(new_n909), .Y(new_n6141));
  INVx1_ASAP7_75t_L         g05885(.A(new_n6141), .Y(new_n6142));
  NAND2xp33_ASAP7_75t_L     g05886(.A(\b[30] ), .B(new_n817), .Y(new_n6143));
  AOI22xp33_ASAP7_75t_L     g05887(.A1(new_n826), .A2(\b[31] ), .B1(new_n823), .B2(new_n3426), .Y(new_n6144));
  AND4x1_ASAP7_75t_L        g05888(.A(new_n6144), .B(new_n6143), .C(new_n6142), .D(\a[14] ), .Y(new_n6145));
  AOI31xp33_ASAP7_75t_L     g05889(.A1(new_n6144), .A2(new_n6143), .A3(new_n6142), .B(\a[14] ), .Y(new_n6146));
  NOR2xp33_ASAP7_75t_L      g05890(.A(new_n6146), .B(new_n6145), .Y(new_n6147));
  NAND3xp33_ASAP7_75t_L     g05891(.A(new_n6140), .B(new_n6136), .C(new_n6147), .Y(new_n6148));
  O2A1O1Ixp33_ASAP7_75t_L   g05892(.A1(new_n5961), .A2(new_n5877), .B(new_n5893), .C(new_n6139), .Y(new_n6149));
  AOI21xp33_ASAP7_75t_L     g05893(.A1(new_n6135), .A2(new_n6132), .B(new_n5962), .Y(new_n6150));
  INVx1_ASAP7_75t_L         g05894(.A(new_n6147), .Y(new_n6151));
  OAI21xp33_ASAP7_75t_L     g05895(.A1(new_n6150), .A2(new_n6149), .B(new_n6151), .Y(new_n6152));
  NAND3xp33_ASAP7_75t_L     g05896(.A(new_n5960), .B(new_n6148), .C(new_n6152), .Y(new_n6153));
  A2O1A1O1Ixp25_ASAP7_75t_L g05897(.A1(new_n5630), .A2(new_n5468), .B(new_n5639), .C(new_n5898), .D(new_n5891), .Y(new_n6154));
  NOR3xp33_ASAP7_75t_L      g05898(.A(new_n6149), .B(new_n6151), .C(new_n6150), .Y(new_n6155));
  AOI21xp33_ASAP7_75t_L     g05899(.A1(new_n6140), .A2(new_n6136), .B(new_n6147), .Y(new_n6156));
  OAI21xp33_ASAP7_75t_L     g05900(.A1(new_n6155), .A2(new_n6156), .B(new_n6154), .Y(new_n6157));
  NAND2xp33_ASAP7_75t_L     g05901(.A(\b[32] ), .B(new_n674), .Y(new_n6158));
  NAND2xp33_ASAP7_75t_L     g05902(.A(\b[33] ), .B(new_n590), .Y(new_n6159));
  AOI22xp33_ASAP7_75t_L     g05903(.A1(new_n600), .A2(\b[34] ), .B1(new_n597), .B2(new_n3833), .Y(new_n6160));
  AND4x1_ASAP7_75t_L        g05904(.A(new_n6160), .B(new_n6159), .C(new_n6158), .D(\a[11] ), .Y(new_n6161));
  AOI31xp33_ASAP7_75t_L     g05905(.A1(new_n6160), .A2(new_n6159), .A3(new_n6158), .B(\a[11] ), .Y(new_n6162));
  NOR2xp33_ASAP7_75t_L      g05906(.A(new_n6162), .B(new_n6161), .Y(new_n6163));
  AND3x1_ASAP7_75t_L        g05907(.A(new_n6157), .B(new_n6153), .C(new_n6163), .Y(new_n6164));
  AOI21xp33_ASAP7_75t_L     g05908(.A1(new_n6157), .A2(new_n6153), .B(new_n6163), .Y(new_n6165));
  MAJIxp5_ASAP7_75t_L       g05909(.A(new_n5708), .B(new_n5918), .C(new_n5912), .Y(new_n6166));
  NOR3xp33_ASAP7_75t_L      g05910(.A(new_n6166), .B(new_n6165), .C(new_n6164), .Y(new_n6167));
  OA21x2_ASAP7_75t_L        g05911(.A1(new_n6164), .A2(new_n6165), .B(new_n6166), .Y(new_n6168));
  NAND2xp33_ASAP7_75t_L     g05912(.A(\b[35] ), .B(new_n480), .Y(new_n6169));
  NAND2xp33_ASAP7_75t_L     g05913(.A(\b[36] ), .B(new_n441), .Y(new_n6170));
  NOR2xp33_ASAP7_75t_L      g05914(.A(new_n4701), .B(new_n667), .Y(new_n6171));
  AOI21xp33_ASAP7_75t_L     g05915(.A1(new_n4709), .A2(new_n448), .B(new_n6171), .Y(new_n6172));
  NAND3xp33_ASAP7_75t_L     g05916(.A(new_n6172), .B(new_n6170), .C(new_n6169), .Y(new_n6173));
  XNOR2x2_ASAP7_75t_L       g05917(.A(\a[8] ), .B(new_n6173), .Y(new_n6174));
  OAI21xp33_ASAP7_75t_L     g05918(.A1(new_n6167), .A2(new_n6168), .B(new_n6174), .Y(new_n6175));
  OR3x1_ASAP7_75t_L         g05919(.A(new_n6168), .B(new_n6174), .C(new_n6167), .Y(new_n6176));
  NAND3xp33_ASAP7_75t_L     g05920(.A(new_n5959), .B(new_n6175), .C(new_n6176), .Y(new_n6177));
  NAND2xp33_ASAP7_75t_L     g05921(.A(new_n6175), .B(new_n6176), .Y(new_n6178));
  A2O1A1Ixp33_ASAP7_75t_L   g05922(.A1(new_n5921), .A2(new_n5700), .B(new_n5922), .C(new_n6178), .Y(new_n6179));
  NAND3xp33_ASAP7_75t_L     g05923(.A(new_n6179), .B(new_n6177), .C(new_n5957), .Y(new_n6180));
  NOR3xp33_ASAP7_75t_L      g05924(.A(new_n6178), .B(new_n5924), .C(new_n5922), .Y(new_n6181));
  AOI21xp33_ASAP7_75t_L     g05925(.A1(new_n6176), .A2(new_n6175), .B(new_n5959), .Y(new_n6182));
  OAI22xp33_ASAP7_75t_L     g05926(.A1(new_n6181), .A2(new_n6182), .B1(new_n5955), .B2(new_n5956), .Y(new_n6183));
  NAND3xp33_ASAP7_75t_L     g05927(.A(new_n5949), .B(new_n6180), .C(new_n6183), .Y(new_n6184));
  A2O1A1O1Ixp25_ASAP7_75t_L g05928(.A1(new_n5445), .A2(new_n5661), .B(new_n5659), .C(new_n5936), .D(new_n5947), .Y(new_n6185));
  INVx1_ASAP7_75t_L         g05929(.A(new_n6180), .Y(new_n6186));
  AOI21xp33_ASAP7_75t_L     g05930(.A1(new_n6179), .A2(new_n6177), .B(new_n5957), .Y(new_n6187));
  OAI21xp33_ASAP7_75t_L     g05931(.A1(new_n6186), .A2(new_n6187), .B(new_n6185), .Y(new_n6188));
  NOR2xp33_ASAP7_75t_L      g05932(.A(new_n5666), .B(new_n277), .Y(new_n6189));
  INVx1_ASAP7_75t_L         g05933(.A(new_n6189), .Y(new_n6190));
  NOR2xp33_ASAP7_75t_L      g05934(.A(new_n5680), .B(new_n261), .Y(new_n6191));
  INVx1_ASAP7_75t_L         g05935(.A(new_n6191), .Y(new_n6192));
  INVx1_ASAP7_75t_L         g05936(.A(new_n5681), .Y(new_n6193));
  NOR2xp33_ASAP7_75t_L      g05937(.A(\b[42] ), .B(\b[43] ), .Y(new_n6194));
  INVx1_ASAP7_75t_L         g05938(.A(\b[43] ), .Y(new_n6195));
  NOR2xp33_ASAP7_75t_L      g05939(.A(new_n5680), .B(new_n6195), .Y(new_n6196));
  NOR2xp33_ASAP7_75t_L      g05940(.A(new_n6194), .B(new_n6196), .Y(new_n6197));
  INVx1_ASAP7_75t_L         g05941(.A(new_n6197), .Y(new_n6198));
  A2O1A1O1Ixp25_ASAP7_75t_L g05942(.A1(new_n5684), .A2(new_n5685), .B(new_n5679), .C(new_n6193), .D(new_n6198), .Y(new_n6199));
  A2O1A1Ixp33_ASAP7_75t_L   g05943(.A1(new_n5685), .A2(new_n5684), .B(new_n5679), .C(new_n6193), .Y(new_n6200));
  NOR2xp33_ASAP7_75t_L      g05944(.A(new_n6197), .B(new_n6200), .Y(new_n6201));
  NOR2xp33_ASAP7_75t_L      g05945(.A(new_n6199), .B(new_n6201), .Y(new_n6202));
  AOI22xp33_ASAP7_75t_L     g05946(.A1(new_n272), .A2(\b[43] ), .B1(new_n269), .B2(new_n6202), .Y(new_n6203));
  AND4x1_ASAP7_75t_L        g05947(.A(new_n6203), .B(new_n6192), .C(new_n6190), .D(\a[2] ), .Y(new_n6204));
  AOI31xp33_ASAP7_75t_L     g05948(.A1(new_n6203), .A2(new_n6192), .A3(new_n6190), .B(\a[2] ), .Y(new_n6205));
  NOR2xp33_ASAP7_75t_L      g05949(.A(new_n6205), .B(new_n6204), .Y(new_n6206));
  NAND3xp33_ASAP7_75t_L     g05950(.A(new_n6184), .B(new_n6188), .C(new_n6206), .Y(new_n6207));
  NAND2xp33_ASAP7_75t_L     g05951(.A(new_n6180), .B(new_n6183), .Y(new_n6208));
  NOR2xp33_ASAP7_75t_L      g05952(.A(new_n6185), .B(new_n6208), .Y(new_n6209));
  AOI21xp33_ASAP7_75t_L     g05953(.A1(new_n6183), .A2(new_n6180), .B(new_n5949), .Y(new_n6210));
  INVx1_ASAP7_75t_L         g05954(.A(new_n6206), .Y(new_n6211));
  OAI21xp33_ASAP7_75t_L     g05955(.A1(new_n6210), .A2(new_n6209), .B(new_n6211), .Y(new_n6212));
  NAND2xp33_ASAP7_75t_L     g05956(.A(new_n6207), .B(new_n6212), .Y(new_n6213));
  MAJIxp5_ASAP7_75t_L       g05957(.A(new_n5944), .B(new_n5691), .C(new_n5941), .Y(new_n6214));
  XOR2x2_ASAP7_75t_L        g05958(.A(new_n6213), .B(new_n6214), .Y(\f[43] ));
  NOR2xp33_ASAP7_75t_L      g05959(.A(new_n5691), .B(new_n5941), .Y(new_n6216));
  NOR3xp33_ASAP7_75t_L      g05960(.A(new_n6209), .B(new_n6210), .C(new_n6206), .Y(new_n6217));
  O2A1O1Ixp33_ASAP7_75t_L   g05961(.A1(new_n6216), .A2(new_n5943), .B(new_n6213), .C(new_n6217), .Y(new_n6218));
  NOR2xp33_ASAP7_75t_L      g05962(.A(\b[43] ), .B(\b[44] ), .Y(new_n6219));
  INVx1_ASAP7_75t_L         g05963(.A(\b[44] ), .Y(new_n6220));
  NOR2xp33_ASAP7_75t_L      g05964(.A(new_n6195), .B(new_n6220), .Y(new_n6221));
  NOR2xp33_ASAP7_75t_L      g05965(.A(new_n6219), .B(new_n6221), .Y(new_n6222));
  A2O1A1Ixp33_ASAP7_75t_L   g05966(.A1(new_n6200), .A2(new_n6197), .B(new_n6196), .C(new_n6222), .Y(new_n6223));
  INVx1_ASAP7_75t_L         g05967(.A(new_n5187), .Y(new_n6224));
  A2O1A1Ixp33_ASAP7_75t_L   g05968(.A1(new_n5189), .A2(new_n6224), .B(new_n5665), .C(new_n5684), .Y(new_n6225));
  A2O1A1O1Ixp25_ASAP7_75t_L g05969(.A1(new_n5682), .A2(new_n6225), .B(new_n5681), .C(new_n6197), .D(new_n6196), .Y(new_n6226));
  INVx1_ASAP7_75t_L         g05970(.A(new_n6222), .Y(new_n6227));
  NAND2xp33_ASAP7_75t_L     g05971(.A(new_n6227), .B(new_n6226), .Y(new_n6228));
  NAND2xp33_ASAP7_75t_L     g05972(.A(new_n6228), .B(new_n6223), .Y(new_n6229));
  NAND2xp33_ASAP7_75t_L     g05973(.A(\b[44] ), .B(new_n272), .Y(new_n6230));
  OAI221xp5_ASAP7_75t_L     g05974(.A1(new_n6195), .A2(new_n261), .B1(new_n292), .B2(new_n6229), .C(new_n6230), .Y(new_n6231));
  AOI21xp33_ASAP7_75t_L     g05975(.A1(new_n291), .A2(\b[42] ), .B(new_n6231), .Y(new_n6232));
  NAND2xp33_ASAP7_75t_L     g05976(.A(\a[2] ), .B(new_n6232), .Y(new_n6233));
  A2O1A1Ixp33_ASAP7_75t_L   g05977(.A1(\b[42] ), .A2(new_n291), .B(new_n6231), .C(new_n265), .Y(new_n6234));
  AND2x2_ASAP7_75t_L        g05978(.A(new_n6234), .B(new_n6233), .Y(new_n6235));
  NAND2xp33_ASAP7_75t_L     g05979(.A(\b[40] ), .B(new_n334), .Y(new_n6236));
  AOI22xp33_ASAP7_75t_L     g05980(.A1(new_n345), .A2(\b[41] ), .B1(new_n342), .B2(new_n5669), .Y(new_n6237));
  NAND2xp33_ASAP7_75t_L     g05981(.A(new_n6236), .B(new_n6237), .Y(new_n6238));
  AOI21xp33_ASAP7_75t_L     g05982(.A1(new_n366), .A2(\b[39] ), .B(new_n6238), .Y(new_n6239));
  NAND2xp33_ASAP7_75t_L     g05983(.A(\a[5] ), .B(new_n6239), .Y(new_n6240));
  A2O1A1Ixp33_ASAP7_75t_L   g05984(.A1(\b[39] ), .A2(new_n366), .B(new_n6238), .C(new_n339), .Y(new_n6241));
  NAND2xp33_ASAP7_75t_L     g05985(.A(new_n6241), .B(new_n6240), .Y(new_n6242));
  INVx1_ASAP7_75t_L         g05986(.A(new_n6242), .Y(new_n6243));
  OAI21xp33_ASAP7_75t_L     g05987(.A1(new_n6164), .A2(new_n6165), .B(new_n6166), .Y(new_n6244));
  OAI21xp33_ASAP7_75t_L     g05988(.A1(new_n6155), .A2(new_n6154), .B(new_n6152), .Y(new_n6245));
  NAND2xp33_ASAP7_75t_L     g05989(.A(\b[30] ), .B(new_n908), .Y(new_n6246));
  NAND2xp33_ASAP7_75t_L     g05990(.A(\b[31] ), .B(new_n817), .Y(new_n6247));
  AOI22xp33_ASAP7_75t_L     g05991(.A1(new_n826), .A2(\b[32] ), .B1(new_n823), .B2(new_n3450), .Y(new_n6248));
  NAND4xp25_ASAP7_75t_L     g05992(.A(new_n6248), .B(\a[14] ), .C(new_n6246), .D(new_n6247), .Y(new_n6249));
  NAND2xp33_ASAP7_75t_L     g05993(.A(new_n6247), .B(new_n6248), .Y(new_n6250));
  A2O1A1Ixp33_ASAP7_75t_L   g05994(.A1(\b[30] ), .A2(new_n908), .B(new_n6250), .C(new_n813), .Y(new_n6251));
  AND2x2_ASAP7_75t_L        g05995(.A(new_n6249), .B(new_n6251), .Y(new_n6252));
  AOI21xp33_ASAP7_75t_L     g05996(.A1(new_n6134), .A2(new_n6133), .B(new_n5968), .Y(new_n6253));
  NOR3xp33_ASAP7_75t_L      g05997(.A(new_n5969), .B(new_n6131), .C(new_n6128), .Y(new_n6254));
  NAND2xp33_ASAP7_75t_L     g05998(.A(new_n6133), .B(new_n6134), .Y(new_n6255));
  NOR2xp33_ASAP7_75t_L      g05999(.A(new_n5968), .B(new_n6255), .Y(new_n6256));
  O2A1O1Ixp33_ASAP7_75t_L   g06000(.A1(new_n6253), .A2(new_n6254), .B(new_n5962), .C(new_n6256), .Y(new_n6257));
  NAND2xp33_ASAP7_75t_L     g06001(.A(\b[27] ), .B(new_n1194), .Y(new_n6258));
  NAND2xp33_ASAP7_75t_L     g06002(.A(\b[28] ), .B(new_n1103), .Y(new_n6259));
  AOI22xp33_ASAP7_75t_L     g06003(.A1(new_n1113), .A2(\b[29] ), .B1(new_n1110), .B2(new_n5472), .Y(new_n6260));
  NAND4xp25_ASAP7_75t_L     g06004(.A(new_n6260), .B(\a[17] ), .C(new_n6258), .D(new_n6259), .Y(new_n6261));
  NAND2xp33_ASAP7_75t_L     g06005(.A(new_n6259), .B(new_n6260), .Y(new_n6262));
  A2O1A1Ixp33_ASAP7_75t_L   g06006(.A1(\b[27] ), .A2(new_n1194), .B(new_n6262), .C(new_n1107), .Y(new_n6263));
  AND2x2_ASAP7_75t_L        g06007(.A(new_n6261), .B(new_n6263), .Y(new_n6264));
  NOR2xp33_ASAP7_75t_L      g06008(.A(new_n6123), .B(new_n6124), .Y(new_n6265));
  MAJIxp5_ASAP7_75t_L       g06009(.A(new_n6130), .B(new_n6125), .C(new_n6265), .Y(new_n6266));
  AOI32xp33_ASAP7_75t_L     g06010(.A1(new_n2483), .A2(new_n2486), .A3(new_n1404), .B1(new_n1406), .B2(\b[26] ), .Y(new_n6267));
  OAI221xp5_ASAP7_75t_L     g06011(.A1(new_n1398), .A2(new_n2180), .B1(new_n2019), .B2(new_n1549), .C(new_n6267), .Y(new_n6268));
  XNOR2x2_ASAP7_75t_L       g06012(.A(\a[20] ), .B(new_n6268), .Y(new_n6269));
  INVx1_ASAP7_75t_L         g06013(.A(new_n6269), .Y(new_n6270));
  NOR3xp33_ASAP7_75t_L      g06014(.A(new_n6104), .B(new_n6089), .C(new_n6091), .Y(new_n6271));
  INVx1_ASAP7_75t_L         g06015(.A(new_n6271), .Y(new_n6272));
  A2O1A1Ixp33_ASAP7_75t_L   g06016(.A1(new_n5856), .A2(new_n6109), .B(new_n6106), .C(new_n6272), .Y(new_n6273));
  NAND2xp33_ASAP7_75t_L     g06017(.A(new_n6056), .B(new_n6049), .Y(new_n6274));
  MAJIxp5_ASAP7_75t_L       g06018(.A(new_n6068), .B(new_n6274), .C(new_n6061), .Y(new_n6275));
  NOR2xp33_ASAP7_75t_L      g06019(.A(new_n952), .B(new_n2932), .Y(new_n6276));
  NAND2xp33_ASAP7_75t_L     g06020(.A(\b[16] ), .B(new_n2706), .Y(new_n6277));
  OAI221xp5_ASAP7_75t_L     g06021(.A1(new_n2708), .A2(new_n1244), .B1(new_n2707), .B2(new_n1251), .C(new_n6277), .Y(new_n6278));
  NOR3xp33_ASAP7_75t_L      g06022(.A(new_n6278), .B(new_n6276), .C(new_n2697), .Y(new_n6279));
  OA21x2_ASAP7_75t_L        g06023(.A1(new_n6276), .A2(new_n6278), .B(new_n2697), .Y(new_n6280));
  NOR2xp33_ASAP7_75t_L      g06024(.A(new_n6279), .B(new_n6280), .Y(new_n6281));
  AOI21xp33_ASAP7_75t_L     g06025(.A1(new_n5971), .A2(new_n6045), .B(new_n6055), .Y(new_n6282));
  NAND2xp33_ASAP7_75t_L     g06026(.A(\b[12] ), .B(new_n3491), .Y(new_n6283));
  NAND2xp33_ASAP7_75t_L     g06027(.A(\b[13] ), .B(new_n3260), .Y(new_n6284));
  AOI32xp33_ASAP7_75t_L     g06028(.A1(new_n877), .A2(new_n874), .A3(new_n3254), .B1(\b[14] ), .B2(new_n3256), .Y(new_n6285));
  AND4x1_ASAP7_75t_L        g06029(.A(new_n6285), .B(new_n6284), .C(new_n6283), .D(\a[32] ), .Y(new_n6286));
  AOI31xp33_ASAP7_75t_L     g06030(.A1(new_n6285), .A2(new_n6284), .A3(new_n6283), .B(\a[32] ), .Y(new_n6287));
  NOR2xp33_ASAP7_75t_L      g06031(.A(new_n6287), .B(new_n6286), .Y(new_n6288));
  INVx1_ASAP7_75t_L         g06032(.A(new_n6288), .Y(new_n6289));
  OAI211xp5_ASAP7_75t_L     g06033(.A1(new_n6019), .A2(new_n6020), .B(new_n6014), .C(new_n6010), .Y(new_n6290));
  INVx1_ASAP7_75t_L         g06034(.A(new_n6290), .Y(new_n6291));
  NOR2xp33_ASAP7_75t_L      g06035(.A(new_n382), .B(new_n4781), .Y(new_n6292));
  INVx1_ASAP7_75t_L         g06036(.A(new_n6292), .Y(new_n6293));
  NAND2xp33_ASAP7_75t_L     g06037(.A(\b[7] ), .B(new_n4548), .Y(new_n6294));
  AOI32xp33_ASAP7_75t_L     g06038(.A1(new_n508), .A2(new_n506), .A3(new_n4542), .B1(\b[8] ), .B2(new_n4544), .Y(new_n6295));
  NAND4xp25_ASAP7_75t_L     g06039(.A(new_n6295), .B(\a[38] ), .C(new_n6293), .D(new_n6294), .Y(new_n6296));
  AOI31xp33_ASAP7_75t_L     g06040(.A1(new_n6295), .A2(new_n6294), .A3(new_n6293), .B(\a[38] ), .Y(new_n6297));
  INVx1_ASAP7_75t_L         g06041(.A(new_n6297), .Y(new_n6298));
  A2O1A1Ixp33_ASAP7_75t_L   g06042(.A1(new_n5753), .A2(new_n6011), .B(new_n6012), .C(new_n6009), .Y(new_n6299));
  NAND2xp33_ASAP7_75t_L     g06043(.A(\b[3] ), .B(new_n5526), .Y(new_n6300));
  NAND2xp33_ASAP7_75t_L     g06044(.A(\b[4] ), .B(new_n5240), .Y(new_n6301));
  AOI22xp33_ASAP7_75t_L     g06045(.A1(new_n5249), .A2(\b[5] ), .B1(new_n5247), .B2(new_n360), .Y(new_n6302));
  NAND4xp25_ASAP7_75t_L     g06046(.A(new_n6302), .B(\a[41] ), .C(new_n6300), .D(new_n6301), .Y(new_n6303));
  OAI221xp5_ASAP7_75t_L     g06047(.A1(new_n5253), .A2(new_n353), .B1(new_n5252), .B2(new_n359), .C(new_n6301), .Y(new_n6304));
  A2O1A1Ixp33_ASAP7_75t_L   g06048(.A1(\b[3] ), .A2(new_n5526), .B(new_n6304), .C(new_n5244), .Y(new_n6305));
  AND3x1_ASAP7_75t_L        g06049(.A(new_n6000), .B(new_n6003), .C(new_n5993), .Y(new_n6306));
  INVx1_ASAP7_75t_L         g06050(.A(new_n5991), .Y(new_n6307));
  NOR3xp33_ASAP7_75t_L      g06051(.A(new_n5998), .B(new_n6307), .C(new_n5990), .Y(new_n6308));
  INVx1_ASAP7_75t_L         g06052(.A(new_n6308), .Y(new_n6309));
  NOR2xp33_ASAP7_75t_L      g06053(.A(new_n258), .B(new_n6309), .Y(new_n6310));
  NAND2xp33_ASAP7_75t_L     g06054(.A(new_n6001), .B(new_n5990), .Y(new_n6311));
  INVx1_ASAP7_75t_L         g06055(.A(new_n6002), .Y(new_n6312));
  NAND2xp33_ASAP7_75t_L     g06056(.A(\b[1] ), .B(new_n5992), .Y(new_n6313));
  OAI221xp5_ASAP7_75t_L     g06057(.A1(new_n6311), .A2(new_n283), .B1(new_n278), .B2(new_n6312), .C(new_n6313), .Y(new_n6314));
  NOR2xp33_ASAP7_75t_L      g06058(.A(new_n6310), .B(new_n6314), .Y(new_n6315));
  A2O1A1Ixp33_ASAP7_75t_L   g06059(.A1(new_n5981), .A2(new_n6306), .B(new_n5996), .C(new_n6315), .Y(new_n6316));
  O2A1O1Ixp33_ASAP7_75t_L   g06060(.A1(new_n258), .A2(new_n5744), .B(new_n6306), .C(new_n5996), .Y(new_n6317));
  A2O1A1Ixp33_ASAP7_75t_L   g06061(.A1(\b[0] ), .A2(new_n6308), .B(new_n6314), .C(new_n6317), .Y(new_n6318));
  NAND4xp25_ASAP7_75t_L     g06062(.A(new_n6318), .B(new_n6303), .C(new_n6305), .D(new_n6316), .Y(new_n6319));
  AOI211xp5_ASAP7_75t_L     g06063(.A1(\b[3] ), .A2(new_n5526), .B(new_n5244), .C(new_n6304), .Y(new_n6320));
  INVx1_ASAP7_75t_L         g06064(.A(new_n6305), .Y(new_n6321));
  NOR2xp33_ASAP7_75t_L      g06065(.A(new_n6311), .B(new_n283), .Y(new_n6322));
  AOI221xp5_ASAP7_75t_L     g06066(.A1(\b[2] ), .A2(new_n6002), .B1(new_n5992), .B2(\b[1] ), .C(new_n6322), .Y(new_n6323));
  OAI21xp33_ASAP7_75t_L     g06067(.A1(new_n258), .A2(new_n6309), .B(new_n6323), .Y(new_n6324));
  O2A1O1Ixp33_ASAP7_75t_L   g06068(.A1(new_n5745), .A2(new_n6004), .B(\a[44] ), .C(new_n6324), .Y(new_n6325));
  A2O1A1Ixp33_ASAP7_75t_L   g06069(.A1(\b[0] ), .A2(new_n5990), .B(new_n6004), .C(\a[44] ), .Y(new_n6326));
  O2A1O1Ixp33_ASAP7_75t_L   g06070(.A1(new_n6309), .A2(new_n258), .B(new_n6323), .C(new_n6326), .Y(new_n6327));
  OAI22xp33_ASAP7_75t_L     g06071(.A1(new_n6321), .A2(new_n6320), .B1(new_n6327), .B2(new_n6325), .Y(new_n6328));
  NAND2xp33_ASAP7_75t_L     g06072(.A(new_n6319), .B(new_n6328), .Y(new_n6329));
  NAND2xp33_ASAP7_75t_L     g06073(.A(new_n6329), .B(new_n6299), .Y(new_n6330));
  O2A1O1Ixp33_ASAP7_75t_L   g06074(.A1(new_n5982), .A2(new_n5762), .B(new_n6006), .C(new_n6013), .Y(new_n6331));
  NAND3xp33_ASAP7_75t_L     g06075(.A(new_n6331), .B(new_n6319), .C(new_n6328), .Y(new_n6332));
  AOI22xp33_ASAP7_75t_L     g06076(.A1(new_n6298), .A2(new_n6296), .B1(new_n6332), .B2(new_n6330), .Y(new_n6333));
  INVx1_ASAP7_75t_L         g06077(.A(new_n6296), .Y(new_n6334));
  AOI21xp33_ASAP7_75t_L     g06078(.A1(new_n6328), .A2(new_n6319), .B(new_n6331), .Y(new_n6335));
  NOR2xp33_ASAP7_75t_L      g06079(.A(new_n6329), .B(new_n6299), .Y(new_n6336));
  NOR4xp25_ASAP7_75t_L      g06080(.A(new_n6336), .B(new_n6335), .C(new_n6334), .D(new_n6297), .Y(new_n6337));
  NOR2xp33_ASAP7_75t_L      g06081(.A(new_n6333), .B(new_n6337), .Y(new_n6338));
  A2O1A1Ixp33_ASAP7_75t_L   g06082(.A1(new_n6027), .A2(new_n6024), .B(new_n6291), .C(new_n6338), .Y(new_n6339));
  AOI21xp33_ASAP7_75t_L     g06083(.A1(new_n6024), .A2(new_n6027), .B(new_n6291), .Y(new_n6340));
  NAND2xp33_ASAP7_75t_L     g06084(.A(new_n6296), .B(new_n6298), .Y(new_n6341));
  OAI21xp33_ASAP7_75t_L     g06085(.A1(new_n6335), .A2(new_n6336), .B(new_n6341), .Y(new_n6342));
  NAND4xp25_ASAP7_75t_L     g06086(.A(new_n6330), .B(new_n6332), .C(new_n6296), .D(new_n6298), .Y(new_n6343));
  NAND2xp33_ASAP7_75t_L     g06087(.A(new_n6343), .B(new_n6342), .Y(new_n6344));
  NAND2xp33_ASAP7_75t_L     g06088(.A(new_n6344), .B(new_n6340), .Y(new_n6345));
  NOR2xp33_ASAP7_75t_L      g06089(.A(new_n559), .B(new_n4986), .Y(new_n6346));
  NAND2xp33_ASAP7_75t_L     g06090(.A(\b[10] ), .B(new_n3874), .Y(new_n6347));
  OAI221xp5_ASAP7_75t_L     g06091(.A1(new_n4115), .A2(new_n695), .B1(new_n4114), .B2(new_n701), .C(new_n6347), .Y(new_n6348));
  OR3x1_ASAP7_75t_L         g06092(.A(new_n6348), .B(new_n3878), .C(new_n6346), .Y(new_n6349));
  A2O1A1Ixp33_ASAP7_75t_L   g06093(.A1(\b[9] ), .A2(new_n4111), .B(new_n6348), .C(new_n3878), .Y(new_n6350));
  AND2x2_ASAP7_75t_L        g06094(.A(new_n6350), .B(new_n6349), .Y(new_n6351));
  NAND3xp33_ASAP7_75t_L     g06095(.A(new_n6351), .B(new_n6345), .C(new_n6339), .Y(new_n6352));
  A2O1A1O1Ixp25_ASAP7_75t_L g06096(.A1(new_n6023), .A2(new_n6022), .B(new_n6029), .C(new_n6290), .D(new_n6344), .Y(new_n6353));
  A2O1A1Ixp33_ASAP7_75t_L   g06097(.A1(new_n6023), .A2(new_n6022), .B(new_n6029), .C(new_n6290), .Y(new_n6354));
  NOR2xp33_ASAP7_75t_L      g06098(.A(new_n6338), .B(new_n6354), .Y(new_n6355));
  NAND2xp33_ASAP7_75t_L     g06099(.A(new_n6350), .B(new_n6349), .Y(new_n6356));
  OAI21xp33_ASAP7_75t_L     g06100(.A1(new_n6355), .A2(new_n6353), .B(new_n6356), .Y(new_n6357));
  NAND2xp33_ASAP7_75t_L     g06101(.A(new_n6039), .B(new_n6040), .Y(new_n6358));
  MAJIxp5_ASAP7_75t_L       g06102(.A(new_n5980), .B(new_n6037), .C(new_n6358), .Y(new_n6359));
  NAND3xp33_ASAP7_75t_L     g06103(.A(new_n6359), .B(new_n6357), .C(new_n6352), .Y(new_n6360));
  NOR3xp33_ASAP7_75t_L      g06104(.A(new_n6353), .B(new_n6356), .C(new_n6355), .Y(new_n6361));
  AOI21xp33_ASAP7_75t_L     g06105(.A1(new_n6345), .A2(new_n6339), .B(new_n6351), .Y(new_n6362));
  A2O1A1Ixp33_ASAP7_75t_L   g06106(.A1(new_n5797), .A2(new_n5786), .B(new_n5799), .C(new_n6038), .Y(new_n6363));
  OAI211xp5_ASAP7_75t_L     g06107(.A1(new_n6361), .A2(new_n6362), .B(new_n6041), .C(new_n6363), .Y(new_n6364));
  AOI21xp33_ASAP7_75t_L     g06108(.A1(new_n6364), .A2(new_n6360), .B(new_n6289), .Y(new_n6365));
  AOI211xp5_ASAP7_75t_L     g06109(.A1(new_n6363), .A2(new_n6041), .B(new_n6361), .C(new_n6362), .Y(new_n6366));
  AOI21xp33_ASAP7_75t_L     g06110(.A1(new_n6357), .A2(new_n6352), .B(new_n6359), .Y(new_n6367));
  NOR3xp33_ASAP7_75t_L      g06111(.A(new_n6366), .B(new_n6367), .C(new_n6288), .Y(new_n6368));
  NOR3xp33_ASAP7_75t_L      g06112(.A(new_n6282), .B(new_n6365), .C(new_n6368), .Y(new_n6369));
  A2O1A1Ixp33_ASAP7_75t_L   g06113(.A1(new_n5804), .A2(new_n5970), .B(new_n6054), .C(new_n6048), .Y(new_n6370));
  NOR2xp33_ASAP7_75t_L      g06114(.A(new_n6368), .B(new_n6365), .Y(new_n6371));
  NOR2xp33_ASAP7_75t_L      g06115(.A(new_n6370), .B(new_n6371), .Y(new_n6372));
  OAI21xp33_ASAP7_75t_L     g06116(.A1(new_n6369), .A2(new_n6372), .B(new_n6281), .Y(new_n6373));
  INVx1_ASAP7_75t_L         g06117(.A(new_n6281), .Y(new_n6374));
  A2O1A1Ixp33_ASAP7_75t_L   g06118(.A1(new_n6045), .A2(new_n5971), .B(new_n6055), .C(new_n6371), .Y(new_n6375));
  OAI21xp33_ASAP7_75t_L     g06119(.A1(new_n6365), .A2(new_n6368), .B(new_n6282), .Y(new_n6376));
  NAND3xp33_ASAP7_75t_L     g06120(.A(new_n6375), .B(new_n6374), .C(new_n6376), .Y(new_n6377));
  NAND3xp33_ASAP7_75t_L     g06121(.A(new_n6275), .B(new_n6373), .C(new_n6377), .Y(new_n6378));
  NOR2xp33_ASAP7_75t_L      g06122(.A(new_n6064), .B(new_n6063), .Y(new_n6379));
  MAJIxp5_ASAP7_75t_L       g06123(.A(new_n6073), .B(new_n6065), .C(new_n6379), .Y(new_n6380));
  AOI21xp33_ASAP7_75t_L     g06124(.A1(new_n6375), .A2(new_n6376), .B(new_n6374), .Y(new_n6381));
  NOR3xp33_ASAP7_75t_L      g06125(.A(new_n6372), .B(new_n6369), .C(new_n6281), .Y(new_n6382));
  OAI21xp33_ASAP7_75t_L     g06126(.A1(new_n6381), .A2(new_n6382), .B(new_n6380), .Y(new_n6383));
  NOR2xp33_ASAP7_75t_L      g06127(.A(new_n1594), .B(new_n2234), .Y(new_n6384));
  AOI221xp5_ASAP7_75t_L     g06128(.A1(new_n2232), .A2(\b[19] ), .B1(new_n2226), .B2(new_n1600), .C(new_n6384), .Y(new_n6385));
  OAI211xp5_ASAP7_75t_L     g06129(.A1(new_n1356), .A2(new_n2387), .B(new_n6385), .C(\a[26] ), .Y(new_n6386));
  INVx1_ASAP7_75t_L         g06130(.A(new_n6386), .Y(new_n6387));
  O2A1O1Ixp33_ASAP7_75t_L   g06131(.A1(new_n1356), .A2(new_n2387), .B(new_n6385), .C(\a[26] ), .Y(new_n6388));
  NOR2xp33_ASAP7_75t_L      g06132(.A(new_n6388), .B(new_n6387), .Y(new_n6389));
  NAND3xp33_ASAP7_75t_L     g06133(.A(new_n6389), .B(new_n6383), .C(new_n6378), .Y(new_n6390));
  NOR3xp33_ASAP7_75t_L      g06134(.A(new_n6380), .B(new_n6381), .C(new_n6382), .Y(new_n6391));
  AOI21xp33_ASAP7_75t_L     g06135(.A1(new_n6377), .A2(new_n6373), .B(new_n6275), .Y(new_n6392));
  INVx1_ASAP7_75t_L         g06136(.A(new_n6388), .Y(new_n6393));
  NAND2xp33_ASAP7_75t_L     g06137(.A(new_n6386), .B(new_n6393), .Y(new_n6394));
  OAI21xp33_ASAP7_75t_L     g06138(.A1(new_n6392), .A2(new_n6391), .B(new_n6394), .Y(new_n6395));
  NOR2xp33_ASAP7_75t_L      g06139(.A(new_n6084), .B(new_n6083), .Y(new_n6396));
  MAJIxp5_ASAP7_75t_L       g06140(.A(new_n6088), .B(new_n6396), .C(new_n6085), .Y(new_n6397));
  NAND3xp33_ASAP7_75t_L     g06141(.A(new_n6397), .B(new_n6395), .C(new_n6390), .Y(new_n6398));
  NAND2xp33_ASAP7_75t_L     g06142(.A(new_n6383), .B(new_n6378), .Y(new_n6399));
  NOR2xp33_ASAP7_75t_L      g06143(.A(new_n6394), .B(new_n6399), .Y(new_n6400));
  AOI21xp33_ASAP7_75t_L     g06144(.A1(new_n6383), .A2(new_n6378), .B(new_n6389), .Y(new_n6401));
  NAND2xp33_ASAP7_75t_L     g06145(.A(new_n6074), .B(new_n6069), .Y(new_n6402));
  MAJIxp5_ASAP7_75t_L       g06146(.A(new_n6090), .B(new_n6402), .C(new_n6079), .Y(new_n6403));
  OAI21xp33_ASAP7_75t_L     g06147(.A1(new_n6401), .A2(new_n6400), .B(new_n6403), .Y(new_n6404));
  AOI32xp33_ASAP7_75t_L     g06148(.A1(new_n1998), .A2(new_n2001), .A3(new_n1764), .B1(new_n1766), .B2(\b[23] ), .Y(new_n6405));
  OAI221xp5_ASAP7_75t_L     g06149(.A1(new_n1758), .A2(new_n1857), .B1(new_n1709), .B2(new_n1911), .C(new_n6405), .Y(new_n6406));
  XNOR2x2_ASAP7_75t_L       g06150(.A(new_n1761), .B(new_n6406), .Y(new_n6407));
  AO21x2_ASAP7_75t_L        g06151(.A1(new_n6404), .A2(new_n6398), .B(new_n6407), .Y(new_n6408));
  NAND3xp33_ASAP7_75t_L     g06152(.A(new_n6398), .B(new_n6404), .C(new_n6407), .Y(new_n6409));
  NAND2xp33_ASAP7_75t_L     g06153(.A(new_n6409), .B(new_n6408), .Y(new_n6410));
  NOR2xp33_ASAP7_75t_L      g06154(.A(new_n6410), .B(new_n6273), .Y(new_n6411));
  A2O1A1O1Ixp25_ASAP7_75t_L g06155(.A1(new_n5602), .A2(new_n5854), .B(new_n5849), .C(new_n5855), .D(new_n6108), .Y(new_n6412));
  AOI21xp33_ASAP7_75t_L     g06156(.A1(new_n6398), .A2(new_n6404), .B(new_n6407), .Y(new_n6413));
  AND3x1_ASAP7_75t_L        g06157(.A(new_n6398), .B(new_n6404), .C(new_n6407), .Y(new_n6414));
  NOR2xp33_ASAP7_75t_L      g06158(.A(new_n6413), .B(new_n6414), .Y(new_n6415));
  O2A1O1Ixp33_ASAP7_75t_L   g06159(.A1(new_n6106), .A2(new_n6412), .B(new_n6272), .C(new_n6415), .Y(new_n6416));
  NOR3xp33_ASAP7_75t_L      g06160(.A(new_n6416), .B(new_n6411), .C(new_n6270), .Y(new_n6417));
  NAND4xp25_ASAP7_75t_L     g06161(.A(new_n6115), .B(new_n6409), .C(new_n6408), .D(new_n6272), .Y(new_n6418));
  A2O1A1Ixp33_ASAP7_75t_L   g06162(.A1(new_n6114), .A2(new_n6113), .B(new_n6271), .C(new_n6410), .Y(new_n6419));
  AOI21xp33_ASAP7_75t_L     g06163(.A1(new_n6419), .A2(new_n6418), .B(new_n6269), .Y(new_n6420));
  NOR3xp33_ASAP7_75t_L      g06164(.A(new_n6266), .B(new_n6417), .C(new_n6420), .Y(new_n6421));
  NOR3xp33_ASAP7_75t_L      g06165(.A(new_n6124), .B(new_n6123), .C(new_n6121), .Y(new_n6422));
  INVx1_ASAP7_75t_L         g06166(.A(new_n6422), .Y(new_n6423));
  A2O1A1Ixp33_ASAP7_75t_L   g06167(.A1(new_n6126), .A2(new_n6122), .B(new_n6127), .C(new_n6423), .Y(new_n6424));
  NAND3xp33_ASAP7_75t_L     g06168(.A(new_n6419), .B(new_n6418), .C(new_n6269), .Y(new_n6425));
  OAI21xp33_ASAP7_75t_L     g06169(.A1(new_n6411), .A2(new_n6416), .B(new_n6270), .Y(new_n6426));
  AOI21xp33_ASAP7_75t_L     g06170(.A1(new_n6426), .A2(new_n6425), .B(new_n6424), .Y(new_n6427));
  OAI21xp33_ASAP7_75t_L     g06171(.A1(new_n6421), .A2(new_n6427), .B(new_n6264), .Y(new_n6428));
  NAND2xp33_ASAP7_75t_L     g06172(.A(new_n6261), .B(new_n6263), .Y(new_n6429));
  NAND3xp33_ASAP7_75t_L     g06173(.A(new_n6424), .B(new_n6425), .C(new_n6426), .Y(new_n6430));
  OAI21xp33_ASAP7_75t_L     g06174(.A1(new_n6420), .A2(new_n6417), .B(new_n6266), .Y(new_n6431));
  NAND3xp33_ASAP7_75t_L     g06175(.A(new_n6430), .B(new_n6429), .C(new_n6431), .Y(new_n6432));
  NAND2xp33_ASAP7_75t_L     g06176(.A(new_n6432), .B(new_n6428), .Y(new_n6433));
  NOR2xp33_ASAP7_75t_L      g06177(.A(new_n6257), .B(new_n6433), .Y(new_n6434));
  MAJIxp5_ASAP7_75t_L       g06178(.A(new_n6138), .B(new_n5968), .C(new_n6255), .Y(new_n6435));
  AOI21xp33_ASAP7_75t_L     g06179(.A1(new_n6432), .A2(new_n6428), .B(new_n6435), .Y(new_n6436));
  OAI21xp33_ASAP7_75t_L     g06180(.A1(new_n6436), .A2(new_n6434), .B(new_n6252), .Y(new_n6437));
  NAND2xp33_ASAP7_75t_L     g06181(.A(new_n6249), .B(new_n6251), .Y(new_n6438));
  NAND3xp33_ASAP7_75t_L     g06182(.A(new_n6435), .B(new_n6428), .C(new_n6432), .Y(new_n6439));
  NAND2xp33_ASAP7_75t_L     g06183(.A(new_n6257), .B(new_n6433), .Y(new_n6440));
  NAND3xp33_ASAP7_75t_L     g06184(.A(new_n6439), .B(new_n6440), .C(new_n6438), .Y(new_n6441));
  NAND3xp33_ASAP7_75t_L     g06185(.A(new_n6245), .B(new_n6437), .C(new_n6441), .Y(new_n6442));
  A2O1A1O1Ixp25_ASAP7_75t_L g06186(.A1(new_n5898), .A2(new_n5909), .B(new_n5891), .C(new_n6148), .D(new_n6156), .Y(new_n6443));
  AOI21xp33_ASAP7_75t_L     g06187(.A1(new_n6439), .A2(new_n6440), .B(new_n6438), .Y(new_n6444));
  NOR3xp33_ASAP7_75t_L      g06188(.A(new_n6434), .B(new_n6436), .C(new_n6252), .Y(new_n6445));
  OAI21xp33_ASAP7_75t_L     g06189(.A1(new_n6444), .A2(new_n6445), .B(new_n6443), .Y(new_n6446));
  NAND2xp33_ASAP7_75t_L     g06190(.A(\b[33] ), .B(new_n674), .Y(new_n6447));
  NAND2xp33_ASAP7_75t_L     g06191(.A(\b[34] ), .B(new_n590), .Y(new_n6448));
  AOI22xp33_ASAP7_75t_L     g06192(.A1(new_n600), .A2(\b[35] ), .B1(new_n597), .B2(new_n5649), .Y(new_n6449));
  AND4x1_ASAP7_75t_L        g06193(.A(new_n6449), .B(new_n6448), .C(new_n6447), .D(\a[11] ), .Y(new_n6450));
  AOI31xp33_ASAP7_75t_L     g06194(.A1(new_n6449), .A2(new_n6448), .A3(new_n6447), .B(\a[11] ), .Y(new_n6451));
  NOR2xp33_ASAP7_75t_L      g06195(.A(new_n6451), .B(new_n6450), .Y(new_n6452));
  NAND3xp33_ASAP7_75t_L     g06196(.A(new_n6442), .B(new_n6446), .C(new_n6452), .Y(new_n6453));
  NOR3xp33_ASAP7_75t_L      g06197(.A(new_n6443), .B(new_n6445), .C(new_n6444), .Y(new_n6454));
  AOI221xp5_ASAP7_75t_L     g06198(.A1(new_n5960), .A2(new_n6148), .B1(new_n6441), .B2(new_n6437), .C(new_n6156), .Y(new_n6455));
  INVx1_ASAP7_75t_L         g06199(.A(new_n6452), .Y(new_n6456));
  OAI21xp33_ASAP7_75t_L     g06200(.A1(new_n6454), .A2(new_n6455), .B(new_n6456), .Y(new_n6457));
  NAND2xp33_ASAP7_75t_L     g06201(.A(new_n6153), .B(new_n6157), .Y(new_n6458));
  INVx1_ASAP7_75t_L         g06202(.A(new_n6458), .Y(new_n6459));
  INVx1_ASAP7_75t_L         g06203(.A(new_n6163), .Y(new_n6460));
  NAND2xp33_ASAP7_75t_L     g06204(.A(new_n6460), .B(new_n6459), .Y(new_n6461));
  NAND4xp25_ASAP7_75t_L     g06205(.A(new_n6244), .B(new_n6461), .C(new_n6457), .D(new_n6453), .Y(new_n6462));
  NAND2xp33_ASAP7_75t_L     g06206(.A(new_n6457), .B(new_n6453), .Y(new_n6463));
  MAJIxp5_ASAP7_75t_L       g06207(.A(new_n5916), .B(new_n5917), .C(new_n5906), .Y(new_n6464));
  MAJIxp5_ASAP7_75t_L       g06208(.A(new_n6464), .B(new_n6458), .C(new_n6163), .Y(new_n6465));
  NAND2xp33_ASAP7_75t_L     g06209(.A(new_n6465), .B(new_n6463), .Y(new_n6466));
  NAND2xp33_ASAP7_75t_L     g06210(.A(\b[36] ), .B(new_n480), .Y(new_n6467));
  NAND2xp33_ASAP7_75t_L     g06211(.A(\b[37] ), .B(new_n441), .Y(new_n6468));
  AOI22xp33_ASAP7_75t_L     g06212(.A1(new_n451), .A2(\b[38] ), .B1(new_n448), .B2(new_n4923), .Y(new_n6469));
  AND4x1_ASAP7_75t_L        g06213(.A(new_n6469), .B(new_n6468), .C(new_n6467), .D(\a[8] ), .Y(new_n6470));
  AOI31xp33_ASAP7_75t_L     g06214(.A1(new_n6469), .A2(new_n6468), .A3(new_n6467), .B(\a[8] ), .Y(new_n6471));
  NOR2xp33_ASAP7_75t_L      g06215(.A(new_n6471), .B(new_n6470), .Y(new_n6472));
  NAND3xp33_ASAP7_75t_L     g06216(.A(new_n6466), .B(new_n6462), .C(new_n6472), .Y(new_n6473));
  AO21x2_ASAP7_75t_L        g06217(.A1(new_n6462), .A2(new_n6466), .B(new_n6472), .Y(new_n6474));
  NOR3xp33_ASAP7_75t_L      g06218(.A(new_n6168), .B(new_n6174), .C(new_n6167), .Y(new_n6475));
  A2O1A1O1Ixp25_ASAP7_75t_L g06219(.A1(new_n5921), .A2(new_n5700), .B(new_n5922), .C(new_n6175), .D(new_n6475), .Y(new_n6476));
  AO21x2_ASAP7_75t_L        g06220(.A1(new_n6473), .A2(new_n6474), .B(new_n6476), .Y(new_n6477));
  NAND3xp33_ASAP7_75t_L     g06221(.A(new_n6476), .B(new_n6474), .C(new_n6473), .Y(new_n6478));
  AOI21xp33_ASAP7_75t_L     g06222(.A1(new_n6477), .A2(new_n6478), .B(new_n6243), .Y(new_n6479));
  AOI21xp33_ASAP7_75t_L     g06223(.A1(new_n6474), .A2(new_n6473), .B(new_n6476), .Y(new_n6480));
  AND3x1_ASAP7_75t_L        g06224(.A(new_n6476), .B(new_n6474), .C(new_n6473), .Y(new_n6481));
  NOR3xp33_ASAP7_75t_L      g06225(.A(new_n6481), .B(new_n6480), .C(new_n6242), .Y(new_n6482));
  NOR2xp33_ASAP7_75t_L      g06226(.A(new_n6479), .B(new_n6482), .Y(new_n6483));
  O2A1O1Ixp33_ASAP7_75t_L   g06227(.A1(new_n6186), .A2(new_n6185), .B(new_n6183), .C(new_n6483), .Y(new_n6484));
  AO21x2_ASAP7_75t_L        g06228(.A1(new_n5661), .A2(new_n5445), .B(new_n5659), .Y(new_n6485));
  A2O1A1O1Ixp25_ASAP7_75t_L g06229(.A1(new_n5936), .A2(new_n6485), .B(new_n5947), .C(new_n6180), .D(new_n6187), .Y(new_n6486));
  AND2x2_ASAP7_75t_L        g06230(.A(new_n6483), .B(new_n6486), .Y(new_n6487));
  NOR3xp33_ASAP7_75t_L      g06231(.A(new_n6487), .B(new_n6235), .C(new_n6484), .Y(new_n6488));
  INVx1_ASAP7_75t_L         g06232(.A(new_n6488), .Y(new_n6489));
  OAI21xp33_ASAP7_75t_L     g06233(.A1(new_n6484), .A2(new_n6487), .B(new_n6235), .Y(new_n6490));
  NAND2xp33_ASAP7_75t_L     g06234(.A(new_n6490), .B(new_n6489), .Y(new_n6491));
  XOR2x2_ASAP7_75t_L        g06235(.A(new_n6491), .B(new_n6218), .Y(\f[44] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g06236(.A1(new_n6213), .A2(new_n6214), .B(new_n6217), .C(new_n6490), .D(new_n6488), .Y(new_n6493));
  NAND2xp33_ASAP7_75t_L     g06237(.A(new_n6446), .B(new_n6442), .Y(new_n6494));
  NOR2xp33_ASAP7_75t_L      g06238(.A(new_n6452), .B(new_n6494), .Y(new_n6495));
  A2O1A1O1Ixp25_ASAP7_75t_L g06239(.A1(new_n6460), .A2(new_n6459), .B(new_n6168), .C(new_n6463), .D(new_n6495), .Y(new_n6496));
  NAND2xp33_ASAP7_75t_L     g06240(.A(\b[34] ), .B(new_n674), .Y(new_n6497));
  NAND2xp33_ASAP7_75t_L     g06241(.A(\b[35] ), .B(new_n590), .Y(new_n6498));
  AOI22xp33_ASAP7_75t_L     g06242(.A1(new_n600), .A2(\b[36] ), .B1(new_n597), .B2(new_n4473), .Y(new_n6499));
  AND4x1_ASAP7_75t_L        g06243(.A(new_n6499), .B(new_n6498), .C(new_n6497), .D(\a[11] ), .Y(new_n6500));
  AOI31xp33_ASAP7_75t_L     g06244(.A1(new_n6499), .A2(new_n6498), .A3(new_n6497), .B(\a[11] ), .Y(new_n6501));
  OAI21xp33_ASAP7_75t_L     g06245(.A1(new_n6444), .A2(new_n6443), .B(new_n6441), .Y(new_n6502));
  NOR3xp33_ASAP7_75t_L      g06246(.A(new_n6427), .B(new_n6264), .C(new_n6421), .Y(new_n6503));
  NAND2xp33_ASAP7_75t_L     g06247(.A(\b[28] ), .B(new_n1194), .Y(new_n6504));
  NAND2xp33_ASAP7_75t_L     g06248(.A(\b[29] ), .B(new_n1103), .Y(new_n6505));
  AOI22xp33_ASAP7_75t_L     g06249(.A1(new_n1113), .A2(\b[30] ), .B1(new_n1110), .B2(new_n3219), .Y(new_n6506));
  NAND4xp25_ASAP7_75t_L     g06250(.A(new_n6506), .B(\a[17] ), .C(new_n6504), .D(new_n6505), .Y(new_n6507));
  NAND2xp33_ASAP7_75t_L     g06251(.A(new_n6505), .B(new_n6506), .Y(new_n6508));
  A2O1A1Ixp33_ASAP7_75t_L   g06252(.A1(\b[28] ), .A2(new_n1194), .B(new_n6508), .C(new_n1107), .Y(new_n6509));
  AND2x2_ASAP7_75t_L        g06253(.A(new_n6507), .B(new_n6509), .Y(new_n6510));
  A2O1A1O1Ixp25_ASAP7_75t_L g06254(.A1(new_n6130), .A2(new_n6129), .B(new_n6422), .C(new_n6425), .D(new_n6420), .Y(new_n6511));
  NOR2xp33_ASAP7_75t_L      g06255(.A(new_n6061), .B(new_n6274), .Y(new_n6512));
  INVx1_ASAP7_75t_L         g06256(.A(new_n6512), .Y(new_n6513));
  A2O1A1Ixp33_ASAP7_75t_L   g06257(.A1(new_n6074), .A2(new_n6513), .B(new_n6381), .C(new_n6377), .Y(new_n6514));
  INVx1_ASAP7_75t_L         g06258(.A(new_n6368), .Y(new_n6515));
  OAI21xp33_ASAP7_75t_L     g06259(.A1(new_n6365), .A2(new_n6282), .B(new_n6515), .Y(new_n6516));
  NOR2xp33_ASAP7_75t_L      g06260(.A(new_n793), .B(new_n3492), .Y(new_n6517));
  INVx1_ASAP7_75t_L         g06261(.A(new_n6517), .Y(new_n6518));
  NAND2xp33_ASAP7_75t_L     g06262(.A(\b[14] ), .B(new_n3260), .Y(new_n6519));
  AOI22xp33_ASAP7_75t_L     g06263(.A1(new_n3256), .A2(\b[15] ), .B1(new_n3254), .B2(new_n959), .Y(new_n6520));
  NAND4xp25_ASAP7_75t_L     g06264(.A(new_n6520), .B(\a[32] ), .C(new_n6518), .D(new_n6519), .Y(new_n6521));
  AOI31xp33_ASAP7_75t_L     g06265(.A1(new_n6520), .A2(new_n6519), .A3(new_n6518), .B(\a[32] ), .Y(new_n6522));
  INVx1_ASAP7_75t_L         g06266(.A(new_n6522), .Y(new_n6523));
  AND2x2_ASAP7_75t_L        g06267(.A(new_n6521), .B(new_n6523), .Y(new_n6524));
  A2O1A1Ixp33_ASAP7_75t_L   g06268(.A1(new_n6363), .A2(new_n6041), .B(new_n6361), .C(new_n6357), .Y(new_n6525));
  NOR2xp33_ASAP7_75t_L      g06269(.A(new_n631), .B(new_n4986), .Y(new_n6526));
  INVx1_ASAP7_75t_L         g06270(.A(new_n6526), .Y(new_n6527));
  NOR2xp33_ASAP7_75t_L      g06271(.A(new_n695), .B(new_n4312), .Y(new_n6528));
  INVx1_ASAP7_75t_L         g06272(.A(new_n6528), .Y(new_n6529));
  AOI22xp33_ASAP7_75t_L     g06273(.A1(new_n3884), .A2(\b[12] ), .B1(new_n3881), .B2(new_n970), .Y(new_n6530));
  AND4x1_ASAP7_75t_L        g06274(.A(new_n6530), .B(new_n6529), .C(new_n6527), .D(\a[35] ), .Y(new_n6531));
  AOI31xp33_ASAP7_75t_L     g06275(.A1(new_n6530), .A2(new_n6529), .A3(new_n6527), .B(\a[35] ), .Y(new_n6532));
  NOR2xp33_ASAP7_75t_L      g06276(.A(new_n6532), .B(new_n6531), .Y(new_n6533));
  NAND3xp33_ASAP7_75t_L     g06277(.A(new_n6341), .B(new_n6330), .C(new_n6332), .Y(new_n6534));
  INVx1_ASAP7_75t_L         g06278(.A(new_n6534), .Y(new_n6535));
  NAND5xp2_ASAP7_75t_L      g06279(.A(new_n6003), .B(new_n6000), .C(new_n5993), .D(new_n5981), .E(\a[44] ), .Y(new_n6536));
  INVx1_ASAP7_75t_L         g06280(.A(\a[45] ), .Y(new_n6537));
  NAND2xp33_ASAP7_75t_L     g06281(.A(\a[44] ), .B(new_n6537), .Y(new_n6538));
  NAND2xp33_ASAP7_75t_L     g06282(.A(\a[45] ), .B(new_n5996), .Y(new_n6539));
  AND2x2_ASAP7_75t_L        g06283(.A(new_n6538), .B(new_n6539), .Y(new_n6540));
  NOR2xp33_ASAP7_75t_L      g06284(.A(new_n258), .B(new_n6540), .Y(new_n6541));
  OAI31xp33_ASAP7_75t_L     g06285(.A1(new_n6536), .A2(new_n6314), .A3(new_n6310), .B(new_n6541), .Y(new_n6542));
  OR4x2_ASAP7_75t_L         g06286(.A(new_n6541), .B(new_n6536), .C(new_n6314), .D(new_n6310), .Y(new_n6543));
  NAND2xp33_ASAP7_75t_L     g06287(.A(new_n6307), .B(new_n5744), .Y(new_n6544));
  NAND2xp33_ASAP7_75t_L     g06288(.A(\b[3] ), .B(new_n6002), .Y(new_n6545));
  OAI221xp5_ASAP7_75t_L     g06289(.A1(new_n278), .A2(new_n6544), .B1(new_n6311), .B2(new_n303), .C(new_n6545), .Y(new_n6546));
  AO211x2_ASAP7_75t_L       g06290(.A1(\b[1] ), .A2(new_n6308), .B(new_n5996), .C(new_n6546), .Y(new_n6547));
  A2O1A1Ixp33_ASAP7_75t_L   g06291(.A1(\b[1] ), .A2(new_n6308), .B(new_n6546), .C(new_n5996), .Y(new_n6548));
  AOI22xp33_ASAP7_75t_L     g06292(.A1(new_n6547), .A2(new_n6548), .B1(new_n6542), .B2(new_n6543), .Y(new_n6549));
  AND4x1_ASAP7_75t_L        g06293(.A(new_n6543), .B(new_n6542), .C(new_n6548), .D(new_n6547), .Y(new_n6550));
  NAND2xp33_ASAP7_75t_L     g06294(.A(\b[5] ), .B(new_n5240), .Y(new_n6551));
  NAND2xp33_ASAP7_75t_L     g06295(.A(\b[6] ), .B(new_n5249), .Y(new_n6552));
  OAI311xp33_ASAP7_75t_L    g06296(.A1(new_n388), .A2(new_n386), .A3(new_n5252), .B1(new_n6552), .C1(new_n6551), .Y(new_n6553));
  AOI211xp5_ASAP7_75t_L     g06297(.A1(\b[4] ), .A2(new_n5526), .B(new_n5244), .C(new_n6553), .Y(new_n6554));
  A2O1A1Ixp33_ASAP7_75t_L   g06298(.A1(\b[4] ), .A2(new_n5526), .B(new_n6553), .C(new_n5244), .Y(new_n6555));
  INVx1_ASAP7_75t_L         g06299(.A(new_n6555), .Y(new_n6556));
  NOR4xp25_ASAP7_75t_L      g06300(.A(new_n6550), .B(new_n6556), .C(new_n6549), .D(new_n6554), .Y(new_n6557));
  AO22x1_ASAP7_75t_L        g06301(.A1(new_n6548), .A2(new_n6547), .B1(new_n6542), .B2(new_n6543), .Y(new_n6558));
  NAND4xp25_ASAP7_75t_L     g06302(.A(new_n6543), .B(new_n6542), .C(new_n6547), .D(new_n6548), .Y(new_n6559));
  INVx1_ASAP7_75t_L         g06303(.A(new_n6554), .Y(new_n6560));
  AOI22xp33_ASAP7_75t_L     g06304(.A1(new_n6560), .A2(new_n6555), .B1(new_n6559), .B2(new_n6558), .Y(new_n6561));
  NOR2xp33_ASAP7_75t_L      g06305(.A(new_n6557), .B(new_n6561), .Y(new_n6562));
  NAND2xp33_ASAP7_75t_L     g06306(.A(new_n6305), .B(new_n6303), .Y(new_n6563));
  NOR2xp33_ASAP7_75t_L      g06307(.A(new_n6325), .B(new_n6327), .Y(new_n6564));
  NAND2xp33_ASAP7_75t_L     g06308(.A(new_n6563), .B(new_n6564), .Y(new_n6565));
  NAND3xp33_ASAP7_75t_L     g06309(.A(new_n6330), .B(new_n6562), .C(new_n6565), .Y(new_n6566));
  NAND4xp25_ASAP7_75t_L     g06310(.A(new_n6558), .B(new_n6555), .C(new_n6560), .D(new_n6559), .Y(new_n6567));
  OAI22xp33_ASAP7_75t_L     g06311(.A1(new_n6550), .A2(new_n6549), .B1(new_n6556), .B2(new_n6554), .Y(new_n6568));
  NAND2xp33_ASAP7_75t_L     g06312(.A(new_n6567), .B(new_n6568), .Y(new_n6569));
  A2O1A1Ixp33_ASAP7_75t_L   g06313(.A1(new_n6564), .A2(new_n6563), .B(new_n6335), .C(new_n6569), .Y(new_n6570));
  NAND2xp33_ASAP7_75t_L     g06314(.A(\b[7] ), .B(new_n4780), .Y(new_n6571));
  NAND2xp33_ASAP7_75t_L     g06315(.A(\b[8] ), .B(new_n4548), .Y(new_n6572));
  AOI32xp33_ASAP7_75t_L     g06316(.A1(new_n765), .A2(new_n977), .A3(new_n4542), .B1(new_n4544), .B2(\b[9] ), .Y(new_n6573));
  NAND4xp25_ASAP7_75t_L     g06317(.A(new_n6573), .B(\a[38] ), .C(new_n6571), .D(new_n6572), .Y(new_n6574));
  INVx1_ASAP7_75t_L         g06318(.A(new_n6574), .Y(new_n6575));
  AOI31xp33_ASAP7_75t_L     g06319(.A1(new_n6573), .A2(new_n6572), .A3(new_n6571), .B(\a[38] ), .Y(new_n6576));
  AOI211xp5_ASAP7_75t_L     g06320(.A1(new_n6566), .A2(new_n6570), .B(new_n6575), .C(new_n6576), .Y(new_n6577));
  A2O1A1Ixp33_ASAP7_75t_L   g06321(.A1(new_n6319), .A2(new_n6328), .B(new_n6331), .C(new_n6565), .Y(new_n6578));
  NOR2xp33_ASAP7_75t_L      g06322(.A(new_n6569), .B(new_n6578), .Y(new_n6579));
  A2O1A1O1Ixp25_ASAP7_75t_L g06323(.A1(new_n6319), .A2(new_n6328), .B(new_n6331), .C(new_n6565), .D(new_n6562), .Y(new_n6580));
  INVx1_ASAP7_75t_L         g06324(.A(new_n6576), .Y(new_n6581));
  AOI211xp5_ASAP7_75t_L     g06325(.A1(new_n6581), .A2(new_n6574), .B(new_n6579), .C(new_n6580), .Y(new_n6582));
  NOR2xp33_ASAP7_75t_L      g06326(.A(new_n6582), .B(new_n6577), .Y(new_n6583));
  A2O1A1Ixp33_ASAP7_75t_L   g06327(.A1(new_n6344), .A2(new_n6354), .B(new_n6535), .C(new_n6583), .Y(new_n6584));
  A2O1A1O1Ixp25_ASAP7_75t_L g06328(.A1(new_n6027), .A2(new_n6024), .B(new_n6291), .C(new_n6344), .D(new_n6535), .Y(new_n6585));
  OAI211xp5_ASAP7_75t_L     g06329(.A1(new_n6579), .A2(new_n6580), .B(new_n6574), .C(new_n6581), .Y(new_n6586));
  OAI211xp5_ASAP7_75t_L     g06330(.A1(new_n6575), .A2(new_n6576), .B(new_n6566), .C(new_n6570), .Y(new_n6587));
  NAND2xp33_ASAP7_75t_L     g06331(.A(new_n6587), .B(new_n6586), .Y(new_n6588));
  NAND2xp33_ASAP7_75t_L     g06332(.A(new_n6588), .B(new_n6585), .Y(new_n6589));
  AOI21xp33_ASAP7_75t_L     g06333(.A1(new_n6584), .A2(new_n6589), .B(new_n6533), .Y(new_n6590));
  OR2x4_ASAP7_75t_L         g06334(.A(new_n6532), .B(new_n6531), .Y(new_n6591));
  NOR2xp33_ASAP7_75t_L      g06335(.A(new_n6588), .B(new_n6585), .Y(new_n6592));
  OAI21xp33_ASAP7_75t_L     g06336(.A1(new_n6338), .A2(new_n6340), .B(new_n6534), .Y(new_n6593));
  NOR2xp33_ASAP7_75t_L      g06337(.A(new_n6593), .B(new_n6583), .Y(new_n6594));
  NOR3xp33_ASAP7_75t_L      g06338(.A(new_n6591), .B(new_n6594), .C(new_n6592), .Y(new_n6595));
  OAI21xp33_ASAP7_75t_L     g06339(.A1(new_n6590), .A2(new_n6595), .B(new_n6525), .Y(new_n6596));
  AOI21xp33_ASAP7_75t_L     g06340(.A1(new_n6359), .A2(new_n6352), .B(new_n6362), .Y(new_n6597));
  OAI21xp33_ASAP7_75t_L     g06341(.A1(new_n6592), .A2(new_n6594), .B(new_n6591), .Y(new_n6598));
  NAND3xp33_ASAP7_75t_L     g06342(.A(new_n6584), .B(new_n6589), .C(new_n6533), .Y(new_n6599));
  NAND3xp33_ASAP7_75t_L     g06343(.A(new_n6597), .B(new_n6598), .C(new_n6599), .Y(new_n6600));
  NAND3xp33_ASAP7_75t_L     g06344(.A(new_n6524), .B(new_n6596), .C(new_n6600), .Y(new_n6601));
  NAND2xp33_ASAP7_75t_L     g06345(.A(new_n6521), .B(new_n6523), .Y(new_n6602));
  AOI21xp33_ASAP7_75t_L     g06346(.A1(new_n6599), .A2(new_n6598), .B(new_n6597), .Y(new_n6603));
  NAND2xp33_ASAP7_75t_L     g06347(.A(new_n6599), .B(new_n6598), .Y(new_n6604));
  NOR2xp33_ASAP7_75t_L      g06348(.A(new_n6525), .B(new_n6604), .Y(new_n6605));
  OAI21xp33_ASAP7_75t_L     g06349(.A1(new_n6603), .A2(new_n6605), .B(new_n6602), .Y(new_n6606));
  NAND3xp33_ASAP7_75t_L     g06350(.A(new_n6516), .B(new_n6601), .C(new_n6606), .Y(new_n6607));
  OAI21xp33_ASAP7_75t_L     g06351(.A1(new_n6367), .A2(new_n6366), .B(new_n6288), .Y(new_n6608));
  A2O1A1O1Ixp25_ASAP7_75t_L g06352(.A1(new_n6045), .A2(new_n5971), .B(new_n6055), .C(new_n6608), .D(new_n6368), .Y(new_n6609));
  NOR3xp33_ASAP7_75t_L      g06353(.A(new_n6605), .B(new_n6603), .C(new_n6602), .Y(new_n6610));
  AOI21xp33_ASAP7_75t_L     g06354(.A1(new_n6600), .A2(new_n6596), .B(new_n6524), .Y(new_n6611));
  OAI21xp33_ASAP7_75t_L     g06355(.A1(new_n6610), .A2(new_n6611), .B(new_n6609), .Y(new_n6612));
  NAND2xp33_ASAP7_75t_L     g06356(.A(\b[16] ), .B(new_n2931), .Y(new_n6613));
  NOR2xp33_ASAP7_75t_L      g06357(.A(new_n1356), .B(new_n2708), .Y(new_n6614));
  AOI221xp5_ASAP7_75t_L     g06358(.A1(new_n2706), .A2(\b[17] ), .B1(new_n2700), .B2(new_n1363), .C(new_n6614), .Y(new_n6615));
  AND3x1_ASAP7_75t_L        g06359(.A(new_n6615), .B(new_n6613), .C(\a[29] ), .Y(new_n6616));
  O2A1O1Ixp33_ASAP7_75t_L   g06360(.A1(new_n1051), .A2(new_n2932), .B(new_n6615), .C(\a[29] ), .Y(new_n6617));
  NOR2xp33_ASAP7_75t_L      g06361(.A(new_n6617), .B(new_n6616), .Y(new_n6618));
  AO21x2_ASAP7_75t_L        g06362(.A1(new_n6612), .A2(new_n6607), .B(new_n6618), .Y(new_n6619));
  NAND3xp33_ASAP7_75t_L     g06363(.A(new_n6607), .B(new_n6612), .C(new_n6618), .Y(new_n6620));
  NAND3xp33_ASAP7_75t_L     g06364(.A(new_n6514), .B(new_n6619), .C(new_n6620), .Y(new_n6621));
  NAND2xp33_ASAP7_75t_L     g06365(.A(new_n6066), .B(new_n6062), .Y(new_n6622));
  A2O1A1O1Ixp25_ASAP7_75t_L g06366(.A1(new_n6073), .A2(new_n6622), .B(new_n6512), .C(new_n6373), .D(new_n6382), .Y(new_n6623));
  AOI21xp33_ASAP7_75t_L     g06367(.A1(new_n6607), .A2(new_n6612), .B(new_n6618), .Y(new_n6624));
  AND3x1_ASAP7_75t_L        g06368(.A(new_n6607), .B(new_n6618), .C(new_n6612), .Y(new_n6625));
  OAI21xp33_ASAP7_75t_L     g06369(.A1(new_n6624), .A2(new_n6625), .B(new_n6623), .Y(new_n6626));
  NAND2xp33_ASAP7_75t_L     g06370(.A(\b[19] ), .B(new_n2386), .Y(new_n6627));
  NAND2xp33_ASAP7_75t_L     g06371(.A(\b[20] ), .B(new_n2232), .Y(new_n6628));
  AOI22xp33_ASAP7_75t_L     g06372(.A1(new_n2228), .A2(\b[21] ), .B1(new_n2226), .B2(new_n1715), .Y(new_n6629));
  AND4x1_ASAP7_75t_L        g06373(.A(new_n6629), .B(new_n6628), .C(new_n6627), .D(\a[26] ), .Y(new_n6630));
  AOI31xp33_ASAP7_75t_L     g06374(.A1(new_n6629), .A2(new_n6628), .A3(new_n6627), .B(\a[26] ), .Y(new_n6631));
  NOR2xp33_ASAP7_75t_L      g06375(.A(new_n6631), .B(new_n6630), .Y(new_n6632));
  NAND3xp33_ASAP7_75t_L     g06376(.A(new_n6621), .B(new_n6626), .C(new_n6632), .Y(new_n6633));
  NOR3xp33_ASAP7_75t_L      g06377(.A(new_n6623), .B(new_n6624), .C(new_n6625), .Y(new_n6634));
  AOI221xp5_ASAP7_75t_L     g06378(.A1(new_n6275), .A2(new_n6373), .B1(new_n6620), .B2(new_n6619), .C(new_n6382), .Y(new_n6635));
  INVx1_ASAP7_75t_L         g06379(.A(new_n6632), .Y(new_n6636));
  OAI21xp33_ASAP7_75t_L     g06380(.A1(new_n6635), .A2(new_n6634), .B(new_n6636), .Y(new_n6637));
  NAND2xp33_ASAP7_75t_L     g06381(.A(new_n6637), .B(new_n6633), .Y(new_n6638));
  NOR2xp33_ASAP7_75t_L      g06382(.A(new_n6392), .B(new_n6391), .Y(new_n6639));
  NAND2xp33_ASAP7_75t_L     g06383(.A(new_n6394), .B(new_n6639), .Y(new_n6640));
  A2O1A1Ixp33_ASAP7_75t_L   g06384(.A1(new_n6395), .A2(new_n6390), .B(new_n6397), .C(new_n6640), .Y(new_n6641));
  NOR2xp33_ASAP7_75t_L      g06385(.A(new_n6638), .B(new_n6641), .Y(new_n6642));
  MAJIxp5_ASAP7_75t_L       g06386(.A(new_n6403), .B(new_n6394), .C(new_n6639), .Y(new_n6643));
  AOI21xp33_ASAP7_75t_L     g06387(.A1(new_n6637), .A2(new_n6633), .B(new_n6643), .Y(new_n6644));
  NAND2xp33_ASAP7_75t_L     g06388(.A(\b[22] ), .B(new_n1910), .Y(new_n6645));
  NAND2xp33_ASAP7_75t_L     g06389(.A(\b[23] ), .B(new_n1770), .Y(new_n6646));
  AOI22xp33_ASAP7_75t_L     g06390(.A1(new_n1766), .A2(\b[24] ), .B1(new_n1764), .B2(new_n2027), .Y(new_n6647));
  NAND4xp25_ASAP7_75t_L     g06391(.A(new_n6647), .B(\a[23] ), .C(new_n6645), .D(new_n6646), .Y(new_n6648));
  NAND2xp33_ASAP7_75t_L     g06392(.A(new_n6646), .B(new_n6647), .Y(new_n6649));
  A2O1A1Ixp33_ASAP7_75t_L   g06393(.A1(\b[22] ), .A2(new_n1910), .B(new_n6649), .C(new_n1761), .Y(new_n6650));
  AND2x2_ASAP7_75t_L        g06394(.A(new_n6648), .B(new_n6650), .Y(new_n6651));
  OAI21xp33_ASAP7_75t_L     g06395(.A1(new_n6644), .A2(new_n6642), .B(new_n6651), .Y(new_n6652));
  NAND3xp33_ASAP7_75t_L     g06396(.A(new_n6643), .B(new_n6637), .C(new_n6633), .Y(new_n6653));
  NAND2xp33_ASAP7_75t_L     g06397(.A(new_n6085), .B(new_n6396), .Y(new_n6654));
  AOI22xp33_ASAP7_75t_L     g06398(.A1(new_n6390), .A2(new_n6395), .B1(new_n6654), .B2(new_n6103), .Y(new_n6655));
  INVx1_ASAP7_75t_L         g06399(.A(new_n6640), .Y(new_n6656));
  OAI21xp33_ASAP7_75t_L     g06400(.A1(new_n6656), .A2(new_n6655), .B(new_n6638), .Y(new_n6657));
  NAND2xp33_ASAP7_75t_L     g06401(.A(new_n6648), .B(new_n6650), .Y(new_n6658));
  NAND3xp33_ASAP7_75t_L     g06402(.A(new_n6653), .B(new_n6657), .C(new_n6658), .Y(new_n6659));
  O2A1O1Ixp33_ASAP7_75t_L   g06403(.A1(new_n6106), .A2(new_n6412), .B(new_n6272), .C(new_n6413), .Y(new_n6660));
  OAI211xp5_ASAP7_75t_L     g06404(.A1(new_n6414), .A2(new_n6660), .B(new_n6652), .C(new_n6659), .Y(new_n6661));
  AOI21xp33_ASAP7_75t_L     g06405(.A1(new_n6653), .A2(new_n6657), .B(new_n6658), .Y(new_n6662));
  NOR3xp33_ASAP7_75t_L      g06406(.A(new_n6651), .B(new_n6642), .C(new_n6644), .Y(new_n6663));
  A2O1A1O1Ixp25_ASAP7_75t_L g06407(.A1(new_n6113), .A2(new_n6114), .B(new_n6271), .C(new_n6408), .D(new_n6414), .Y(new_n6664));
  OAI21xp33_ASAP7_75t_L     g06408(.A1(new_n6662), .A2(new_n6663), .B(new_n6664), .Y(new_n6665));
  NOR2xp33_ASAP7_75t_L      g06409(.A(new_n2180), .B(new_n1549), .Y(new_n6666));
  INVx1_ASAP7_75t_L         g06410(.A(new_n6666), .Y(new_n6667));
  NAND2xp33_ASAP7_75t_L     g06411(.A(\b[26] ), .B(new_n1410), .Y(new_n6668));
  AOI22xp33_ASAP7_75t_L     g06412(.A1(new_n1406), .A2(\b[27] ), .B1(new_n1404), .B2(new_n2657), .Y(new_n6669));
  AND4x1_ASAP7_75t_L        g06413(.A(new_n6669), .B(new_n6668), .C(new_n6667), .D(\a[20] ), .Y(new_n6670));
  AOI31xp33_ASAP7_75t_L     g06414(.A1(new_n6669), .A2(new_n6668), .A3(new_n6667), .B(\a[20] ), .Y(new_n6671));
  NOR2xp33_ASAP7_75t_L      g06415(.A(new_n6671), .B(new_n6670), .Y(new_n6672));
  NAND3xp33_ASAP7_75t_L     g06416(.A(new_n6661), .B(new_n6672), .C(new_n6665), .Y(new_n6673));
  NOR3xp33_ASAP7_75t_L      g06417(.A(new_n6664), .B(new_n6663), .C(new_n6662), .Y(new_n6674));
  AOI211xp5_ASAP7_75t_L     g06418(.A1(new_n6652), .A2(new_n6659), .B(new_n6414), .C(new_n6660), .Y(new_n6675));
  INVx1_ASAP7_75t_L         g06419(.A(new_n6672), .Y(new_n6676));
  OAI21xp33_ASAP7_75t_L     g06420(.A1(new_n6674), .A2(new_n6675), .B(new_n6676), .Y(new_n6677));
  AOI21xp33_ASAP7_75t_L     g06421(.A1(new_n6677), .A2(new_n6673), .B(new_n6511), .Y(new_n6678));
  OAI21xp33_ASAP7_75t_L     g06422(.A1(new_n6417), .A2(new_n6266), .B(new_n6426), .Y(new_n6679));
  NAND2xp33_ASAP7_75t_L     g06423(.A(new_n6677), .B(new_n6673), .Y(new_n6680));
  NOR2xp33_ASAP7_75t_L      g06424(.A(new_n6680), .B(new_n6679), .Y(new_n6681));
  NOR3xp33_ASAP7_75t_L      g06425(.A(new_n6681), .B(new_n6678), .C(new_n6510), .Y(new_n6682));
  NAND2xp33_ASAP7_75t_L     g06426(.A(new_n6507), .B(new_n6509), .Y(new_n6683));
  NAND2xp33_ASAP7_75t_L     g06427(.A(new_n6680), .B(new_n6679), .Y(new_n6684));
  NAND3xp33_ASAP7_75t_L     g06428(.A(new_n6511), .B(new_n6673), .C(new_n6677), .Y(new_n6685));
  AOI21xp33_ASAP7_75t_L     g06429(.A1(new_n6684), .A2(new_n6685), .B(new_n6683), .Y(new_n6686));
  NOR2xp33_ASAP7_75t_L      g06430(.A(new_n6686), .B(new_n6682), .Y(new_n6687));
  A2O1A1Ixp33_ASAP7_75t_L   g06431(.A1(new_n6428), .A2(new_n6435), .B(new_n6503), .C(new_n6687), .Y(new_n6688));
  A2O1A1O1Ixp25_ASAP7_75t_L g06432(.A1(new_n5962), .A2(new_n6139), .B(new_n6256), .C(new_n6428), .D(new_n6503), .Y(new_n6689));
  NAND3xp33_ASAP7_75t_L     g06433(.A(new_n6684), .B(new_n6683), .C(new_n6685), .Y(new_n6690));
  OAI21xp33_ASAP7_75t_L     g06434(.A1(new_n6678), .A2(new_n6681), .B(new_n6510), .Y(new_n6691));
  NAND2xp33_ASAP7_75t_L     g06435(.A(new_n6690), .B(new_n6691), .Y(new_n6692));
  NAND2xp33_ASAP7_75t_L     g06436(.A(new_n6689), .B(new_n6692), .Y(new_n6693));
  NAND2xp33_ASAP7_75t_L     g06437(.A(new_n823), .B(new_n3813), .Y(new_n6694));
  OAI221xp5_ASAP7_75t_L     g06438(.A1(new_n912), .A2(new_n3807), .B1(new_n3443), .B2(new_n994), .C(new_n6694), .Y(new_n6695));
  AOI21xp33_ASAP7_75t_L     g06439(.A1(new_n908), .A2(\b[31] ), .B(new_n6695), .Y(new_n6696));
  NAND2xp33_ASAP7_75t_L     g06440(.A(\a[14] ), .B(new_n6696), .Y(new_n6697));
  A2O1A1Ixp33_ASAP7_75t_L   g06441(.A1(\b[31] ), .A2(new_n908), .B(new_n6695), .C(new_n813), .Y(new_n6698));
  AND4x1_ASAP7_75t_L        g06442(.A(new_n6688), .B(new_n6698), .C(new_n6693), .D(new_n6697), .Y(new_n6699));
  NAND2xp33_ASAP7_75t_L     g06443(.A(new_n6698), .B(new_n6697), .Y(new_n6700));
  INVx1_ASAP7_75t_L         g06444(.A(new_n6700), .Y(new_n6701));
  AOI21xp33_ASAP7_75t_L     g06445(.A1(new_n6693), .A2(new_n6688), .B(new_n6701), .Y(new_n6702));
  OAI21xp33_ASAP7_75t_L     g06446(.A1(new_n6699), .A2(new_n6702), .B(new_n6502), .Y(new_n6703));
  A2O1A1O1Ixp25_ASAP7_75t_L g06447(.A1(new_n6148), .A2(new_n5960), .B(new_n6156), .C(new_n6437), .D(new_n6445), .Y(new_n6704));
  XOR2x2_ASAP7_75t_L        g06448(.A(new_n6689), .B(new_n6692), .Y(new_n6705));
  NAND2xp33_ASAP7_75t_L     g06449(.A(new_n6701), .B(new_n6705), .Y(new_n6706));
  XNOR2x2_ASAP7_75t_L       g06450(.A(new_n6689), .B(new_n6692), .Y(new_n6707));
  NAND2xp33_ASAP7_75t_L     g06451(.A(new_n6700), .B(new_n6707), .Y(new_n6708));
  NAND3xp33_ASAP7_75t_L     g06452(.A(new_n6706), .B(new_n6708), .C(new_n6704), .Y(new_n6709));
  OAI211xp5_ASAP7_75t_L     g06453(.A1(new_n6500), .A2(new_n6501), .B(new_n6709), .C(new_n6703), .Y(new_n6710));
  NOR2xp33_ASAP7_75t_L      g06454(.A(new_n6501), .B(new_n6500), .Y(new_n6711));
  AOI21xp33_ASAP7_75t_L     g06455(.A1(new_n6706), .A2(new_n6708), .B(new_n6704), .Y(new_n6712));
  NOR3xp33_ASAP7_75t_L      g06456(.A(new_n6702), .B(new_n6502), .C(new_n6699), .Y(new_n6713));
  OAI21xp33_ASAP7_75t_L     g06457(.A1(new_n6713), .A2(new_n6712), .B(new_n6711), .Y(new_n6714));
  NAND2xp33_ASAP7_75t_L     g06458(.A(new_n6714), .B(new_n6710), .Y(new_n6715));
  NAND2xp33_ASAP7_75t_L     g06459(.A(new_n6715), .B(new_n6496), .Y(new_n6716));
  AOI22xp33_ASAP7_75t_L     g06460(.A1(new_n6453), .A2(new_n6457), .B1(new_n6461), .B2(new_n6244), .Y(new_n6717));
  OAI211xp5_ASAP7_75t_L     g06461(.A1(new_n6495), .A2(new_n6717), .B(new_n6710), .C(new_n6714), .Y(new_n6718));
  NOR2xp33_ASAP7_75t_L      g06462(.A(new_n4701), .B(new_n481), .Y(new_n6719));
  INVx1_ASAP7_75t_L         g06463(.A(new_n6719), .Y(new_n6720));
  NAND2xp33_ASAP7_75t_L     g06464(.A(\b[38] ), .B(new_n441), .Y(new_n6721));
  AOI22xp33_ASAP7_75t_L     g06465(.A1(new_n451), .A2(\b[39] ), .B1(new_n448), .B2(new_n5174), .Y(new_n6722));
  AND4x1_ASAP7_75t_L        g06466(.A(new_n6722), .B(new_n6721), .C(new_n6720), .D(\a[8] ), .Y(new_n6723));
  AOI31xp33_ASAP7_75t_L     g06467(.A1(new_n6722), .A2(new_n6721), .A3(new_n6720), .B(\a[8] ), .Y(new_n6724));
  NOR2xp33_ASAP7_75t_L      g06468(.A(new_n6724), .B(new_n6723), .Y(new_n6725));
  NAND3xp33_ASAP7_75t_L     g06469(.A(new_n6716), .B(new_n6718), .C(new_n6725), .Y(new_n6726));
  AOI211xp5_ASAP7_75t_L     g06470(.A1(new_n6710), .A2(new_n6714), .B(new_n6495), .C(new_n6717), .Y(new_n6727));
  O2A1O1Ixp33_ASAP7_75t_L   g06471(.A1(new_n6494), .A2(new_n6452), .B(new_n6466), .C(new_n6715), .Y(new_n6728));
  INVx1_ASAP7_75t_L         g06472(.A(new_n6725), .Y(new_n6729));
  OAI21xp33_ASAP7_75t_L     g06473(.A1(new_n6727), .A2(new_n6728), .B(new_n6729), .Y(new_n6730));
  OAI211xp5_ASAP7_75t_L     g06474(.A1(new_n6470), .A2(new_n6471), .B(new_n6466), .C(new_n6462), .Y(new_n6731));
  NAND4xp25_ASAP7_75t_L     g06475(.A(new_n6477), .B(new_n6731), .C(new_n6730), .D(new_n6726), .Y(new_n6732));
  NOR3xp33_ASAP7_75t_L      g06476(.A(new_n6728), .B(new_n6729), .C(new_n6727), .Y(new_n6733));
  AOI21xp33_ASAP7_75t_L     g06477(.A1(new_n6716), .A2(new_n6718), .B(new_n6725), .Y(new_n6734));
  NAND2xp33_ASAP7_75t_L     g06478(.A(new_n6462), .B(new_n6466), .Y(new_n6735));
  MAJIxp5_ASAP7_75t_L       g06479(.A(new_n6476), .B(new_n6472), .C(new_n6735), .Y(new_n6736));
  OAI21xp33_ASAP7_75t_L     g06480(.A1(new_n6734), .A2(new_n6733), .B(new_n6736), .Y(new_n6737));
  NOR2xp33_ASAP7_75t_L      g06481(.A(new_n5186), .B(new_n365), .Y(new_n6738));
  INVx1_ASAP7_75t_L         g06482(.A(new_n6738), .Y(new_n6739));
  NAND2xp33_ASAP7_75t_L     g06483(.A(\b[41] ), .B(new_n334), .Y(new_n6740));
  AOI22xp33_ASAP7_75t_L     g06484(.A1(new_n345), .A2(\b[42] ), .B1(new_n342), .B2(new_n5688), .Y(new_n6741));
  AND4x1_ASAP7_75t_L        g06485(.A(new_n6741), .B(new_n6740), .C(new_n6739), .D(\a[5] ), .Y(new_n6742));
  AOI31xp33_ASAP7_75t_L     g06486(.A1(new_n6741), .A2(new_n6740), .A3(new_n6739), .B(\a[5] ), .Y(new_n6743));
  NOR2xp33_ASAP7_75t_L      g06487(.A(new_n6743), .B(new_n6742), .Y(new_n6744));
  NAND3xp33_ASAP7_75t_L     g06488(.A(new_n6732), .B(new_n6737), .C(new_n6744), .Y(new_n6745));
  NOR3xp33_ASAP7_75t_L      g06489(.A(new_n6736), .B(new_n6733), .C(new_n6734), .Y(new_n6746));
  AOI22xp33_ASAP7_75t_L     g06490(.A1(new_n6726), .A2(new_n6730), .B1(new_n6731), .B2(new_n6477), .Y(new_n6747));
  INVx1_ASAP7_75t_L         g06491(.A(new_n6744), .Y(new_n6748));
  OAI21xp33_ASAP7_75t_L     g06492(.A1(new_n6746), .A2(new_n6747), .B(new_n6748), .Y(new_n6749));
  NAND2xp33_ASAP7_75t_L     g06493(.A(new_n6745), .B(new_n6749), .Y(new_n6750));
  NAND3xp33_ASAP7_75t_L     g06494(.A(new_n6477), .B(new_n6242), .C(new_n6478), .Y(new_n6751));
  OAI21xp33_ASAP7_75t_L     g06495(.A1(new_n6483), .A2(new_n6486), .B(new_n6751), .Y(new_n6752));
  XOR2x2_ASAP7_75t_L        g06496(.A(new_n6750), .B(new_n6752), .Y(new_n6753));
  INVx1_ASAP7_75t_L         g06497(.A(new_n6221), .Y(new_n6754));
  NOR2xp33_ASAP7_75t_L      g06498(.A(\b[44] ), .B(\b[45] ), .Y(new_n6755));
  INVx1_ASAP7_75t_L         g06499(.A(\b[45] ), .Y(new_n6756));
  NOR2xp33_ASAP7_75t_L      g06500(.A(new_n6220), .B(new_n6756), .Y(new_n6757));
  NOR2xp33_ASAP7_75t_L      g06501(.A(new_n6755), .B(new_n6757), .Y(new_n6758));
  INVx1_ASAP7_75t_L         g06502(.A(new_n6758), .Y(new_n6759));
  O2A1O1Ixp33_ASAP7_75t_L   g06503(.A1(new_n6227), .A2(new_n6226), .B(new_n6754), .C(new_n6759), .Y(new_n6760));
  A2O1A1O1Ixp25_ASAP7_75t_L g06504(.A1(new_n6197), .A2(new_n6200), .B(new_n6196), .C(new_n6222), .D(new_n6221), .Y(new_n6761));
  NAND2xp33_ASAP7_75t_L     g06505(.A(new_n6759), .B(new_n6761), .Y(new_n6762));
  INVx1_ASAP7_75t_L         g06506(.A(new_n6762), .Y(new_n6763));
  NOR2xp33_ASAP7_75t_L      g06507(.A(new_n6760), .B(new_n6763), .Y(new_n6764));
  AOI22xp33_ASAP7_75t_L     g06508(.A1(new_n272), .A2(\b[45] ), .B1(new_n269), .B2(new_n6764), .Y(new_n6765));
  OAI221xp5_ASAP7_75t_L     g06509(.A1(new_n261), .A2(new_n6220), .B1(new_n6195), .B2(new_n277), .C(new_n6765), .Y(new_n6766));
  XNOR2x2_ASAP7_75t_L       g06510(.A(new_n265), .B(new_n6766), .Y(new_n6767));
  NOR2xp33_ASAP7_75t_L      g06511(.A(new_n6767), .B(new_n6753), .Y(new_n6768));
  INVx1_ASAP7_75t_L         g06512(.A(new_n6768), .Y(new_n6769));
  NAND2xp33_ASAP7_75t_L     g06513(.A(new_n6767), .B(new_n6753), .Y(new_n6770));
  AND2x2_ASAP7_75t_L        g06514(.A(new_n6770), .B(new_n6769), .Y(new_n6771));
  XNOR2x2_ASAP7_75t_L       g06515(.A(new_n6493), .B(new_n6771), .Y(\f[45] ));
  NAND2xp33_ASAP7_75t_L     g06516(.A(\b[42] ), .B(new_n334), .Y(new_n6773));
  AOI22xp33_ASAP7_75t_L     g06517(.A1(new_n345), .A2(\b[43] ), .B1(new_n342), .B2(new_n6202), .Y(new_n6774));
  NAND2xp33_ASAP7_75t_L     g06518(.A(new_n6773), .B(new_n6774), .Y(new_n6775));
  AOI211xp5_ASAP7_75t_L     g06519(.A1(\b[41] ), .A2(new_n366), .B(new_n339), .C(new_n6775), .Y(new_n6776));
  INVx1_ASAP7_75t_L         g06520(.A(new_n6775), .Y(new_n6777));
  O2A1O1Ixp33_ASAP7_75t_L   g06521(.A1(new_n5666), .A2(new_n365), .B(new_n6777), .C(\a[5] ), .Y(new_n6778));
  NOR2xp33_ASAP7_75t_L      g06522(.A(new_n6776), .B(new_n6778), .Y(new_n6779));
  NOR3xp33_ASAP7_75t_L      g06523(.A(new_n6728), .B(new_n6725), .C(new_n6727), .Y(new_n6780));
  O2A1O1Ixp33_ASAP7_75t_L   g06524(.A1(new_n6734), .A2(new_n6733), .B(new_n6736), .C(new_n6780), .Y(new_n6781));
  OAI21xp33_ASAP7_75t_L     g06525(.A1(new_n6686), .A2(new_n6689), .B(new_n6690), .Y(new_n6782));
  NAND2xp33_ASAP7_75t_L     g06526(.A(new_n6665), .B(new_n6661), .Y(new_n6783));
  NOR2xp33_ASAP7_75t_L      g06527(.A(new_n6672), .B(new_n6783), .Y(new_n6784));
  NOR2xp33_ASAP7_75t_L      g06528(.A(new_n2852), .B(new_n1412), .Y(new_n6785));
  INVx1_ASAP7_75t_L         g06529(.A(new_n6785), .Y(new_n6786));
  OAI221xp5_ASAP7_75t_L     g06530(.A1(new_n2650), .A2(new_n1398), .B1(new_n1411), .B2(new_n5212), .C(new_n6786), .Y(new_n6787));
  INVx1_ASAP7_75t_L         g06531(.A(new_n6787), .Y(new_n6788));
  OAI211xp5_ASAP7_75t_L     g06532(.A1(new_n2477), .A2(new_n1549), .B(new_n6788), .C(\a[20] ), .Y(new_n6789));
  A2O1A1Ixp33_ASAP7_75t_L   g06533(.A1(\b[26] ), .A2(new_n1548), .B(new_n6787), .C(new_n1401), .Y(new_n6790));
  AND2x2_ASAP7_75t_L        g06534(.A(new_n6790), .B(new_n6789), .Y(new_n6791));
  NOR2xp33_ASAP7_75t_L      g06535(.A(new_n6592), .B(new_n6594), .Y(new_n6792));
  NAND2xp33_ASAP7_75t_L     g06536(.A(\b[11] ), .B(new_n4111), .Y(new_n6793));
  NAND2xp33_ASAP7_75t_L     g06537(.A(\b[12] ), .B(new_n3874), .Y(new_n6794));
  AOI22xp33_ASAP7_75t_L     g06538(.A1(new_n3884), .A2(\b[13] ), .B1(new_n3881), .B2(new_n800), .Y(new_n6795));
  AND4x1_ASAP7_75t_L        g06539(.A(new_n6795), .B(new_n6794), .C(new_n6793), .D(\a[35] ), .Y(new_n6796));
  AOI31xp33_ASAP7_75t_L     g06540(.A1(new_n6795), .A2(new_n6794), .A3(new_n6793), .B(\a[35] ), .Y(new_n6797));
  NOR2xp33_ASAP7_75t_L      g06541(.A(new_n6797), .B(new_n6796), .Y(new_n6798));
  INVx1_ASAP7_75t_L         g06542(.A(new_n6798), .Y(new_n6799));
  A2O1A1O1Ixp25_ASAP7_75t_L g06543(.A1(new_n6344), .A2(new_n6354), .B(new_n6535), .C(new_n6586), .D(new_n6582), .Y(new_n6800));
  INVx1_ASAP7_75t_L         g06544(.A(new_n6541), .Y(new_n6801));
  NOR3xp33_ASAP7_75t_L      g06545(.A(new_n6324), .B(new_n6801), .C(new_n6536), .Y(new_n6802));
  NOR2xp33_ASAP7_75t_L      g06546(.A(new_n278), .B(new_n6309), .Y(new_n6803));
  NOR2xp33_ASAP7_75t_L      g06547(.A(new_n299), .B(new_n6544), .Y(new_n6804));
  OAI32xp33_ASAP7_75t_L     g06548(.A1(new_n325), .A2(new_n327), .A3(new_n6311), .B1(new_n6312), .B2(new_n323), .Y(new_n6805));
  NOR4xp25_ASAP7_75t_L      g06549(.A(new_n6805), .B(new_n5996), .C(new_n6803), .D(new_n6804), .Y(new_n6806));
  INVx1_ASAP7_75t_L         g06550(.A(new_n6806), .Y(new_n6807));
  OAI31xp33_ASAP7_75t_L     g06551(.A1(new_n6805), .A2(new_n6804), .A3(new_n6803), .B(new_n5996), .Y(new_n6808));
  NAND2xp33_ASAP7_75t_L     g06552(.A(\a[47] ), .B(new_n6541), .Y(new_n6809));
  NAND2xp33_ASAP7_75t_L     g06553(.A(new_n6539), .B(new_n6538), .Y(new_n6810));
  XNOR2x2_ASAP7_75t_L       g06554(.A(\a[46] ), .B(\a[45] ), .Y(new_n6811));
  NOR2xp33_ASAP7_75t_L      g06555(.A(new_n6811), .B(new_n6810), .Y(new_n6812));
  NAND2xp33_ASAP7_75t_L     g06556(.A(\b[0] ), .B(new_n6812), .Y(new_n6813));
  INVx1_ASAP7_75t_L         g06557(.A(\a[46] ), .Y(new_n6814));
  NAND2xp33_ASAP7_75t_L     g06558(.A(\a[47] ), .B(new_n6814), .Y(new_n6815));
  INVx1_ASAP7_75t_L         g06559(.A(\a[47] ), .Y(new_n6816));
  NAND2xp33_ASAP7_75t_L     g06560(.A(\a[46] ), .B(new_n6816), .Y(new_n6817));
  AND2x2_ASAP7_75t_L        g06561(.A(new_n6815), .B(new_n6817), .Y(new_n6818));
  NOR2xp33_ASAP7_75t_L      g06562(.A(new_n6540), .B(new_n6818), .Y(new_n6819));
  NAND2xp33_ASAP7_75t_L     g06563(.A(new_n271), .B(new_n6819), .Y(new_n6820));
  NAND2xp33_ASAP7_75t_L     g06564(.A(new_n6817), .B(new_n6815), .Y(new_n6821));
  NOR2xp33_ASAP7_75t_L      g06565(.A(new_n6821), .B(new_n6540), .Y(new_n6822));
  NAND2xp33_ASAP7_75t_L     g06566(.A(\b[1] ), .B(new_n6822), .Y(new_n6823));
  NAND3xp33_ASAP7_75t_L     g06567(.A(new_n6820), .B(new_n6823), .C(new_n6813), .Y(new_n6824));
  XOR2x2_ASAP7_75t_L        g06568(.A(new_n6809), .B(new_n6824), .Y(new_n6825));
  NAND3xp33_ASAP7_75t_L     g06569(.A(new_n6807), .B(new_n6825), .C(new_n6808), .Y(new_n6826));
  INVx1_ASAP7_75t_L         g06570(.A(new_n6808), .Y(new_n6827));
  XNOR2x2_ASAP7_75t_L       g06571(.A(new_n6809), .B(new_n6824), .Y(new_n6828));
  OAI21xp33_ASAP7_75t_L     g06572(.A1(new_n6806), .A2(new_n6827), .B(new_n6828), .Y(new_n6829));
  OAI211xp5_ASAP7_75t_L     g06573(.A1(new_n6802), .A2(new_n6549), .B(new_n6826), .C(new_n6829), .Y(new_n6830));
  NOR2xp33_ASAP7_75t_L      g06574(.A(new_n6536), .B(new_n6324), .Y(new_n6831));
  NAND2xp33_ASAP7_75t_L     g06575(.A(new_n6548), .B(new_n6547), .Y(new_n6832));
  MAJIxp5_ASAP7_75t_L       g06576(.A(new_n6832), .B(new_n6541), .C(new_n6831), .Y(new_n6833));
  NOR3xp33_ASAP7_75t_L      g06577(.A(new_n6827), .B(new_n6828), .C(new_n6806), .Y(new_n6834));
  AOI21xp33_ASAP7_75t_L     g06578(.A1(new_n6807), .A2(new_n6808), .B(new_n6825), .Y(new_n6835));
  OAI21xp33_ASAP7_75t_L     g06579(.A1(new_n6834), .A2(new_n6835), .B(new_n6833), .Y(new_n6836));
  NAND2xp33_ASAP7_75t_L     g06580(.A(\b[6] ), .B(new_n5240), .Y(new_n6837));
  AOI32xp33_ASAP7_75t_L     g06581(.A1(new_n424), .A2(new_n426), .A3(new_n5247), .B1(new_n5249), .B2(\b[7] ), .Y(new_n6838));
  OAI211xp5_ASAP7_75t_L     g06582(.A1(new_n353), .A2(new_n5521), .B(new_n6838), .C(new_n6837), .Y(new_n6839));
  NOR2xp33_ASAP7_75t_L      g06583(.A(new_n5244), .B(new_n6839), .Y(new_n6840));
  INVx1_ASAP7_75t_L         g06584(.A(new_n6840), .Y(new_n6841));
  NAND2xp33_ASAP7_75t_L     g06585(.A(new_n5244), .B(new_n6839), .Y(new_n6842));
  NAND4xp25_ASAP7_75t_L     g06586(.A(new_n6841), .B(new_n6830), .C(new_n6836), .D(new_n6842), .Y(new_n6843));
  NOR3xp33_ASAP7_75t_L      g06587(.A(new_n6833), .B(new_n6834), .C(new_n6835), .Y(new_n6844));
  AOI211xp5_ASAP7_75t_L     g06588(.A1(new_n6829), .A2(new_n6826), .B(new_n6549), .C(new_n6802), .Y(new_n6845));
  INVx1_ASAP7_75t_L         g06589(.A(new_n6842), .Y(new_n6846));
  OAI22xp33_ASAP7_75t_L     g06590(.A1(new_n6844), .A2(new_n6845), .B1(new_n6846), .B2(new_n6840), .Y(new_n6847));
  NAND2xp33_ASAP7_75t_L     g06591(.A(new_n6843), .B(new_n6847), .Y(new_n6848));
  AOI211xp5_ASAP7_75t_L     g06592(.A1(new_n6560), .A2(new_n6555), .B(new_n6549), .C(new_n6550), .Y(new_n6849));
  INVx1_ASAP7_75t_L         g06593(.A(new_n6849), .Y(new_n6850));
  A2O1A1Ixp33_ASAP7_75t_L   g06594(.A1(new_n6330), .A2(new_n6565), .B(new_n6562), .C(new_n6850), .Y(new_n6851));
  NOR2xp33_ASAP7_75t_L      g06595(.A(new_n6848), .B(new_n6851), .Y(new_n6852));
  O2A1O1Ixp33_ASAP7_75t_L   g06596(.A1(new_n6557), .A2(new_n6561), .B(new_n6578), .C(new_n6849), .Y(new_n6853));
  AOI21xp33_ASAP7_75t_L     g06597(.A1(new_n6847), .A2(new_n6843), .B(new_n6853), .Y(new_n6854));
  NOR2xp33_ASAP7_75t_L      g06598(.A(new_n503), .B(new_n4781), .Y(new_n6855));
  INVx1_ASAP7_75t_L         g06599(.A(new_n6855), .Y(new_n6856));
  NAND2xp33_ASAP7_75t_L     g06600(.A(\b[9] ), .B(new_n4548), .Y(new_n6857));
  AOI22xp33_ASAP7_75t_L     g06601(.A1(new_n4544), .A2(\b[10] ), .B1(new_n4542), .B2(new_n852), .Y(new_n6858));
  NAND4xp25_ASAP7_75t_L     g06602(.A(new_n6858), .B(\a[38] ), .C(new_n6856), .D(new_n6857), .Y(new_n6859));
  AOI31xp33_ASAP7_75t_L     g06603(.A1(new_n6858), .A2(new_n6857), .A3(new_n6856), .B(\a[38] ), .Y(new_n6860));
  INVx1_ASAP7_75t_L         g06604(.A(new_n6860), .Y(new_n6861));
  OAI211xp5_ASAP7_75t_L     g06605(.A1(new_n6854), .A2(new_n6852), .B(new_n6859), .C(new_n6861), .Y(new_n6862));
  NAND3xp33_ASAP7_75t_L     g06606(.A(new_n6853), .B(new_n6847), .C(new_n6843), .Y(new_n6863));
  A2O1A1Ixp33_ASAP7_75t_L   g06607(.A1(new_n6569), .A2(new_n6578), .B(new_n6849), .C(new_n6848), .Y(new_n6864));
  NAND2xp33_ASAP7_75t_L     g06608(.A(new_n6859), .B(new_n6861), .Y(new_n6865));
  NAND3xp33_ASAP7_75t_L     g06609(.A(new_n6865), .B(new_n6863), .C(new_n6864), .Y(new_n6866));
  AND3x1_ASAP7_75t_L        g06610(.A(new_n6800), .B(new_n6866), .C(new_n6862), .Y(new_n6867));
  AOI21xp33_ASAP7_75t_L     g06611(.A1(new_n6866), .A2(new_n6862), .B(new_n6800), .Y(new_n6868));
  NOR3xp33_ASAP7_75t_L      g06612(.A(new_n6799), .B(new_n6867), .C(new_n6868), .Y(new_n6869));
  NAND3xp33_ASAP7_75t_L     g06613(.A(new_n6800), .B(new_n6866), .C(new_n6862), .Y(new_n6870));
  AO21x2_ASAP7_75t_L        g06614(.A1(new_n6866), .A2(new_n6862), .B(new_n6800), .Y(new_n6871));
  AOI21xp33_ASAP7_75t_L     g06615(.A1(new_n6871), .A2(new_n6870), .B(new_n6798), .Y(new_n6872));
  NOR2xp33_ASAP7_75t_L      g06616(.A(new_n6872), .B(new_n6869), .Y(new_n6873));
  A2O1A1Ixp33_ASAP7_75t_L   g06617(.A1(new_n6792), .A2(new_n6591), .B(new_n6603), .C(new_n6873), .Y(new_n6874));
  NAND2xp33_ASAP7_75t_L     g06618(.A(new_n6589), .B(new_n6584), .Y(new_n6875));
  NOR2xp33_ASAP7_75t_L      g06619(.A(new_n6533), .B(new_n6875), .Y(new_n6876));
  O2A1O1Ixp33_ASAP7_75t_L   g06620(.A1(new_n6590), .A2(new_n6595), .B(new_n6525), .C(new_n6876), .Y(new_n6877));
  NAND3xp33_ASAP7_75t_L     g06621(.A(new_n6871), .B(new_n6870), .C(new_n6798), .Y(new_n6878));
  OAI21xp33_ASAP7_75t_L     g06622(.A1(new_n6868), .A2(new_n6867), .B(new_n6799), .Y(new_n6879));
  NAND2xp33_ASAP7_75t_L     g06623(.A(new_n6878), .B(new_n6879), .Y(new_n6880));
  NAND2xp33_ASAP7_75t_L     g06624(.A(new_n6880), .B(new_n6877), .Y(new_n6881));
  NAND2xp33_ASAP7_75t_L     g06625(.A(\b[14] ), .B(new_n3491), .Y(new_n6882));
  NAND2xp33_ASAP7_75t_L     g06626(.A(\b[15] ), .B(new_n3260), .Y(new_n6883));
  AOI22xp33_ASAP7_75t_L     g06627(.A1(new_n3256), .A2(\b[16] ), .B1(new_n3254), .B2(new_n1058), .Y(new_n6884));
  NAND4xp25_ASAP7_75t_L     g06628(.A(new_n6884), .B(\a[32] ), .C(new_n6882), .D(new_n6883), .Y(new_n6885));
  NAND2xp33_ASAP7_75t_L     g06629(.A(new_n6883), .B(new_n6884), .Y(new_n6886));
  A2O1A1Ixp33_ASAP7_75t_L   g06630(.A1(\b[14] ), .A2(new_n3491), .B(new_n6886), .C(new_n3251), .Y(new_n6887));
  NAND2xp33_ASAP7_75t_L     g06631(.A(new_n6885), .B(new_n6887), .Y(new_n6888));
  INVx1_ASAP7_75t_L         g06632(.A(new_n6888), .Y(new_n6889));
  NAND3xp33_ASAP7_75t_L     g06633(.A(new_n6889), .B(new_n6881), .C(new_n6874), .Y(new_n6890));
  O2A1O1Ixp33_ASAP7_75t_L   g06634(.A1(new_n6533), .A2(new_n6875), .B(new_n6596), .C(new_n6880), .Y(new_n6891));
  MAJIxp5_ASAP7_75t_L       g06635(.A(new_n6597), .B(new_n6533), .C(new_n6875), .Y(new_n6892));
  NOR2xp33_ASAP7_75t_L      g06636(.A(new_n6892), .B(new_n6873), .Y(new_n6893));
  OAI21xp33_ASAP7_75t_L     g06637(.A1(new_n6891), .A2(new_n6893), .B(new_n6888), .Y(new_n6894));
  NAND3xp33_ASAP7_75t_L     g06638(.A(new_n6602), .B(new_n6596), .C(new_n6600), .Y(new_n6895));
  OAI21xp33_ASAP7_75t_L     g06639(.A1(new_n6610), .A2(new_n6611), .B(new_n6516), .Y(new_n6896));
  NAND4xp25_ASAP7_75t_L     g06640(.A(new_n6896), .B(new_n6890), .C(new_n6894), .D(new_n6895), .Y(new_n6897));
  NOR3xp33_ASAP7_75t_L      g06641(.A(new_n6893), .B(new_n6891), .C(new_n6888), .Y(new_n6898));
  AOI21xp33_ASAP7_75t_L     g06642(.A1(new_n6874), .A2(new_n6881), .B(new_n6889), .Y(new_n6899));
  NAND2xp33_ASAP7_75t_L     g06643(.A(new_n6596), .B(new_n6600), .Y(new_n6900));
  MAJIxp5_ASAP7_75t_L       g06644(.A(new_n6609), .B(new_n6524), .C(new_n6900), .Y(new_n6901));
  OAI21xp33_ASAP7_75t_L     g06645(.A1(new_n6898), .A2(new_n6899), .B(new_n6901), .Y(new_n6902));
  NOR2xp33_ASAP7_75t_L      g06646(.A(new_n1244), .B(new_n2932), .Y(new_n6903));
  NAND2xp33_ASAP7_75t_L     g06647(.A(\b[18] ), .B(new_n2706), .Y(new_n6904));
  OAI221xp5_ASAP7_75t_L     g06648(.A1(new_n2708), .A2(new_n1493), .B1(new_n2707), .B2(new_n2793), .C(new_n6904), .Y(new_n6905));
  OR3x1_ASAP7_75t_L         g06649(.A(new_n6905), .B(new_n2697), .C(new_n6903), .Y(new_n6906));
  A2O1A1Ixp33_ASAP7_75t_L   g06650(.A1(\b[17] ), .A2(new_n2931), .B(new_n6905), .C(new_n2697), .Y(new_n6907));
  NAND4xp25_ASAP7_75t_L     g06651(.A(new_n6897), .B(new_n6902), .C(new_n6907), .D(new_n6906), .Y(new_n6908));
  NOR3xp33_ASAP7_75t_L      g06652(.A(new_n6899), .B(new_n6901), .C(new_n6898), .Y(new_n6909));
  AOI22xp33_ASAP7_75t_L     g06653(.A1(new_n6890), .A2(new_n6894), .B1(new_n6895), .B2(new_n6896), .Y(new_n6910));
  NAND2xp33_ASAP7_75t_L     g06654(.A(new_n6907), .B(new_n6906), .Y(new_n6911));
  OAI21xp33_ASAP7_75t_L     g06655(.A1(new_n6909), .A2(new_n6910), .B(new_n6911), .Y(new_n6912));
  A2O1A1O1Ixp25_ASAP7_75t_L g06656(.A1(new_n6373), .A2(new_n6275), .B(new_n6382), .C(new_n6620), .D(new_n6624), .Y(new_n6913));
  NAND3xp33_ASAP7_75t_L     g06657(.A(new_n6913), .B(new_n6912), .C(new_n6908), .Y(new_n6914));
  AO21x2_ASAP7_75t_L        g06658(.A1(new_n6908), .A2(new_n6912), .B(new_n6913), .Y(new_n6915));
  NAND2xp33_ASAP7_75t_L     g06659(.A(\b[20] ), .B(new_n2386), .Y(new_n6916));
  NAND2xp33_ASAP7_75t_L     g06660(.A(\b[21] ), .B(new_n2232), .Y(new_n6917));
  AOI32xp33_ASAP7_75t_L     g06661(.A1(new_n1862), .A2(new_n1860), .A3(new_n2226), .B1(\b[22] ), .B2(new_n2228), .Y(new_n6918));
  NAND4xp25_ASAP7_75t_L     g06662(.A(new_n6918), .B(\a[26] ), .C(new_n6916), .D(new_n6917), .Y(new_n6919));
  NAND2xp33_ASAP7_75t_L     g06663(.A(new_n6917), .B(new_n6918), .Y(new_n6920));
  A2O1A1Ixp33_ASAP7_75t_L   g06664(.A1(\b[20] ), .A2(new_n2386), .B(new_n6920), .C(new_n2223), .Y(new_n6921));
  AND2x2_ASAP7_75t_L        g06665(.A(new_n6919), .B(new_n6921), .Y(new_n6922));
  NAND3xp33_ASAP7_75t_L     g06666(.A(new_n6915), .B(new_n6922), .C(new_n6914), .Y(new_n6923));
  AND3x1_ASAP7_75t_L        g06667(.A(new_n6913), .B(new_n6912), .C(new_n6908), .Y(new_n6924));
  AOI21xp33_ASAP7_75t_L     g06668(.A1(new_n6912), .A2(new_n6908), .B(new_n6913), .Y(new_n6925));
  NAND2xp33_ASAP7_75t_L     g06669(.A(new_n6919), .B(new_n6921), .Y(new_n6926));
  OAI21xp33_ASAP7_75t_L     g06670(.A1(new_n6925), .A2(new_n6924), .B(new_n6926), .Y(new_n6927));
  NAND2xp33_ASAP7_75t_L     g06671(.A(new_n6923), .B(new_n6927), .Y(new_n6928));
  NAND2xp33_ASAP7_75t_L     g06672(.A(new_n6626), .B(new_n6621), .Y(new_n6929));
  MAJIxp5_ASAP7_75t_L       g06673(.A(new_n6643), .B(new_n6929), .C(new_n6632), .Y(new_n6930));
  NOR2xp33_ASAP7_75t_L      g06674(.A(new_n6928), .B(new_n6930), .Y(new_n6931));
  NOR3xp33_ASAP7_75t_L      g06675(.A(new_n6924), .B(new_n6925), .C(new_n6926), .Y(new_n6932));
  AOI21xp33_ASAP7_75t_L     g06676(.A1(new_n6915), .A2(new_n6914), .B(new_n6922), .Y(new_n6933));
  NOR2xp33_ASAP7_75t_L      g06677(.A(new_n6933), .B(new_n6932), .Y(new_n6934));
  NOR2xp33_ASAP7_75t_L      g06678(.A(new_n6632), .B(new_n6929), .Y(new_n6935));
  INVx1_ASAP7_75t_L         g06679(.A(new_n6935), .Y(new_n6936));
  AOI21xp33_ASAP7_75t_L     g06680(.A1(new_n6657), .A2(new_n6936), .B(new_n6934), .Y(new_n6937));
  NOR2xp33_ASAP7_75t_L      g06681(.A(new_n1995), .B(new_n1911), .Y(new_n6938));
  NAND2xp33_ASAP7_75t_L     g06682(.A(\b[24] ), .B(new_n1770), .Y(new_n6939));
  OAI221xp5_ASAP7_75t_L     g06683(.A1(new_n1772), .A2(new_n2180), .B1(new_n1771), .B2(new_n2187), .C(new_n6939), .Y(new_n6940));
  OR3x1_ASAP7_75t_L         g06684(.A(new_n6940), .B(new_n1761), .C(new_n6938), .Y(new_n6941));
  A2O1A1Ixp33_ASAP7_75t_L   g06685(.A1(\b[23] ), .A2(new_n1910), .B(new_n6940), .C(new_n1761), .Y(new_n6942));
  NAND2xp33_ASAP7_75t_L     g06686(.A(new_n6942), .B(new_n6941), .Y(new_n6943));
  NOR3xp33_ASAP7_75t_L      g06687(.A(new_n6931), .B(new_n6937), .C(new_n6943), .Y(new_n6944));
  AOI21xp33_ASAP7_75t_L     g06688(.A1(new_n6641), .A2(new_n6638), .B(new_n6935), .Y(new_n6945));
  NAND2xp33_ASAP7_75t_L     g06689(.A(new_n6934), .B(new_n6945), .Y(new_n6946));
  A2O1A1Ixp33_ASAP7_75t_L   g06690(.A1(new_n6638), .A2(new_n6641), .B(new_n6935), .C(new_n6928), .Y(new_n6947));
  AND2x2_ASAP7_75t_L        g06691(.A(new_n6942), .B(new_n6941), .Y(new_n6948));
  AOI21xp33_ASAP7_75t_L     g06692(.A1(new_n6946), .A2(new_n6947), .B(new_n6948), .Y(new_n6949));
  A2O1A1Ixp33_ASAP7_75t_L   g06693(.A1(new_n6114), .A2(new_n6113), .B(new_n6271), .C(new_n6408), .Y(new_n6950));
  A2O1A1Ixp33_ASAP7_75t_L   g06694(.A1(new_n6950), .A2(new_n6409), .B(new_n6662), .C(new_n6659), .Y(new_n6951));
  OAI21xp33_ASAP7_75t_L     g06695(.A1(new_n6949), .A2(new_n6944), .B(new_n6951), .Y(new_n6952));
  NAND3xp33_ASAP7_75t_L     g06696(.A(new_n6946), .B(new_n6947), .C(new_n6948), .Y(new_n6953));
  OAI21xp33_ASAP7_75t_L     g06697(.A1(new_n6937), .A2(new_n6931), .B(new_n6943), .Y(new_n6954));
  A2O1A1O1Ixp25_ASAP7_75t_L g06698(.A1(new_n6408), .A2(new_n6273), .B(new_n6414), .C(new_n6652), .D(new_n6663), .Y(new_n6955));
  NAND3xp33_ASAP7_75t_L     g06699(.A(new_n6955), .B(new_n6954), .C(new_n6953), .Y(new_n6956));
  AOI21xp33_ASAP7_75t_L     g06700(.A1(new_n6956), .A2(new_n6952), .B(new_n6791), .Y(new_n6957));
  NAND2xp33_ASAP7_75t_L     g06701(.A(new_n6790), .B(new_n6789), .Y(new_n6958));
  AOI21xp33_ASAP7_75t_L     g06702(.A1(new_n6954), .A2(new_n6953), .B(new_n6955), .Y(new_n6959));
  NOR3xp33_ASAP7_75t_L      g06703(.A(new_n6951), .B(new_n6949), .C(new_n6944), .Y(new_n6960));
  NOR3xp33_ASAP7_75t_L      g06704(.A(new_n6959), .B(new_n6960), .C(new_n6958), .Y(new_n6961));
  NOR2xp33_ASAP7_75t_L      g06705(.A(new_n6961), .B(new_n6957), .Y(new_n6962));
  A2O1A1Ixp33_ASAP7_75t_L   g06706(.A1(new_n6680), .A2(new_n6679), .B(new_n6784), .C(new_n6962), .Y(new_n6963));
  AOI21xp33_ASAP7_75t_L     g06707(.A1(new_n6679), .A2(new_n6680), .B(new_n6784), .Y(new_n6964));
  OAI21xp33_ASAP7_75t_L     g06708(.A1(new_n6960), .A2(new_n6959), .B(new_n6958), .Y(new_n6965));
  NAND3xp33_ASAP7_75t_L     g06709(.A(new_n6956), .B(new_n6791), .C(new_n6952), .Y(new_n6966));
  NAND2xp33_ASAP7_75t_L     g06710(.A(new_n6965), .B(new_n6966), .Y(new_n6967));
  NAND2xp33_ASAP7_75t_L     g06711(.A(new_n6967), .B(new_n6964), .Y(new_n6968));
  AOI22xp33_ASAP7_75t_L     g06712(.A1(new_n1113), .A2(\b[31] ), .B1(new_n1110), .B2(new_n3426), .Y(new_n6969));
  OAI221xp5_ASAP7_75t_L     g06713(.A1(new_n1298), .A2(new_n3212), .B1(new_n2871), .B2(new_n1195), .C(new_n6969), .Y(new_n6970));
  XNOR2x2_ASAP7_75t_L       g06714(.A(\a[17] ), .B(new_n6970), .Y(new_n6971));
  NAND3xp33_ASAP7_75t_L     g06715(.A(new_n6963), .B(new_n6968), .C(new_n6971), .Y(new_n6972));
  O2A1O1Ixp33_ASAP7_75t_L   g06716(.A1(new_n6783), .A2(new_n6672), .B(new_n6684), .C(new_n6967), .Y(new_n6973));
  MAJIxp5_ASAP7_75t_L       g06717(.A(new_n6511), .B(new_n6783), .C(new_n6672), .Y(new_n6974));
  NOR2xp33_ASAP7_75t_L      g06718(.A(new_n6974), .B(new_n6962), .Y(new_n6975));
  XNOR2x2_ASAP7_75t_L       g06719(.A(new_n1107), .B(new_n6970), .Y(new_n6976));
  OAI21xp33_ASAP7_75t_L     g06720(.A1(new_n6975), .A2(new_n6973), .B(new_n6976), .Y(new_n6977));
  NAND3xp33_ASAP7_75t_L     g06721(.A(new_n6782), .B(new_n6972), .C(new_n6977), .Y(new_n6978));
  A2O1A1O1Ixp25_ASAP7_75t_L g06722(.A1(new_n6428), .A2(new_n6435), .B(new_n6503), .C(new_n6691), .D(new_n6682), .Y(new_n6979));
  NOR3xp33_ASAP7_75t_L      g06723(.A(new_n6973), .B(new_n6975), .C(new_n6976), .Y(new_n6980));
  AOI21xp33_ASAP7_75t_L     g06724(.A1(new_n6963), .A2(new_n6968), .B(new_n6971), .Y(new_n6981));
  OAI21xp33_ASAP7_75t_L     g06725(.A1(new_n6980), .A2(new_n6981), .B(new_n6979), .Y(new_n6982));
  NAND2xp33_ASAP7_75t_L     g06726(.A(\b[33] ), .B(new_n817), .Y(new_n6983));
  AOI22xp33_ASAP7_75t_L     g06727(.A1(new_n826), .A2(\b[34] ), .B1(new_n823), .B2(new_n3833), .Y(new_n6984));
  NAND2xp33_ASAP7_75t_L     g06728(.A(new_n6983), .B(new_n6984), .Y(new_n6985));
  AOI211xp5_ASAP7_75t_L     g06729(.A1(\b[32] ), .A2(new_n908), .B(new_n813), .C(new_n6985), .Y(new_n6986));
  INVx1_ASAP7_75t_L         g06730(.A(new_n6985), .Y(new_n6987));
  O2A1O1Ixp33_ASAP7_75t_L   g06731(.A1(new_n3443), .A2(new_n909), .B(new_n6987), .C(\a[14] ), .Y(new_n6988));
  NOR2xp33_ASAP7_75t_L      g06732(.A(new_n6986), .B(new_n6988), .Y(new_n6989));
  NAND3xp33_ASAP7_75t_L     g06733(.A(new_n6989), .B(new_n6978), .C(new_n6982), .Y(new_n6990));
  AOI21xp33_ASAP7_75t_L     g06734(.A1(new_n6982), .A2(new_n6978), .B(new_n6989), .Y(new_n6991));
  INVx1_ASAP7_75t_L         g06735(.A(new_n6991), .Y(new_n6992));
  MAJIxp5_ASAP7_75t_L       g06736(.A(new_n6502), .B(new_n6705), .C(new_n6700), .Y(new_n6993));
  NAND3xp33_ASAP7_75t_L     g06737(.A(new_n6993), .B(new_n6992), .C(new_n6990), .Y(new_n6994));
  AND3x1_ASAP7_75t_L        g06738(.A(new_n6989), .B(new_n6982), .C(new_n6978), .Y(new_n6995));
  MAJIxp5_ASAP7_75t_L       g06739(.A(new_n6704), .B(new_n6707), .C(new_n6701), .Y(new_n6996));
  OAI21xp33_ASAP7_75t_L     g06740(.A1(new_n6995), .A2(new_n6991), .B(new_n6996), .Y(new_n6997));
  NOR2xp33_ASAP7_75t_L      g06741(.A(new_n4701), .B(new_n676), .Y(new_n6998));
  AOI221xp5_ASAP7_75t_L     g06742(.A1(new_n590), .A2(\b[36] ), .B1(new_n597), .B2(new_n4709), .C(new_n6998), .Y(new_n6999));
  OA211x2_ASAP7_75t_L       g06743(.A1(new_n1620), .A2(new_n4053), .B(new_n6999), .C(\a[11] ), .Y(new_n7000));
  O2A1O1Ixp33_ASAP7_75t_L   g06744(.A1(new_n4053), .A2(new_n1620), .B(new_n6999), .C(\a[11] ), .Y(new_n7001));
  NOR2xp33_ASAP7_75t_L      g06745(.A(new_n7001), .B(new_n7000), .Y(new_n7002));
  NAND3xp33_ASAP7_75t_L     g06746(.A(new_n6994), .B(new_n6997), .C(new_n7002), .Y(new_n7003));
  NAND2xp33_ASAP7_75t_L     g06747(.A(new_n6997), .B(new_n6994), .Y(new_n7004));
  OAI21xp33_ASAP7_75t_L     g06748(.A1(new_n7000), .A2(new_n7001), .B(new_n7004), .Y(new_n7005));
  NOR3xp33_ASAP7_75t_L      g06749(.A(new_n6712), .B(new_n6713), .C(new_n6711), .Y(new_n7006));
  A2O1A1O1Ixp25_ASAP7_75t_L g06750(.A1(new_n6465), .A2(new_n6463), .B(new_n6495), .C(new_n6714), .D(new_n7006), .Y(new_n7007));
  AND3x1_ASAP7_75t_L        g06751(.A(new_n7005), .B(new_n7007), .C(new_n7003), .Y(new_n7008));
  AOI21xp33_ASAP7_75t_L     g06752(.A1(new_n7005), .A2(new_n7003), .B(new_n7007), .Y(new_n7009));
  NAND2xp33_ASAP7_75t_L     g06753(.A(\b[38] ), .B(new_n480), .Y(new_n7010));
  NAND2xp33_ASAP7_75t_L     g06754(.A(\b[39] ), .B(new_n441), .Y(new_n7011));
  AOI22xp33_ASAP7_75t_L     g06755(.A1(new_n451), .A2(\b[40] ), .B1(new_n448), .B2(new_n5194), .Y(new_n7012));
  AND4x1_ASAP7_75t_L        g06756(.A(new_n7012), .B(new_n7011), .C(new_n7010), .D(\a[8] ), .Y(new_n7013));
  AOI31xp33_ASAP7_75t_L     g06757(.A1(new_n7012), .A2(new_n7011), .A3(new_n7010), .B(\a[8] ), .Y(new_n7014));
  NOR2xp33_ASAP7_75t_L      g06758(.A(new_n7014), .B(new_n7013), .Y(new_n7015));
  NOR3xp33_ASAP7_75t_L      g06759(.A(new_n7008), .B(new_n7009), .C(new_n7015), .Y(new_n7016));
  NAND3xp33_ASAP7_75t_L     g06760(.A(new_n7005), .B(new_n7003), .C(new_n7007), .Y(new_n7017));
  AO21x2_ASAP7_75t_L        g06761(.A1(new_n7003), .A2(new_n7005), .B(new_n7007), .Y(new_n7018));
  INVx1_ASAP7_75t_L         g06762(.A(new_n7015), .Y(new_n7019));
  AOI21xp33_ASAP7_75t_L     g06763(.A1(new_n7018), .A2(new_n7017), .B(new_n7019), .Y(new_n7020));
  OAI21xp33_ASAP7_75t_L     g06764(.A1(new_n7016), .A2(new_n7020), .B(new_n6781), .Y(new_n7021));
  NAND2xp33_ASAP7_75t_L     g06765(.A(new_n6726), .B(new_n6730), .Y(new_n7022));
  NOR2xp33_ASAP7_75t_L      g06766(.A(new_n7020), .B(new_n7016), .Y(new_n7023));
  A2O1A1Ixp33_ASAP7_75t_L   g06767(.A1(new_n6736), .A2(new_n7022), .B(new_n6780), .C(new_n7023), .Y(new_n7024));
  NAND3xp33_ASAP7_75t_L     g06768(.A(new_n7024), .B(new_n7021), .C(new_n6779), .Y(new_n7025));
  AO21x2_ASAP7_75t_L        g06769(.A1(new_n7021), .A2(new_n7024), .B(new_n6779), .Y(new_n7026));
  NOR3xp33_ASAP7_75t_L      g06770(.A(new_n6747), .B(new_n6744), .C(new_n6746), .Y(new_n7027));
  AOI21xp33_ASAP7_75t_L     g06771(.A1(new_n6752), .A2(new_n6750), .B(new_n7027), .Y(new_n7028));
  AND3x1_ASAP7_75t_L        g06772(.A(new_n7028), .B(new_n7026), .C(new_n7025), .Y(new_n7029));
  AOI21xp33_ASAP7_75t_L     g06773(.A1(new_n7026), .A2(new_n7025), .B(new_n7028), .Y(new_n7030));
  NOR2xp33_ASAP7_75t_L      g06774(.A(new_n7030), .B(new_n7029), .Y(new_n7031));
  NOR2xp33_ASAP7_75t_L      g06775(.A(\b[45] ), .B(\b[46] ), .Y(new_n7032));
  INVx1_ASAP7_75t_L         g06776(.A(\b[46] ), .Y(new_n7033));
  NOR2xp33_ASAP7_75t_L      g06777(.A(new_n6756), .B(new_n7033), .Y(new_n7034));
  NOR2xp33_ASAP7_75t_L      g06778(.A(new_n7032), .B(new_n7034), .Y(new_n7035));
  A2O1A1Ixp33_ASAP7_75t_L   g06779(.A1(\b[45] ), .A2(\b[44] ), .B(new_n6760), .C(new_n7035), .Y(new_n7036));
  INVx1_ASAP7_75t_L         g06780(.A(new_n7036), .Y(new_n7037));
  INVx1_ASAP7_75t_L         g06781(.A(new_n6757), .Y(new_n7038));
  A2O1A1Ixp33_ASAP7_75t_L   g06782(.A1(new_n6223), .A2(new_n6754), .B(new_n6755), .C(new_n7038), .Y(new_n7039));
  NOR2xp33_ASAP7_75t_L      g06783(.A(new_n7035), .B(new_n7039), .Y(new_n7040));
  NOR2xp33_ASAP7_75t_L      g06784(.A(new_n7037), .B(new_n7040), .Y(new_n7041));
  AOI22xp33_ASAP7_75t_L     g06785(.A1(new_n272), .A2(\b[46] ), .B1(new_n269), .B2(new_n7041), .Y(new_n7042));
  OAI221xp5_ASAP7_75t_L     g06786(.A1(new_n261), .A2(new_n6756), .B1(new_n6220), .B2(new_n277), .C(new_n7042), .Y(new_n7043));
  XNOR2x2_ASAP7_75t_L       g06787(.A(new_n265), .B(new_n7043), .Y(new_n7044));
  XNOR2x2_ASAP7_75t_L       g06788(.A(new_n7044), .B(new_n7031), .Y(new_n7045));
  O2A1O1Ixp33_ASAP7_75t_L   g06789(.A1(new_n6493), .A2(new_n6768), .B(new_n6770), .C(new_n7045), .Y(new_n7046));
  INVx1_ASAP7_75t_L         g06790(.A(new_n7045), .Y(new_n7047));
  OAI21xp33_ASAP7_75t_L     g06791(.A1(new_n6768), .A2(new_n6493), .B(new_n6770), .Y(new_n7048));
  NOR2xp33_ASAP7_75t_L      g06792(.A(new_n7048), .B(new_n7047), .Y(new_n7049));
  NOR2xp33_ASAP7_75t_L      g06793(.A(new_n7046), .B(new_n7049), .Y(\f[46] ));
  NAND2xp33_ASAP7_75t_L     g06794(.A(new_n7021), .B(new_n7024), .Y(new_n7051));
  MAJIxp5_ASAP7_75t_L       g06795(.A(new_n7028), .B(new_n6779), .C(new_n7051), .Y(new_n7052));
  NAND2xp33_ASAP7_75t_L     g06796(.A(\b[42] ), .B(new_n366), .Y(new_n7053));
  NAND2xp33_ASAP7_75t_L     g06797(.A(\b[43] ), .B(new_n334), .Y(new_n7054));
  INVx1_ASAP7_75t_L         g06798(.A(new_n6229), .Y(new_n7055));
  AOI22xp33_ASAP7_75t_L     g06799(.A1(new_n345), .A2(\b[44] ), .B1(new_n342), .B2(new_n7055), .Y(new_n7056));
  AND4x1_ASAP7_75t_L        g06800(.A(new_n7056), .B(new_n7054), .C(new_n7053), .D(\a[5] ), .Y(new_n7057));
  AOI31xp33_ASAP7_75t_L     g06801(.A1(new_n7056), .A2(new_n7054), .A3(new_n7053), .B(\a[5] ), .Y(new_n7058));
  NOR2xp33_ASAP7_75t_L      g06802(.A(new_n7058), .B(new_n7057), .Y(new_n7059));
  INVx1_ASAP7_75t_L         g06803(.A(new_n7059), .Y(new_n7060));
  OAI21xp33_ASAP7_75t_L     g06804(.A1(new_n6980), .A2(new_n6979), .B(new_n6977), .Y(new_n7061));
  NAND2xp33_ASAP7_75t_L     g06805(.A(\b[30] ), .B(new_n1194), .Y(new_n7062));
  NAND2xp33_ASAP7_75t_L     g06806(.A(\b[31] ), .B(new_n1103), .Y(new_n7063));
  AOI22xp33_ASAP7_75t_L     g06807(.A1(new_n1113), .A2(\b[32] ), .B1(new_n1110), .B2(new_n3450), .Y(new_n7064));
  AND4x1_ASAP7_75t_L        g06808(.A(new_n7064), .B(new_n7063), .C(new_n7062), .D(\a[17] ), .Y(new_n7065));
  AOI31xp33_ASAP7_75t_L     g06809(.A1(new_n7064), .A2(new_n7063), .A3(new_n7062), .B(\a[17] ), .Y(new_n7066));
  NOR2xp33_ASAP7_75t_L      g06810(.A(new_n7066), .B(new_n7065), .Y(new_n7067));
  NOR2xp33_ASAP7_75t_L      g06811(.A(new_n6960), .B(new_n6959), .Y(new_n7068));
  MAJIxp5_ASAP7_75t_L       g06812(.A(new_n6974), .B(new_n6958), .C(new_n7068), .Y(new_n7069));
  NAND2xp33_ASAP7_75t_L     g06813(.A(\b[28] ), .B(new_n1410), .Y(new_n7070));
  OAI221xp5_ASAP7_75t_L     g06814(.A1(new_n1412), .A2(new_n2871), .B1(new_n1411), .B2(new_n2881), .C(new_n7070), .Y(new_n7071));
  AOI21xp33_ASAP7_75t_L     g06815(.A1(new_n1548), .A2(\b[27] ), .B(new_n7071), .Y(new_n7072));
  NAND2xp33_ASAP7_75t_L     g06816(.A(\a[20] ), .B(new_n7072), .Y(new_n7073));
  A2O1A1Ixp33_ASAP7_75t_L   g06817(.A1(\b[27] ), .A2(new_n1548), .B(new_n7071), .C(new_n1401), .Y(new_n7074));
  NAND2xp33_ASAP7_75t_L     g06818(.A(new_n7074), .B(new_n7073), .Y(new_n7075));
  INVx1_ASAP7_75t_L         g06819(.A(new_n7075), .Y(new_n7076));
  NOR2xp33_ASAP7_75t_L      g06820(.A(new_n6937), .B(new_n6931), .Y(new_n7077));
  MAJIxp5_ASAP7_75t_L       g06821(.A(new_n6951), .B(new_n6943), .C(new_n7077), .Y(new_n7078));
  AOI22xp33_ASAP7_75t_L     g06822(.A1(new_n1766), .A2(\b[26] ), .B1(new_n1764), .B2(new_n2888), .Y(new_n7079));
  OAI221xp5_ASAP7_75t_L     g06823(.A1(new_n1758), .A2(new_n2180), .B1(new_n2019), .B2(new_n1911), .C(new_n7079), .Y(new_n7080));
  XNOR2x2_ASAP7_75t_L       g06824(.A(new_n1761), .B(new_n7080), .Y(new_n7081));
  NOR3xp33_ASAP7_75t_L      g06825(.A(new_n6924), .B(new_n6922), .C(new_n6925), .Y(new_n7082));
  INVx1_ASAP7_75t_L         g06826(.A(new_n7082), .Y(new_n7083));
  OAI21xp33_ASAP7_75t_L     g06827(.A1(new_n6934), .A2(new_n6945), .B(new_n7083), .Y(new_n7084));
  NAND3xp33_ASAP7_75t_L     g06828(.A(new_n6897), .B(new_n6911), .C(new_n6902), .Y(new_n7085));
  A2O1A1Ixp33_ASAP7_75t_L   g06829(.A1(new_n6908), .A2(new_n6912), .B(new_n6913), .C(new_n7085), .Y(new_n7086));
  XNOR2x2_ASAP7_75t_L       g06830(.A(new_n6892), .B(new_n6880), .Y(new_n7087));
  MAJIxp5_ASAP7_75t_L       g06831(.A(new_n6901), .B(new_n6888), .C(new_n7087), .Y(new_n7088));
  NAND2xp33_ASAP7_75t_L     g06832(.A(\b[16] ), .B(new_n3260), .Y(new_n7089));
  OAI221xp5_ASAP7_75t_L     g06833(.A1(new_n3262), .A2(new_n1244), .B1(new_n3261), .B2(new_n1251), .C(new_n7089), .Y(new_n7090));
  INVx1_ASAP7_75t_L         g06834(.A(new_n7090), .Y(new_n7091));
  OAI211xp5_ASAP7_75t_L     g06835(.A1(new_n952), .A2(new_n3492), .B(new_n7091), .C(\a[32] ), .Y(new_n7092));
  A2O1A1Ixp33_ASAP7_75t_L   g06836(.A1(\b[15] ), .A2(new_n3491), .B(new_n7090), .C(new_n3251), .Y(new_n7093));
  NAND2xp33_ASAP7_75t_L     g06837(.A(new_n7093), .B(new_n7092), .Y(new_n7094));
  A2O1A1O1Ixp25_ASAP7_75t_L g06838(.A1(new_n6525), .A2(new_n6604), .B(new_n6876), .C(new_n6878), .D(new_n6872), .Y(new_n7095));
  NAND2xp33_ASAP7_75t_L     g06839(.A(new_n6830), .B(new_n6836), .Y(new_n7096));
  NOR2xp33_ASAP7_75t_L      g06840(.A(new_n6840), .B(new_n6846), .Y(new_n7097));
  NOR2xp33_ASAP7_75t_L      g06841(.A(new_n7096), .B(new_n7097), .Y(new_n7098));
  NOR2xp33_ASAP7_75t_L      g06842(.A(new_n382), .B(new_n5521), .Y(new_n7099));
  INVx1_ASAP7_75t_L         g06843(.A(new_n7099), .Y(new_n7100));
  NAND2xp33_ASAP7_75t_L     g06844(.A(\b[7] ), .B(new_n5240), .Y(new_n7101));
  AOI32xp33_ASAP7_75t_L     g06845(.A1(new_n508), .A2(new_n506), .A3(new_n5247), .B1(\b[8] ), .B2(new_n5249), .Y(new_n7102));
  NAND4xp25_ASAP7_75t_L     g06846(.A(new_n7102), .B(\a[41] ), .C(new_n7100), .D(new_n7101), .Y(new_n7103));
  AOI31xp33_ASAP7_75t_L     g06847(.A1(new_n7102), .A2(new_n7101), .A3(new_n7100), .B(\a[41] ), .Y(new_n7104));
  INVx1_ASAP7_75t_L         g06848(.A(new_n7104), .Y(new_n7105));
  INVx1_ASAP7_75t_L         g06849(.A(new_n6802), .Y(new_n7106));
  A2O1A1Ixp33_ASAP7_75t_L   g06850(.A1(new_n6558), .A2(new_n7106), .B(new_n6834), .C(new_n6829), .Y(new_n7107));
  NAND2xp33_ASAP7_75t_L     g06851(.A(\b[3] ), .B(new_n6308), .Y(new_n7108));
  NAND2xp33_ASAP7_75t_L     g06852(.A(\b[4] ), .B(new_n5992), .Y(new_n7109));
  AOI22xp33_ASAP7_75t_L     g06853(.A1(new_n6002), .A2(\b[5] ), .B1(new_n5999), .B2(new_n360), .Y(new_n7110));
  NAND4xp25_ASAP7_75t_L     g06854(.A(new_n7110), .B(\a[44] ), .C(new_n7108), .D(new_n7109), .Y(new_n7111));
  OAI221xp5_ASAP7_75t_L     g06855(.A1(new_n6312), .A2(new_n353), .B1(new_n6311), .B2(new_n359), .C(new_n7109), .Y(new_n7112));
  A2O1A1Ixp33_ASAP7_75t_L   g06856(.A1(\b[3] ), .A2(new_n6308), .B(new_n7112), .C(new_n5996), .Y(new_n7113));
  AND3x1_ASAP7_75t_L        g06857(.A(new_n6820), .B(new_n6823), .C(new_n6813), .Y(new_n7114));
  NAND3xp33_ASAP7_75t_L     g06858(.A(new_n6540), .B(new_n6811), .C(new_n6821), .Y(new_n7115));
  NOR2xp33_ASAP7_75t_L      g06859(.A(new_n258), .B(new_n7115), .Y(new_n7116));
  NAND2xp33_ASAP7_75t_L     g06860(.A(new_n6821), .B(new_n6810), .Y(new_n7117));
  INVx1_ASAP7_75t_L         g06861(.A(new_n6822), .Y(new_n7118));
  NAND2xp33_ASAP7_75t_L     g06862(.A(\b[1] ), .B(new_n6812), .Y(new_n7119));
  OAI221xp5_ASAP7_75t_L     g06863(.A1(new_n7117), .A2(new_n283), .B1(new_n278), .B2(new_n7118), .C(new_n7119), .Y(new_n7120));
  NOR2xp33_ASAP7_75t_L      g06864(.A(new_n7116), .B(new_n7120), .Y(new_n7121));
  A2O1A1Ixp33_ASAP7_75t_L   g06865(.A1(new_n6801), .A2(new_n7114), .B(new_n6816), .C(new_n7121), .Y(new_n7122));
  O2A1O1Ixp33_ASAP7_75t_L   g06866(.A1(new_n258), .A2(new_n6540), .B(new_n7114), .C(new_n6816), .Y(new_n7123));
  INVx1_ASAP7_75t_L         g06867(.A(new_n7115), .Y(new_n7124));
  A2O1A1Ixp33_ASAP7_75t_L   g06868(.A1(\b[0] ), .A2(new_n7124), .B(new_n7120), .C(new_n7123), .Y(new_n7125));
  NAND4xp25_ASAP7_75t_L     g06869(.A(new_n7125), .B(new_n7111), .C(new_n7113), .D(new_n7122), .Y(new_n7126));
  AOI211xp5_ASAP7_75t_L     g06870(.A1(\b[3] ), .A2(new_n6308), .B(new_n5996), .C(new_n7112), .Y(new_n7127));
  INVx1_ASAP7_75t_L         g06871(.A(new_n7113), .Y(new_n7128));
  NOR2xp33_ASAP7_75t_L      g06872(.A(new_n7117), .B(new_n283), .Y(new_n7129));
  AOI221xp5_ASAP7_75t_L     g06873(.A1(\b[2] ), .A2(new_n6822), .B1(new_n6812), .B2(\b[1] ), .C(new_n7129), .Y(new_n7130));
  OAI21xp33_ASAP7_75t_L     g06874(.A1(new_n258), .A2(new_n7115), .B(new_n7130), .Y(new_n7131));
  O2A1O1Ixp33_ASAP7_75t_L   g06875(.A1(new_n6541), .A2(new_n6824), .B(\a[47] ), .C(new_n7131), .Y(new_n7132));
  A2O1A1Ixp33_ASAP7_75t_L   g06876(.A1(\b[0] ), .A2(new_n6810), .B(new_n6824), .C(\a[47] ), .Y(new_n7133));
  O2A1O1Ixp33_ASAP7_75t_L   g06877(.A1(new_n7115), .A2(new_n258), .B(new_n7130), .C(new_n7133), .Y(new_n7134));
  OAI22xp33_ASAP7_75t_L     g06878(.A1(new_n7128), .A2(new_n7127), .B1(new_n7134), .B2(new_n7132), .Y(new_n7135));
  NAND2xp33_ASAP7_75t_L     g06879(.A(new_n7126), .B(new_n7135), .Y(new_n7136));
  NAND2xp33_ASAP7_75t_L     g06880(.A(new_n7136), .B(new_n7107), .Y(new_n7137));
  O2A1O1Ixp33_ASAP7_75t_L   g06881(.A1(new_n6802), .A2(new_n6549), .B(new_n6826), .C(new_n6835), .Y(new_n7138));
  NAND3xp33_ASAP7_75t_L     g06882(.A(new_n7138), .B(new_n7126), .C(new_n7135), .Y(new_n7139));
  AOI22xp33_ASAP7_75t_L     g06883(.A1(new_n7105), .A2(new_n7103), .B1(new_n7139), .B2(new_n7137), .Y(new_n7140));
  INVx1_ASAP7_75t_L         g06884(.A(new_n7103), .Y(new_n7141));
  AOI21xp33_ASAP7_75t_L     g06885(.A1(new_n7135), .A2(new_n7126), .B(new_n7138), .Y(new_n7142));
  NOR2xp33_ASAP7_75t_L      g06886(.A(new_n7136), .B(new_n7107), .Y(new_n7143));
  NOR4xp25_ASAP7_75t_L      g06887(.A(new_n7143), .B(new_n7142), .C(new_n7141), .D(new_n7104), .Y(new_n7144));
  NOR2xp33_ASAP7_75t_L      g06888(.A(new_n7140), .B(new_n7144), .Y(new_n7145));
  A2O1A1Ixp33_ASAP7_75t_L   g06889(.A1(new_n6851), .A2(new_n6848), .B(new_n7098), .C(new_n7145), .Y(new_n7146));
  AOI21xp33_ASAP7_75t_L     g06890(.A1(new_n6851), .A2(new_n6848), .B(new_n7098), .Y(new_n7147));
  OAI22xp33_ASAP7_75t_L     g06891(.A1(new_n7143), .A2(new_n7142), .B1(new_n7104), .B2(new_n7141), .Y(new_n7148));
  NAND4xp25_ASAP7_75t_L     g06892(.A(new_n7137), .B(new_n7139), .C(new_n7103), .D(new_n7105), .Y(new_n7149));
  NAND2xp33_ASAP7_75t_L     g06893(.A(new_n7149), .B(new_n7148), .Y(new_n7150));
  NAND2xp33_ASAP7_75t_L     g06894(.A(new_n7150), .B(new_n7147), .Y(new_n7151));
  NOR2xp33_ASAP7_75t_L      g06895(.A(new_n559), .B(new_n4781), .Y(new_n7152));
  INVx1_ASAP7_75t_L         g06896(.A(new_n7152), .Y(new_n7153));
  NAND2xp33_ASAP7_75t_L     g06897(.A(\b[10] ), .B(new_n4548), .Y(new_n7154));
  AOI32xp33_ASAP7_75t_L     g06898(.A1(new_n700), .A2(new_n698), .A3(new_n4542), .B1(\b[11] ), .B2(new_n4544), .Y(new_n7155));
  AND4x1_ASAP7_75t_L        g06899(.A(new_n7155), .B(new_n7154), .C(new_n7153), .D(\a[38] ), .Y(new_n7156));
  AOI31xp33_ASAP7_75t_L     g06900(.A1(new_n7155), .A2(new_n7154), .A3(new_n7153), .B(\a[38] ), .Y(new_n7157));
  NOR2xp33_ASAP7_75t_L      g06901(.A(new_n7157), .B(new_n7156), .Y(new_n7158));
  NAND3xp33_ASAP7_75t_L     g06902(.A(new_n7146), .B(new_n7151), .C(new_n7158), .Y(new_n7159));
  OAI211xp5_ASAP7_75t_L     g06903(.A1(new_n6840), .A2(new_n6846), .B(new_n6836), .C(new_n6830), .Y(new_n7160));
  A2O1A1O1Ixp25_ASAP7_75t_L g06904(.A1(new_n6847), .A2(new_n6843), .B(new_n6853), .C(new_n7160), .D(new_n7150), .Y(new_n7161));
  A2O1A1Ixp33_ASAP7_75t_L   g06905(.A1(new_n6847), .A2(new_n6843), .B(new_n6853), .C(new_n7160), .Y(new_n7162));
  NOR2xp33_ASAP7_75t_L      g06906(.A(new_n7145), .B(new_n7162), .Y(new_n7163));
  INVx1_ASAP7_75t_L         g06907(.A(new_n7158), .Y(new_n7164));
  OAI21xp33_ASAP7_75t_L     g06908(.A1(new_n7163), .A2(new_n7161), .B(new_n7164), .Y(new_n7165));
  AOI21xp33_ASAP7_75t_L     g06909(.A1(new_n6864), .A2(new_n6863), .B(new_n6865), .Y(new_n7166));
  OAI21xp33_ASAP7_75t_L     g06910(.A1(new_n7166), .A2(new_n6800), .B(new_n6866), .Y(new_n7167));
  NAND3xp33_ASAP7_75t_L     g06911(.A(new_n7167), .B(new_n7165), .C(new_n7159), .Y(new_n7168));
  NOR3xp33_ASAP7_75t_L      g06912(.A(new_n7161), .B(new_n7163), .C(new_n7164), .Y(new_n7169));
  AOI21xp33_ASAP7_75t_L     g06913(.A1(new_n7146), .A2(new_n7151), .B(new_n7158), .Y(new_n7170));
  A2O1A1Ixp33_ASAP7_75t_L   g06914(.A1(new_n6593), .A2(new_n6586), .B(new_n6582), .C(new_n6862), .Y(new_n7171));
  OAI211xp5_ASAP7_75t_L     g06915(.A1(new_n7169), .A2(new_n7170), .B(new_n7171), .C(new_n6866), .Y(new_n7172));
  NAND2xp33_ASAP7_75t_L     g06916(.A(\b[12] ), .B(new_n4111), .Y(new_n7173));
  NAND2xp33_ASAP7_75t_L     g06917(.A(\b[13] ), .B(new_n3874), .Y(new_n7174));
  AOI32xp33_ASAP7_75t_L     g06918(.A1(new_n877), .A2(new_n874), .A3(new_n3881), .B1(\b[14] ), .B2(new_n3884), .Y(new_n7175));
  AND4x1_ASAP7_75t_L        g06919(.A(new_n7175), .B(new_n7174), .C(new_n7173), .D(\a[35] ), .Y(new_n7176));
  AOI31xp33_ASAP7_75t_L     g06920(.A1(new_n7175), .A2(new_n7174), .A3(new_n7173), .B(\a[35] ), .Y(new_n7177));
  NOR2xp33_ASAP7_75t_L      g06921(.A(new_n7177), .B(new_n7176), .Y(new_n7178));
  NAND3xp33_ASAP7_75t_L     g06922(.A(new_n7168), .B(new_n7172), .C(new_n7178), .Y(new_n7179));
  AOI211xp5_ASAP7_75t_L     g06923(.A1(new_n7171), .A2(new_n6866), .B(new_n7169), .C(new_n7170), .Y(new_n7180));
  AOI21xp33_ASAP7_75t_L     g06924(.A1(new_n7165), .A2(new_n7159), .B(new_n7167), .Y(new_n7181));
  INVx1_ASAP7_75t_L         g06925(.A(new_n7178), .Y(new_n7182));
  OAI21xp33_ASAP7_75t_L     g06926(.A1(new_n7181), .A2(new_n7180), .B(new_n7182), .Y(new_n7183));
  AOI21xp33_ASAP7_75t_L     g06927(.A1(new_n7183), .A2(new_n7179), .B(new_n7095), .Y(new_n7184));
  NAND2xp33_ASAP7_75t_L     g06928(.A(new_n6591), .B(new_n6792), .Y(new_n7185));
  A2O1A1Ixp33_ASAP7_75t_L   g06929(.A1(new_n6596), .A2(new_n7185), .B(new_n6869), .C(new_n6879), .Y(new_n7186));
  NAND2xp33_ASAP7_75t_L     g06930(.A(new_n7179), .B(new_n7183), .Y(new_n7187));
  NOR2xp33_ASAP7_75t_L      g06931(.A(new_n7187), .B(new_n7186), .Y(new_n7188));
  OAI21xp33_ASAP7_75t_L     g06932(.A1(new_n7184), .A2(new_n7188), .B(new_n7094), .Y(new_n7189));
  NAND2xp33_ASAP7_75t_L     g06933(.A(new_n7187), .B(new_n7186), .Y(new_n7190));
  NAND3xp33_ASAP7_75t_L     g06934(.A(new_n7095), .B(new_n7179), .C(new_n7183), .Y(new_n7191));
  NAND4xp25_ASAP7_75t_L     g06935(.A(new_n7190), .B(new_n7191), .C(new_n7092), .D(new_n7093), .Y(new_n7192));
  NAND2xp33_ASAP7_75t_L     g06936(.A(new_n7189), .B(new_n7192), .Y(new_n7193));
  NOR2xp33_ASAP7_75t_L      g06937(.A(new_n7088), .B(new_n7193), .Y(new_n7194));
  NOR3xp33_ASAP7_75t_L      g06938(.A(new_n6889), .B(new_n6891), .C(new_n6893), .Y(new_n7195));
  AOI211xp5_ASAP7_75t_L     g06939(.A1(new_n7189), .A2(new_n7192), .B(new_n7195), .C(new_n6910), .Y(new_n7196));
  NOR2xp33_ASAP7_75t_L      g06940(.A(new_n1594), .B(new_n2708), .Y(new_n7197));
  AOI221xp5_ASAP7_75t_L     g06941(.A1(new_n2706), .A2(\b[19] ), .B1(new_n2700), .B2(new_n1600), .C(new_n7197), .Y(new_n7198));
  OA211x2_ASAP7_75t_L       g06942(.A1(new_n2932), .A2(new_n1356), .B(new_n7198), .C(\a[29] ), .Y(new_n7199));
  O2A1O1Ixp33_ASAP7_75t_L   g06943(.A1(new_n1356), .A2(new_n2932), .B(new_n7198), .C(\a[29] ), .Y(new_n7200));
  OAI22xp33_ASAP7_75t_L     g06944(.A1(new_n7196), .A2(new_n7194), .B1(new_n7200), .B2(new_n7199), .Y(new_n7201));
  OAI211xp5_ASAP7_75t_L     g06945(.A1(new_n7195), .A2(new_n6910), .B(new_n7189), .C(new_n7192), .Y(new_n7202));
  NAND2xp33_ASAP7_75t_L     g06946(.A(new_n7088), .B(new_n7193), .Y(new_n7203));
  NOR2xp33_ASAP7_75t_L      g06947(.A(new_n7200), .B(new_n7199), .Y(new_n7204));
  NAND3xp33_ASAP7_75t_L     g06948(.A(new_n7202), .B(new_n7204), .C(new_n7203), .Y(new_n7205));
  AOI21xp33_ASAP7_75t_L     g06949(.A1(new_n7201), .A2(new_n7205), .B(new_n7086), .Y(new_n7206));
  AND3x1_ASAP7_75t_L        g06950(.A(new_n7086), .B(new_n7201), .C(new_n7205), .Y(new_n7207));
  NOR2xp33_ASAP7_75t_L      g06951(.A(new_n1709), .B(new_n2387), .Y(new_n7208));
  NAND2xp33_ASAP7_75t_L     g06952(.A(\b[22] ), .B(new_n2232), .Y(new_n7209));
  OAI221xp5_ASAP7_75t_L     g06953(.A1(new_n2234), .A2(new_n1995), .B1(new_n2233), .B2(new_n4860), .C(new_n7209), .Y(new_n7210));
  NOR3xp33_ASAP7_75t_L      g06954(.A(new_n7210), .B(new_n7208), .C(new_n2223), .Y(new_n7211));
  OA21x2_ASAP7_75t_L        g06955(.A1(new_n7208), .A2(new_n7210), .B(new_n2223), .Y(new_n7212));
  NOR2xp33_ASAP7_75t_L      g06956(.A(new_n7211), .B(new_n7212), .Y(new_n7213));
  OAI21xp33_ASAP7_75t_L     g06957(.A1(new_n7206), .A2(new_n7207), .B(new_n7213), .Y(new_n7214));
  AO21x2_ASAP7_75t_L        g06958(.A1(new_n7205), .A2(new_n7201), .B(new_n7086), .Y(new_n7215));
  NAND3xp33_ASAP7_75t_L     g06959(.A(new_n7086), .B(new_n7201), .C(new_n7205), .Y(new_n7216));
  OR2x4_ASAP7_75t_L         g06960(.A(new_n7211), .B(new_n7212), .Y(new_n7217));
  NAND3xp33_ASAP7_75t_L     g06961(.A(new_n7217), .B(new_n7215), .C(new_n7216), .Y(new_n7218));
  NAND2xp33_ASAP7_75t_L     g06962(.A(new_n7214), .B(new_n7218), .Y(new_n7219));
  NOR2xp33_ASAP7_75t_L      g06963(.A(new_n7219), .B(new_n7084), .Y(new_n7220));
  AOI21xp33_ASAP7_75t_L     g06964(.A1(new_n7215), .A2(new_n7216), .B(new_n7217), .Y(new_n7221));
  NOR3xp33_ASAP7_75t_L      g06965(.A(new_n7207), .B(new_n7213), .C(new_n7206), .Y(new_n7222));
  NOR2xp33_ASAP7_75t_L      g06966(.A(new_n7221), .B(new_n7222), .Y(new_n7223));
  O2A1O1Ixp33_ASAP7_75t_L   g06967(.A1(new_n6934), .A2(new_n6945), .B(new_n7083), .C(new_n7223), .Y(new_n7224));
  NOR3xp33_ASAP7_75t_L      g06968(.A(new_n7224), .B(new_n7081), .C(new_n7220), .Y(new_n7225));
  XNOR2x2_ASAP7_75t_L       g06969(.A(\a[23] ), .B(new_n7080), .Y(new_n7226));
  A2O1A1O1Ixp25_ASAP7_75t_L g06970(.A1(new_n6641), .A2(new_n6638), .B(new_n6935), .C(new_n6928), .D(new_n7082), .Y(new_n7227));
  NAND2xp33_ASAP7_75t_L     g06971(.A(new_n7227), .B(new_n7223), .Y(new_n7228));
  A2O1A1Ixp33_ASAP7_75t_L   g06972(.A1(new_n6930), .A2(new_n6928), .B(new_n7082), .C(new_n7219), .Y(new_n7229));
  AOI21xp33_ASAP7_75t_L     g06973(.A1(new_n7229), .A2(new_n7228), .B(new_n7226), .Y(new_n7230));
  NOR3xp33_ASAP7_75t_L      g06974(.A(new_n7078), .B(new_n7225), .C(new_n7230), .Y(new_n7231));
  NAND2xp33_ASAP7_75t_L     g06975(.A(new_n6953), .B(new_n6954), .Y(new_n7232));
  NAND2xp33_ASAP7_75t_L     g06976(.A(new_n6947), .B(new_n6946), .Y(new_n7233));
  NOR2xp33_ASAP7_75t_L      g06977(.A(new_n6948), .B(new_n7233), .Y(new_n7234));
  NAND3xp33_ASAP7_75t_L     g06978(.A(new_n7229), .B(new_n7226), .C(new_n7228), .Y(new_n7235));
  OAI21xp33_ASAP7_75t_L     g06979(.A1(new_n7220), .A2(new_n7224), .B(new_n7081), .Y(new_n7236));
  AOI221xp5_ASAP7_75t_L     g06980(.A1(new_n7232), .A2(new_n6951), .B1(new_n7235), .B2(new_n7236), .C(new_n7234), .Y(new_n7237));
  OAI21xp33_ASAP7_75t_L     g06981(.A1(new_n7237), .A2(new_n7231), .B(new_n7076), .Y(new_n7238));
  MAJIxp5_ASAP7_75t_L       g06982(.A(new_n6955), .B(new_n7233), .C(new_n6948), .Y(new_n7239));
  NAND3xp33_ASAP7_75t_L     g06983(.A(new_n7239), .B(new_n7235), .C(new_n7236), .Y(new_n7240));
  OAI21xp33_ASAP7_75t_L     g06984(.A1(new_n7225), .A2(new_n7230), .B(new_n7078), .Y(new_n7241));
  NAND3xp33_ASAP7_75t_L     g06985(.A(new_n7240), .B(new_n7075), .C(new_n7241), .Y(new_n7242));
  NAND2xp33_ASAP7_75t_L     g06986(.A(new_n7238), .B(new_n7242), .Y(new_n7243));
  NOR2xp33_ASAP7_75t_L      g06987(.A(new_n7069), .B(new_n7243), .Y(new_n7244));
  NOR3xp33_ASAP7_75t_L      g06988(.A(new_n6959), .B(new_n6791), .C(new_n6960), .Y(new_n7245));
  AOI221xp5_ASAP7_75t_L     g06989(.A1(new_n6974), .A2(new_n6967), .B1(new_n7238), .B2(new_n7242), .C(new_n7245), .Y(new_n7246));
  OAI21xp33_ASAP7_75t_L     g06990(.A1(new_n7246), .A2(new_n7244), .B(new_n7067), .Y(new_n7247));
  INVx1_ASAP7_75t_L         g06991(.A(new_n7067), .Y(new_n7248));
  INVx1_ASAP7_75t_L         g06992(.A(new_n7245), .Y(new_n7249));
  A2O1A1Ixp33_ASAP7_75t_L   g06993(.A1(new_n6965), .A2(new_n6966), .B(new_n6964), .C(new_n7249), .Y(new_n7250));
  NAND3xp33_ASAP7_75t_L     g06994(.A(new_n7250), .B(new_n7238), .C(new_n7242), .Y(new_n7251));
  NAND2xp33_ASAP7_75t_L     g06995(.A(new_n7069), .B(new_n7243), .Y(new_n7252));
  NAND3xp33_ASAP7_75t_L     g06996(.A(new_n7251), .B(new_n7248), .C(new_n7252), .Y(new_n7253));
  NAND3xp33_ASAP7_75t_L     g06997(.A(new_n7061), .B(new_n7247), .C(new_n7253), .Y(new_n7254));
  INVx1_ASAP7_75t_L         g06998(.A(new_n6256), .Y(new_n7255));
  OAI21xp33_ASAP7_75t_L     g06999(.A1(new_n6253), .A2(new_n6254), .B(new_n5962), .Y(new_n7256));
  AOI21xp33_ASAP7_75t_L     g07000(.A1(new_n6430), .A2(new_n6431), .B(new_n6429), .Y(new_n7257));
  A2O1A1Ixp33_ASAP7_75t_L   g07001(.A1(new_n7256), .A2(new_n7255), .B(new_n7257), .C(new_n6432), .Y(new_n7258));
  A2O1A1O1Ixp25_ASAP7_75t_L g07002(.A1(new_n6687), .A2(new_n7258), .B(new_n6682), .C(new_n6972), .D(new_n6981), .Y(new_n7259));
  AOI21xp33_ASAP7_75t_L     g07003(.A1(new_n7251), .A2(new_n7252), .B(new_n7248), .Y(new_n7260));
  NOR3xp33_ASAP7_75t_L      g07004(.A(new_n7244), .B(new_n7246), .C(new_n7067), .Y(new_n7261));
  OAI21xp33_ASAP7_75t_L     g07005(.A1(new_n7260), .A2(new_n7261), .B(new_n7259), .Y(new_n7262));
  NAND2xp33_ASAP7_75t_L     g07006(.A(\b[33] ), .B(new_n908), .Y(new_n7263));
  NAND2xp33_ASAP7_75t_L     g07007(.A(\b[34] ), .B(new_n817), .Y(new_n7264));
  AOI22xp33_ASAP7_75t_L     g07008(.A1(new_n826), .A2(\b[35] ), .B1(new_n823), .B2(new_n5649), .Y(new_n7265));
  AND4x1_ASAP7_75t_L        g07009(.A(new_n7265), .B(new_n7264), .C(new_n7263), .D(\a[14] ), .Y(new_n7266));
  AOI31xp33_ASAP7_75t_L     g07010(.A1(new_n7265), .A2(new_n7264), .A3(new_n7263), .B(\a[14] ), .Y(new_n7267));
  NOR2xp33_ASAP7_75t_L      g07011(.A(new_n7267), .B(new_n7266), .Y(new_n7268));
  NAND3xp33_ASAP7_75t_L     g07012(.A(new_n7254), .B(new_n7262), .C(new_n7268), .Y(new_n7269));
  NOR3xp33_ASAP7_75t_L      g07013(.A(new_n7259), .B(new_n7260), .C(new_n7261), .Y(new_n7270));
  AOI221xp5_ASAP7_75t_L     g07014(.A1(new_n6782), .A2(new_n6972), .B1(new_n7247), .B2(new_n7253), .C(new_n6981), .Y(new_n7271));
  INVx1_ASAP7_75t_L         g07015(.A(new_n7268), .Y(new_n7272));
  OAI21xp33_ASAP7_75t_L     g07016(.A1(new_n7271), .A2(new_n7270), .B(new_n7272), .Y(new_n7273));
  NAND2xp33_ASAP7_75t_L     g07017(.A(new_n7269), .B(new_n7273), .Y(new_n7274));
  NAND2xp33_ASAP7_75t_L     g07018(.A(new_n6982), .B(new_n6978), .Y(new_n7275));
  MAJIxp5_ASAP7_75t_L       g07019(.A(new_n6993), .B(new_n7275), .C(new_n6989), .Y(new_n7276));
  NOR2xp33_ASAP7_75t_L      g07020(.A(new_n7276), .B(new_n7274), .Y(new_n7277));
  OAI211xp5_ASAP7_75t_L     g07021(.A1(new_n6986), .A2(new_n6988), .B(new_n6978), .C(new_n6982), .Y(new_n7278));
  AOI22xp33_ASAP7_75t_L     g07022(.A1(new_n7269), .A2(new_n7273), .B1(new_n7278), .B2(new_n6997), .Y(new_n7279));
  NAND2xp33_ASAP7_75t_L     g07023(.A(\b[36] ), .B(new_n674), .Y(new_n7280));
  NAND2xp33_ASAP7_75t_L     g07024(.A(\b[37] ), .B(new_n590), .Y(new_n7281));
  AOI22xp33_ASAP7_75t_L     g07025(.A1(new_n600), .A2(\b[38] ), .B1(new_n597), .B2(new_n4923), .Y(new_n7282));
  NAND4xp25_ASAP7_75t_L     g07026(.A(new_n7282), .B(\a[11] ), .C(new_n7280), .D(new_n7281), .Y(new_n7283));
  NAND2xp33_ASAP7_75t_L     g07027(.A(new_n7281), .B(new_n7282), .Y(new_n7284));
  A2O1A1Ixp33_ASAP7_75t_L   g07028(.A1(\b[36] ), .A2(new_n674), .B(new_n7284), .C(new_n594), .Y(new_n7285));
  NAND2xp33_ASAP7_75t_L     g07029(.A(new_n7283), .B(new_n7285), .Y(new_n7286));
  NOR3xp33_ASAP7_75t_L      g07030(.A(new_n7279), .B(new_n7277), .C(new_n7286), .Y(new_n7287));
  OA21x2_ASAP7_75t_L        g07031(.A1(new_n7277), .A2(new_n7279), .B(new_n7286), .Y(new_n7288));
  MAJIxp5_ASAP7_75t_L       g07032(.A(new_n7007), .B(new_n7004), .C(new_n7002), .Y(new_n7289));
  NOR3xp33_ASAP7_75t_L      g07033(.A(new_n7289), .B(new_n7288), .C(new_n7287), .Y(new_n7290));
  OA21x2_ASAP7_75t_L        g07034(.A1(new_n7287), .A2(new_n7288), .B(new_n7289), .Y(new_n7291));
  NAND2xp33_ASAP7_75t_L     g07035(.A(\b[39] ), .B(new_n480), .Y(new_n7292));
  NAND2xp33_ASAP7_75t_L     g07036(.A(\b[40] ), .B(new_n441), .Y(new_n7293));
  AOI22xp33_ASAP7_75t_L     g07037(.A1(new_n451), .A2(\b[41] ), .B1(new_n448), .B2(new_n5669), .Y(new_n7294));
  AND4x1_ASAP7_75t_L        g07038(.A(new_n7294), .B(new_n7293), .C(new_n7292), .D(\a[8] ), .Y(new_n7295));
  AOI31xp33_ASAP7_75t_L     g07039(.A1(new_n7294), .A2(new_n7293), .A3(new_n7292), .B(\a[8] ), .Y(new_n7296));
  NOR2xp33_ASAP7_75t_L      g07040(.A(new_n7296), .B(new_n7295), .Y(new_n7297));
  NOR3xp33_ASAP7_75t_L      g07041(.A(new_n7291), .B(new_n7297), .C(new_n7290), .Y(new_n7298));
  INVx1_ASAP7_75t_L         g07042(.A(new_n7298), .Y(new_n7299));
  OAI21xp33_ASAP7_75t_L     g07043(.A1(new_n7290), .A2(new_n7291), .B(new_n7297), .Y(new_n7300));
  INVx1_ASAP7_75t_L         g07044(.A(new_n6780), .Y(new_n7301));
  NAND3xp33_ASAP7_75t_L     g07045(.A(new_n7018), .B(new_n7019), .C(new_n7017), .Y(new_n7302));
  A2O1A1Ixp33_ASAP7_75t_L   g07046(.A1(new_n6737), .A2(new_n7301), .B(new_n7020), .C(new_n7302), .Y(new_n7303));
  NAND3xp33_ASAP7_75t_L     g07047(.A(new_n7299), .B(new_n7303), .C(new_n7300), .Y(new_n7304));
  INVx1_ASAP7_75t_L         g07048(.A(new_n7300), .Y(new_n7305));
  OAI21xp33_ASAP7_75t_L     g07049(.A1(new_n7009), .A2(new_n7008), .B(new_n7015), .Y(new_n7306));
  A2O1A1O1Ixp25_ASAP7_75t_L g07050(.A1(new_n6736), .A2(new_n7022), .B(new_n6780), .C(new_n7306), .D(new_n7016), .Y(new_n7307));
  OAI21xp33_ASAP7_75t_L     g07051(.A1(new_n7298), .A2(new_n7305), .B(new_n7307), .Y(new_n7308));
  AOI21xp33_ASAP7_75t_L     g07052(.A1(new_n7304), .A2(new_n7308), .B(new_n7060), .Y(new_n7309));
  NOR3xp33_ASAP7_75t_L      g07053(.A(new_n7307), .B(new_n7305), .C(new_n7298), .Y(new_n7310));
  AOI21xp33_ASAP7_75t_L     g07054(.A1(new_n7299), .A2(new_n7300), .B(new_n7303), .Y(new_n7311));
  NOR3xp33_ASAP7_75t_L      g07055(.A(new_n7310), .B(new_n7311), .C(new_n7059), .Y(new_n7312));
  NOR2xp33_ASAP7_75t_L      g07056(.A(new_n7309), .B(new_n7312), .Y(new_n7313));
  XNOR2x2_ASAP7_75t_L       g07057(.A(new_n7313), .B(new_n7052), .Y(new_n7314));
  NOR2xp33_ASAP7_75t_L      g07058(.A(\b[46] ), .B(\b[47] ), .Y(new_n7315));
  INVx1_ASAP7_75t_L         g07059(.A(\b[47] ), .Y(new_n7316));
  NOR2xp33_ASAP7_75t_L      g07060(.A(new_n7033), .B(new_n7316), .Y(new_n7317));
  NOR2xp33_ASAP7_75t_L      g07061(.A(new_n7315), .B(new_n7317), .Y(new_n7318));
  A2O1A1Ixp33_ASAP7_75t_L   g07062(.A1(new_n7039), .A2(new_n7035), .B(new_n7034), .C(new_n7318), .Y(new_n7319));
  O2A1O1Ixp33_ASAP7_75t_L   g07063(.A1(new_n6757), .A2(new_n6760), .B(new_n7035), .C(new_n7034), .Y(new_n7320));
  OAI21xp33_ASAP7_75t_L     g07064(.A1(new_n7315), .A2(new_n7317), .B(new_n7320), .Y(new_n7321));
  NAND2xp33_ASAP7_75t_L     g07065(.A(new_n7321), .B(new_n7319), .Y(new_n7322));
  INVx1_ASAP7_75t_L         g07066(.A(new_n7322), .Y(new_n7323));
  AOI22xp33_ASAP7_75t_L     g07067(.A1(new_n272), .A2(\b[47] ), .B1(new_n269), .B2(new_n7323), .Y(new_n7324));
  OAI221xp5_ASAP7_75t_L     g07068(.A1(new_n261), .A2(new_n7033), .B1(new_n6756), .B2(new_n277), .C(new_n7324), .Y(new_n7325));
  XNOR2x2_ASAP7_75t_L       g07069(.A(\a[2] ), .B(new_n7325), .Y(new_n7326));
  XOR2x2_ASAP7_75t_L        g07070(.A(new_n7326), .B(new_n7314), .Y(new_n7327));
  MAJIxp5_ASAP7_75t_L       g07071(.A(new_n7048), .B(new_n7031), .C(new_n7044), .Y(new_n7328));
  XNOR2x2_ASAP7_75t_L       g07072(.A(new_n7328), .B(new_n7327), .Y(\f[47] ));
  A2O1A1Ixp33_ASAP7_75t_L   g07073(.A1(new_n7044), .A2(new_n7031), .B(new_n7046), .C(new_n7327), .Y(new_n7330));
  INVx1_ASAP7_75t_L         g07074(.A(new_n7317), .Y(new_n7331));
  NOR2xp33_ASAP7_75t_L      g07075(.A(\b[47] ), .B(\b[48] ), .Y(new_n7332));
  INVx1_ASAP7_75t_L         g07076(.A(\b[48] ), .Y(new_n7333));
  NOR2xp33_ASAP7_75t_L      g07077(.A(new_n7316), .B(new_n7333), .Y(new_n7334));
  NOR2xp33_ASAP7_75t_L      g07078(.A(new_n7332), .B(new_n7334), .Y(new_n7335));
  INVx1_ASAP7_75t_L         g07079(.A(new_n7335), .Y(new_n7336));
  O2A1O1Ixp33_ASAP7_75t_L   g07080(.A1(new_n7315), .A2(new_n7320), .B(new_n7331), .C(new_n7336), .Y(new_n7337));
  A2O1A1O1Ixp25_ASAP7_75t_L g07081(.A1(new_n7035), .A2(new_n7039), .B(new_n7034), .C(new_n7318), .D(new_n7317), .Y(new_n7338));
  NAND2xp33_ASAP7_75t_L     g07082(.A(new_n7336), .B(new_n7338), .Y(new_n7339));
  INVx1_ASAP7_75t_L         g07083(.A(new_n7339), .Y(new_n7340));
  NOR2xp33_ASAP7_75t_L      g07084(.A(new_n7337), .B(new_n7340), .Y(new_n7341));
  AOI22xp33_ASAP7_75t_L     g07085(.A1(new_n272), .A2(\b[48] ), .B1(new_n269), .B2(new_n7341), .Y(new_n7342));
  OAI221xp5_ASAP7_75t_L     g07086(.A1(new_n261), .A2(new_n7316), .B1(new_n7033), .B2(new_n277), .C(new_n7342), .Y(new_n7343));
  XNOR2x2_ASAP7_75t_L       g07087(.A(\a[2] ), .B(new_n7343), .Y(new_n7344));
  NOR2xp33_ASAP7_75t_L      g07088(.A(new_n6779), .B(new_n7051), .Y(new_n7345));
  O2A1O1Ixp33_ASAP7_75t_L   g07089(.A1(new_n7345), .A2(new_n7030), .B(new_n7313), .C(new_n7312), .Y(new_n7346));
  NOR3xp33_ASAP7_75t_L      g07090(.A(new_n7270), .B(new_n7271), .C(new_n7268), .Y(new_n7347));
  AOI21xp33_ASAP7_75t_L     g07091(.A1(new_n7274), .A2(new_n7276), .B(new_n7347), .Y(new_n7348));
  NAND2xp33_ASAP7_75t_L     g07092(.A(\b[34] ), .B(new_n908), .Y(new_n7349));
  NAND2xp33_ASAP7_75t_L     g07093(.A(\b[35] ), .B(new_n817), .Y(new_n7350));
  AOI22xp33_ASAP7_75t_L     g07094(.A1(new_n826), .A2(\b[36] ), .B1(new_n823), .B2(new_n4473), .Y(new_n7351));
  AND4x1_ASAP7_75t_L        g07095(.A(new_n7351), .B(new_n7350), .C(new_n7349), .D(\a[14] ), .Y(new_n7352));
  AOI31xp33_ASAP7_75t_L     g07096(.A1(new_n7351), .A2(new_n7350), .A3(new_n7349), .B(\a[14] ), .Y(new_n7353));
  NOR2xp33_ASAP7_75t_L      g07097(.A(new_n7353), .B(new_n7352), .Y(new_n7354));
  INVx1_ASAP7_75t_L         g07098(.A(new_n7354), .Y(new_n7355));
  A2O1A1O1Ixp25_ASAP7_75t_L g07099(.A1(new_n6972), .A2(new_n6782), .B(new_n6981), .C(new_n7247), .D(new_n7261), .Y(new_n7356));
  NOR3xp33_ASAP7_75t_L      g07100(.A(new_n7076), .B(new_n7231), .C(new_n7237), .Y(new_n7357));
  NOR2xp33_ASAP7_75t_L      g07101(.A(new_n2852), .B(new_n1549), .Y(new_n7358));
  INVx1_ASAP7_75t_L         g07102(.A(new_n7358), .Y(new_n7359));
  NAND2xp33_ASAP7_75t_L     g07103(.A(\b[29] ), .B(new_n1410), .Y(new_n7360));
  AOI22xp33_ASAP7_75t_L     g07104(.A1(new_n1406), .A2(\b[30] ), .B1(new_n1404), .B2(new_n3219), .Y(new_n7361));
  AND4x1_ASAP7_75t_L        g07105(.A(new_n7361), .B(new_n7360), .C(new_n7359), .D(\a[20] ), .Y(new_n7362));
  AOI31xp33_ASAP7_75t_L     g07106(.A1(new_n7361), .A2(new_n7360), .A3(new_n7359), .B(\a[20] ), .Y(new_n7363));
  NOR2xp33_ASAP7_75t_L      g07107(.A(new_n7363), .B(new_n7362), .Y(new_n7364));
  A2O1A1O1Ixp25_ASAP7_75t_L g07108(.A1(new_n6951), .A2(new_n7232), .B(new_n7234), .C(new_n7235), .D(new_n7230), .Y(new_n7365));
  NAND3xp33_ASAP7_75t_L     g07109(.A(new_n7168), .B(new_n7172), .C(new_n7182), .Y(new_n7366));
  A2O1A1Ixp33_ASAP7_75t_L   g07110(.A1(new_n7179), .A2(new_n7183), .B(new_n7095), .C(new_n7366), .Y(new_n7367));
  NOR2xp33_ASAP7_75t_L      g07111(.A(new_n793), .B(new_n4986), .Y(new_n7368));
  NAND2xp33_ASAP7_75t_L     g07112(.A(\b[14] ), .B(new_n3874), .Y(new_n7369));
  OAI221xp5_ASAP7_75t_L     g07113(.A1(new_n4115), .A2(new_n952), .B1(new_n4114), .B2(new_n2573), .C(new_n7369), .Y(new_n7370));
  OR3x1_ASAP7_75t_L         g07114(.A(new_n7370), .B(new_n3878), .C(new_n7368), .Y(new_n7371));
  A2O1A1Ixp33_ASAP7_75t_L   g07115(.A1(\b[13] ), .A2(new_n4111), .B(new_n7370), .C(new_n3878), .Y(new_n7372));
  NAND2xp33_ASAP7_75t_L     g07116(.A(new_n7372), .B(new_n7371), .Y(new_n7373));
  A2O1A1Ixp33_ASAP7_75t_L   g07117(.A1(new_n7171), .A2(new_n6866), .B(new_n7169), .C(new_n7165), .Y(new_n7374));
  NOR2xp33_ASAP7_75t_L      g07118(.A(new_n631), .B(new_n4781), .Y(new_n7375));
  INVx1_ASAP7_75t_L         g07119(.A(new_n7375), .Y(new_n7376));
  NOR2xp33_ASAP7_75t_L      g07120(.A(new_n695), .B(new_n4536), .Y(new_n7377));
  INVx1_ASAP7_75t_L         g07121(.A(new_n7377), .Y(new_n7378));
  AOI22xp33_ASAP7_75t_L     g07122(.A1(new_n4544), .A2(\b[12] ), .B1(new_n4542), .B2(new_n970), .Y(new_n7379));
  AND4x1_ASAP7_75t_L        g07123(.A(new_n7379), .B(new_n7378), .C(new_n7376), .D(\a[38] ), .Y(new_n7380));
  AOI31xp33_ASAP7_75t_L     g07124(.A1(new_n7379), .A2(new_n7378), .A3(new_n7376), .B(\a[38] ), .Y(new_n7381));
  NOR2xp33_ASAP7_75t_L      g07125(.A(new_n7381), .B(new_n7380), .Y(new_n7382));
  AOI211xp5_ASAP7_75t_L     g07126(.A1(new_n7105), .A2(new_n7103), .B(new_n7142), .C(new_n7143), .Y(new_n7383));
  NAND5xp2_ASAP7_75t_L      g07127(.A(new_n6823), .B(new_n6820), .C(new_n6813), .D(new_n6801), .E(\a[47] ), .Y(new_n7384));
  INVx1_ASAP7_75t_L         g07128(.A(\a[48] ), .Y(new_n7385));
  NAND2xp33_ASAP7_75t_L     g07129(.A(\a[47] ), .B(new_n7385), .Y(new_n7386));
  NAND2xp33_ASAP7_75t_L     g07130(.A(\a[48] ), .B(new_n6816), .Y(new_n7387));
  AND2x2_ASAP7_75t_L        g07131(.A(new_n7386), .B(new_n7387), .Y(new_n7388));
  NOR2xp33_ASAP7_75t_L      g07132(.A(new_n258), .B(new_n7388), .Y(new_n7389));
  OAI31xp33_ASAP7_75t_L     g07133(.A1(new_n7384), .A2(new_n7120), .A3(new_n7116), .B(new_n7389), .Y(new_n7390));
  OR4x2_ASAP7_75t_L         g07134(.A(new_n7389), .B(new_n7384), .C(new_n7120), .D(new_n7116), .Y(new_n7391));
  INVx1_ASAP7_75t_L         g07135(.A(new_n6812), .Y(new_n7392));
  NAND2xp33_ASAP7_75t_L     g07136(.A(\b[3] ), .B(new_n6822), .Y(new_n7393));
  OAI221xp5_ASAP7_75t_L     g07137(.A1(new_n278), .A2(new_n7392), .B1(new_n7117), .B2(new_n303), .C(new_n7393), .Y(new_n7394));
  INVx1_ASAP7_75t_L         g07138(.A(new_n7394), .Y(new_n7395));
  OAI211xp5_ASAP7_75t_L     g07139(.A1(new_n276), .A2(new_n7115), .B(new_n7395), .C(\a[47] ), .Y(new_n7396));
  A2O1A1Ixp33_ASAP7_75t_L   g07140(.A1(\b[1] ), .A2(new_n7124), .B(new_n7394), .C(new_n6816), .Y(new_n7397));
  AO22x1_ASAP7_75t_L        g07141(.A1(new_n7390), .A2(new_n7391), .B1(new_n7397), .B2(new_n7396), .Y(new_n7398));
  NAND4xp25_ASAP7_75t_L     g07142(.A(new_n7396), .B(new_n7391), .C(new_n7390), .D(new_n7397), .Y(new_n7399));
  NAND2xp33_ASAP7_75t_L     g07143(.A(\b[4] ), .B(new_n6308), .Y(new_n7400));
  NAND2xp33_ASAP7_75t_L     g07144(.A(\b[5] ), .B(new_n5992), .Y(new_n7401));
  AOI22xp33_ASAP7_75t_L     g07145(.A1(new_n6002), .A2(\b[6] ), .B1(new_n5999), .B2(new_n389), .Y(new_n7402));
  NAND4xp25_ASAP7_75t_L     g07146(.A(new_n7402), .B(\a[44] ), .C(new_n7400), .D(new_n7401), .Y(new_n7403));
  OAI221xp5_ASAP7_75t_L     g07147(.A1(new_n6312), .A2(new_n382), .B1(new_n6311), .B2(new_n540), .C(new_n7401), .Y(new_n7404));
  A2O1A1Ixp33_ASAP7_75t_L   g07148(.A1(\b[4] ), .A2(new_n6308), .B(new_n7404), .C(new_n5996), .Y(new_n7405));
  NAND4xp25_ASAP7_75t_L     g07149(.A(new_n7398), .B(new_n7405), .C(new_n7403), .D(new_n7399), .Y(new_n7406));
  AOI22xp33_ASAP7_75t_L     g07150(.A1(new_n7391), .A2(new_n7390), .B1(new_n7397), .B2(new_n7396), .Y(new_n7407));
  AND4x1_ASAP7_75t_L        g07151(.A(new_n7391), .B(new_n7396), .C(new_n7390), .D(new_n7397), .Y(new_n7408));
  AOI211xp5_ASAP7_75t_L     g07152(.A1(\b[4] ), .A2(new_n6308), .B(new_n5996), .C(new_n7404), .Y(new_n7409));
  AOI31xp33_ASAP7_75t_L     g07153(.A1(new_n7402), .A2(new_n7401), .A3(new_n7400), .B(\a[44] ), .Y(new_n7410));
  OAI22xp33_ASAP7_75t_L     g07154(.A1(new_n7409), .A2(new_n7410), .B1(new_n7407), .B2(new_n7408), .Y(new_n7411));
  NAND2xp33_ASAP7_75t_L     g07155(.A(new_n7113), .B(new_n7111), .Y(new_n7412));
  NOR2xp33_ASAP7_75t_L      g07156(.A(new_n7132), .B(new_n7134), .Y(new_n7413));
  NAND2xp33_ASAP7_75t_L     g07157(.A(new_n7412), .B(new_n7413), .Y(new_n7414));
  NAND4xp25_ASAP7_75t_L     g07158(.A(new_n7137), .B(new_n7414), .C(new_n7411), .D(new_n7406), .Y(new_n7415));
  NAND2xp33_ASAP7_75t_L     g07159(.A(new_n7406), .B(new_n7411), .Y(new_n7416));
  A2O1A1Ixp33_ASAP7_75t_L   g07160(.A1(new_n7413), .A2(new_n7412), .B(new_n7142), .C(new_n7416), .Y(new_n7417));
  NAND2xp33_ASAP7_75t_L     g07161(.A(\b[7] ), .B(new_n5526), .Y(new_n7418));
  NAND2xp33_ASAP7_75t_L     g07162(.A(\b[8] ), .B(new_n5240), .Y(new_n7419));
  AOI22xp33_ASAP7_75t_L     g07163(.A1(new_n5249), .A2(\b[9] ), .B1(new_n5247), .B2(new_n566), .Y(new_n7420));
  NAND4xp25_ASAP7_75t_L     g07164(.A(new_n7420), .B(\a[41] ), .C(new_n7418), .D(new_n7419), .Y(new_n7421));
  INVx1_ASAP7_75t_L         g07165(.A(new_n7421), .Y(new_n7422));
  OAI221xp5_ASAP7_75t_L     g07166(.A1(new_n5253), .A2(new_n559), .B1(new_n5252), .B2(new_n978), .C(new_n7419), .Y(new_n7423));
  A2O1A1Ixp33_ASAP7_75t_L   g07167(.A1(\b[7] ), .A2(new_n5526), .B(new_n7423), .C(new_n5244), .Y(new_n7424));
  INVx1_ASAP7_75t_L         g07168(.A(new_n7424), .Y(new_n7425));
  AOI211xp5_ASAP7_75t_L     g07169(.A1(new_n7415), .A2(new_n7417), .B(new_n7422), .C(new_n7425), .Y(new_n7426));
  A2O1A1Ixp33_ASAP7_75t_L   g07170(.A1(new_n7126), .A2(new_n7135), .B(new_n7138), .C(new_n7414), .Y(new_n7427));
  NOR2xp33_ASAP7_75t_L      g07171(.A(new_n7416), .B(new_n7427), .Y(new_n7428));
  AOI22xp33_ASAP7_75t_L     g07172(.A1(new_n7406), .A2(new_n7411), .B1(new_n7414), .B2(new_n7137), .Y(new_n7429));
  AOI211xp5_ASAP7_75t_L     g07173(.A1(new_n7424), .A2(new_n7421), .B(new_n7428), .C(new_n7429), .Y(new_n7430));
  NOR2xp33_ASAP7_75t_L      g07174(.A(new_n7430), .B(new_n7426), .Y(new_n7431));
  A2O1A1Ixp33_ASAP7_75t_L   g07175(.A1(new_n7150), .A2(new_n7162), .B(new_n7383), .C(new_n7431), .Y(new_n7432));
  A2O1A1O1Ixp25_ASAP7_75t_L g07176(.A1(new_n6851), .A2(new_n6848), .B(new_n7098), .C(new_n7150), .D(new_n7383), .Y(new_n7433));
  OAI211xp5_ASAP7_75t_L     g07177(.A1(new_n7428), .A2(new_n7429), .B(new_n7421), .C(new_n7424), .Y(new_n7434));
  OAI211xp5_ASAP7_75t_L     g07178(.A1(new_n7422), .A2(new_n7425), .B(new_n7415), .C(new_n7417), .Y(new_n7435));
  NAND2xp33_ASAP7_75t_L     g07179(.A(new_n7435), .B(new_n7434), .Y(new_n7436));
  NAND2xp33_ASAP7_75t_L     g07180(.A(new_n7436), .B(new_n7433), .Y(new_n7437));
  AOI21xp33_ASAP7_75t_L     g07181(.A1(new_n7432), .A2(new_n7437), .B(new_n7382), .Y(new_n7438));
  OR2x4_ASAP7_75t_L         g07182(.A(new_n7381), .B(new_n7380), .Y(new_n7439));
  NOR2xp33_ASAP7_75t_L      g07183(.A(new_n7436), .B(new_n7433), .Y(new_n7440));
  INVx1_ASAP7_75t_L         g07184(.A(new_n7383), .Y(new_n7441));
  A2O1A1Ixp33_ASAP7_75t_L   g07185(.A1(new_n7148), .A2(new_n7149), .B(new_n7147), .C(new_n7441), .Y(new_n7442));
  NOR2xp33_ASAP7_75t_L      g07186(.A(new_n7431), .B(new_n7442), .Y(new_n7443));
  NOR3xp33_ASAP7_75t_L      g07187(.A(new_n7439), .B(new_n7443), .C(new_n7440), .Y(new_n7444));
  OAI21xp33_ASAP7_75t_L     g07188(.A1(new_n7438), .A2(new_n7444), .B(new_n7374), .Y(new_n7445));
  AOI21xp33_ASAP7_75t_L     g07189(.A1(new_n7167), .A2(new_n7159), .B(new_n7170), .Y(new_n7446));
  OAI21xp33_ASAP7_75t_L     g07190(.A1(new_n7440), .A2(new_n7443), .B(new_n7439), .Y(new_n7447));
  NAND3xp33_ASAP7_75t_L     g07191(.A(new_n7432), .B(new_n7437), .C(new_n7382), .Y(new_n7448));
  NAND3xp33_ASAP7_75t_L     g07192(.A(new_n7446), .B(new_n7447), .C(new_n7448), .Y(new_n7449));
  NAND3xp33_ASAP7_75t_L     g07193(.A(new_n7449), .B(new_n7445), .C(new_n7373), .Y(new_n7450));
  AND2x2_ASAP7_75t_L        g07194(.A(new_n7372), .B(new_n7371), .Y(new_n7451));
  AOI21xp33_ASAP7_75t_L     g07195(.A1(new_n7448), .A2(new_n7447), .B(new_n7446), .Y(new_n7452));
  NOR3xp33_ASAP7_75t_L      g07196(.A(new_n7374), .B(new_n7438), .C(new_n7444), .Y(new_n7453));
  OAI21xp33_ASAP7_75t_L     g07197(.A1(new_n7452), .A2(new_n7453), .B(new_n7451), .Y(new_n7454));
  NAND3xp33_ASAP7_75t_L     g07198(.A(new_n7367), .B(new_n7450), .C(new_n7454), .Y(new_n7455));
  INVx1_ASAP7_75t_L         g07199(.A(new_n7366), .Y(new_n7456));
  A2O1A1O1Ixp25_ASAP7_75t_L g07200(.A1(new_n6892), .A2(new_n6873), .B(new_n6872), .C(new_n7187), .D(new_n7456), .Y(new_n7457));
  NAND2xp33_ASAP7_75t_L     g07201(.A(new_n7450), .B(new_n7454), .Y(new_n7458));
  NAND2xp33_ASAP7_75t_L     g07202(.A(new_n7458), .B(new_n7457), .Y(new_n7459));
  AOI22xp33_ASAP7_75t_L     g07203(.A1(new_n3256), .A2(\b[18] ), .B1(new_n3254), .B2(new_n1363), .Y(new_n7460));
  OAI221xp5_ASAP7_75t_L     g07204(.A1(new_n3248), .A2(new_n1244), .B1(new_n1051), .B2(new_n3492), .C(new_n7460), .Y(new_n7461));
  XNOR2x2_ASAP7_75t_L       g07205(.A(\a[32] ), .B(new_n7461), .Y(new_n7462));
  NAND3xp33_ASAP7_75t_L     g07206(.A(new_n7459), .B(new_n7455), .C(new_n7462), .Y(new_n7463));
  NAND2xp33_ASAP7_75t_L     g07207(.A(new_n7172), .B(new_n7168), .Y(new_n7464));
  O2A1O1Ixp33_ASAP7_75t_L   g07208(.A1(new_n7464), .A2(new_n7178), .B(new_n7190), .C(new_n7458), .Y(new_n7465));
  AOI21xp33_ASAP7_75t_L     g07209(.A1(new_n7454), .A2(new_n7450), .B(new_n7367), .Y(new_n7466));
  XNOR2x2_ASAP7_75t_L       g07210(.A(new_n3251), .B(new_n7461), .Y(new_n7467));
  OAI21xp33_ASAP7_75t_L     g07211(.A1(new_n7465), .A2(new_n7466), .B(new_n7467), .Y(new_n7468));
  NAND2xp33_ASAP7_75t_L     g07212(.A(new_n7468), .B(new_n7463), .Y(new_n7469));
  NAND3xp33_ASAP7_75t_L     g07213(.A(new_n7191), .B(new_n7190), .C(new_n7094), .Y(new_n7470));
  A2O1A1Ixp33_ASAP7_75t_L   g07214(.A1(new_n7189), .A2(new_n7192), .B(new_n7088), .C(new_n7470), .Y(new_n7471));
  NOR2xp33_ASAP7_75t_L      g07215(.A(new_n7471), .B(new_n7469), .Y(new_n7472));
  NOR3xp33_ASAP7_75t_L      g07216(.A(new_n7466), .B(new_n7465), .C(new_n7467), .Y(new_n7473));
  AOI21xp33_ASAP7_75t_L     g07217(.A1(new_n7459), .A2(new_n7455), .B(new_n7462), .Y(new_n7474));
  OAI21xp33_ASAP7_75t_L     g07218(.A1(new_n7473), .A2(new_n7474), .B(new_n7471), .Y(new_n7475));
  INVx1_ASAP7_75t_L         g07219(.A(new_n7475), .Y(new_n7476));
  NAND2xp33_ASAP7_75t_L     g07220(.A(\b[19] ), .B(new_n2931), .Y(new_n7477));
  NAND2xp33_ASAP7_75t_L     g07221(.A(\b[20] ), .B(new_n2706), .Y(new_n7478));
  AOI22xp33_ASAP7_75t_L     g07222(.A1(new_n2702), .A2(\b[21] ), .B1(new_n2700), .B2(new_n1715), .Y(new_n7479));
  NAND4xp25_ASAP7_75t_L     g07223(.A(new_n7479), .B(\a[29] ), .C(new_n7477), .D(new_n7478), .Y(new_n7480));
  NAND2xp33_ASAP7_75t_L     g07224(.A(new_n7478), .B(new_n7479), .Y(new_n7481));
  A2O1A1Ixp33_ASAP7_75t_L   g07225(.A1(\b[19] ), .A2(new_n2931), .B(new_n7481), .C(new_n2697), .Y(new_n7482));
  NAND2xp33_ASAP7_75t_L     g07226(.A(new_n7480), .B(new_n7482), .Y(new_n7483));
  NOR3xp33_ASAP7_75t_L      g07227(.A(new_n7476), .B(new_n7472), .C(new_n7483), .Y(new_n7484));
  AO21x2_ASAP7_75t_L        g07228(.A1(new_n7192), .A2(new_n7189), .B(new_n7088), .Y(new_n7485));
  NAND4xp25_ASAP7_75t_L     g07229(.A(new_n7485), .B(new_n7463), .C(new_n7468), .D(new_n7470), .Y(new_n7486));
  INVx1_ASAP7_75t_L         g07230(.A(new_n7483), .Y(new_n7487));
  AOI21xp33_ASAP7_75t_L     g07231(.A1(new_n7486), .A2(new_n7475), .B(new_n7487), .Y(new_n7488));
  AOI21xp33_ASAP7_75t_L     g07232(.A1(new_n7202), .A2(new_n7203), .B(new_n7204), .Y(new_n7489));
  AO21x2_ASAP7_75t_L        g07233(.A1(new_n7205), .A2(new_n7086), .B(new_n7489), .Y(new_n7490));
  NOR3xp33_ASAP7_75t_L      g07234(.A(new_n7490), .B(new_n7484), .C(new_n7488), .Y(new_n7491));
  NAND3xp33_ASAP7_75t_L     g07235(.A(new_n7487), .B(new_n7475), .C(new_n7486), .Y(new_n7492));
  OAI21xp33_ASAP7_75t_L     g07236(.A1(new_n7472), .A2(new_n7476), .B(new_n7483), .Y(new_n7493));
  AOI21xp33_ASAP7_75t_L     g07237(.A1(new_n7086), .A2(new_n7205), .B(new_n7489), .Y(new_n7494));
  AOI21xp33_ASAP7_75t_L     g07238(.A1(new_n7493), .A2(new_n7492), .B(new_n7494), .Y(new_n7495));
  NAND2xp33_ASAP7_75t_L     g07239(.A(\b[22] ), .B(new_n2386), .Y(new_n7496));
  NAND2xp33_ASAP7_75t_L     g07240(.A(\b[23] ), .B(new_n2232), .Y(new_n7497));
  AOI22xp33_ASAP7_75t_L     g07241(.A1(new_n2228), .A2(\b[24] ), .B1(new_n2226), .B2(new_n2027), .Y(new_n7498));
  NAND4xp25_ASAP7_75t_L     g07242(.A(new_n7498), .B(\a[26] ), .C(new_n7496), .D(new_n7497), .Y(new_n7499));
  NAND2xp33_ASAP7_75t_L     g07243(.A(new_n7497), .B(new_n7498), .Y(new_n7500));
  A2O1A1Ixp33_ASAP7_75t_L   g07244(.A1(\b[22] ), .A2(new_n2386), .B(new_n7500), .C(new_n2223), .Y(new_n7501));
  AND2x2_ASAP7_75t_L        g07245(.A(new_n7499), .B(new_n7501), .Y(new_n7502));
  OAI21xp33_ASAP7_75t_L     g07246(.A1(new_n7495), .A2(new_n7491), .B(new_n7502), .Y(new_n7503));
  NAND3xp33_ASAP7_75t_L     g07247(.A(new_n7493), .B(new_n7494), .C(new_n7492), .Y(new_n7504));
  OAI21xp33_ASAP7_75t_L     g07248(.A1(new_n7488), .A2(new_n7484), .B(new_n7490), .Y(new_n7505));
  NAND2xp33_ASAP7_75t_L     g07249(.A(new_n7499), .B(new_n7501), .Y(new_n7506));
  NAND3xp33_ASAP7_75t_L     g07250(.A(new_n7505), .B(new_n7504), .C(new_n7506), .Y(new_n7507));
  O2A1O1Ixp33_ASAP7_75t_L   g07251(.A1(new_n6934), .A2(new_n6945), .B(new_n7083), .C(new_n7221), .Y(new_n7508));
  OAI211xp5_ASAP7_75t_L     g07252(.A1(new_n7222), .A2(new_n7508), .B(new_n7503), .C(new_n7507), .Y(new_n7509));
  AOI21xp33_ASAP7_75t_L     g07253(.A1(new_n7505), .A2(new_n7504), .B(new_n7506), .Y(new_n7510));
  NOR3xp33_ASAP7_75t_L      g07254(.A(new_n7491), .B(new_n7502), .C(new_n7495), .Y(new_n7511));
  A2O1A1O1Ixp25_ASAP7_75t_L g07255(.A1(new_n6928), .A2(new_n6930), .B(new_n7082), .C(new_n7214), .D(new_n7222), .Y(new_n7512));
  OAI21xp33_ASAP7_75t_L     g07256(.A1(new_n7510), .A2(new_n7511), .B(new_n7512), .Y(new_n7513));
  NOR2xp33_ASAP7_75t_L      g07257(.A(new_n2180), .B(new_n1911), .Y(new_n7514));
  INVx1_ASAP7_75t_L         g07258(.A(new_n7514), .Y(new_n7515));
  NAND2xp33_ASAP7_75t_L     g07259(.A(\b[26] ), .B(new_n1770), .Y(new_n7516));
  AOI22xp33_ASAP7_75t_L     g07260(.A1(new_n1766), .A2(\b[27] ), .B1(new_n1764), .B2(new_n2657), .Y(new_n7517));
  AND4x1_ASAP7_75t_L        g07261(.A(new_n7517), .B(new_n7516), .C(new_n7515), .D(\a[23] ), .Y(new_n7518));
  AOI31xp33_ASAP7_75t_L     g07262(.A1(new_n7517), .A2(new_n7516), .A3(new_n7515), .B(\a[23] ), .Y(new_n7519));
  NOR2xp33_ASAP7_75t_L      g07263(.A(new_n7519), .B(new_n7518), .Y(new_n7520));
  NAND3xp33_ASAP7_75t_L     g07264(.A(new_n7509), .B(new_n7513), .C(new_n7520), .Y(new_n7521));
  NOR3xp33_ASAP7_75t_L      g07265(.A(new_n7512), .B(new_n7511), .C(new_n7510), .Y(new_n7522));
  AOI211xp5_ASAP7_75t_L     g07266(.A1(new_n7503), .A2(new_n7507), .B(new_n7222), .C(new_n7508), .Y(new_n7523));
  INVx1_ASAP7_75t_L         g07267(.A(new_n7520), .Y(new_n7524));
  OAI21xp33_ASAP7_75t_L     g07268(.A1(new_n7523), .A2(new_n7522), .B(new_n7524), .Y(new_n7525));
  AOI21xp33_ASAP7_75t_L     g07269(.A1(new_n7525), .A2(new_n7521), .B(new_n7365), .Y(new_n7526));
  NAND2xp33_ASAP7_75t_L     g07270(.A(new_n6943), .B(new_n7077), .Y(new_n7527));
  A2O1A1Ixp33_ASAP7_75t_L   g07271(.A1(new_n6952), .A2(new_n7527), .B(new_n7225), .C(new_n7236), .Y(new_n7528));
  NAND2xp33_ASAP7_75t_L     g07272(.A(new_n7521), .B(new_n7525), .Y(new_n7529));
  NOR2xp33_ASAP7_75t_L      g07273(.A(new_n7528), .B(new_n7529), .Y(new_n7530));
  NOR3xp33_ASAP7_75t_L      g07274(.A(new_n7530), .B(new_n7526), .C(new_n7364), .Y(new_n7531));
  INVx1_ASAP7_75t_L         g07275(.A(new_n7364), .Y(new_n7532));
  NAND2xp33_ASAP7_75t_L     g07276(.A(new_n7528), .B(new_n7529), .Y(new_n7533));
  NAND3xp33_ASAP7_75t_L     g07277(.A(new_n7365), .B(new_n7521), .C(new_n7525), .Y(new_n7534));
  AOI21xp33_ASAP7_75t_L     g07278(.A1(new_n7533), .A2(new_n7534), .B(new_n7532), .Y(new_n7535));
  NOR2xp33_ASAP7_75t_L      g07279(.A(new_n7535), .B(new_n7531), .Y(new_n7536));
  A2O1A1Ixp33_ASAP7_75t_L   g07280(.A1(new_n7238), .A2(new_n7250), .B(new_n7357), .C(new_n7536), .Y(new_n7537));
  A2O1A1O1Ixp25_ASAP7_75t_L g07281(.A1(new_n6974), .A2(new_n6967), .B(new_n7245), .C(new_n7238), .D(new_n7357), .Y(new_n7538));
  OAI21xp33_ASAP7_75t_L     g07282(.A1(new_n7531), .A2(new_n7535), .B(new_n7538), .Y(new_n7539));
  NAND2xp33_ASAP7_75t_L     g07283(.A(\b[32] ), .B(new_n1103), .Y(new_n7540));
  AOI22xp33_ASAP7_75t_L     g07284(.A1(new_n1113), .A2(\b[33] ), .B1(new_n1110), .B2(new_n3813), .Y(new_n7541));
  NAND2xp33_ASAP7_75t_L     g07285(.A(new_n7540), .B(new_n7541), .Y(new_n7542));
  AOI211xp5_ASAP7_75t_L     g07286(.A1(\b[31] ), .A2(new_n1194), .B(new_n1107), .C(new_n7542), .Y(new_n7543));
  INVx1_ASAP7_75t_L         g07287(.A(new_n7542), .Y(new_n7544));
  O2A1O1Ixp33_ASAP7_75t_L   g07288(.A1(new_n3419), .A2(new_n1195), .B(new_n7544), .C(\a[17] ), .Y(new_n7545));
  NOR2xp33_ASAP7_75t_L      g07289(.A(new_n7543), .B(new_n7545), .Y(new_n7546));
  NAND3xp33_ASAP7_75t_L     g07290(.A(new_n7537), .B(new_n7539), .C(new_n7546), .Y(new_n7547));
  AO21x2_ASAP7_75t_L        g07291(.A1(new_n7539), .A2(new_n7537), .B(new_n7546), .Y(new_n7548));
  AO21x2_ASAP7_75t_L        g07292(.A1(new_n7547), .A2(new_n7548), .B(new_n7356), .Y(new_n7549));
  NAND3xp33_ASAP7_75t_L     g07293(.A(new_n7356), .B(new_n7548), .C(new_n7547), .Y(new_n7550));
  NAND3xp33_ASAP7_75t_L     g07294(.A(new_n7549), .B(new_n7355), .C(new_n7550), .Y(new_n7551));
  AOI21xp33_ASAP7_75t_L     g07295(.A1(new_n7548), .A2(new_n7547), .B(new_n7356), .Y(new_n7552));
  AND3x1_ASAP7_75t_L        g07296(.A(new_n7356), .B(new_n7548), .C(new_n7547), .Y(new_n7553));
  OAI21xp33_ASAP7_75t_L     g07297(.A1(new_n7552), .A2(new_n7553), .B(new_n7354), .Y(new_n7554));
  NAND2xp33_ASAP7_75t_L     g07298(.A(new_n7551), .B(new_n7554), .Y(new_n7555));
  NAND2xp33_ASAP7_75t_L     g07299(.A(new_n7555), .B(new_n7348), .Y(new_n7556));
  NOR3xp33_ASAP7_75t_L      g07300(.A(new_n7553), .B(new_n7354), .C(new_n7552), .Y(new_n7557));
  AOI21xp33_ASAP7_75t_L     g07301(.A1(new_n7549), .A2(new_n7550), .B(new_n7355), .Y(new_n7558));
  NOR2xp33_ASAP7_75t_L      g07302(.A(new_n7558), .B(new_n7557), .Y(new_n7559));
  A2O1A1Ixp33_ASAP7_75t_L   g07303(.A1(new_n7276), .A2(new_n7274), .B(new_n7347), .C(new_n7559), .Y(new_n7560));
  NAND2xp33_ASAP7_75t_L     g07304(.A(\b[38] ), .B(new_n590), .Y(new_n7561));
  AOI22xp33_ASAP7_75t_L     g07305(.A1(new_n600), .A2(\b[39] ), .B1(new_n597), .B2(new_n5174), .Y(new_n7562));
  NAND2xp33_ASAP7_75t_L     g07306(.A(new_n7561), .B(new_n7562), .Y(new_n7563));
  AOI211xp5_ASAP7_75t_L     g07307(.A1(\b[37] ), .A2(new_n674), .B(new_n594), .C(new_n7563), .Y(new_n7564));
  INVx1_ASAP7_75t_L         g07308(.A(new_n7564), .Y(new_n7565));
  A2O1A1Ixp33_ASAP7_75t_L   g07309(.A1(\b[37] ), .A2(new_n674), .B(new_n7563), .C(new_n594), .Y(new_n7566));
  AND2x2_ASAP7_75t_L        g07310(.A(new_n7566), .B(new_n7565), .Y(new_n7567));
  NAND3xp33_ASAP7_75t_L     g07311(.A(new_n7560), .B(new_n7556), .C(new_n7567), .Y(new_n7568));
  AOI221xp5_ASAP7_75t_L     g07312(.A1(new_n7274), .A2(new_n7276), .B1(new_n7551), .B2(new_n7554), .C(new_n7347), .Y(new_n7569));
  NOR2xp33_ASAP7_75t_L      g07313(.A(new_n7555), .B(new_n7348), .Y(new_n7570));
  NAND2xp33_ASAP7_75t_L     g07314(.A(new_n7566), .B(new_n7565), .Y(new_n7571));
  OAI21xp33_ASAP7_75t_L     g07315(.A1(new_n7569), .A2(new_n7570), .B(new_n7571), .Y(new_n7572));
  NOR2xp33_ASAP7_75t_L      g07316(.A(new_n7277), .B(new_n7279), .Y(new_n7573));
  MAJIxp5_ASAP7_75t_L       g07317(.A(new_n7289), .B(new_n7573), .C(new_n7286), .Y(new_n7574));
  NAND3xp33_ASAP7_75t_L     g07318(.A(new_n7574), .B(new_n7572), .C(new_n7568), .Y(new_n7575));
  NAND2xp33_ASAP7_75t_L     g07319(.A(new_n7572), .B(new_n7568), .Y(new_n7576));
  AOI211xp5_ASAP7_75t_L     g07320(.A1(new_n7285), .A2(new_n7283), .B(new_n7277), .C(new_n7279), .Y(new_n7577));
  OAI21xp33_ASAP7_75t_L     g07321(.A1(new_n7577), .A2(new_n7291), .B(new_n7576), .Y(new_n7578));
  AND2x2_ASAP7_75t_L        g07322(.A(new_n7575), .B(new_n7578), .Y(new_n7579));
  NAND2xp33_ASAP7_75t_L     g07323(.A(\b[42] ), .B(new_n451), .Y(new_n7580));
  OAI221xp5_ASAP7_75t_L     g07324(.A1(new_n5666), .A2(new_n529), .B1(new_n482), .B2(new_n5687), .C(new_n7580), .Y(new_n7581));
  AOI21xp33_ASAP7_75t_L     g07325(.A1(new_n480), .A2(\b[40] ), .B(new_n7581), .Y(new_n7582));
  NAND2xp33_ASAP7_75t_L     g07326(.A(\a[8] ), .B(new_n7582), .Y(new_n7583));
  A2O1A1Ixp33_ASAP7_75t_L   g07327(.A1(\b[40] ), .A2(new_n480), .B(new_n7581), .C(new_n445), .Y(new_n7584));
  NAND2xp33_ASAP7_75t_L     g07328(.A(new_n7584), .B(new_n7583), .Y(new_n7585));
  INVx1_ASAP7_75t_L         g07329(.A(new_n7585), .Y(new_n7586));
  NAND2xp33_ASAP7_75t_L     g07330(.A(new_n7586), .B(new_n7579), .Y(new_n7587));
  NAND2xp33_ASAP7_75t_L     g07331(.A(new_n7575), .B(new_n7578), .Y(new_n7588));
  NAND2xp33_ASAP7_75t_L     g07332(.A(new_n7585), .B(new_n7588), .Y(new_n7589));
  OAI21xp33_ASAP7_75t_L     g07333(.A1(new_n7305), .A2(new_n7307), .B(new_n7299), .Y(new_n7590));
  NAND3xp33_ASAP7_75t_L     g07334(.A(new_n7587), .B(new_n7590), .C(new_n7589), .Y(new_n7591));
  NOR2xp33_ASAP7_75t_L      g07335(.A(new_n7585), .B(new_n7588), .Y(new_n7592));
  NOR2xp33_ASAP7_75t_L      g07336(.A(new_n7586), .B(new_n7579), .Y(new_n7593));
  NOR2xp33_ASAP7_75t_L      g07337(.A(new_n6727), .B(new_n6728), .Y(new_n7594));
  MAJx2_ASAP7_75t_L         g07338(.A(new_n6736), .B(new_n6729), .C(new_n7594), .Y(new_n7595));
  A2O1A1O1Ixp25_ASAP7_75t_L g07339(.A1(new_n7306), .A2(new_n7595), .B(new_n7016), .C(new_n7300), .D(new_n7298), .Y(new_n7596));
  OAI21xp33_ASAP7_75t_L     g07340(.A1(new_n7592), .A2(new_n7593), .B(new_n7596), .Y(new_n7597));
  NAND2xp33_ASAP7_75t_L     g07341(.A(\b[43] ), .B(new_n366), .Y(new_n7598));
  NAND2xp33_ASAP7_75t_L     g07342(.A(\b[44] ), .B(new_n334), .Y(new_n7599));
  AOI22xp33_ASAP7_75t_L     g07343(.A1(new_n345), .A2(\b[45] ), .B1(new_n342), .B2(new_n6764), .Y(new_n7600));
  AND4x1_ASAP7_75t_L        g07344(.A(new_n7600), .B(new_n7599), .C(new_n7598), .D(\a[5] ), .Y(new_n7601));
  AOI31xp33_ASAP7_75t_L     g07345(.A1(new_n7600), .A2(new_n7599), .A3(new_n7598), .B(\a[5] ), .Y(new_n7602));
  NOR2xp33_ASAP7_75t_L      g07346(.A(new_n7602), .B(new_n7601), .Y(new_n7603));
  AOI21xp33_ASAP7_75t_L     g07347(.A1(new_n7597), .A2(new_n7591), .B(new_n7603), .Y(new_n7604));
  NAND3xp33_ASAP7_75t_L     g07348(.A(new_n7597), .B(new_n7591), .C(new_n7603), .Y(new_n7605));
  INVx1_ASAP7_75t_L         g07349(.A(new_n7605), .Y(new_n7606));
  NOR3xp33_ASAP7_75t_L      g07350(.A(new_n7346), .B(new_n7604), .C(new_n7606), .Y(new_n7607));
  INVx1_ASAP7_75t_L         g07351(.A(new_n7604), .Y(new_n7608));
  AOI221xp5_ASAP7_75t_L     g07352(.A1(new_n7313), .A2(new_n7052), .B1(new_n7605), .B2(new_n7608), .C(new_n7312), .Y(new_n7609));
  OAI21xp33_ASAP7_75t_L     g07353(.A1(new_n7607), .A2(new_n7609), .B(new_n7344), .Y(new_n7610));
  NOR3xp33_ASAP7_75t_L      g07354(.A(new_n7609), .B(new_n7607), .C(new_n7344), .Y(new_n7611));
  INVx1_ASAP7_75t_L         g07355(.A(new_n7611), .Y(new_n7612));
  NAND2xp33_ASAP7_75t_L     g07356(.A(new_n7610), .B(new_n7612), .Y(new_n7613));
  O2A1O1Ixp33_ASAP7_75t_L   g07357(.A1(new_n7314), .A2(new_n7326), .B(new_n7330), .C(new_n7613), .Y(new_n7614));
  MAJIxp5_ASAP7_75t_L       g07358(.A(new_n7328), .B(new_n7314), .C(new_n7326), .Y(new_n7615));
  AOI21xp33_ASAP7_75t_L     g07359(.A1(new_n7612), .A2(new_n7610), .B(new_n7615), .Y(new_n7616));
  NOR2xp33_ASAP7_75t_L      g07360(.A(new_n7616), .B(new_n7614), .Y(\f[48] ));
  INVx1_ASAP7_75t_L         g07361(.A(new_n7615), .Y(new_n7618));
  OAI21xp33_ASAP7_75t_L     g07362(.A1(new_n7526), .A2(new_n7530), .B(new_n7364), .Y(new_n7619));
  A2O1A1O1Ixp25_ASAP7_75t_L g07363(.A1(new_n7238), .A2(new_n7250), .B(new_n7357), .C(new_n7619), .D(new_n7531), .Y(new_n7620));
  NAND2xp33_ASAP7_75t_L     g07364(.A(new_n7513), .B(new_n7509), .Y(new_n7621));
  NOR2xp33_ASAP7_75t_L      g07365(.A(new_n7520), .B(new_n7621), .Y(new_n7622));
  NOR2xp33_ASAP7_75t_L      g07366(.A(new_n2477), .B(new_n1911), .Y(new_n7623));
  NAND2xp33_ASAP7_75t_L     g07367(.A(\b[27] ), .B(new_n1770), .Y(new_n7624));
  OAI221xp5_ASAP7_75t_L     g07368(.A1(new_n1772), .A2(new_n2852), .B1(new_n1771), .B2(new_n5212), .C(new_n7624), .Y(new_n7625));
  OR3x1_ASAP7_75t_L         g07369(.A(new_n7625), .B(new_n1761), .C(new_n7623), .Y(new_n7626));
  A2O1A1Ixp33_ASAP7_75t_L   g07370(.A1(\b[26] ), .A2(new_n1910), .B(new_n7625), .C(new_n1761), .Y(new_n7627));
  AND2x2_ASAP7_75t_L        g07371(.A(new_n7627), .B(new_n7626), .Y(new_n7628));
  NOR2xp33_ASAP7_75t_L      g07372(.A(new_n7440), .B(new_n7443), .Y(new_n7629));
  NAND2xp33_ASAP7_75t_L     g07373(.A(new_n7439), .B(new_n7629), .Y(new_n7630));
  A2O1A1Ixp33_ASAP7_75t_L   g07374(.A1(new_n7447), .A2(new_n7448), .B(new_n7446), .C(new_n7630), .Y(new_n7631));
  NAND2xp33_ASAP7_75t_L     g07375(.A(\b[11] ), .B(new_n4780), .Y(new_n7632));
  NAND2xp33_ASAP7_75t_L     g07376(.A(\b[12] ), .B(new_n4548), .Y(new_n7633));
  AOI22xp33_ASAP7_75t_L     g07377(.A1(new_n4544), .A2(\b[13] ), .B1(new_n4542), .B2(new_n800), .Y(new_n7634));
  AND4x1_ASAP7_75t_L        g07378(.A(new_n7634), .B(new_n7633), .C(new_n7632), .D(\a[38] ), .Y(new_n7635));
  AOI31xp33_ASAP7_75t_L     g07379(.A1(new_n7634), .A2(new_n7633), .A3(new_n7632), .B(\a[38] ), .Y(new_n7636));
  NOR2xp33_ASAP7_75t_L      g07380(.A(new_n7636), .B(new_n7635), .Y(new_n7637));
  A2O1A1O1Ixp25_ASAP7_75t_L g07381(.A1(new_n7150), .A2(new_n7162), .B(new_n7383), .C(new_n7434), .D(new_n7430), .Y(new_n7638));
  INVx1_ASAP7_75t_L         g07382(.A(new_n7389), .Y(new_n7639));
  NOR3xp33_ASAP7_75t_L      g07383(.A(new_n7131), .B(new_n7639), .C(new_n7384), .Y(new_n7640));
  NOR2xp33_ASAP7_75t_L      g07384(.A(new_n278), .B(new_n7115), .Y(new_n7641));
  NOR2xp33_ASAP7_75t_L      g07385(.A(new_n299), .B(new_n7392), .Y(new_n7642));
  OAI32xp33_ASAP7_75t_L     g07386(.A1(new_n325), .A2(new_n327), .A3(new_n7117), .B1(new_n7118), .B2(new_n323), .Y(new_n7643));
  NOR4xp25_ASAP7_75t_L      g07387(.A(new_n7643), .B(new_n6816), .C(new_n7641), .D(new_n7642), .Y(new_n7644));
  NOR3xp33_ASAP7_75t_L      g07388(.A(new_n7643), .B(new_n7642), .C(new_n7641), .Y(new_n7645));
  NOR2xp33_ASAP7_75t_L      g07389(.A(\a[47] ), .B(new_n7645), .Y(new_n7646));
  NAND2xp33_ASAP7_75t_L     g07390(.A(new_n7387), .B(new_n7386), .Y(new_n7647));
  XNOR2x2_ASAP7_75t_L       g07391(.A(\a[49] ), .B(\a[48] ), .Y(new_n7648));
  NOR2xp33_ASAP7_75t_L      g07392(.A(new_n7648), .B(new_n7647), .Y(new_n7649));
  NAND2xp33_ASAP7_75t_L     g07393(.A(\b[0] ), .B(new_n7649), .Y(new_n7650));
  INVx1_ASAP7_75t_L         g07394(.A(\a[49] ), .Y(new_n7651));
  NAND2xp33_ASAP7_75t_L     g07395(.A(\a[50] ), .B(new_n7651), .Y(new_n7652));
  INVx1_ASAP7_75t_L         g07396(.A(\a[50] ), .Y(new_n7653));
  NAND2xp33_ASAP7_75t_L     g07397(.A(\a[49] ), .B(new_n7653), .Y(new_n7654));
  AND2x2_ASAP7_75t_L        g07398(.A(new_n7652), .B(new_n7654), .Y(new_n7655));
  NOR2xp33_ASAP7_75t_L      g07399(.A(new_n7388), .B(new_n7655), .Y(new_n7656));
  NAND2xp33_ASAP7_75t_L     g07400(.A(new_n271), .B(new_n7656), .Y(new_n7657));
  NAND2xp33_ASAP7_75t_L     g07401(.A(new_n7654), .B(new_n7652), .Y(new_n7658));
  NOR2xp33_ASAP7_75t_L      g07402(.A(new_n7658), .B(new_n7388), .Y(new_n7659));
  NAND2xp33_ASAP7_75t_L     g07403(.A(\b[1] ), .B(new_n7659), .Y(new_n7660));
  NAND3xp33_ASAP7_75t_L     g07404(.A(new_n7657), .B(new_n7660), .C(new_n7650), .Y(new_n7661));
  NAND3xp33_ASAP7_75t_L     g07405(.A(new_n7661), .B(new_n7389), .C(\a[50] ), .Y(new_n7662));
  NAND2xp33_ASAP7_75t_L     g07406(.A(\a[50] ), .B(new_n7389), .Y(new_n7663));
  AND3x1_ASAP7_75t_L        g07407(.A(new_n7657), .B(new_n7660), .C(new_n7650), .Y(new_n7664));
  NAND2xp33_ASAP7_75t_L     g07408(.A(new_n7663), .B(new_n7664), .Y(new_n7665));
  AO211x2_ASAP7_75t_L       g07409(.A1(new_n7665), .A2(new_n7662), .B(new_n7644), .C(new_n7646), .Y(new_n7666));
  XNOR2x2_ASAP7_75t_L       g07410(.A(new_n7663), .B(new_n7661), .Y(new_n7667));
  OAI21xp33_ASAP7_75t_L     g07411(.A1(new_n7644), .A2(new_n7646), .B(new_n7667), .Y(new_n7668));
  OAI211xp5_ASAP7_75t_L     g07412(.A1(new_n7640), .A2(new_n7407), .B(new_n7666), .C(new_n7668), .Y(new_n7669));
  INVx1_ASAP7_75t_L         g07413(.A(new_n7640), .Y(new_n7670));
  NOR3xp33_ASAP7_75t_L      g07414(.A(new_n7646), .B(new_n7667), .C(new_n7644), .Y(new_n7671));
  OA21x2_ASAP7_75t_L        g07415(.A1(new_n7644), .A2(new_n7646), .B(new_n7667), .Y(new_n7672));
  OAI211xp5_ASAP7_75t_L     g07416(.A1(new_n7671), .A2(new_n7672), .B(new_n7398), .C(new_n7670), .Y(new_n7673));
  NAND2xp33_ASAP7_75t_L     g07417(.A(\b[6] ), .B(new_n5992), .Y(new_n7674));
  AOI32xp33_ASAP7_75t_L     g07418(.A1(new_n424), .A2(new_n426), .A3(new_n5999), .B1(new_n6002), .B2(\b[7] ), .Y(new_n7675));
  OAI211xp5_ASAP7_75t_L     g07419(.A1(new_n353), .A2(new_n6309), .B(new_n7675), .C(new_n7674), .Y(new_n7676));
  NOR2xp33_ASAP7_75t_L      g07420(.A(new_n5996), .B(new_n7676), .Y(new_n7677));
  INVx1_ASAP7_75t_L         g07421(.A(new_n7677), .Y(new_n7678));
  NAND2xp33_ASAP7_75t_L     g07422(.A(new_n5996), .B(new_n7676), .Y(new_n7679));
  NAND4xp25_ASAP7_75t_L     g07423(.A(new_n7673), .B(new_n7669), .C(new_n7678), .D(new_n7679), .Y(new_n7680));
  AO22x1_ASAP7_75t_L        g07424(.A1(new_n7679), .A2(new_n7678), .B1(new_n7669), .B2(new_n7673), .Y(new_n7681));
  NAND2xp33_ASAP7_75t_L     g07425(.A(new_n7680), .B(new_n7681), .Y(new_n7682));
  AOI211xp5_ASAP7_75t_L     g07426(.A1(new_n7405), .A2(new_n7403), .B(new_n7407), .C(new_n7408), .Y(new_n7683));
  AO21x2_ASAP7_75t_L        g07427(.A1(new_n7416), .A2(new_n7427), .B(new_n7683), .Y(new_n7684));
  NOR2xp33_ASAP7_75t_L      g07428(.A(new_n7684), .B(new_n7682), .Y(new_n7685));
  AOI21xp33_ASAP7_75t_L     g07429(.A1(new_n7427), .A2(new_n7416), .B(new_n7683), .Y(new_n7686));
  AOI21xp33_ASAP7_75t_L     g07430(.A1(new_n7681), .A2(new_n7680), .B(new_n7686), .Y(new_n7687));
  NAND2xp33_ASAP7_75t_L     g07431(.A(\b[8] ), .B(new_n5526), .Y(new_n7688));
  NAND2xp33_ASAP7_75t_L     g07432(.A(\b[9] ), .B(new_n5240), .Y(new_n7689));
  AOI22xp33_ASAP7_75t_L     g07433(.A1(new_n5249), .A2(\b[10] ), .B1(new_n5247), .B2(new_n852), .Y(new_n7690));
  NAND4xp25_ASAP7_75t_L     g07434(.A(new_n7690), .B(\a[41] ), .C(new_n7688), .D(new_n7689), .Y(new_n7691));
  INVx1_ASAP7_75t_L         g07435(.A(new_n7691), .Y(new_n7692));
  AOI31xp33_ASAP7_75t_L     g07436(.A1(new_n7690), .A2(new_n7689), .A3(new_n7688), .B(\a[41] ), .Y(new_n7693));
  NOR2xp33_ASAP7_75t_L      g07437(.A(new_n7693), .B(new_n7692), .Y(new_n7694));
  OAI21xp33_ASAP7_75t_L     g07438(.A1(new_n7687), .A2(new_n7685), .B(new_n7694), .Y(new_n7695));
  NAND3xp33_ASAP7_75t_L     g07439(.A(new_n7686), .B(new_n7681), .C(new_n7680), .Y(new_n7696));
  A2O1A1Ixp33_ASAP7_75t_L   g07440(.A1(new_n7416), .A2(new_n7427), .B(new_n7683), .C(new_n7682), .Y(new_n7697));
  INVx1_ASAP7_75t_L         g07441(.A(new_n7693), .Y(new_n7698));
  NAND2xp33_ASAP7_75t_L     g07442(.A(new_n7691), .B(new_n7698), .Y(new_n7699));
  NAND3xp33_ASAP7_75t_L     g07443(.A(new_n7697), .B(new_n7699), .C(new_n7696), .Y(new_n7700));
  NAND3xp33_ASAP7_75t_L     g07444(.A(new_n7638), .B(new_n7700), .C(new_n7695), .Y(new_n7701));
  AO21x2_ASAP7_75t_L        g07445(.A1(new_n7700), .A2(new_n7695), .B(new_n7638), .Y(new_n7702));
  NAND3xp33_ASAP7_75t_L     g07446(.A(new_n7702), .B(new_n7701), .C(new_n7637), .Y(new_n7703));
  INVx1_ASAP7_75t_L         g07447(.A(new_n7637), .Y(new_n7704));
  AND3x1_ASAP7_75t_L        g07448(.A(new_n7638), .B(new_n7700), .C(new_n7695), .Y(new_n7705));
  AOI21xp33_ASAP7_75t_L     g07449(.A1(new_n7700), .A2(new_n7695), .B(new_n7638), .Y(new_n7706));
  OAI21xp33_ASAP7_75t_L     g07450(.A1(new_n7706), .A2(new_n7705), .B(new_n7704), .Y(new_n7707));
  NAND3xp33_ASAP7_75t_L     g07451(.A(new_n7631), .B(new_n7703), .C(new_n7707), .Y(new_n7708));
  NAND2xp33_ASAP7_75t_L     g07452(.A(new_n7437), .B(new_n7432), .Y(new_n7709));
  NOR2xp33_ASAP7_75t_L      g07453(.A(new_n7382), .B(new_n7709), .Y(new_n7710));
  O2A1O1Ixp33_ASAP7_75t_L   g07454(.A1(new_n7438), .A2(new_n7444), .B(new_n7374), .C(new_n7710), .Y(new_n7711));
  NAND2xp33_ASAP7_75t_L     g07455(.A(new_n7703), .B(new_n7707), .Y(new_n7712));
  NAND2xp33_ASAP7_75t_L     g07456(.A(new_n7712), .B(new_n7711), .Y(new_n7713));
  NAND2xp33_ASAP7_75t_L     g07457(.A(\b[14] ), .B(new_n4111), .Y(new_n7714));
  NAND2xp33_ASAP7_75t_L     g07458(.A(\b[15] ), .B(new_n3874), .Y(new_n7715));
  AOI22xp33_ASAP7_75t_L     g07459(.A1(new_n3884), .A2(\b[16] ), .B1(new_n3881), .B2(new_n1058), .Y(new_n7716));
  NAND4xp25_ASAP7_75t_L     g07460(.A(new_n7716), .B(\a[35] ), .C(new_n7714), .D(new_n7715), .Y(new_n7717));
  NAND2xp33_ASAP7_75t_L     g07461(.A(new_n7715), .B(new_n7716), .Y(new_n7718));
  A2O1A1Ixp33_ASAP7_75t_L   g07462(.A1(\b[14] ), .A2(new_n4111), .B(new_n7718), .C(new_n3878), .Y(new_n7719));
  AND2x2_ASAP7_75t_L        g07463(.A(new_n7717), .B(new_n7719), .Y(new_n7720));
  NAND3xp33_ASAP7_75t_L     g07464(.A(new_n7708), .B(new_n7713), .C(new_n7720), .Y(new_n7721));
  O2A1O1Ixp33_ASAP7_75t_L   g07465(.A1(new_n7382), .A2(new_n7709), .B(new_n7445), .C(new_n7712), .Y(new_n7722));
  AOI21xp33_ASAP7_75t_L     g07466(.A1(new_n7707), .A2(new_n7703), .B(new_n7631), .Y(new_n7723));
  NAND2xp33_ASAP7_75t_L     g07467(.A(new_n7717), .B(new_n7719), .Y(new_n7724));
  OAI21xp33_ASAP7_75t_L     g07468(.A1(new_n7722), .A2(new_n7723), .B(new_n7724), .Y(new_n7725));
  NOR3xp33_ASAP7_75t_L      g07469(.A(new_n7451), .B(new_n7453), .C(new_n7452), .Y(new_n7726));
  A2O1A1O1Ixp25_ASAP7_75t_L g07470(.A1(new_n7187), .A2(new_n7186), .B(new_n7456), .C(new_n7454), .D(new_n7726), .Y(new_n7727));
  NAND3xp33_ASAP7_75t_L     g07471(.A(new_n7727), .B(new_n7725), .C(new_n7721), .Y(new_n7728));
  AO21x2_ASAP7_75t_L        g07472(.A1(new_n7721), .A2(new_n7725), .B(new_n7727), .Y(new_n7729));
  NAND2xp33_ASAP7_75t_L     g07473(.A(\b[17] ), .B(new_n3491), .Y(new_n7730));
  NAND2xp33_ASAP7_75t_L     g07474(.A(\b[18] ), .B(new_n3260), .Y(new_n7731));
  AOI22xp33_ASAP7_75t_L     g07475(.A1(new_n3256), .A2(\b[19] ), .B1(new_n3254), .B2(new_n1499), .Y(new_n7732));
  NAND4xp25_ASAP7_75t_L     g07476(.A(new_n7732), .B(\a[32] ), .C(new_n7730), .D(new_n7731), .Y(new_n7733));
  OAI221xp5_ASAP7_75t_L     g07477(.A1(new_n3262), .A2(new_n1493), .B1(new_n3261), .B2(new_n2793), .C(new_n7731), .Y(new_n7734));
  A2O1A1Ixp33_ASAP7_75t_L   g07478(.A1(\b[17] ), .A2(new_n3491), .B(new_n7734), .C(new_n3251), .Y(new_n7735));
  AND2x2_ASAP7_75t_L        g07479(.A(new_n7733), .B(new_n7735), .Y(new_n7736));
  NAND3xp33_ASAP7_75t_L     g07480(.A(new_n7729), .B(new_n7728), .C(new_n7736), .Y(new_n7737));
  AND3x1_ASAP7_75t_L        g07481(.A(new_n7727), .B(new_n7725), .C(new_n7721), .Y(new_n7738));
  AOI21xp33_ASAP7_75t_L     g07482(.A1(new_n7725), .A2(new_n7721), .B(new_n7727), .Y(new_n7739));
  NAND2xp33_ASAP7_75t_L     g07483(.A(new_n7733), .B(new_n7735), .Y(new_n7740));
  OAI21xp33_ASAP7_75t_L     g07484(.A1(new_n7739), .A2(new_n7738), .B(new_n7740), .Y(new_n7741));
  NOR2xp33_ASAP7_75t_L      g07485(.A(new_n7465), .B(new_n7466), .Y(new_n7742));
  NAND2xp33_ASAP7_75t_L     g07486(.A(new_n7467), .B(new_n7742), .Y(new_n7743));
  AND4x1_ASAP7_75t_L        g07487(.A(new_n7475), .B(new_n7743), .C(new_n7737), .D(new_n7741), .Y(new_n7744));
  MAJIxp5_ASAP7_75t_L       g07488(.A(new_n7471), .B(new_n7467), .C(new_n7742), .Y(new_n7745));
  AOI21xp33_ASAP7_75t_L     g07489(.A1(new_n7741), .A2(new_n7737), .B(new_n7745), .Y(new_n7746));
  NOR2xp33_ASAP7_75t_L      g07490(.A(new_n1594), .B(new_n2932), .Y(new_n7747));
  NAND2xp33_ASAP7_75t_L     g07491(.A(\b[21] ), .B(new_n2706), .Y(new_n7748));
  OAI221xp5_ASAP7_75t_L     g07492(.A1(new_n2708), .A2(new_n1857), .B1(new_n2707), .B2(new_n1863), .C(new_n7748), .Y(new_n7749));
  OR3x1_ASAP7_75t_L         g07493(.A(new_n7749), .B(new_n2697), .C(new_n7747), .Y(new_n7750));
  A2O1A1Ixp33_ASAP7_75t_L   g07494(.A1(\b[20] ), .A2(new_n2931), .B(new_n7749), .C(new_n2697), .Y(new_n7751));
  NAND2xp33_ASAP7_75t_L     g07495(.A(new_n7751), .B(new_n7750), .Y(new_n7752));
  NOR3xp33_ASAP7_75t_L      g07496(.A(new_n7744), .B(new_n7746), .C(new_n7752), .Y(new_n7753));
  NAND3xp33_ASAP7_75t_L     g07497(.A(new_n7745), .B(new_n7741), .C(new_n7737), .Y(new_n7754));
  NAND2xp33_ASAP7_75t_L     g07498(.A(new_n7737), .B(new_n7741), .Y(new_n7755));
  INVx1_ASAP7_75t_L         g07499(.A(new_n7743), .Y(new_n7756));
  A2O1A1Ixp33_ASAP7_75t_L   g07500(.A1(new_n7469), .A2(new_n7471), .B(new_n7756), .C(new_n7755), .Y(new_n7757));
  AND2x2_ASAP7_75t_L        g07501(.A(new_n7751), .B(new_n7750), .Y(new_n7758));
  AOI21xp33_ASAP7_75t_L     g07502(.A1(new_n7757), .A2(new_n7754), .B(new_n7758), .Y(new_n7759));
  NAND2xp33_ASAP7_75t_L     g07503(.A(new_n7475), .B(new_n7486), .Y(new_n7760));
  MAJIxp5_ASAP7_75t_L       g07504(.A(new_n7494), .B(new_n7487), .C(new_n7760), .Y(new_n7761));
  NOR3xp33_ASAP7_75t_L      g07505(.A(new_n7761), .B(new_n7759), .C(new_n7753), .Y(new_n7762));
  NAND3xp33_ASAP7_75t_L     g07506(.A(new_n7757), .B(new_n7754), .C(new_n7758), .Y(new_n7763));
  OAI21xp33_ASAP7_75t_L     g07507(.A1(new_n7746), .A2(new_n7744), .B(new_n7752), .Y(new_n7764));
  NOR2xp33_ASAP7_75t_L      g07508(.A(new_n7472), .B(new_n7476), .Y(new_n7765));
  NAND2xp33_ASAP7_75t_L     g07509(.A(new_n7483), .B(new_n7765), .Y(new_n7766));
  AOI22xp33_ASAP7_75t_L     g07510(.A1(new_n7763), .A2(new_n7764), .B1(new_n7766), .B2(new_n7505), .Y(new_n7767));
  NAND2xp33_ASAP7_75t_L     g07511(.A(\b[23] ), .B(new_n2386), .Y(new_n7768));
  NAND2xp33_ASAP7_75t_L     g07512(.A(\b[24] ), .B(new_n2232), .Y(new_n7769));
  AOI22xp33_ASAP7_75t_L     g07513(.A1(new_n2228), .A2(\b[25] ), .B1(new_n2226), .B2(new_n2188), .Y(new_n7770));
  AND4x1_ASAP7_75t_L        g07514(.A(new_n7770), .B(new_n7769), .C(new_n7768), .D(\a[26] ), .Y(new_n7771));
  AOI31xp33_ASAP7_75t_L     g07515(.A1(new_n7770), .A2(new_n7769), .A3(new_n7768), .B(\a[26] ), .Y(new_n7772));
  OR2x4_ASAP7_75t_L         g07516(.A(new_n7772), .B(new_n7771), .Y(new_n7773));
  NOR3xp33_ASAP7_75t_L      g07517(.A(new_n7773), .B(new_n7767), .C(new_n7762), .Y(new_n7774));
  NAND4xp25_ASAP7_75t_L     g07518(.A(new_n7505), .B(new_n7766), .C(new_n7764), .D(new_n7763), .Y(new_n7775));
  OAI21xp33_ASAP7_75t_L     g07519(.A1(new_n7759), .A2(new_n7753), .B(new_n7761), .Y(new_n7776));
  NOR2xp33_ASAP7_75t_L      g07520(.A(new_n7772), .B(new_n7771), .Y(new_n7777));
  AOI21xp33_ASAP7_75t_L     g07521(.A1(new_n7775), .A2(new_n7776), .B(new_n7777), .Y(new_n7778));
  A2O1A1Ixp33_ASAP7_75t_L   g07522(.A1(new_n6930), .A2(new_n6928), .B(new_n7082), .C(new_n7214), .Y(new_n7779));
  A2O1A1Ixp33_ASAP7_75t_L   g07523(.A1(new_n7779), .A2(new_n7218), .B(new_n7510), .C(new_n7507), .Y(new_n7780));
  OAI21xp33_ASAP7_75t_L     g07524(.A1(new_n7774), .A2(new_n7778), .B(new_n7780), .Y(new_n7781));
  NAND3xp33_ASAP7_75t_L     g07525(.A(new_n7775), .B(new_n7776), .C(new_n7777), .Y(new_n7782));
  OAI21xp33_ASAP7_75t_L     g07526(.A1(new_n7762), .A2(new_n7767), .B(new_n7773), .Y(new_n7783));
  A2O1A1O1Ixp25_ASAP7_75t_L g07527(.A1(new_n7214), .A2(new_n7084), .B(new_n7222), .C(new_n7503), .D(new_n7511), .Y(new_n7784));
  NAND3xp33_ASAP7_75t_L     g07528(.A(new_n7784), .B(new_n7783), .C(new_n7782), .Y(new_n7785));
  AOI21xp33_ASAP7_75t_L     g07529(.A1(new_n7785), .A2(new_n7781), .B(new_n7628), .Y(new_n7786));
  NAND2xp33_ASAP7_75t_L     g07530(.A(new_n7627), .B(new_n7626), .Y(new_n7787));
  AOI21xp33_ASAP7_75t_L     g07531(.A1(new_n7783), .A2(new_n7782), .B(new_n7784), .Y(new_n7788));
  NOR3xp33_ASAP7_75t_L      g07532(.A(new_n7780), .B(new_n7778), .C(new_n7774), .Y(new_n7789));
  NOR3xp33_ASAP7_75t_L      g07533(.A(new_n7789), .B(new_n7788), .C(new_n7787), .Y(new_n7790));
  NOR2xp33_ASAP7_75t_L      g07534(.A(new_n7786), .B(new_n7790), .Y(new_n7791));
  A2O1A1Ixp33_ASAP7_75t_L   g07535(.A1(new_n7529), .A2(new_n7528), .B(new_n7622), .C(new_n7791), .Y(new_n7792));
  AOI21xp33_ASAP7_75t_L     g07536(.A1(new_n7529), .A2(new_n7528), .B(new_n7622), .Y(new_n7793));
  OAI21xp33_ASAP7_75t_L     g07537(.A1(new_n7788), .A2(new_n7789), .B(new_n7787), .Y(new_n7794));
  NAND3xp33_ASAP7_75t_L     g07538(.A(new_n7785), .B(new_n7781), .C(new_n7628), .Y(new_n7795));
  NAND2xp33_ASAP7_75t_L     g07539(.A(new_n7795), .B(new_n7794), .Y(new_n7796));
  NAND2xp33_ASAP7_75t_L     g07540(.A(new_n7796), .B(new_n7793), .Y(new_n7797));
  NAND2xp33_ASAP7_75t_L     g07541(.A(\b[29] ), .B(new_n1548), .Y(new_n7798));
  NAND2xp33_ASAP7_75t_L     g07542(.A(\b[30] ), .B(new_n1410), .Y(new_n7799));
  AOI22xp33_ASAP7_75t_L     g07543(.A1(new_n1406), .A2(\b[31] ), .B1(new_n1404), .B2(new_n3426), .Y(new_n7800));
  AND4x1_ASAP7_75t_L        g07544(.A(new_n7800), .B(new_n7799), .C(new_n7798), .D(\a[20] ), .Y(new_n7801));
  AOI31xp33_ASAP7_75t_L     g07545(.A1(new_n7800), .A2(new_n7799), .A3(new_n7798), .B(\a[20] ), .Y(new_n7802));
  NOR2xp33_ASAP7_75t_L      g07546(.A(new_n7802), .B(new_n7801), .Y(new_n7803));
  AOI21xp33_ASAP7_75t_L     g07547(.A1(new_n7792), .A2(new_n7797), .B(new_n7803), .Y(new_n7804));
  O2A1O1Ixp33_ASAP7_75t_L   g07548(.A1(new_n7621), .A2(new_n7520), .B(new_n7533), .C(new_n7796), .Y(new_n7805));
  NAND3xp33_ASAP7_75t_L     g07549(.A(new_n7509), .B(new_n7513), .C(new_n7524), .Y(new_n7806));
  A2O1A1Ixp33_ASAP7_75t_L   g07550(.A1(new_n7521), .A2(new_n7525), .B(new_n7365), .C(new_n7806), .Y(new_n7807));
  NOR2xp33_ASAP7_75t_L      g07551(.A(new_n7807), .B(new_n7791), .Y(new_n7808));
  INVx1_ASAP7_75t_L         g07552(.A(new_n7803), .Y(new_n7809));
  NOR3xp33_ASAP7_75t_L      g07553(.A(new_n7805), .B(new_n7808), .C(new_n7809), .Y(new_n7810));
  OAI21xp33_ASAP7_75t_L     g07554(.A1(new_n7804), .A2(new_n7810), .B(new_n7620), .Y(new_n7811));
  NAND3xp33_ASAP7_75t_L     g07555(.A(new_n7533), .B(new_n7534), .C(new_n7532), .Y(new_n7812));
  OAI21xp33_ASAP7_75t_L     g07556(.A1(new_n7535), .A2(new_n7538), .B(new_n7812), .Y(new_n7813));
  OAI21xp33_ASAP7_75t_L     g07557(.A1(new_n7808), .A2(new_n7805), .B(new_n7809), .Y(new_n7814));
  NAND3xp33_ASAP7_75t_L     g07558(.A(new_n7792), .B(new_n7803), .C(new_n7797), .Y(new_n7815));
  NAND3xp33_ASAP7_75t_L     g07559(.A(new_n7813), .B(new_n7814), .C(new_n7815), .Y(new_n7816));
  NAND2xp33_ASAP7_75t_L     g07560(.A(\b[32] ), .B(new_n1194), .Y(new_n7817));
  NAND2xp33_ASAP7_75t_L     g07561(.A(\b[33] ), .B(new_n1103), .Y(new_n7818));
  AOI22xp33_ASAP7_75t_L     g07562(.A1(new_n1113), .A2(\b[34] ), .B1(new_n1110), .B2(new_n3833), .Y(new_n7819));
  NAND4xp25_ASAP7_75t_L     g07563(.A(new_n7819), .B(\a[17] ), .C(new_n7817), .D(new_n7818), .Y(new_n7820));
  NAND2xp33_ASAP7_75t_L     g07564(.A(new_n7818), .B(new_n7819), .Y(new_n7821));
  A2O1A1Ixp33_ASAP7_75t_L   g07565(.A1(\b[32] ), .A2(new_n1194), .B(new_n7821), .C(new_n1107), .Y(new_n7822));
  NAND2xp33_ASAP7_75t_L     g07566(.A(new_n7820), .B(new_n7822), .Y(new_n7823));
  INVx1_ASAP7_75t_L         g07567(.A(new_n7823), .Y(new_n7824));
  NAND3xp33_ASAP7_75t_L     g07568(.A(new_n7824), .B(new_n7816), .C(new_n7811), .Y(new_n7825));
  AOI21xp33_ASAP7_75t_L     g07569(.A1(new_n7815), .A2(new_n7814), .B(new_n7813), .Y(new_n7826));
  NOR3xp33_ASAP7_75t_L      g07570(.A(new_n7620), .B(new_n7804), .C(new_n7810), .Y(new_n7827));
  OAI21xp33_ASAP7_75t_L     g07571(.A1(new_n7826), .A2(new_n7827), .B(new_n7823), .Y(new_n7828));
  OAI211xp5_ASAP7_75t_L     g07572(.A1(new_n7543), .A2(new_n7545), .B(new_n7537), .C(new_n7539), .Y(new_n7829));
  NAND4xp25_ASAP7_75t_L     g07573(.A(new_n7549), .B(new_n7829), .C(new_n7828), .D(new_n7825), .Y(new_n7830));
  NAND2xp33_ASAP7_75t_L     g07574(.A(new_n7825), .B(new_n7828), .Y(new_n7831));
  NAND2xp33_ASAP7_75t_L     g07575(.A(new_n7539), .B(new_n7537), .Y(new_n7832));
  MAJIxp5_ASAP7_75t_L       g07576(.A(new_n7356), .B(new_n7546), .C(new_n7832), .Y(new_n7833));
  NAND2xp33_ASAP7_75t_L     g07577(.A(new_n7833), .B(new_n7831), .Y(new_n7834));
  NAND2xp33_ASAP7_75t_L     g07578(.A(\b[36] ), .B(new_n817), .Y(new_n7835));
  NOR2xp33_ASAP7_75t_L      g07579(.A(new_n4701), .B(new_n912), .Y(new_n7836));
  AOI21xp33_ASAP7_75t_L     g07580(.A1(new_n4709), .A2(new_n823), .B(new_n7836), .Y(new_n7837));
  NAND2xp33_ASAP7_75t_L     g07581(.A(new_n7835), .B(new_n7837), .Y(new_n7838));
  AOI211xp5_ASAP7_75t_L     g07582(.A1(\b[35] ), .A2(new_n908), .B(new_n813), .C(new_n7838), .Y(new_n7839));
  AND2x2_ASAP7_75t_L        g07583(.A(new_n7835), .B(new_n7837), .Y(new_n7840));
  O2A1O1Ixp33_ASAP7_75t_L   g07584(.A1(new_n4053), .A2(new_n909), .B(new_n7840), .C(\a[14] ), .Y(new_n7841));
  NOR2xp33_ASAP7_75t_L      g07585(.A(new_n7839), .B(new_n7841), .Y(new_n7842));
  NAND3xp33_ASAP7_75t_L     g07586(.A(new_n7842), .B(new_n7830), .C(new_n7834), .Y(new_n7843));
  AO21x2_ASAP7_75t_L        g07587(.A1(new_n7830), .A2(new_n7834), .B(new_n7842), .Y(new_n7844));
  A2O1A1O1Ixp25_ASAP7_75t_L g07588(.A1(new_n7276), .A2(new_n7274), .B(new_n7347), .C(new_n7554), .D(new_n7557), .Y(new_n7845));
  NAND3xp33_ASAP7_75t_L     g07589(.A(new_n7845), .B(new_n7844), .C(new_n7843), .Y(new_n7846));
  AO21x2_ASAP7_75t_L        g07590(.A1(new_n7843), .A2(new_n7844), .B(new_n7845), .Y(new_n7847));
  NAND2xp33_ASAP7_75t_L     g07591(.A(\b[38] ), .B(new_n674), .Y(new_n7848));
  NAND2xp33_ASAP7_75t_L     g07592(.A(\b[39] ), .B(new_n590), .Y(new_n7849));
  AOI22xp33_ASAP7_75t_L     g07593(.A1(new_n600), .A2(\b[40] ), .B1(new_n597), .B2(new_n5194), .Y(new_n7850));
  NAND4xp25_ASAP7_75t_L     g07594(.A(new_n7850), .B(\a[11] ), .C(new_n7848), .D(new_n7849), .Y(new_n7851));
  NAND2xp33_ASAP7_75t_L     g07595(.A(new_n7849), .B(new_n7850), .Y(new_n7852));
  A2O1A1Ixp33_ASAP7_75t_L   g07596(.A1(\b[38] ), .A2(new_n674), .B(new_n7852), .C(new_n594), .Y(new_n7853));
  AND2x2_ASAP7_75t_L        g07597(.A(new_n7851), .B(new_n7853), .Y(new_n7854));
  NAND3xp33_ASAP7_75t_L     g07598(.A(new_n7847), .B(new_n7846), .C(new_n7854), .Y(new_n7855));
  AND3x1_ASAP7_75t_L        g07599(.A(new_n7845), .B(new_n7844), .C(new_n7843), .Y(new_n7856));
  AOI21xp33_ASAP7_75t_L     g07600(.A1(new_n7844), .A2(new_n7843), .B(new_n7845), .Y(new_n7857));
  NAND2xp33_ASAP7_75t_L     g07601(.A(new_n7851), .B(new_n7853), .Y(new_n7858));
  OAI21xp33_ASAP7_75t_L     g07602(.A1(new_n7857), .A2(new_n7856), .B(new_n7858), .Y(new_n7859));
  NAND3xp33_ASAP7_75t_L     g07603(.A(new_n7560), .B(new_n7556), .C(new_n7571), .Y(new_n7860));
  NAND4xp25_ASAP7_75t_L     g07604(.A(new_n7578), .B(new_n7860), .C(new_n7859), .D(new_n7855), .Y(new_n7861));
  NAND2xp33_ASAP7_75t_L     g07605(.A(new_n7855), .B(new_n7859), .Y(new_n7862));
  NAND2xp33_ASAP7_75t_L     g07606(.A(new_n7556), .B(new_n7560), .Y(new_n7863));
  MAJIxp5_ASAP7_75t_L       g07607(.A(new_n7574), .B(new_n7863), .C(new_n7567), .Y(new_n7864));
  NAND2xp33_ASAP7_75t_L     g07608(.A(new_n7862), .B(new_n7864), .Y(new_n7865));
  NOR2xp33_ASAP7_75t_L      g07609(.A(new_n5666), .B(new_n481), .Y(new_n7866));
  INVx1_ASAP7_75t_L         g07610(.A(new_n7866), .Y(new_n7867));
  NAND2xp33_ASAP7_75t_L     g07611(.A(\b[42] ), .B(new_n441), .Y(new_n7868));
  AOI22xp33_ASAP7_75t_L     g07612(.A1(new_n451), .A2(\b[43] ), .B1(new_n448), .B2(new_n6202), .Y(new_n7869));
  AND4x1_ASAP7_75t_L        g07613(.A(new_n7869), .B(new_n7868), .C(new_n7867), .D(\a[8] ), .Y(new_n7870));
  AOI31xp33_ASAP7_75t_L     g07614(.A1(new_n7869), .A2(new_n7868), .A3(new_n7867), .B(\a[8] ), .Y(new_n7871));
  NOR2xp33_ASAP7_75t_L      g07615(.A(new_n7871), .B(new_n7870), .Y(new_n7872));
  NAND3xp33_ASAP7_75t_L     g07616(.A(new_n7861), .B(new_n7865), .C(new_n7872), .Y(new_n7873));
  NOR2xp33_ASAP7_75t_L      g07617(.A(new_n7862), .B(new_n7864), .Y(new_n7874));
  NOR3xp33_ASAP7_75t_L      g07618(.A(new_n7856), .B(new_n7857), .C(new_n7858), .Y(new_n7875));
  AOI21xp33_ASAP7_75t_L     g07619(.A1(new_n7847), .A2(new_n7846), .B(new_n7854), .Y(new_n7876));
  NOR2xp33_ASAP7_75t_L      g07620(.A(new_n7876), .B(new_n7875), .Y(new_n7877));
  AOI21xp33_ASAP7_75t_L     g07621(.A1(new_n7578), .A2(new_n7860), .B(new_n7877), .Y(new_n7878));
  INVx1_ASAP7_75t_L         g07622(.A(new_n7872), .Y(new_n7879));
  OAI21xp33_ASAP7_75t_L     g07623(.A1(new_n7874), .A2(new_n7878), .B(new_n7879), .Y(new_n7880));
  NOR2xp33_ASAP7_75t_L      g07624(.A(new_n7586), .B(new_n7588), .Y(new_n7881));
  O2A1O1Ixp33_ASAP7_75t_L   g07625(.A1(new_n7592), .A2(new_n7593), .B(new_n7590), .C(new_n7881), .Y(new_n7882));
  NAND3xp33_ASAP7_75t_L     g07626(.A(new_n7882), .B(new_n7880), .C(new_n7873), .Y(new_n7883));
  NAND2xp33_ASAP7_75t_L     g07627(.A(new_n7873), .B(new_n7880), .Y(new_n7884));
  MAJIxp5_ASAP7_75t_L       g07628(.A(new_n7596), .B(new_n7586), .C(new_n7588), .Y(new_n7885));
  NAND2xp33_ASAP7_75t_L     g07629(.A(new_n7885), .B(new_n7884), .Y(new_n7886));
  INVx1_ASAP7_75t_L         g07630(.A(new_n7041), .Y(new_n7887));
  NAND2xp33_ASAP7_75t_L     g07631(.A(\b[46] ), .B(new_n345), .Y(new_n7888));
  OAI221xp5_ASAP7_75t_L     g07632(.A1(new_n6756), .A2(new_n406), .B1(new_n367), .B2(new_n7887), .C(new_n7888), .Y(new_n7889));
  AOI21xp33_ASAP7_75t_L     g07633(.A1(new_n366), .A2(\b[44] ), .B(new_n7889), .Y(new_n7890));
  NAND2xp33_ASAP7_75t_L     g07634(.A(\a[5] ), .B(new_n7890), .Y(new_n7891));
  A2O1A1Ixp33_ASAP7_75t_L   g07635(.A1(\b[44] ), .A2(new_n366), .B(new_n7889), .C(new_n339), .Y(new_n7892));
  NAND2xp33_ASAP7_75t_L     g07636(.A(new_n7892), .B(new_n7891), .Y(new_n7893));
  INVx1_ASAP7_75t_L         g07637(.A(new_n7893), .Y(new_n7894));
  NAND3xp33_ASAP7_75t_L     g07638(.A(new_n7883), .B(new_n7886), .C(new_n7894), .Y(new_n7895));
  INVx1_ASAP7_75t_L         g07639(.A(new_n7895), .Y(new_n7896));
  AOI21xp33_ASAP7_75t_L     g07640(.A1(new_n7883), .A2(new_n7886), .B(new_n7894), .Y(new_n7897));
  A2O1A1O1Ixp25_ASAP7_75t_L g07641(.A1(new_n7313), .A2(new_n7052), .B(new_n7312), .C(new_n7605), .D(new_n7604), .Y(new_n7898));
  INVx1_ASAP7_75t_L         g07642(.A(new_n7898), .Y(new_n7899));
  NOR3xp33_ASAP7_75t_L      g07643(.A(new_n7899), .B(new_n7896), .C(new_n7897), .Y(new_n7900));
  INVx1_ASAP7_75t_L         g07644(.A(new_n7897), .Y(new_n7901));
  AOI21xp33_ASAP7_75t_L     g07645(.A1(new_n7901), .A2(new_n7895), .B(new_n7898), .Y(new_n7902));
  NAND2xp33_ASAP7_75t_L     g07646(.A(\b[47] ), .B(new_n291), .Y(new_n7903));
  NAND2xp33_ASAP7_75t_L     g07647(.A(\b[48] ), .B(new_n380), .Y(new_n7904));
  INVx1_ASAP7_75t_L         g07648(.A(new_n7334), .Y(new_n7905));
  NOR2xp33_ASAP7_75t_L      g07649(.A(\b[48] ), .B(\b[49] ), .Y(new_n7906));
  INVx1_ASAP7_75t_L         g07650(.A(\b[49] ), .Y(new_n7907));
  NOR2xp33_ASAP7_75t_L      g07651(.A(new_n7333), .B(new_n7907), .Y(new_n7908));
  NOR2xp33_ASAP7_75t_L      g07652(.A(new_n7906), .B(new_n7908), .Y(new_n7909));
  INVx1_ASAP7_75t_L         g07653(.A(new_n7909), .Y(new_n7910));
  A2O1A1O1Ixp25_ASAP7_75t_L g07654(.A1(new_n7331), .A2(new_n7319), .B(new_n7332), .C(new_n7905), .D(new_n7910), .Y(new_n7911));
  A2O1A1Ixp33_ASAP7_75t_L   g07655(.A1(new_n7319), .A2(new_n7331), .B(new_n7332), .C(new_n7905), .Y(new_n7912));
  NOR2xp33_ASAP7_75t_L      g07656(.A(new_n7909), .B(new_n7912), .Y(new_n7913));
  NOR2xp33_ASAP7_75t_L      g07657(.A(new_n7911), .B(new_n7913), .Y(new_n7914));
  AOI22xp33_ASAP7_75t_L     g07658(.A1(new_n272), .A2(\b[49] ), .B1(new_n269), .B2(new_n7914), .Y(new_n7915));
  NAND4xp25_ASAP7_75t_L     g07659(.A(new_n7915), .B(\a[2] ), .C(new_n7903), .D(new_n7904), .Y(new_n7916));
  NAND2xp33_ASAP7_75t_L     g07660(.A(new_n7904), .B(new_n7915), .Y(new_n7917));
  A2O1A1Ixp33_ASAP7_75t_L   g07661(.A1(\b[47] ), .A2(new_n291), .B(new_n7917), .C(new_n265), .Y(new_n7918));
  AND2x2_ASAP7_75t_L        g07662(.A(new_n7916), .B(new_n7918), .Y(new_n7919));
  OAI21xp33_ASAP7_75t_L     g07663(.A1(new_n7902), .A2(new_n7900), .B(new_n7919), .Y(new_n7920));
  NOR3xp33_ASAP7_75t_L      g07664(.A(new_n7900), .B(new_n7902), .C(new_n7919), .Y(new_n7921));
  INVx1_ASAP7_75t_L         g07665(.A(new_n7921), .Y(new_n7922));
  NAND2xp33_ASAP7_75t_L     g07666(.A(new_n7920), .B(new_n7922), .Y(new_n7923));
  O2A1O1Ixp33_ASAP7_75t_L   g07667(.A1(new_n7618), .A2(new_n7613), .B(new_n7612), .C(new_n7923), .Y(new_n7924));
  AOI211xp5_ASAP7_75t_L     g07668(.A1(new_n7922), .A2(new_n7920), .B(new_n7611), .C(new_n7614), .Y(new_n7925));
  NOR2xp33_ASAP7_75t_L      g07669(.A(new_n7924), .B(new_n7925), .Y(\f[49] ));
  NAND2xp33_ASAP7_75t_L     g07670(.A(\b[45] ), .B(new_n366), .Y(new_n7927));
  NAND2xp33_ASAP7_75t_L     g07671(.A(\b[46] ), .B(new_n334), .Y(new_n7928));
  AOI22xp33_ASAP7_75t_L     g07672(.A1(new_n345), .A2(\b[47] ), .B1(new_n342), .B2(new_n7323), .Y(new_n7929));
  AND4x1_ASAP7_75t_L        g07673(.A(new_n7929), .B(new_n7928), .C(new_n7927), .D(\a[5] ), .Y(new_n7930));
  AOI31xp33_ASAP7_75t_L     g07674(.A1(new_n7929), .A2(new_n7928), .A3(new_n7927), .B(\a[5] ), .Y(new_n7931));
  NOR2xp33_ASAP7_75t_L      g07675(.A(new_n7931), .B(new_n7930), .Y(new_n7932));
  NOR2xp33_ASAP7_75t_L      g07676(.A(new_n7874), .B(new_n7878), .Y(new_n7933));
  MAJIxp5_ASAP7_75t_L       g07677(.A(new_n7885), .B(new_n7933), .C(new_n7879), .Y(new_n7934));
  OAI21xp33_ASAP7_75t_L     g07678(.A1(new_n7810), .A2(new_n7620), .B(new_n7814), .Y(new_n7935));
  NAND2xp33_ASAP7_75t_L     g07679(.A(\b[30] ), .B(new_n1548), .Y(new_n7936));
  NAND2xp33_ASAP7_75t_L     g07680(.A(\b[31] ), .B(new_n1410), .Y(new_n7937));
  AOI22xp33_ASAP7_75t_L     g07681(.A1(new_n1406), .A2(\b[32] ), .B1(new_n1404), .B2(new_n3450), .Y(new_n7938));
  AND4x1_ASAP7_75t_L        g07682(.A(new_n7938), .B(new_n7937), .C(new_n7936), .D(\a[20] ), .Y(new_n7939));
  AOI31xp33_ASAP7_75t_L     g07683(.A1(new_n7938), .A2(new_n7937), .A3(new_n7936), .B(\a[20] ), .Y(new_n7940));
  NOR2xp33_ASAP7_75t_L      g07684(.A(new_n7940), .B(new_n7939), .Y(new_n7941));
  NOR3xp33_ASAP7_75t_L      g07685(.A(new_n7789), .B(new_n7788), .C(new_n7628), .Y(new_n7942));
  AOI21xp33_ASAP7_75t_L     g07686(.A1(new_n7796), .A2(new_n7807), .B(new_n7942), .Y(new_n7943));
  NAND2xp33_ASAP7_75t_L     g07687(.A(\b[27] ), .B(new_n1910), .Y(new_n7944));
  NAND2xp33_ASAP7_75t_L     g07688(.A(\b[28] ), .B(new_n1770), .Y(new_n7945));
  AOI22xp33_ASAP7_75t_L     g07689(.A1(new_n1766), .A2(\b[29] ), .B1(new_n1764), .B2(new_n5472), .Y(new_n7946));
  NAND4xp25_ASAP7_75t_L     g07690(.A(new_n7946), .B(\a[23] ), .C(new_n7944), .D(new_n7945), .Y(new_n7947));
  AOI31xp33_ASAP7_75t_L     g07691(.A1(new_n7946), .A2(new_n7945), .A3(new_n7944), .B(\a[23] ), .Y(new_n7948));
  INVx1_ASAP7_75t_L         g07692(.A(new_n7948), .Y(new_n7949));
  AND2x2_ASAP7_75t_L        g07693(.A(new_n7947), .B(new_n7949), .Y(new_n7950));
  NOR2xp33_ASAP7_75t_L      g07694(.A(new_n7762), .B(new_n7767), .Y(new_n7951));
  MAJIxp5_ASAP7_75t_L       g07695(.A(new_n7780), .B(new_n7773), .C(new_n7951), .Y(new_n7952));
  NAND2xp33_ASAP7_75t_L     g07696(.A(\b[24] ), .B(new_n2386), .Y(new_n7953));
  NAND2xp33_ASAP7_75t_L     g07697(.A(\b[25] ), .B(new_n2232), .Y(new_n7954));
  AOI22xp33_ASAP7_75t_L     g07698(.A1(new_n2228), .A2(\b[26] ), .B1(new_n2226), .B2(new_n2888), .Y(new_n7955));
  NAND4xp25_ASAP7_75t_L     g07699(.A(new_n7955), .B(\a[26] ), .C(new_n7953), .D(new_n7954), .Y(new_n7956));
  AOI31xp33_ASAP7_75t_L     g07700(.A1(new_n7955), .A2(new_n7954), .A3(new_n7953), .B(\a[26] ), .Y(new_n7957));
  INVx1_ASAP7_75t_L         g07701(.A(new_n7957), .Y(new_n7958));
  NAND2xp33_ASAP7_75t_L     g07702(.A(new_n7956), .B(new_n7958), .Y(new_n7959));
  NOR2xp33_ASAP7_75t_L      g07703(.A(new_n7487), .B(new_n7760), .Y(new_n7960));
  O2A1O1Ixp33_ASAP7_75t_L   g07704(.A1(new_n7484), .A2(new_n7488), .B(new_n7490), .C(new_n7960), .Y(new_n7961));
  NOR3xp33_ASAP7_75t_L      g07705(.A(new_n7744), .B(new_n7746), .C(new_n7758), .Y(new_n7962));
  INVx1_ASAP7_75t_L         g07706(.A(new_n7962), .Y(new_n7963));
  A2O1A1Ixp33_ASAP7_75t_L   g07707(.A1(new_n7764), .A2(new_n7763), .B(new_n7961), .C(new_n7963), .Y(new_n7964));
  NOR3xp33_ASAP7_75t_L      g07708(.A(new_n7738), .B(new_n7739), .C(new_n7736), .Y(new_n7965));
  A2O1A1O1Ixp25_ASAP7_75t_L g07709(.A1(new_n7471), .A2(new_n7469), .B(new_n7756), .C(new_n7755), .D(new_n7965), .Y(new_n7966));
  NAND3xp33_ASAP7_75t_L     g07710(.A(new_n7708), .B(new_n7713), .C(new_n7724), .Y(new_n7967));
  A2O1A1Ixp33_ASAP7_75t_L   g07711(.A1(new_n7725), .A2(new_n7721), .B(new_n7727), .C(new_n7967), .Y(new_n7968));
  NAND2xp33_ASAP7_75t_L     g07712(.A(\b[16] ), .B(new_n3874), .Y(new_n7969));
  OAI221xp5_ASAP7_75t_L     g07713(.A1(new_n4115), .A2(new_n1244), .B1(new_n4114), .B2(new_n1251), .C(new_n7969), .Y(new_n7970));
  INVx1_ASAP7_75t_L         g07714(.A(new_n7970), .Y(new_n7971));
  OAI211xp5_ASAP7_75t_L     g07715(.A1(new_n952), .A2(new_n4986), .B(new_n7971), .C(\a[35] ), .Y(new_n7972));
  A2O1A1Ixp33_ASAP7_75t_L   g07716(.A1(\b[15] ), .A2(new_n4111), .B(new_n7970), .C(new_n3878), .Y(new_n7973));
  NAND2xp33_ASAP7_75t_L     g07717(.A(new_n7973), .B(new_n7972), .Y(new_n7974));
  NAND2xp33_ASAP7_75t_L     g07718(.A(new_n7448), .B(new_n7447), .Y(new_n7975));
  AOI21xp33_ASAP7_75t_L     g07719(.A1(new_n7702), .A2(new_n7701), .B(new_n7637), .Y(new_n7976));
  A2O1A1O1Ixp25_ASAP7_75t_L g07720(.A1(new_n7374), .A2(new_n7975), .B(new_n7710), .C(new_n7703), .D(new_n7976), .Y(new_n7977));
  INVx1_ASAP7_75t_L         g07721(.A(new_n7679), .Y(new_n7978));
  OAI211xp5_ASAP7_75t_L     g07722(.A1(new_n7677), .A2(new_n7978), .B(new_n7673), .C(new_n7669), .Y(new_n7979));
  INVx1_ASAP7_75t_L         g07723(.A(new_n7979), .Y(new_n7980));
  NOR2xp33_ASAP7_75t_L      g07724(.A(new_n382), .B(new_n6309), .Y(new_n7981));
  NAND2xp33_ASAP7_75t_L     g07725(.A(\b[7] ), .B(new_n5992), .Y(new_n7982));
  OAI221xp5_ASAP7_75t_L     g07726(.A1(new_n6312), .A2(new_n503), .B1(new_n6311), .B2(new_n509), .C(new_n7982), .Y(new_n7983));
  NOR3xp33_ASAP7_75t_L      g07727(.A(new_n7983), .B(new_n7981), .C(new_n5996), .Y(new_n7984));
  OA21x2_ASAP7_75t_L        g07728(.A1(new_n7981), .A2(new_n7983), .B(new_n5996), .Y(new_n7985));
  O2A1O1Ixp33_ASAP7_75t_L   g07729(.A1(new_n7640), .A2(new_n7407), .B(new_n7666), .C(new_n7672), .Y(new_n7986));
  NAND2xp33_ASAP7_75t_L     g07730(.A(\b[4] ), .B(new_n6812), .Y(new_n7987));
  OAI221xp5_ASAP7_75t_L     g07731(.A1(new_n7118), .A2(new_n353), .B1(new_n7117), .B2(new_n359), .C(new_n7987), .Y(new_n7988));
  AOI211xp5_ASAP7_75t_L     g07732(.A1(\b[3] ), .A2(new_n7124), .B(new_n6816), .C(new_n7988), .Y(new_n7989));
  INVx1_ASAP7_75t_L         g07733(.A(new_n7989), .Y(new_n7990));
  A2O1A1Ixp33_ASAP7_75t_L   g07734(.A1(\b[3] ), .A2(new_n7124), .B(new_n7988), .C(new_n6816), .Y(new_n7991));
  INVx1_ASAP7_75t_L         g07735(.A(new_n7648), .Y(new_n7992));
  NOR3xp33_ASAP7_75t_L      g07736(.A(new_n7655), .B(new_n7992), .C(new_n7647), .Y(new_n7993));
  INVx1_ASAP7_75t_L         g07737(.A(new_n7993), .Y(new_n7994));
  NOR2xp33_ASAP7_75t_L      g07738(.A(new_n258), .B(new_n7994), .Y(new_n7995));
  NAND2xp33_ASAP7_75t_L     g07739(.A(new_n7658), .B(new_n7647), .Y(new_n7996));
  NAND2xp33_ASAP7_75t_L     g07740(.A(new_n7647), .B(new_n7655), .Y(new_n7997));
  NAND2xp33_ASAP7_75t_L     g07741(.A(\b[1] ), .B(new_n7649), .Y(new_n7998));
  OAI221xp5_ASAP7_75t_L     g07742(.A1(new_n7996), .A2(new_n283), .B1(new_n278), .B2(new_n7997), .C(new_n7998), .Y(new_n7999));
  NOR2xp33_ASAP7_75t_L      g07743(.A(new_n7999), .B(new_n7995), .Y(new_n8000));
  A2O1A1Ixp33_ASAP7_75t_L   g07744(.A1(new_n7639), .A2(new_n7664), .B(new_n7653), .C(new_n8000), .Y(new_n8001));
  O2A1O1Ixp33_ASAP7_75t_L   g07745(.A1(new_n258), .A2(new_n7388), .B(new_n7664), .C(new_n7653), .Y(new_n8002));
  A2O1A1Ixp33_ASAP7_75t_L   g07746(.A1(\b[0] ), .A2(new_n7993), .B(new_n7999), .C(new_n8002), .Y(new_n8003));
  NAND4xp25_ASAP7_75t_L     g07747(.A(new_n7990), .B(new_n8003), .C(new_n8001), .D(new_n7991), .Y(new_n8004));
  INVx1_ASAP7_75t_L         g07748(.A(new_n7991), .Y(new_n8005));
  INVx1_ASAP7_75t_L         g07749(.A(new_n8001), .Y(new_n8006));
  A2O1A1Ixp33_ASAP7_75t_L   g07750(.A1(\b[0] ), .A2(new_n7647), .B(new_n7661), .C(\a[50] ), .Y(new_n8007));
  INVx1_ASAP7_75t_L         g07751(.A(new_n7999), .Y(new_n8008));
  O2A1O1Ixp33_ASAP7_75t_L   g07752(.A1(new_n7994), .A2(new_n258), .B(new_n8008), .C(new_n8007), .Y(new_n8009));
  OAI22xp33_ASAP7_75t_L     g07753(.A1(new_n8006), .A2(new_n8009), .B1(new_n7989), .B2(new_n8005), .Y(new_n8010));
  AOI21xp33_ASAP7_75t_L     g07754(.A1(new_n8010), .A2(new_n8004), .B(new_n7986), .Y(new_n8011));
  A2O1A1Ixp33_ASAP7_75t_L   g07755(.A1(new_n7398), .A2(new_n7670), .B(new_n7671), .C(new_n7668), .Y(new_n8012));
  NAND2xp33_ASAP7_75t_L     g07756(.A(new_n8004), .B(new_n8010), .Y(new_n8013));
  NOR2xp33_ASAP7_75t_L      g07757(.A(new_n8013), .B(new_n8012), .Y(new_n8014));
  OAI22xp33_ASAP7_75t_L     g07758(.A1(new_n8011), .A2(new_n8014), .B1(new_n7984), .B2(new_n7985), .Y(new_n8015));
  INVx1_ASAP7_75t_L         g07759(.A(new_n7984), .Y(new_n8016));
  A2O1A1Ixp33_ASAP7_75t_L   g07760(.A1(\b[6] ), .A2(new_n6308), .B(new_n7983), .C(new_n5996), .Y(new_n8017));
  NAND2xp33_ASAP7_75t_L     g07761(.A(new_n8013), .B(new_n8012), .Y(new_n8018));
  NAND3xp33_ASAP7_75t_L     g07762(.A(new_n7986), .B(new_n8004), .C(new_n8010), .Y(new_n8019));
  NAND4xp25_ASAP7_75t_L     g07763(.A(new_n8019), .B(new_n8016), .C(new_n8018), .D(new_n8017), .Y(new_n8020));
  AND2x2_ASAP7_75t_L        g07764(.A(new_n8020), .B(new_n8015), .Y(new_n8021));
  A2O1A1Ixp33_ASAP7_75t_L   g07765(.A1(new_n7684), .A2(new_n7682), .B(new_n7980), .C(new_n8021), .Y(new_n8022));
  O2A1O1Ixp33_ASAP7_75t_L   g07766(.A1(new_n7683), .A2(new_n7429), .B(new_n7682), .C(new_n7980), .Y(new_n8023));
  NAND2xp33_ASAP7_75t_L     g07767(.A(new_n8020), .B(new_n8015), .Y(new_n8024));
  NAND2xp33_ASAP7_75t_L     g07768(.A(new_n8024), .B(new_n8023), .Y(new_n8025));
  NOR2xp33_ASAP7_75t_L      g07769(.A(new_n559), .B(new_n5521), .Y(new_n8026));
  NAND2xp33_ASAP7_75t_L     g07770(.A(\b[10] ), .B(new_n5240), .Y(new_n8027));
  OAI221xp5_ASAP7_75t_L     g07771(.A1(new_n5253), .A2(new_n695), .B1(new_n5252), .B2(new_n701), .C(new_n8027), .Y(new_n8028));
  OR3x1_ASAP7_75t_L         g07772(.A(new_n8028), .B(new_n5244), .C(new_n8026), .Y(new_n8029));
  A2O1A1Ixp33_ASAP7_75t_L   g07773(.A1(\b[9] ), .A2(new_n5526), .B(new_n8028), .C(new_n5244), .Y(new_n8030));
  AND2x2_ASAP7_75t_L        g07774(.A(new_n8030), .B(new_n8029), .Y(new_n8031));
  NAND3xp33_ASAP7_75t_L     g07775(.A(new_n8031), .B(new_n8022), .C(new_n8025), .Y(new_n8032));
  A2O1A1O1Ixp25_ASAP7_75t_L g07776(.A1(new_n7681), .A2(new_n7680), .B(new_n7686), .C(new_n7979), .D(new_n8024), .Y(new_n8033));
  A2O1A1Ixp33_ASAP7_75t_L   g07777(.A1(new_n7681), .A2(new_n7680), .B(new_n7686), .C(new_n7979), .Y(new_n8034));
  NOR2xp33_ASAP7_75t_L      g07778(.A(new_n8034), .B(new_n8021), .Y(new_n8035));
  NAND2xp33_ASAP7_75t_L     g07779(.A(new_n8030), .B(new_n8029), .Y(new_n8036));
  OAI21xp33_ASAP7_75t_L     g07780(.A1(new_n8033), .A2(new_n8035), .B(new_n8036), .Y(new_n8037));
  AOI21xp33_ASAP7_75t_L     g07781(.A1(new_n7697), .A2(new_n7696), .B(new_n7699), .Y(new_n8038));
  OAI21xp33_ASAP7_75t_L     g07782(.A1(new_n8038), .A2(new_n7638), .B(new_n7700), .Y(new_n8039));
  NAND3xp33_ASAP7_75t_L     g07783(.A(new_n8039), .B(new_n8037), .C(new_n8032), .Y(new_n8040));
  NOR3xp33_ASAP7_75t_L      g07784(.A(new_n8035), .B(new_n8033), .C(new_n8036), .Y(new_n8041));
  AOI21xp33_ASAP7_75t_L     g07785(.A1(new_n8022), .A2(new_n8025), .B(new_n8031), .Y(new_n8042));
  A2O1A1Ixp33_ASAP7_75t_L   g07786(.A1(new_n7442), .A2(new_n7434), .B(new_n7430), .C(new_n7695), .Y(new_n8043));
  OAI211xp5_ASAP7_75t_L     g07787(.A1(new_n8041), .A2(new_n8042), .B(new_n7700), .C(new_n8043), .Y(new_n8044));
  NAND2xp33_ASAP7_75t_L     g07788(.A(\b[12] ), .B(new_n4780), .Y(new_n8045));
  NAND2xp33_ASAP7_75t_L     g07789(.A(\b[13] ), .B(new_n4548), .Y(new_n8046));
  AOI32xp33_ASAP7_75t_L     g07790(.A1(new_n877), .A2(new_n874), .A3(new_n4542), .B1(\b[14] ), .B2(new_n4544), .Y(new_n8047));
  AND4x1_ASAP7_75t_L        g07791(.A(new_n8047), .B(new_n8046), .C(new_n8045), .D(\a[38] ), .Y(new_n8048));
  AOI31xp33_ASAP7_75t_L     g07792(.A1(new_n8047), .A2(new_n8046), .A3(new_n8045), .B(\a[38] ), .Y(new_n8049));
  NOR2xp33_ASAP7_75t_L      g07793(.A(new_n8049), .B(new_n8048), .Y(new_n8050));
  NAND3xp33_ASAP7_75t_L     g07794(.A(new_n8044), .B(new_n8040), .C(new_n8050), .Y(new_n8051));
  AOI211xp5_ASAP7_75t_L     g07795(.A1(new_n8043), .A2(new_n7700), .B(new_n8041), .C(new_n8042), .Y(new_n8052));
  AOI21xp33_ASAP7_75t_L     g07796(.A1(new_n8037), .A2(new_n8032), .B(new_n8039), .Y(new_n8053));
  INVx1_ASAP7_75t_L         g07797(.A(new_n8050), .Y(new_n8054));
  OAI21xp33_ASAP7_75t_L     g07798(.A1(new_n8053), .A2(new_n8052), .B(new_n8054), .Y(new_n8055));
  AOI21xp33_ASAP7_75t_L     g07799(.A1(new_n8055), .A2(new_n8051), .B(new_n7977), .Y(new_n8056));
  INVx1_ASAP7_75t_L         g07800(.A(new_n7703), .Y(new_n8057));
  A2O1A1Ixp33_ASAP7_75t_L   g07801(.A1(new_n7445), .A2(new_n7630), .B(new_n8057), .C(new_n7707), .Y(new_n8058));
  NAND2xp33_ASAP7_75t_L     g07802(.A(new_n8051), .B(new_n8055), .Y(new_n8059));
  NOR2xp33_ASAP7_75t_L      g07803(.A(new_n8059), .B(new_n8058), .Y(new_n8060));
  OAI21xp33_ASAP7_75t_L     g07804(.A1(new_n8056), .A2(new_n8060), .B(new_n7974), .Y(new_n8061));
  AND2x2_ASAP7_75t_L        g07805(.A(new_n7973), .B(new_n7972), .Y(new_n8062));
  NAND2xp33_ASAP7_75t_L     g07806(.A(new_n8059), .B(new_n8058), .Y(new_n8063));
  NAND3xp33_ASAP7_75t_L     g07807(.A(new_n7977), .B(new_n8051), .C(new_n8055), .Y(new_n8064));
  NAND3xp33_ASAP7_75t_L     g07808(.A(new_n8062), .B(new_n8063), .C(new_n8064), .Y(new_n8065));
  NAND3xp33_ASAP7_75t_L     g07809(.A(new_n7968), .B(new_n8061), .C(new_n8065), .Y(new_n8066));
  NOR3xp33_ASAP7_75t_L      g07810(.A(new_n7723), .B(new_n7722), .C(new_n7724), .Y(new_n8067));
  AOI21xp33_ASAP7_75t_L     g07811(.A1(new_n7708), .A2(new_n7713), .B(new_n7720), .Y(new_n8068));
  NOR2xp33_ASAP7_75t_L      g07812(.A(new_n8068), .B(new_n8067), .Y(new_n8069));
  AOI21xp33_ASAP7_75t_L     g07813(.A1(new_n8063), .A2(new_n8064), .B(new_n8062), .Y(new_n8070));
  NOR3xp33_ASAP7_75t_L      g07814(.A(new_n8060), .B(new_n8056), .C(new_n7974), .Y(new_n8071));
  OAI221xp5_ASAP7_75t_L     g07815(.A1(new_n8071), .A2(new_n8070), .B1(new_n7727), .B2(new_n8069), .C(new_n7967), .Y(new_n8072));
  NAND2xp33_ASAP7_75t_L     g07816(.A(\b[18] ), .B(new_n3491), .Y(new_n8073));
  NOR2xp33_ASAP7_75t_L      g07817(.A(new_n1493), .B(new_n3248), .Y(new_n8074));
  AOI221xp5_ASAP7_75t_L     g07818(.A1(new_n3256), .A2(\b[20] ), .B1(new_n3254), .B2(new_n1600), .C(new_n8074), .Y(new_n8075));
  AND3x1_ASAP7_75t_L        g07819(.A(new_n8075), .B(new_n8073), .C(\a[32] ), .Y(new_n8076));
  O2A1O1Ixp33_ASAP7_75t_L   g07820(.A1(new_n1356), .A2(new_n3492), .B(new_n8075), .C(\a[32] ), .Y(new_n8077));
  NOR2xp33_ASAP7_75t_L      g07821(.A(new_n8077), .B(new_n8076), .Y(new_n8078));
  AO21x2_ASAP7_75t_L        g07822(.A1(new_n8066), .A2(new_n8072), .B(new_n8078), .Y(new_n8079));
  NAND3xp33_ASAP7_75t_L     g07823(.A(new_n8072), .B(new_n8066), .C(new_n8078), .Y(new_n8080));
  NAND2xp33_ASAP7_75t_L     g07824(.A(new_n8080), .B(new_n8079), .Y(new_n8081));
  NAND2xp33_ASAP7_75t_L     g07825(.A(new_n8081), .B(new_n7966), .Y(new_n8082));
  MAJx2_ASAP7_75t_L         g07826(.A(new_n7471), .B(new_n7467), .C(new_n7742), .Y(new_n8083));
  AOI21xp33_ASAP7_75t_L     g07827(.A1(new_n8072), .A2(new_n8066), .B(new_n8078), .Y(new_n8084));
  AND3x1_ASAP7_75t_L        g07828(.A(new_n8072), .B(new_n8066), .C(new_n8078), .Y(new_n8085));
  NOR2xp33_ASAP7_75t_L      g07829(.A(new_n8084), .B(new_n8085), .Y(new_n8086));
  A2O1A1Ixp33_ASAP7_75t_L   g07830(.A1(new_n8083), .A2(new_n7755), .B(new_n7965), .C(new_n8086), .Y(new_n8087));
  NAND2xp33_ASAP7_75t_L     g07831(.A(\b[22] ), .B(new_n2706), .Y(new_n8088));
  OAI221xp5_ASAP7_75t_L     g07832(.A1(new_n2708), .A2(new_n1995), .B1(new_n2707), .B2(new_n4860), .C(new_n8088), .Y(new_n8089));
  AOI21xp33_ASAP7_75t_L     g07833(.A1(new_n2931), .A2(\b[21] ), .B(new_n8089), .Y(new_n8090));
  NAND2xp33_ASAP7_75t_L     g07834(.A(\a[29] ), .B(new_n8090), .Y(new_n8091));
  A2O1A1Ixp33_ASAP7_75t_L   g07835(.A1(\b[21] ), .A2(new_n2931), .B(new_n8089), .C(new_n2697), .Y(new_n8092));
  NAND2xp33_ASAP7_75t_L     g07836(.A(new_n8092), .B(new_n8091), .Y(new_n8093));
  AOI21xp33_ASAP7_75t_L     g07837(.A1(new_n8087), .A2(new_n8082), .B(new_n8093), .Y(new_n8094));
  INVx1_ASAP7_75t_L         g07838(.A(new_n7965), .Y(new_n8095));
  A2O1A1Ixp33_ASAP7_75t_L   g07839(.A1(new_n7741), .A2(new_n7737), .B(new_n7745), .C(new_n8095), .Y(new_n8096));
  NOR2xp33_ASAP7_75t_L      g07840(.A(new_n8096), .B(new_n8086), .Y(new_n8097));
  NOR2xp33_ASAP7_75t_L      g07841(.A(new_n8081), .B(new_n7966), .Y(new_n8098));
  AND2x2_ASAP7_75t_L        g07842(.A(new_n8092), .B(new_n8091), .Y(new_n8099));
  NOR3xp33_ASAP7_75t_L      g07843(.A(new_n8098), .B(new_n8097), .C(new_n8099), .Y(new_n8100));
  NOR3xp33_ASAP7_75t_L      g07844(.A(new_n7964), .B(new_n8094), .C(new_n8100), .Y(new_n8101));
  O2A1O1Ixp33_ASAP7_75t_L   g07845(.A1(new_n7753), .A2(new_n7759), .B(new_n7761), .C(new_n7962), .Y(new_n8102));
  OAI21xp33_ASAP7_75t_L     g07846(.A1(new_n8097), .A2(new_n8098), .B(new_n8099), .Y(new_n8103));
  NAND3xp33_ASAP7_75t_L     g07847(.A(new_n8087), .B(new_n8082), .C(new_n8093), .Y(new_n8104));
  AOI21xp33_ASAP7_75t_L     g07848(.A1(new_n8104), .A2(new_n8103), .B(new_n8102), .Y(new_n8105));
  NOR3xp33_ASAP7_75t_L      g07849(.A(new_n8101), .B(new_n8105), .C(new_n7959), .Y(new_n8106));
  AND2x2_ASAP7_75t_L        g07850(.A(new_n7956), .B(new_n7958), .Y(new_n8107));
  NAND3xp33_ASAP7_75t_L     g07851(.A(new_n8102), .B(new_n8103), .C(new_n8104), .Y(new_n8108));
  OAI21xp33_ASAP7_75t_L     g07852(.A1(new_n8094), .A2(new_n8100), .B(new_n7964), .Y(new_n8109));
  AOI21xp33_ASAP7_75t_L     g07853(.A1(new_n8109), .A2(new_n8108), .B(new_n8107), .Y(new_n8110));
  NOR3xp33_ASAP7_75t_L      g07854(.A(new_n7952), .B(new_n8106), .C(new_n8110), .Y(new_n8111));
  NAND2xp33_ASAP7_75t_L     g07855(.A(new_n7776), .B(new_n7775), .Y(new_n8112));
  MAJIxp5_ASAP7_75t_L       g07856(.A(new_n7784), .B(new_n8112), .C(new_n7777), .Y(new_n8113));
  NAND3xp33_ASAP7_75t_L     g07857(.A(new_n8109), .B(new_n8107), .C(new_n8108), .Y(new_n8114));
  OAI21xp33_ASAP7_75t_L     g07858(.A1(new_n8105), .A2(new_n8101), .B(new_n7959), .Y(new_n8115));
  AOI21xp33_ASAP7_75t_L     g07859(.A1(new_n8115), .A2(new_n8114), .B(new_n8113), .Y(new_n8116));
  OAI21xp33_ASAP7_75t_L     g07860(.A1(new_n8116), .A2(new_n8111), .B(new_n7950), .Y(new_n8117));
  NAND2xp33_ASAP7_75t_L     g07861(.A(new_n7947), .B(new_n7949), .Y(new_n8118));
  NAND3xp33_ASAP7_75t_L     g07862(.A(new_n8113), .B(new_n8114), .C(new_n8115), .Y(new_n8119));
  OAI21xp33_ASAP7_75t_L     g07863(.A1(new_n8110), .A2(new_n8106), .B(new_n7952), .Y(new_n8120));
  NAND3xp33_ASAP7_75t_L     g07864(.A(new_n8119), .B(new_n8118), .C(new_n8120), .Y(new_n8121));
  NAND2xp33_ASAP7_75t_L     g07865(.A(new_n8121), .B(new_n8117), .Y(new_n8122));
  NOR2xp33_ASAP7_75t_L      g07866(.A(new_n7943), .B(new_n8122), .Y(new_n8123));
  AOI221xp5_ASAP7_75t_L     g07867(.A1(new_n7807), .A2(new_n7796), .B1(new_n8121), .B2(new_n8117), .C(new_n7942), .Y(new_n8124));
  OAI21xp33_ASAP7_75t_L     g07868(.A1(new_n8124), .A2(new_n8123), .B(new_n7941), .Y(new_n8125));
  INVx1_ASAP7_75t_L         g07869(.A(new_n7941), .Y(new_n8126));
  INVx1_ASAP7_75t_L         g07870(.A(new_n7942), .Y(new_n8127));
  OAI21xp33_ASAP7_75t_L     g07871(.A1(new_n7793), .A2(new_n7791), .B(new_n8127), .Y(new_n8128));
  NAND3xp33_ASAP7_75t_L     g07872(.A(new_n8128), .B(new_n8117), .C(new_n8121), .Y(new_n8129));
  INVx1_ASAP7_75t_L         g07873(.A(new_n8124), .Y(new_n8130));
  NAND3xp33_ASAP7_75t_L     g07874(.A(new_n8130), .B(new_n8129), .C(new_n8126), .Y(new_n8131));
  NAND3xp33_ASAP7_75t_L     g07875(.A(new_n7935), .B(new_n8125), .C(new_n8131), .Y(new_n8132));
  INVx1_ASAP7_75t_L         g07876(.A(new_n7238), .Y(new_n8133));
  OAI21xp33_ASAP7_75t_L     g07877(.A1(new_n8133), .A2(new_n7069), .B(new_n7242), .Y(new_n8134));
  A2O1A1O1Ixp25_ASAP7_75t_L g07878(.A1(new_n7536), .A2(new_n8134), .B(new_n7531), .C(new_n7815), .D(new_n7804), .Y(new_n8135));
  AOI21xp33_ASAP7_75t_L     g07879(.A1(new_n8130), .A2(new_n8129), .B(new_n8126), .Y(new_n8136));
  NOR3xp33_ASAP7_75t_L      g07880(.A(new_n8123), .B(new_n8124), .C(new_n7941), .Y(new_n8137));
  OAI21xp33_ASAP7_75t_L     g07881(.A1(new_n8136), .A2(new_n8137), .B(new_n8135), .Y(new_n8138));
  NAND2xp33_ASAP7_75t_L     g07882(.A(\b[33] ), .B(new_n1194), .Y(new_n8139));
  NAND2xp33_ASAP7_75t_L     g07883(.A(\b[34] ), .B(new_n1103), .Y(new_n8140));
  AOI22xp33_ASAP7_75t_L     g07884(.A1(new_n1113), .A2(\b[35] ), .B1(new_n1110), .B2(new_n5649), .Y(new_n8141));
  NAND4xp25_ASAP7_75t_L     g07885(.A(new_n8141), .B(\a[17] ), .C(new_n8139), .D(new_n8140), .Y(new_n8142));
  NAND2xp33_ASAP7_75t_L     g07886(.A(new_n8140), .B(new_n8141), .Y(new_n8143));
  A2O1A1Ixp33_ASAP7_75t_L   g07887(.A1(\b[33] ), .A2(new_n1194), .B(new_n8143), .C(new_n1107), .Y(new_n8144));
  AND2x2_ASAP7_75t_L        g07888(.A(new_n8142), .B(new_n8144), .Y(new_n8145));
  NAND3xp33_ASAP7_75t_L     g07889(.A(new_n8145), .B(new_n8132), .C(new_n8138), .Y(new_n8146));
  NOR3xp33_ASAP7_75t_L      g07890(.A(new_n8135), .B(new_n8136), .C(new_n8137), .Y(new_n8147));
  AOI21xp33_ASAP7_75t_L     g07891(.A1(new_n8131), .A2(new_n8125), .B(new_n7935), .Y(new_n8148));
  NAND2xp33_ASAP7_75t_L     g07892(.A(new_n8142), .B(new_n8144), .Y(new_n8149));
  OAI21xp33_ASAP7_75t_L     g07893(.A1(new_n8147), .A2(new_n8148), .B(new_n8149), .Y(new_n8150));
  AND2x2_ASAP7_75t_L        g07894(.A(new_n8150), .B(new_n8146), .Y(new_n8151));
  NOR3xp33_ASAP7_75t_L      g07895(.A(new_n7827), .B(new_n7823), .C(new_n7826), .Y(new_n8152));
  AOI21xp33_ASAP7_75t_L     g07896(.A1(new_n7816), .A2(new_n7811), .B(new_n7824), .Y(new_n8153));
  NOR3xp33_ASAP7_75t_L      g07897(.A(new_n7827), .B(new_n7824), .C(new_n7826), .Y(new_n8154));
  O2A1O1Ixp33_ASAP7_75t_L   g07898(.A1(new_n8152), .A2(new_n8153), .B(new_n7833), .C(new_n8154), .Y(new_n8155));
  NAND2xp33_ASAP7_75t_L     g07899(.A(new_n8155), .B(new_n8151), .Y(new_n8156));
  NAND2xp33_ASAP7_75t_L     g07900(.A(new_n8150), .B(new_n8146), .Y(new_n8157));
  A2O1A1Ixp33_ASAP7_75t_L   g07901(.A1(new_n7831), .A2(new_n7833), .B(new_n8154), .C(new_n8157), .Y(new_n8158));
  INVx1_ASAP7_75t_L         g07902(.A(new_n4922), .Y(new_n8159));
  NAND2xp33_ASAP7_75t_L     g07903(.A(new_n4918), .B(new_n8159), .Y(new_n8160));
  NAND2xp33_ASAP7_75t_L     g07904(.A(\b[37] ), .B(new_n817), .Y(new_n8161));
  OAI221xp5_ASAP7_75t_L     g07905(.A1(new_n912), .A2(new_n4915), .B1(new_n911), .B2(new_n8160), .C(new_n8161), .Y(new_n8162));
  AOI21xp33_ASAP7_75t_L     g07906(.A1(new_n908), .A2(\b[36] ), .B(new_n8162), .Y(new_n8163));
  NAND2xp33_ASAP7_75t_L     g07907(.A(\a[14] ), .B(new_n8163), .Y(new_n8164));
  A2O1A1Ixp33_ASAP7_75t_L   g07908(.A1(\b[36] ), .A2(new_n908), .B(new_n8162), .C(new_n813), .Y(new_n8165));
  AND2x2_ASAP7_75t_L        g07909(.A(new_n8165), .B(new_n8164), .Y(new_n8166));
  NAND3xp33_ASAP7_75t_L     g07910(.A(new_n8156), .B(new_n8166), .C(new_n8158), .Y(new_n8167));
  NOR2xp33_ASAP7_75t_L      g07911(.A(new_n8153), .B(new_n8152), .Y(new_n8168));
  MAJx2_ASAP7_75t_L         g07912(.A(new_n7356), .B(new_n7832), .C(new_n7546), .Y(new_n8169));
  INVx1_ASAP7_75t_L         g07913(.A(new_n8154), .Y(new_n8170));
  OAI21xp33_ASAP7_75t_L     g07914(.A1(new_n8168), .A2(new_n8169), .B(new_n8170), .Y(new_n8171));
  NOR2xp33_ASAP7_75t_L      g07915(.A(new_n8157), .B(new_n8171), .Y(new_n8172));
  AOI21xp33_ASAP7_75t_L     g07916(.A1(new_n8150), .A2(new_n8146), .B(new_n8155), .Y(new_n8173));
  NAND2xp33_ASAP7_75t_L     g07917(.A(new_n8165), .B(new_n8164), .Y(new_n8174));
  OAI21xp33_ASAP7_75t_L     g07918(.A1(new_n8173), .A2(new_n8172), .B(new_n8174), .Y(new_n8175));
  NAND2xp33_ASAP7_75t_L     g07919(.A(new_n7834), .B(new_n7830), .Y(new_n8176));
  INVx1_ASAP7_75t_L         g07920(.A(new_n8176), .Y(new_n8177));
  OAI21xp33_ASAP7_75t_L     g07921(.A1(new_n7839), .A2(new_n7841), .B(new_n8177), .Y(new_n8178));
  NAND4xp25_ASAP7_75t_L     g07922(.A(new_n7847), .B(new_n8178), .C(new_n8175), .D(new_n8167), .Y(new_n8179));
  NOR3xp33_ASAP7_75t_L      g07923(.A(new_n8172), .B(new_n8173), .C(new_n8174), .Y(new_n8180));
  AOI21xp33_ASAP7_75t_L     g07924(.A1(new_n8156), .A2(new_n8158), .B(new_n8166), .Y(new_n8181));
  MAJIxp5_ASAP7_75t_L       g07925(.A(new_n7845), .B(new_n7842), .C(new_n8176), .Y(new_n8182));
  OAI21xp33_ASAP7_75t_L     g07926(.A1(new_n8180), .A2(new_n8181), .B(new_n8182), .Y(new_n8183));
  NAND2xp33_ASAP7_75t_L     g07927(.A(\b[39] ), .B(new_n674), .Y(new_n8184));
  NAND2xp33_ASAP7_75t_L     g07928(.A(\b[40] ), .B(new_n590), .Y(new_n8185));
  AOI22xp33_ASAP7_75t_L     g07929(.A1(new_n600), .A2(\b[41] ), .B1(new_n597), .B2(new_n5669), .Y(new_n8186));
  AND4x1_ASAP7_75t_L        g07930(.A(new_n8186), .B(new_n8185), .C(new_n8184), .D(\a[11] ), .Y(new_n8187));
  AOI31xp33_ASAP7_75t_L     g07931(.A1(new_n8186), .A2(new_n8185), .A3(new_n8184), .B(\a[11] ), .Y(new_n8188));
  NOR2xp33_ASAP7_75t_L      g07932(.A(new_n8188), .B(new_n8187), .Y(new_n8189));
  NAND3xp33_ASAP7_75t_L     g07933(.A(new_n8179), .B(new_n8183), .C(new_n8189), .Y(new_n8190));
  NOR3xp33_ASAP7_75t_L      g07934(.A(new_n8182), .B(new_n8181), .C(new_n8180), .Y(new_n8191));
  OA21x2_ASAP7_75t_L        g07935(.A1(new_n8180), .A2(new_n8181), .B(new_n8182), .Y(new_n8192));
  INVx1_ASAP7_75t_L         g07936(.A(new_n8189), .Y(new_n8193));
  OAI21xp33_ASAP7_75t_L     g07937(.A1(new_n8191), .A2(new_n8192), .B(new_n8193), .Y(new_n8194));
  NAND2xp33_ASAP7_75t_L     g07938(.A(new_n8190), .B(new_n8194), .Y(new_n8195));
  NOR3xp33_ASAP7_75t_L      g07939(.A(new_n7856), .B(new_n7857), .C(new_n7854), .Y(new_n8196));
  INVx1_ASAP7_75t_L         g07940(.A(new_n8196), .Y(new_n8197));
  A2O1A1Ixp33_ASAP7_75t_L   g07941(.A1(new_n7578), .A2(new_n7860), .B(new_n7877), .C(new_n8197), .Y(new_n8198));
  NOR2xp33_ASAP7_75t_L      g07942(.A(new_n8195), .B(new_n8198), .Y(new_n8199));
  AOI21xp33_ASAP7_75t_L     g07943(.A1(new_n7864), .A2(new_n7862), .B(new_n8196), .Y(new_n8200));
  AOI21xp33_ASAP7_75t_L     g07944(.A1(new_n8194), .A2(new_n8190), .B(new_n8200), .Y(new_n8201));
  NAND2xp33_ASAP7_75t_L     g07945(.A(\b[42] ), .B(new_n480), .Y(new_n8202));
  NAND2xp33_ASAP7_75t_L     g07946(.A(\b[43] ), .B(new_n441), .Y(new_n8203));
  AOI22xp33_ASAP7_75t_L     g07947(.A1(new_n451), .A2(\b[44] ), .B1(new_n448), .B2(new_n7055), .Y(new_n8204));
  AND4x1_ASAP7_75t_L        g07948(.A(new_n8204), .B(new_n8203), .C(new_n8202), .D(\a[8] ), .Y(new_n8205));
  AOI31xp33_ASAP7_75t_L     g07949(.A1(new_n8204), .A2(new_n8203), .A3(new_n8202), .B(\a[8] ), .Y(new_n8206));
  NOR2xp33_ASAP7_75t_L      g07950(.A(new_n8206), .B(new_n8205), .Y(new_n8207));
  NOR3xp33_ASAP7_75t_L      g07951(.A(new_n8199), .B(new_n8201), .C(new_n8207), .Y(new_n8208));
  NAND3xp33_ASAP7_75t_L     g07952(.A(new_n8200), .B(new_n8194), .C(new_n8190), .Y(new_n8209));
  A2O1A1Ixp33_ASAP7_75t_L   g07953(.A1(new_n7862), .A2(new_n7864), .B(new_n8196), .C(new_n8195), .Y(new_n8210));
  AOI211xp5_ASAP7_75t_L     g07954(.A1(new_n8209), .A2(new_n8210), .B(new_n8205), .C(new_n8206), .Y(new_n8211));
  OAI21xp33_ASAP7_75t_L     g07955(.A1(new_n8208), .A2(new_n8211), .B(new_n7934), .Y(new_n8212));
  NOR3xp33_ASAP7_75t_L      g07956(.A(new_n7878), .B(new_n7872), .C(new_n7874), .Y(new_n8213));
  NOR2xp33_ASAP7_75t_L      g07957(.A(new_n8208), .B(new_n8211), .Y(new_n8214));
  A2O1A1Ixp33_ASAP7_75t_L   g07958(.A1(new_n7885), .A2(new_n7884), .B(new_n8213), .C(new_n8214), .Y(new_n8215));
  NAND3xp33_ASAP7_75t_L     g07959(.A(new_n8215), .B(new_n8212), .C(new_n7932), .Y(new_n8216));
  INVx1_ASAP7_75t_L         g07960(.A(new_n7932), .Y(new_n8217));
  OAI211xp5_ASAP7_75t_L     g07961(.A1(new_n8205), .A2(new_n8206), .B(new_n8209), .C(new_n8210), .Y(new_n8218));
  OAI21xp33_ASAP7_75t_L     g07962(.A1(new_n8201), .A2(new_n8199), .B(new_n8207), .Y(new_n8219));
  AOI221xp5_ASAP7_75t_L     g07963(.A1(new_n7884), .A2(new_n7885), .B1(new_n8218), .B2(new_n8219), .C(new_n8213), .Y(new_n8220));
  NOR3xp33_ASAP7_75t_L      g07964(.A(new_n7934), .B(new_n8208), .C(new_n8211), .Y(new_n8221));
  OAI21xp33_ASAP7_75t_L     g07965(.A1(new_n8220), .A2(new_n8221), .B(new_n8217), .Y(new_n8222));
  NAND2xp33_ASAP7_75t_L     g07966(.A(new_n8222), .B(new_n8216), .Y(new_n8223));
  XNOR2x2_ASAP7_75t_L       g07967(.A(new_n7885), .B(new_n7884), .Y(new_n8224));
  MAJIxp5_ASAP7_75t_L       g07968(.A(new_n7898), .B(new_n8224), .C(new_n7894), .Y(new_n8225));
  XNOR2x2_ASAP7_75t_L       g07969(.A(new_n8225), .B(new_n8223), .Y(new_n8226));
  NOR2xp33_ASAP7_75t_L      g07970(.A(\b[49] ), .B(\b[50] ), .Y(new_n8227));
  INVx1_ASAP7_75t_L         g07971(.A(\b[50] ), .Y(new_n8228));
  NOR2xp33_ASAP7_75t_L      g07972(.A(new_n7907), .B(new_n8228), .Y(new_n8229));
  NOR2xp33_ASAP7_75t_L      g07973(.A(new_n8227), .B(new_n8229), .Y(new_n8230));
  A2O1A1Ixp33_ASAP7_75t_L   g07974(.A1(new_n7912), .A2(new_n7909), .B(new_n7908), .C(new_n8230), .Y(new_n8231));
  O2A1O1Ixp33_ASAP7_75t_L   g07975(.A1(new_n7334), .A2(new_n7337), .B(new_n7909), .C(new_n7908), .Y(new_n8232));
  OAI21xp33_ASAP7_75t_L     g07976(.A1(new_n8227), .A2(new_n8229), .B(new_n8232), .Y(new_n8233));
  NAND2xp33_ASAP7_75t_L     g07977(.A(new_n8233), .B(new_n8231), .Y(new_n8234));
  INVx1_ASAP7_75t_L         g07978(.A(new_n8234), .Y(new_n8235));
  AOI22xp33_ASAP7_75t_L     g07979(.A1(new_n272), .A2(\b[50] ), .B1(new_n269), .B2(new_n8235), .Y(new_n8236));
  OAI221xp5_ASAP7_75t_L     g07980(.A1(new_n261), .A2(new_n7907), .B1(new_n7333), .B2(new_n277), .C(new_n8236), .Y(new_n8237));
  XNOR2x2_ASAP7_75t_L       g07981(.A(\a[2] ), .B(new_n8237), .Y(new_n8238));
  INVx1_ASAP7_75t_L         g07982(.A(new_n8238), .Y(new_n8239));
  XNOR2x2_ASAP7_75t_L       g07983(.A(new_n8239), .B(new_n8226), .Y(new_n8240));
  A2O1A1O1Ixp25_ASAP7_75t_L g07984(.A1(new_n7610), .A2(new_n7615), .B(new_n7611), .C(new_n7920), .D(new_n7921), .Y(new_n8241));
  INVx1_ASAP7_75t_L         g07985(.A(new_n8241), .Y(new_n8242));
  AND2x2_ASAP7_75t_L        g07986(.A(new_n8242), .B(new_n8240), .Y(new_n8243));
  NOR2xp33_ASAP7_75t_L      g07987(.A(new_n8242), .B(new_n8240), .Y(new_n8244));
  NOR2xp33_ASAP7_75t_L      g07988(.A(new_n8244), .B(new_n8243), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g07989(.A(new_n8241), .B(new_n8226), .C(new_n8238), .Y(new_n8246));
  INVx1_ASAP7_75t_L         g07990(.A(new_n8229), .Y(new_n8247));
  NOR2xp33_ASAP7_75t_L      g07991(.A(\b[50] ), .B(\b[51] ), .Y(new_n8248));
  INVx1_ASAP7_75t_L         g07992(.A(\b[51] ), .Y(new_n8249));
  NOR2xp33_ASAP7_75t_L      g07993(.A(new_n8228), .B(new_n8249), .Y(new_n8250));
  NOR2xp33_ASAP7_75t_L      g07994(.A(new_n8248), .B(new_n8250), .Y(new_n8251));
  INVx1_ASAP7_75t_L         g07995(.A(new_n8251), .Y(new_n8252));
  O2A1O1Ixp33_ASAP7_75t_L   g07996(.A1(new_n8227), .A2(new_n8232), .B(new_n8247), .C(new_n8252), .Y(new_n8253));
  A2O1A1O1Ixp25_ASAP7_75t_L g07997(.A1(new_n7909), .A2(new_n7912), .B(new_n7908), .C(new_n8230), .D(new_n8229), .Y(new_n8254));
  NAND2xp33_ASAP7_75t_L     g07998(.A(new_n8252), .B(new_n8254), .Y(new_n8255));
  INVx1_ASAP7_75t_L         g07999(.A(new_n8255), .Y(new_n8256));
  NOR2xp33_ASAP7_75t_L      g08000(.A(new_n8253), .B(new_n8256), .Y(new_n8257));
  NOR2xp33_ASAP7_75t_L      g08001(.A(new_n8249), .B(new_n632), .Y(new_n8258));
  AOI221xp5_ASAP7_75t_L     g08002(.A1(new_n380), .A2(\b[50] ), .B1(new_n269), .B2(new_n8257), .C(new_n8258), .Y(new_n8259));
  OA211x2_ASAP7_75t_L       g08003(.A1(new_n277), .A2(new_n7907), .B(new_n8259), .C(\a[2] ), .Y(new_n8260));
  O2A1O1Ixp33_ASAP7_75t_L   g08004(.A1(new_n7907), .A2(new_n277), .B(new_n8259), .C(\a[2] ), .Y(new_n8261));
  NOR2xp33_ASAP7_75t_L      g08005(.A(new_n8261), .B(new_n8260), .Y(new_n8262));
  NOR3xp33_ASAP7_75t_L      g08006(.A(new_n8221), .B(new_n8220), .C(new_n8217), .Y(new_n8263));
  AOI21xp33_ASAP7_75t_L     g08007(.A1(new_n8215), .A2(new_n8212), .B(new_n7932), .Y(new_n8264));
  NOR3xp33_ASAP7_75t_L      g08008(.A(new_n8221), .B(new_n8220), .C(new_n7932), .Y(new_n8265));
  O2A1O1Ixp33_ASAP7_75t_L   g08009(.A1(new_n8263), .A2(new_n8264), .B(new_n8225), .C(new_n8265), .Y(new_n8266));
  NAND2xp33_ASAP7_75t_L     g08010(.A(\b[47] ), .B(new_n334), .Y(new_n8267));
  AOI22xp33_ASAP7_75t_L     g08011(.A1(new_n345), .A2(\b[48] ), .B1(new_n342), .B2(new_n7341), .Y(new_n8268));
  NAND2xp33_ASAP7_75t_L     g08012(.A(new_n8267), .B(new_n8268), .Y(new_n8269));
  INVx1_ASAP7_75t_L         g08013(.A(new_n8269), .Y(new_n8270));
  OAI211xp5_ASAP7_75t_L     g08014(.A1(new_n7033), .A2(new_n365), .B(new_n8270), .C(\a[5] ), .Y(new_n8271));
  A2O1A1Ixp33_ASAP7_75t_L   g08015(.A1(\b[46] ), .A2(new_n366), .B(new_n8269), .C(new_n339), .Y(new_n8272));
  NAND2xp33_ASAP7_75t_L     g08016(.A(new_n8272), .B(new_n8271), .Y(new_n8273));
  NOR3xp33_ASAP7_75t_L      g08017(.A(new_n8145), .B(new_n8148), .C(new_n8147), .Y(new_n8274));
  INVx1_ASAP7_75t_L         g08018(.A(new_n8274), .Y(new_n8275));
  NAND2xp33_ASAP7_75t_L     g08019(.A(\b[34] ), .B(new_n1194), .Y(new_n8276));
  NAND2xp33_ASAP7_75t_L     g08020(.A(\b[35] ), .B(new_n1103), .Y(new_n8277));
  AOI22xp33_ASAP7_75t_L     g08021(.A1(new_n1113), .A2(\b[36] ), .B1(new_n1110), .B2(new_n4473), .Y(new_n8278));
  AND4x1_ASAP7_75t_L        g08022(.A(new_n8278), .B(new_n8277), .C(new_n8276), .D(\a[17] ), .Y(new_n8279));
  AOI31xp33_ASAP7_75t_L     g08023(.A1(new_n8278), .A2(new_n8277), .A3(new_n8276), .B(\a[17] ), .Y(new_n8280));
  NOR2xp33_ASAP7_75t_L      g08024(.A(new_n8280), .B(new_n8279), .Y(new_n8281));
  A2O1A1O1Ixp25_ASAP7_75t_L g08025(.A1(new_n7813), .A2(new_n7815), .B(new_n7804), .C(new_n8125), .D(new_n8137), .Y(new_n8282));
  NOR3xp33_ASAP7_75t_L      g08026(.A(new_n8111), .B(new_n8116), .C(new_n7950), .Y(new_n8283));
  A2O1A1O1Ixp25_ASAP7_75t_L g08027(.A1(new_n7807), .A2(new_n7796), .B(new_n7942), .C(new_n8117), .D(new_n8283), .Y(new_n8284));
  NAND2xp33_ASAP7_75t_L     g08028(.A(\b[28] ), .B(new_n1910), .Y(new_n8285));
  NAND2xp33_ASAP7_75t_L     g08029(.A(\b[29] ), .B(new_n1770), .Y(new_n8286));
  AOI22xp33_ASAP7_75t_L     g08030(.A1(new_n1766), .A2(\b[30] ), .B1(new_n1764), .B2(new_n3219), .Y(new_n8287));
  AND4x1_ASAP7_75t_L        g08031(.A(new_n8287), .B(new_n8286), .C(new_n8285), .D(\a[23] ), .Y(new_n8288));
  AOI31xp33_ASAP7_75t_L     g08032(.A1(new_n8287), .A2(new_n8286), .A3(new_n8285), .B(\a[23] ), .Y(new_n8289));
  NOR2xp33_ASAP7_75t_L      g08033(.A(new_n8289), .B(new_n8288), .Y(new_n8290));
  NAND2xp33_ASAP7_75t_L     g08034(.A(new_n7782), .B(new_n7783), .Y(new_n8291));
  NOR2xp33_ASAP7_75t_L      g08035(.A(new_n7777), .B(new_n8112), .Y(new_n8292));
  A2O1A1O1Ixp25_ASAP7_75t_L g08036(.A1(new_n7780), .A2(new_n8291), .B(new_n8292), .C(new_n8114), .D(new_n8110), .Y(new_n8293));
  NAND2xp33_ASAP7_75t_L     g08037(.A(new_n8065), .B(new_n8061), .Y(new_n8294));
  NOR3xp33_ASAP7_75t_L      g08038(.A(new_n8060), .B(new_n8062), .C(new_n8056), .Y(new_n8295));
  NOR2xp33_ASAP7_75t_L      g08039(.A(new_n1356), .B(new_n4115), .Y(new_n8296));
  AOI221xp5_ASAP7_75t_L     g08040(.A1(new_n3874), .A2(\b[17] ), .B1(new_n3881), .B2(new_n1363), .C(new_n8296), .Y(new_n8297));
  OAI21xp33_ASAP7_75t_L     g08041(.A1(new_n1051), .A2(new_n4986), .B(new_n8297), .Y(new_n8298));
  NOR2xp33_ASAP7_75t_L      g08042(.A(new_n3878), .B(new_n8298), .Y(new_n8299));
  O2A1O1Ixp33_ASAP7_75t_L   g08043(.A1(new_n1051), .A2(new_n4986), .B(new_n8297), .C(\a[35] ), .Y(new_n8300));
  NOR2xp33_ASAP7_75t_L      g08044(.A(new_n8300), .B(new_n8299), .Y(new_n8301));
  NAND2xp33_ASAP7_75t_L     g08045(.A(new_n8040), .B(new_n8044), .Y(new_n8302));
  NAND2xp33_ASAP7_75t_L     g08046(.A(\b[13] ), .B(new_n4780), .Y(new_n8303));
  NAND2xp33_ASAP7_75t_L     g08047(.A(\b[14] ), .B(new_n4548), .Y(new_n8304));
  AOI22xp33_ASAP7_75t_L     g08048(.A1(new_n4544), .A2(\b[15] ), .B1(new_n4542), .B2(new_n959), .Y(new_n8305));
  AND4x1_ASAP7_75t_L        g08049(.A(new_n8305), .B(new_n8304), .C(new_n8303), .D(\a[38] ), .Y(new_n8306));
  AOI31xp33_ASAP7_75t_L     g08050(.A1(new_n8305), .A2(new_n8304), .A3(new_n8303), .B(\a[38] ), .Y(new_n8307));
  A2O1A1Ixp33_ASAP7_75t_L   g08051(.A1(new_n8043), .A2(new_n7700), .B(new_n8041), .C(new_n8037), .Y(new_n8308));
  NOR2xp33_ASAP7_75t_L      g08052(.A(new_n631), .B(new_n5521), .Y(new_n8309));
  INVx1_ASAP7_75t_L         g08053(.A(new_n8309), .Y(new_n8310));
  NAND2xp33_ASAP7_75t_L     g08054(.A(\b[11] ), .B(new_n5240), .Y(new_n8311));
  AOI32xp33_ASAP7_75t_L     g08055(.A1(new_n771), .A2(new_n774), .A3(new_n5247), .B1(new_n5249), .B2(\b[12] ), .Y(new_n8312));
  AND4x1_ASAP7_75t_L        g08056(.A(new_n8312), .B(new_n8311), .C(new_n8310), .D(\a[41] ), .Y(new_n8313));
  AOI31xp33_ASAP7_75t_L     g08057(.A1(new_n8312), .A2(new_n8311), .A3(new_n8310), .B(\a[41] ), .Y(new_n8314));
  NOR2xp33_ASAP7_75t_L      g08058(.A(new_n8314), .B(new_n8313), .Y(new_n8315));
  AOI211xp5_ASAP7_75t_L     g08059(.A1(new_n8016), .A2(new_n8017), .B(new_n8011), .C(new_n8014), .Y(new_n8316));
  NAND5xp2_ASAP7_75t_L      g08060(.A(new_n7660), .B(new_n7657), .C(new_n7650), .D(new_n7639), .E(\a[50] ), .Y(new_n8317));
  INVx1_ASAP7_75t_L         g08061(.A(\a[51] ), .Y(new_n8318));
  NAND2xp33_ASAP7_75t_L     g08062(.A(\a[50] ), .B(new_n8318), .Y(new_n8319));
  NAND2xp33_ASAP7_75t_L     g08063(.A(\a[51] ), .B(new_n7653), .Y(new_n8320));
  AND2x2_ASAP7_75t_L        g08064(.A(new_n8319), .B(new_n8320), .Y(new_n8321));
  NOR2xp33_ASAP7_75t_L      g08065(.A(new_n258), .B(new_n8321), .Y(new_n8322));
  OAI31xp33_ASAP7_75t_L     g08066(.A1(new_n8317), .A2(new_n7999), .A3(new_n7995), .B(new_n8322), .Y(new_n8323));
  INVx1_ASAP7_75t_L         g08067(.A(new_n8322), .Y(new_n8324));
  NAND5xp2_ASAP7_75t_L      g08068(.A(\a[50] ), .B(new_n8000), .C(new_n8324), .D(new_n7664), .E(new_n7639), .Y(new_n8325));
  NAND2xp33_ASAP7_75t_L     g08069(.A(new_n7992), .B(new_n7388), .Y(new_n8326));
  NAND2xp33_ASAP7_75t_L     g08070(.A(\b[3] ), .B(new_n7659), .Y(new_n8327));
  OAI221xp5_ASAP7_75t_L     g08071(.A1(new_n278), .A2(new_n8326), .B1(new_n7996), .B2(new_n303), .C(new_n8327), .Y(new_n8328));
  AO211x2_ASAP7_75t_L       g08072(.A1(\b[1] ), .A2(new_n7993), .B(new_n7653), .C(new_n8328), .Y(new_n8329));
  A2O1A1Ixp33_ASAP7_75t_L   g08073(.A1(\b[1] ), .A2(new_n7993), .B(new_n8328), .C(new_n7653), .Y(new_n8330));
  AO22x1_ASAP7_75t_L        g08074(.A1(new_n8330), .A2(new_n8329), .B1(new_n8323), .B2(new_n8325), .Y(new_n8331));
  NAND4xp25_ASAP7_75t_L     g08075(.A(new_n8325), .B(new_n8323), .C(new_n8329), .D(new_n8330), .Y(new_n8332));
  NAND2xp33_ASAP7_75t_L     g08076(.A(\b[4] ), .B(new_n7124), .Y(new_n8333));
  NAND2xp33_ASAP7_75t_L     g08077(.A(\b[5] ), .B(new_n6812), .Y(new_n8334));
  AOI22xp33_ASAP7_75t_L     g08078(.A1(new_n6822), .A2(\b[6] ), .B1(new_n6819), .B2(new_n389), .Y(new_n8335));
  NAND4xp25_ASAP7_75t_L     g08079(.A(new_n8335), .B(\a[47] ), .C(new_n8333), .D(new_n8334), .Y(new_n8336));
  OAI221xp5_ASAP7_75t_L     g08080(.A1(new_n7118), .A2(new_n382), .B1(new_n7117), .B2(new_n540), .C(new_n8334), .Y(new_n8337));
  A2O1A1Ixp33_ASAP7_75t_L   g08081(.A1(\b[4] ), .A2(new_n7124), .B(new_n8337), .C(new_n6816), .Y(new_n8338));
  AND4x1_ASAP7_75t_L        g08082(.A(new_n8331), .B(new_n8338), .C(new_n8332), .D(new_n8336), .Y(new_n8339));
  AOI22xp33_ASAP7_75t_L     g08083(.A1(new_n8338), .A2(new_n8336), .B1(new_n8332), .B2(new_n8331), .Y(new_n8340));
  NOR2xp33_ASAP7_75t_L      g08084(.A(new_n8340), .B(new_n8339), .Y(new_n8341));
  NAND2xp33_ASAP7_75t_L     g08085(.A(new_n7991), .B(new_n7990), .Y(new_n8342));
  NOR2xp33_ASAP7_75t_L      g08086(.A(new_n8009), .B(new_n8006), .Y(new_n8343));
  MAJIxp5_ASAP7_75t_L       g08087(.A(new_n8012), .B(new_n8343), .C(new_n8342), .Y(new_n8344));
  NAND2xp33_ASAP7_75t_L     g08088(.A(new_n8341), .B(new_n8344), .Y(new_n8345));
  NAND4xp25_ASAP7_75t_L     g08089(.A(new_n8331), .B(new_n8338), .C(new_n8336), .D(new_n8332), .Y(new_n8346));
  AO22x1_ASAP7_75t_L        g08090(.A1(new_n8336), .A2(new_n8338), .B1(new_n8332), .B2(new_n8331), .Y(new_n8347));
  NAND2xp33_ASAP7_75t_L     g08091(.A(new_n8346), .B(new_n8347), .Y(new_n8348));
  A2O1A1Ixp33_ASAP7_75t_L   g08092(.A1(new_n8343), .A2(new_n8342), .B(new_n8011), .C(new_n8348), .Y(new_n8349));
  NAND2xp33_ASAP7_75t_L     g08093(.A(\b[8] ), .B(new_n5992), .Y(new_n8350));
  OAI221xp5_ASAP7_75t_L     g08094(.A1(new_n6312), .A2(new_n559), .B1(new_n6311), .B2(new_n978), .C(new_n8350), .Y(new_n8351));
  AOI211xp5_ASAP7_75t_L     g08095(.A1(\b[7] ), .A2(new_n6308), .B(new_n5996), .C(new_n8351), .Y(new_n8352));
  A2O1A1Ixp33_ASAP7_75t_L   g08096(.A1(\b[7] ), .A2(new_n6308), .B(new_n8351), .C(new_n5996), .Y(new_n8353));
  INVx1_ASAP7_75t_L         g08097(.A(new_n8353), .Y(new_n8354));
  AOI211xp5_ASAP7_75t_L     g08098(.A1(new_n8349), .A2(new_n8345), .B(new_n8352), .C(new_n8354), .Y(new_n8355));
  NAND2xp33_ASAP7_75t_L     g08099(.A(new_n8343), .B(new_n8342), .Y(new_n8356));
  A2O1A1Ixp33_ASAP7_75t_L   g08100(.A1(new_n8004), .A2(new_n8010), .B(new_n7986), .C(new_n8356), .Y(new_n8357));
  NOR2xp33_ASAP7_75t_L      g08101(.A(new_n8357), .B(new_n8348), .Y(new_n8358));
  NOR2xp33_ASAP7_75t_L      g08102(.A(new_n8341), .B(new_n8344), .Y(new_n8359));
  INVx1_ASAP7_75t_L         g08103(.A(new_n8352), .Y(new_n8360));
  AOI211xp5_ASAP7_75t_L     g08104(.A1(new_n8360), .A2(new_n8353), .B(new_n8359), .C(new_n8358), .Y(new_n8361));
  NOR2xp33_ASAP7_75t_L      g08105(.A(new_n8361), .B(new_n8355), .Y(new_n8362));
  A2O1A1Ixp33_ASAP7_75t_L   g08106(.A1(new_n8024), .A2(new_n8034), .B(new_n8316), .C(new_n8362), .Y(new_n8363));
  O2A1O1Ixp33_ASAP7_75t_L   g08107(.A1(new_n7980), .A2(new_n7687), .B(new_n8024), .C(new_n8316), .Y(new_n8364));
  OAI211xp5_ASAP7_75t_L     g08108(.A1(new_n8359), .A2(new_n8358), .B(new_n8360), .C(new_n8353), .Y(new_n8365));
  OAI211xp5_ASAP7_75t_L     g08109(.A1(new_n8352), .A2(new_n8354), .B(new_n8349), .C(new_n8345), .Y(new_n8366));
  NAND2xp33_ASAP7_75t_L     g08110(.A(new_n8366), .B(new_n8365), .Y(new_n8367));
  NAND2xp33_ASAP7_75t_L     g08111(.A(new_n8364), .B(new_n8367), .Y(new_n8368));
  AOI21xp33_ASAP7_75t_L     g08112(.A1(new_n8363), .A2(new_n8368), .B(new_n8315), .Y(new_n8369));
  INVx1_ASAP7_75t_L         g08113(.A(new_n8315), .Y(new_n8370));
  NOR2xp33_ASAP7_75t_L      g08114(.A(new_n8364), .B(new_n8367), .Y(new_n8371));
  AO21x2_ASAP7_75t_L        g08115(.A1(new_n8024), .A2(new_n8034), .B(new_n8316), .Y(new_n8372));
  NOR2xp33_ASAP7_75t_L      g08116(.A(new_n8372), .B(new_n8362), .Y(new_n8373));
  NOR3xp33_ASAP7_75t_L      g08117(.A(new_n8373), .B(new_n8370), .C(new_n8371), .Y(new_n8374));
  OAI21xp33_ASAP7_75t_L     g08118(.A1(new_n8369), .A2(new_n8374), .B(new_n8308), .Y(new_n8375));
  A2O1A1Ixp33_ASAP7_75t_L   g08119(.A1(new_n6851), .A2(new_n6848), .B(new_n7098), .C(new_n7150), .Y(new_n8376));
  A2O1A1Ixp33_ASAP7_75t_L   g08120(.A1(new_n8376), .A2(new_n7441), .B(new_n7426), .C(new_n7435), .Y(new_n8377));
  NOR3xp33_ASAP7_75t_L      g08121(.A(new_n7685), .B(new_n7694), .C(new_n7687), .Y(new_n8378));
  A2O1A1O1Ixp25_ASAP7_75t_L g08122(.A1(new_n7695), .A2(new_n8377), .B(new_n8378), .C(new_n8032), .D(new_n8042), .Y(new_n8379));
  OAI21xp33_ASAP7_75t_L     g08123(.A1(new_n8371), .A2(new_n8373), .B(new_n8370), .Y(new_n8380));
  NAND3xp33_ASAP7_75t_L     g08124(.A(new_n8363), .B(new_n8315), .C(new_n8368), .Y(new_n8381));
  NAND3xp33_ASAP7_75t_L     g08125(.A(new_n8379), .B(new_n8380), .C(new_n8381), .Y(new_n8382));
  OAI211xp5_ASAP7_75t_L     g08126(.A1(new_n8306), .A2(new_n8307), .B(new_n8382), .C(new_n8375), .Y(new_n8383));
  NOR2xp33_ASAP7_75t_L      g08127(.A(new_n8307), .B(new_n8306), .Y(new_n8384));
  AOI21xp33_ASAP7_75t_L     g08128(.A1(new_n8381), .A2(new_n8380), .B(new_n8379), .Y(new_n8385));
  NOR3xp33_ASAP7_75t_L      g08129(.A(new_n8308), .B(new_n8369), .C(new_n8374), .Y(new_n8386));
  OAI21xp33_ASAP7_75t_L     g08130(.A1(new_n8385), .A2(new_n8386), .B(new_n8384), .Y(new_n8387));
  NAND2xp33_ASAP7_75t_L     g08131(.A(new_n8383), .B(new_n8387), .Y(new_n8388));
  O2A1O1Ixp33_ASAP7_75t_L   g08132(.A1(new_n8302), .A2(new_n8050), .B(new_n8063), .C(new_n8388), .Y(new_n8389));
  NAND3xp33_ASAP7_75t_L     g08133(.A(new_n8044), .B(new_n8040), .C(new_n8054), .Y(new_n8390));
  A2O1A1Ixp33_ASAP7_75t_L   g08134(.A1(new_n8051), .A2(new_n8055), .B(new_n7977), .C(new_n8390), .Y(new_n8391));
  AOI21xp33_ASAP7_75t_L     g08135(.A1(new_n8387), .A2(new_n8383), .B(new_n8391), .Y(new_n8392));
  NOR3xp33_ASAP7_75t_L      g08136(.A(new_n8389), .B(new_n8392), .C(new_n8301), .Y(new_n8393));
  XNOR2x2_ASAP7_75t_L       g08137(.A(new_n3878), .B(new_n8298), .Y(new_n8394));
  NAND3xp33_ASAP7_75t_L     g08138(.A(new_n8391), .B(new_n8383), .C(new_n8387), .Y(new_n8395));
  NAND3xp33_ASAP7_75t_L     g08139(.A(new_n8388), .B(new_n8063), .C(new_n8390), .Y(new_n8396));
  AOI21xp33_ASAP7_75t_L     g08140(.A1(new_n8396), .A2(new_n8395), .B(new_n8394), .Y(new_n8397));
  NOR2xp33_ASAP7_75t_L      g08141(.A(new_n8397), .B(new_n8393), .Y(new_n8398));
  A2O1A1Ixp33_ASAP7_75t_L   g08142(.A1(new_n8294), .A2(new_n7968), .B(new_n8295), .C(new_n8398), .Y(new_n8399));
  O2A1O1Ixp33_ASAP7_75t_L   g08143(.A1(new_n8070), .A2(new_n8071), .B(new_n7968), .C(new_n8295), .Y(new_n8400));
  OAI21xp33_ASAP7_75t_L     g08144(.A1(new_n8393), .A2(new_n8397), .B(new_n8400), .Y(new_n8401));
  NAND2xp33_ASAP7_75t_L     g08145(.A(\b[19] ), .B(new_n3491), .Y(new_n8402));
  NAND2xp33_ASAP7_75t_L     g08146(.A(\b[20] ), .B(new_n3260), .Y(new_n8403));
  AOI22xp33_ASAP7_75t_L     g08147(.A1(new_n3256), .A2(\b[21] ), .B1(new_n3254), .B2(new_n1715), .Y(new_n8404));
  NAND4xp25_ASAP7_75t_L     g08148(.A(new_n8404), .B(\a[32] ), .C(new_n8402), .D(new_n8403), .Y(new_n8405));
  NAND2xp33_ASAP7_75t_L     g08149(.A(new_n8403), .B(new_n8404), .Y(new_n8406));
  A2O1A1Ixp33_ASAP7_75t_L   g08150(.A1(\b[19] ), .A2(new_n3491), .B(new_n8406), .C(new_n3251), .Y(new_n8407));
  AND2x2_ASAP7_75t_L        g08151(.A(new_n8405), .B(new_n8407), .Y(new_n8408));
  NAND3xp33_ASAP7_75t_L     g08152(.A(new_n8399), .B(new_n8401), .C(new_n8408), .Y(new_n8409));
  AO21x2_ASAP7_75t_L        g08153(.A1(new_n8401), .A2(new_n8399), .B(new_n8408), .Y(new_n8410));
  A2O1A1O1Ixp25_ASAP7_75t_L g08154(.A1(new_n7755), .A2(new_n8083), .B(new_n7965), .C(new_n8080), .D(new_n8084), .Y(new_n8411));
  AND3x1_ASAP7_75t_L        g08155(.A(new_n8411), .B(new_n8410), .C(new_n8409), .Y(new_n8412));
  AOI21xp33_ASAP7_75t_L     g08156(.A1(new_n8410), .A2(new_n8409), .B(new_n8411), .Y(new_n8413));
  NAND2xp33_ASAP7_75t_L     g08157(.A(\b[22] ), .B(new_n2931), .Y(new_n8414));
  NAND2xp33_ASAP7_75t_L     g08158(.A(\b[23] ), .B(new_n2706), .Y(new_n8415));
  AOI22xp33_ASAP7_75t_L     g08159(.A1(new_n2702), .A2(\b[24] ), .B1(new_n2700), .B2(new_n2027), .Y(new_n8416));
  NAND4xp25_ASAP7_75t_L     g08160(.A(new_n8416), .B(\a[29] ), .C(new_n8414), .D(new_n8415), .Y(new_n8417));
  NAND2xp33_ASAP7_75t_L     g08161(.A(new_n8415), .B(new_n8416), .Y(new_n8418));
  A2O1A1Ixp33_ASAP7_75t_L   g08162(.A1(\b[22] ), .A2(new_n2931), .B(new_n8418), .C(new_n2697), .Y(new_n8419));
  NAND2xp33_ASAP7_75t_L     g08163(.A(new_n8417), .B(new_n8419), .Y(new_n8420));
  INVx1_ASAP7_75t_L         g08164(.A(new_n8420), .Y(new_n8421));
  OAI21xp33_ASAP7_75t_L     g08165(.A1(new_n8413), .A2(new_n8412), .B(new_n8421), .Y(new_n8422));
  NAND3xp33_ASAP7_75t_L     g08166(.A(new_n8411), .B(new_n8410), .C(new_n8409), .Y(new_n8423));
  AND3x1_ASAP7_75t_L        g08167(.A(new_n8399), .B(new_n8408), .C(new_n8401), .Y(new_n8424));
  AOI21xp33_ASAP7_75t_L     g08168(.A1(new_n8399), .A2(new_n8401), .B(new_n8408), .Y(new_n8425));
  A2O1A1Ixp33_ASAP7_75t_L   g08169(.A1(new_n7757), .A2(new_n8095), .B(new_n8085), .C(new_n8079), .Y(new_n8426));
  OAI21xp33_ASAP7_75t_L     g08170(.A1(new_n8424), .A2(new_n8425), .B(new_n8426), .Y(new_n8427));
  NAND3xp33_ASAP7_75t_L     g08171(.A(new_n8427), .B(new_n8423), .C(new_n8420), .Y(new_n8428));
  A2O1A1Ixp33_ASAP7_75t_L   g08172(.A1(new_n7776), .A2(new_n7963), .B(new_n8094), .C(new_n8104), .Y(new_n8429));
  NAND3xp33_ASAP7_75t_L     g08173(.A(new_n8429), .B(new_n8428), .C(new_n8422), .Y(new_n8430));
  AOI21xp33_ASAP7_75t_L     g08174(.A1(new_n8427), .A2(new_n8423), .B(new_n8420), .Y(new_n8431));
  NOR3xp33_ASAP7_75t_L      g08175(.A(new_n8412), .B(new_n8413), .C(new_n8421), .Y(new_n8432));
  NAND2xp33_ASAP7_75t_L     g08176(.A(new_n7764), .B(new_n7763), .Y(new_n8433));
  A2O1A1O1Ixp25_ASAP7_75t_L g08177(.A1(new_n7761), .A2(new_n8433), .B(new_n7962), .C(new_n8103), .D(new_n8100), .Y(new_n8434));
  OAI21xp33_ASAP7_75t_L     g08178(.A1(new_n8431), .A2(new_n8432), .B(new_n8434), .Y(new_n8435));
  NAND2xp33_ASAP7_75t_L     g08179(.A(\b[25] ), .B(new_n2386), .Y(new_n8436));
  NAND2xp33_ASAP7_75t_L     g08180(.A(\b[26] ), .B(new_n2232), .Y(new_n8437));
  AOI22xp33_ASAP7_75t_L     g08181(.A1(new_n2228), .A2(\b[27] ), .B1(new_n2226), .B2(new_n2657), .Y(new_n8438));
  NAND4xp25_ASAP7_75t_L     g08182(.A(new_n8438), .B(\a[26] ), .C(new_n8436), .D(new_n8437), .Y(new_n8439));
  NAND2xp33_ASAP7_75t_L     g08183(.A(new_n8437), .B(new_n8438), .Y(new_n8440));
  A2O1A1Ixp33_ASAP7_75t_L   g08184(.A1(\b[25] ), .A2(new_n2386), .B(new_n8440), .C(new_n2223), .Y(new_n8441));
  NAND2xp33_ASAP7_75t_L     g08185(.A(new_n8439), .B(new_n8441), .Y(new_n8442));
  INVx1_ASAP7_75t_L         g08186(.A(new_n8442), .Y(new_n8443));
  NAND3xp33_ASAP7_75t_L     g08187(.A(new_n8430), .B(new_n8443), .C(new_n8435), .Y(new_n8444));
  NOR3xp33_ASAP7_75t_L      g08188(.A(new_n8434), .B(new_n8432), .C(new_n8431), .Y(new_n8445));
  AOI21xp33_ASAP7_75t_L     g08189(.A1(new_n8428), .A2(new_n8422), .B(new_n8429), .Y(new_n8446));
  OAI21xp33_ASAP7_75t_L     g08190(.A1(new_n8445), .A2(new_n8446), .B(new_n8442), .Y(new_n8447));
  AOI21xp33_ASAP7_75t_L     g08191(.A1(new_n8447), .A2(new_n8444), .B(new_n8293), .Y(new_n8448));
  INVx1_ASAP7_75t_L         g08192(.A(new_n8292), .Y(new_n8449));
  A2O1A1Ixp33_ASAP7_75t_L   g08193(.A1(new_n7781), .A2(new_n8449), .B(new_n8106), .C(new_n8115), .Y(new_n8450));
  NAND2xp33_ASAP7_75t_L     g08194(.A(new_n8444), .B(new_n8447), .Y(new_n8451));
  NOR2xp33_ASAP7_75t_L      g08195(.A(new_n8450), .B(new_n8451), .Y(new_n8452));
  NOR3xp33_ASAP7_75t_L      g08196(.A(new_n8452), .B(new_n8448), .C(new_n8290), .Y(new_n8453));
  INVx1_ASAP7_75t_L         g08197(.A(new_n8290), .Y(new_n8454));
  A2O1A1Ixp33_ASAP7_75t_L   g08198(.A1(new_n8114), .A2(new_n8113), .B(new_n8110), .C(new_n8451), .Y(new_n8455));
  NOR3xp33_ASAP7_75t_L      g08199(.A(new_n8446), .B(new_n8445), .C(new_n8442), .Y(new_n8456));
  AOI21xp33_ASAP7_75t_L     g08200(.A1(new_n8430), .A2(new_n8435), .B(new_n8443), .Y(new_n8457));
  NOR2xp33_ASAP7_75t_L      g08201(.A(new_n8457), .B(new_n8456), .Y(new_n8458));
  NAND2xp33_ASAP7_75t_L     g08202(.A(new_n8293), .B(new_n8458), .Y(new_n8459));
  AOI21xp33_ASAP7_75t_L     g08203(.A1(new_n8455), .A2(new_n8459), .B(new_n8454), .Y(new_n8460));
  OR3x1_ASAP7_75t_L         g08204(.A(new_n8284), .B(new_n8460), .C(new_n8453), .Y(new_n8461));
  OAI21xp33_ASAP7_75t_L     g08205(.A1(new_n8453), .A2(new_n8460), .B(new_n8284), .Y(new_n8462));
  NAND2xp33_ASAP7_75t_L     g08206(.A(\b[32] ), .B(new_n1410), .Y(new_n8463));
  AOI22xp33_ASAP7_75t_L     g08207(.A1(new_n1406), .A2(\b[33] ), .B1(new_n1404), .B2(new_n3813), .Y(new_n8464));
  NAND2xp33_ASAP7_75t_L     g08208(.A(new_n8463), .B(new_n8464), .Y(new_n8465));
  AOI211xp5_ASAP7_75t_L     g08209(.A1(\b[31] ), .A2(new_n1548), .B(new_n1401), .C(new_n8465), .Y(new_n8466));
  INVx1_ASAP7_75t_L         g08210(.A(new_n8465), .Y(new_n8467));
  O2A1O1Ixp33_ASAP7_75t_L   g08211(.A1(new_n3419), .A2(new_n1549), .B(new_n8467), .C(\a[20] ), .Y(new_n8468));
  NOR2xp33_ASAP7_75t_L      g08212(.A(new_n8466), .B(new_n8468), .Y(new_n8469));
  NAND3xp33_ASAP7_75t_L     g08213(.A(new_n8461), .B(new_n8469), .C(new_n8462), .Y(new_n8470));
  NOR3xp33_ASAP7_75t_L      g08214(.A(new_n8284), .B(new_n8460), .C(new_n8453), .Y(new_n8471));
  OA21x2_ASAP7_75t_L        g08215(.A1(new_n8453), .A2(new_n8460), .B(new_n8284), .Y(new_n8472));
  OR2x4_ASAP7_75t_L         g08216(.A(new_n8466), .B(new_n8468), .Y(new_n8473));
  OAI21xp33_ASAP7_75t_L     g08217(.A1(new_n8471), .A2(new_n8472), .B(new_n8473), .Y(new_n8474));
  AOI21xp33_ASAP7_75t_L     g08218(.A1(new_n8474), .A2(new_n8470), .B(new_n8282), .Y(new_n8475));
  AND3x1_ASAP7_75t_L        g08219(.A(new_n8282), .B(new_n8474), .C(new_n8470), .Y(new_n8476));
  NOR3xp33_ASAP7_75t_L      g08220(.A(new_n8476), .B(new_n8475), .C(new_n8281), .Y(new_n8477));
  INVx1_ASAP7_75t_L         g08221(.A(new_n8281), .Y(new_n8478));
  OAI21xp33_ASAP7_75t_L     g08222(.A1(new_n8136), .A2(new_n8135), .B(new_n8131), .Y(new_n8479));
  NOR3xp33_ASAP7_75t_L      g08223(.A(new_n8473), .B(new_n8472), .C(new_n8471), .Y(new_n8480));
  AOI21xp33_ASAP7_75t_L     g08224(.A1(new_n8461), .A2(new_n8462), .B(new_n8469), .Y(new_n8481));
  OAI21xp33_ASAP7_75t_L     g08225(.A1(new_n8480), .A2(new_n8481), .B(new_n8479), .Y(new_n8482));
  NAND3xp33_ASAP7_75t_L     g08226(.A(new_n8282), .B(new_n8470), .C(new_n8474), .Y(new_n8483));
  AOI21xp33_ASAP7_75t_L     g08227(.A1(new_n8482), .A2(new_n8483), .B(new_n8478), .Y(new_n8484));
  OAI221xp5_ASAP7_75t_L     g08228(.A1(new_n8484), .A2(new_n8477), .B1(new_n8155), .B2(new_n8151), .C(new_n8275), .Y(new_n8485));
  A2O1A1Ixp33_ASAP7_75t_L   g08229(.A1(new_n8150), .A2(new_n8146), .B(new_n8155), .C(new_n8275), .Y(new_n8486));
  NOR2xp33_ASAP7_75t_L      g08230(.A(new_n8484), .B(new_n8477), .Y(new_n8487));
  NAND2xp33_ASAP7_75t_L     g08231(.A(new_n8487), .B(new_n8486), .Y(new_n8488));
  NAND2xp33_ASAP7_75t_L     g08232(.A(\b[37] ), .B(new_n908), .Y(new_n8489));
  NAND2xp33_ASAP7_75t_L     g08233(.A(\b[38] ), .B(new_n817), .Y(new_n8490));
  AOI22xp33_ASAP7_75t_L     g08234(.A1(new_n826), .A2(\b[39] ), .B1(new_n823), .B2(new_n5174), .Y(new_n8491));
  AND4x1_ASAP7_75t_L        g08235(.A(new_n8491), .B(new_n8490), .C(new_n8489), .D(\a[14] ), .Y(new_n8492));
  AOI31xp33_ASAP7_75t_L     g08236(.A1(new_n8491), .A2(new_n8490), .A3(new_n8489), .B(\a[14] ), .Y(new_n8493));
  NOR2xp33_ASAP7_75t_L      g08237(.A(new_n8493), .B(new_n8492), .Y(new_n8494));
  NAND3xp33_ASAP7_75t_L     g08238(.A(new_n8488), .B(new_n8485), .C(new_n8494), .Y(new_n8495));
  NAND3xp33_ASAP7_75t_L     g08239(.A(new_n8482), .B(new_n8478), .C(new_n8483), .Y(new_n8496));
  OAI21xp33_ASAP7_75t_L     g08240(.A1(new_n8475), .A2(new_n8476), .B(new_n8281), .Y(new_n8497));
  AOI221xp5_ASAP7_75t_L     g08241(.A1(new_n8497), .A2(new_n8496), .B1(new_n8157), .B2(new_n8171), .C(new_n8274), .Y(new_n8498));
  NAND2xp33_ASAP7_75t_L     g08242(.A(new_n8496), .B(new_n8497), .Y(new_n8499));
  O2A1O1Ixp33_ASAP7_75t_L   g08243(.A1(new_n8151), .A2(new_n8155), .B(new_n8275), .C(new_n8499), .Y(new_n8500));
  INVx1_ASAP7_75t_L         g08244(.A(new_n8494), .Y(new_n8501));
  OAI21xp33_ASAP7_75t_L     g08245(.A1(new_n8498), .A2(new_n8500), .B(new_n8501), .Y(new_n8502));
  NOR2xp33_ASAP7_75t_L      g08246(.A(new_n8173), .B(new_n8172), .Y(new_n8503));
  NAND2xp33_ASAP7_75t_L     g08247(.A(new_n8174), .B(new_n8503), .Y(new_n8504));
  AND4x1_ASAP7_75t_L        g08248(.A(new_n8183), .B(new_n8504), .C(new_n8495), .D(new_n8502), .Y(new_n8505));
  MAJIxp5_ASAP7_75t_L       g08249(.A(new_n8182), .B(new_n8174), .C(new_n8503), .Y(new_n8506));
  AOI21xp33_ASAP7_75t_L     g08250(.A1(new_n8502), .A2(new_n8495), .B(new_n8506), .Y(new_n8507));
  NOR2xp33_ASAP7_75t_L      g08251(.A(new_n5186), .B(new_n1620), .Y(new_n8508));
  INVx1_ASAP7_75t_L         g08252(.A(new_n8508), .Y(new_n8509));
  NAND2xp33_ASAP7_75t_L     g08253(.A(\b[41] ), .B(new_n590), .Y(new_n8510));
  AOI22xp33_ASAP7_75t_L     g08254(.A1(new_n600), .A2(\b[42] ), .B1(new_n597), .B2(new_n5688), .Y(new_n8511));
  AND4x1_ASAP7_75t_L        g08255(.A(new_n8511), .B(new_n8510), .C(new_n8509), .D(\a[11] ), .Y(new_n8512));
  AOI31xp33_ASAP7_75t_L     g08256(.A1(new_n8511), .A2(new_n8510), .A3(new_n8509), .B(\a[11] ), .Y(new_n8513));
  NOR2xp33_ASAP7_75t_L      g08257(.A(new_n8513), .B(new_n8512), .Y(new_n8514));
  OAI21xp33_ASAP7_75t_L     g08258(.A1(new_n8507), .A2(new_n8505), .B(new_n8514), .Y(new_n8515));
  NAND3xp33_ASAP7_75t_L     g08259(.A(new_n8506), .B(new_n8502), .C(new_n8495), .Y(new_n8516));
  NAND2xp33_ASAP7_75t_L     g08260(.A(new_n8495), .B(new_n8502), .Y(new_n8517));
  INVx1_ASAP7_75t_L         g08261(.A(new_n8504), .Y(new_n8518));
  OAI21xp33_ASAP7_75t_L     g08262(.A1(new_n8518), .A2(new_n8192), .B(new_n8517), .Y(new_n8519));
  INVx1_ASAP7_75t_L         g08263(.A(new_n8514), .Y(new_n8520));
  NAND3xp33_ASAP7_75t_L     g08264(.A(new_n8519), .B(new_n8520), .C(new_n8516), .Y(new_n8521));
  NAND2xp33_ASAP7_75t_L     g08265(.A(new_n8515), .B(new_n8521), .Y(new_n8522));
  NAND2xp33_ASAP7_75t_L     g08266(.A(new_n8183), .B(new_n8179), .Y(new_n8523));
  NOR2xp33_ASAP7_75t_L      g08267(.A(new_n8189), .B(new_n8523), .Y(new_n8524));
  INVx1_ASAP7_75t_L         g08268(.A(new_n8524), .Y(new_n8525));
  AOI21xp33_ASAP7_75t_L     g08269(.A1(new_n8210), .A2(new_n8525), .B(new_n8522), .Y(new_n8526));
  AOI21xp33_ASAP7_75t_L     g08270(.A1(new_n8519), .A2(new_n8516), .B(new_n8520), .Y(new_n8527));
  NOR3xp33_ASAP7_75t_L      g08271(.A(new_n8505), .B(new_n8507), .C(new_n8514), .Y(new_n8528));
  NOR2xp33_ASAP7_75t_L      g08272(.A(new_n8528), .B(new_n8527), .Y(new_n8529));
  MAJIxp5_ASAP7_75t_L       g08273(.A(new_n8200), .B(new_n8523), .C(new_n8189), .Y(new_n8530));
  NOR2xp33_ASAP7_75t_L      g08274(.A(new_n8529), .B(new_n8530), .Y(new_n8531));
  NAND2xp33_ASAP7_75t_L     g08275(.A(\b[43] ), .B(new_n480), .Y(new_n8532));
  NAND2xp33_ASAP7_75t_L     g08276(.A(\b[44] ), .B(new_n441), .Y(new_n8533));
  AOI22xp33_ASAP7_75t_L     g08277(.A1(new_n451), .A2(\b[45] ), .B1(new_n448), .B2(new_n6764), .Y(new_n8534));
  AND4x1_ASAP7_75t_L        g08278(.A(new_n8534), .B(new_n8533), .C(new_n8532), .D(\a[8] ), .Y(new_n8535));
  AOI31xp33_ASAP7_75t_L     g08279(.A1(new_n8534), .A2(new_n8533), .A3(new_n8532), .B(\a[8] ), .Y(new_n8536));
  NOR2xp33_ASAP7_75t_L      g08280(.A(new_n8536), .B(new_n8535), .Y(new_n8537));
  INVx1_ASAP7_75t_L         g08281(.A(new_n8537), .Y(new_n8538));
  NOR3xp33_ASAP7_75t_L      g08282(.A(new_n8526), .B(new_n8531), .C(new_n8538), .Y(new_n8539));
  NAND2xp33_ASAP7_75t_L     g08283(.A(new_n8529), .B(new_n8530), .Y(new_n8540));
  AO221x2_ASAP7_75t_L       g08284(.A1(new_n8521), .A2(new_n8515), .B1(new_n8198), .B2(new_n8195), .C(new_n8524), .Y(new_n8541));
  AOI21xp33_ASAP7_75t_L     g08285(.A1(new_n8540), .A2(new_n8541), .B(new_n8537), .Y(new_n8542));
  OAI21xp33_ASAP7_75t_L     g08286(.A1(new_n8211), .A2(new_n7934), .B(new_n8218), .Y(new_n8543));
  OAI21xp33_ASAP7_75t_L     g08287(.A1(new_n8539), .A2(new_n8542), .B(new_n8543), .Y(new_n8544));
  NOR2xp33_ASAP7_75t_L      g08288(.A(new_n8542), .B(new_n8539), .Y(new_n8545));
  A2O1A1O1Ixp25_ASAP7_75t_L g08289(.A1(new_n7885), .A2(new_n7884), .B(new_n8213), .C(new_n8219), .D(new_n8208), .Y(new_n8546));
  NAND2xp33_ASAP7_75t_L     g08290(.A(new_n8546), .B(new_n8545), .Y(new_n8547));
  AOI21xp33_ASAP7_75t_L     g08291(.A1(new_n8547), .A2(new_n8544), .B(new_n8273), .Y(new_n8548));
  INVx1_ASAP7_75t_L         g08292(.A(new_n8273), .Y(new_n8549));
  INVx1_ASAP7_75t_L         g08293(.A(new_n8544), .Y(new_n8550));
  NAND3xp33_ASAP7_75t_L     g08294(.A(new_n8540), .B(new_n8541), .C(new_n8537), .Y(new_n8551));
  OAI21xp33_ASAP7_75t_L     g08295(.A1(new_n8531), .A2(new_n8526), .B(new_n8538), .Y(new_n8552));
  NAND2xp33_ASAP7_75t_L     g08296(.A(new_n8551), .B(new_n8552), .Y(new_n8553));
  NOR2xp33_ASAP7_75t_L      g08297(.A(new_n8543), .B(new_n8553), .Y(new_n8554));
  NOR3xp33_ASAP7_75t_L      g08298(.A(new_n8550), .B(new_n8549), .C(new_n8554), .Y(new_n8555));
  NOR3xp33_ASAP7_75t_L      g08299(.A(new_n8266), .B(new_n8548), .C(new_n8555), .Y(new_n8556));
  INVx1_ASAP7_75t_L         g08300(.A(new_n8266), .Y(new_n8557));
  OAI21xp33_ASAP7_75t_L     g08301(.A1(new_n8554), .A2(new_n8550), .B(new_n8549), .Y(new_n8558));
  NAND3xp33_ASAP7_75t_L     g08302(.A(new_n8547), .B(new_n8544), .C(new_n8273), .Y(new_n8559));
  AOI21xp33_ASAP7_75t_L     g08303(.A1(new_n8559), .A2(new_n8558), .B(new_n8557), .Y(new_n8560));
  NOR3xp33_ASAP7_75t_L      g08304(.A(new_n8560), .B(new_n8556), .C(new_n8262), .Y(new_n8561));
  INVx1_ASAP7_75t_L         g08305(.A(new_n8561), .Y(new_n8562));
  OAI21xp33_ASAP7_75t_L     g08306(.A1(new_n8556), .A2(new_n8560), .B(new_n8262), .Y(new_n8563));
  NAND2xp33_ASAP7_75t_L     g08307(.A(new_n8563), .B(new_n8562), .Y(new_n8564));
  XNOR2x2_ASAP7_75t_L       g08308(.A(new_n8246), .B(new_n8564), .Y(\f[51] ));
  INVx1_ASAP7_75t_L         g08309(.A(new_n8226), .Y(new_n8566));
  A2O1A1O1Ixp25_ASAP7_75t_L g08310(.A1(new_n8239), .A2(new_n8566), .B(new_n8243), .C(new_n8563), .D(new_n8561), .Y(new_n8567));
  NOR2xp33_ASAP7_75t_L      g08311(.A(\b[51] ), .B(\b[52] ), .Y(new_n8568));
  INVx1_ASAP7_75t_L         g08312(.A(\b[52] ), .Y(new_n8569));
  NOR2xp33_ASAP7_75t_L      g08313(.A(new_n8249), .B(new_n8569), .Y(new_n8570));
  NOR2xp33_ASAP7_75t_L      g08314(.A(new_n8568), .B(new_n8570), .Y(new_n8571));
  A2O1A1Ixp33_ASAP7_75t_L   g08315(.A1(\b[51] ), .A2(\b[50] ), .B(new_n8253), .C(new_n8571), .Y(new_n8572));
  INVx1_ASAP7_75t_L         g08316(.A(new_n8250), .Y(new_n8573));
  A2O1A1Ixp33_ASAP7_75t_L   g08317(.A1(new_n8231), .A2(new_n8247), .B(new_n8248), .C(new_n8573), .Y(new_n8574));
  NOR2xp33_ASAP7_75t_L      g08318(.A(new_n8571), .B(new_n8574), .Y(new_n8575));
  INVx1_ASAP7_75t_L         g08319(.A(new_n8575), .Y(new_n8576));
  AND2x2_ASAP7_75t_L        g08320(.A(new_n8572), .B(new_n8576), .Y(new_n8577));
  NOR2xp33_ASAP7_75t_L      g08321(.A(new_n8569), .B(new_n632), .Y(new_n8578));
  AOI221xp5_ASAP7_75t_L     g08322(.A1(new_n380), .A2(\b[51] ), .B1(new_n269), .B2(new_n8577), .C(new_n8578), .Y(new_n8579));
  OA211x2_ASAP7_75t_L       g08323(.A1(new_n277), .A2(new_n8228), .B(new_n8579), .C(\a[2] ), .Y(new_n8580));
  O2A1O1Ixp33_ASAP7_75t_L   g08324(.A1(new_n8228), .A2(new_n277), .B(new_n8579), .C(\a[2] ), .Y(new_n8581));
  NOR2xp33_ASAP7_75t_L      g08325(.A(new_n8581), .B(new_n8580), .Y(new_n8582));
  A2O1A1O1Ixp25_ASAP7_75t_L g08326(.A1(new_n8225), .A2(new_n8223), .B(new_n8265), .C(new_n8558), .D(new_n8555), .Y(new_n8583));
  NAND3xp33_ASAP7_75t_L     g08327(.A(new_n8540), .B(new_n8541), .C(new_n8538), .Y(new_n8584));
  NAND2xp33_ASAP7_75t_L     g08328(.A(\b[45] ), .B(new_n441), .Y(new_n8585));
  OAI221xp5_ASAP7_75t_L     g08329(.A1(new_n667), .A2(new_n7033), .B1(new_n482), .B2(new_n7887), .C(new_n8585), .Y(new_n8586));
  AOI21xp33_ASAP7_75t_L     g08330(.A1(new_n480), .A2(\b[44] ), .B(new_n8586), .Y(new_n8587));
  NAND2xp33_ASAP7_75t_L     g08331(.A(\a[8] ), .B(new_n8587), .Y(new_n8588));
  A2O1A1Ixp33_ASAP7_75t_L   g08332(.A1(\b[44] ), .A2(new_n480), .B(new_n8586), .C(new_n445), .Y(new_n8589));
  NAND2xp33_ASAP7_75t_L     g08333(.A(new_n8589), .B(new_n8588), .Y(new_n8590));
  INVx1_ASAP7_75t_L         g08334(.A(new_n8590), .Y(new_n8591));
  A2O1A1O1Ixp25_ASAP7_75t_L g08335(.A1(new_n8195), .A2(new_n8198), .B(new_n8524), .C(new_n8515), .D(new_n8528), .Y(new_n8592));
  NAND3xp33_ASAP7_75t_L     g08336(.A(new_n8430), .B(new_n8435), .C(new_n8442), .Y(new_n8593));
  NOR2xp33_ASAP7_75t_L      g08337(.A(new_n2852), .B(new_n2234), .Y(new_n8594));
  AOI221xp5_ASAP7_75t_L     g08338(.A1(new_n2232), .A2(\b[27] ), .B1(new_n2226), .B2(new_n2858), .C(new_n8594), .Y(new_n8595));
  OAI211xp5_ASAP7_75t_L     g08339(.A1(new_n2477), .A2(new_n2387), .B(new_n8595), .C(\a[26] ), .Y(new_n8596));
  INVx1_ASAP7_75t_L         g08340(.A(new_n8595), .Y(new_n8597));
  A2O1A1Ixp33_ASAP7_75t_L   g08341(.A1(\b[26] ), .A2(new_n2386), .B(new_n8597), .C(new_n2223), .Y(new_n8598));
  AND2x2_ASAP7_75t_L        g08342(.A(new_n8596), .B(new_n8598), .Y(new_n8599));
  A2O1A1O1Ixp25_ASAP7_75t_L g08343(.A1(new_n8103), .A2(new_n7964), .B(new_n8100), .C(new_n8422), .D(new_n8432), .Y(new_n8600));
  NOR2xp33_ASAP7_75t_L      g08344(.A(new_n8425), .B(new_n8424), .Y(new_n8601));
  NAND2xp33_ASAP7_75t_L     g08345(.A(new_n8401), .B(new_n8399), .Y(new_n8602));
  AO21x2_ASAP7_75t_L        g08346(.A1(new_n8407), .A2(new_n8405), .B(new_n8602), .Y(new_n8603));
  NOR2xp33_ASAP7_75t_L      g08347(.A(new_n1594), .B(new_n3492), .Y(new_n8604));
  NAND2xp33_ASAP7_75t_L     g08348(.A(\b[21] ), .B(new_n3260), .Y(new_n8605));
  OAI221xp5_ASAP7_75t_L     g08349(.A1(new_n3262), .A2(new_n1857), .B1(new_n3261), .B2(new_n1863), .C(new_n8605), .Y(new_n8606));
  OR3x1_ASAP7_75t_L         g08350(.A(new_n8606), .B(new_n3251), .C(new_n8604), .Y(new_n8607));
  A2O1A1Ixp33_ASAP7_75t_L   g08351(.A1(\b[20] ), .A2(new_n3491), .B(new_n8606), .C(new_n3251), .Y(new_n8608));
  AND2x2_ASAP7_75t_L        g08352(.A(new_n8608), .B(new_n8607), .Y(new_n8609));
  OAI21xp33_ASAP7_75t_L     g08353(.A1(new_n8392), .A2(new_n8389), .B(new_n8301), .Y(new_n8610));
  A2O1A1O1Ixp25_ASAP7_75t_L g08354(.A1(new_n7968), .A2(new_n8294), .B(new_n8295), .C(new_n8610), .D(new_n8393), .Y(new_n8611));
  NOR3xp33_ASAP7_75t_L      g08355(.A(new_n8373), .B(new_n8371), .C(new_n8315), .Y(new_n8612));
  INVx1_ASAP7_75t_L         g08356(.A(new_n8612), .Y(new_n8613));
  A2O1A1Ixp33_ASAP7_75t_L   g08357(.A1(new_n8380), .A2(new_n8381), .B(new_n8379), .C(new_n8613), .Y(new_n8614));
  NOR2xp33_ASAP7_75t_L      g08358(.A(new_n695), .B(new_n5521), .Y(new_n8615));
  INVx1_ASAP7_75t_L         g08359(.A(new_n8615), .Y(new_n8616));
  NAND2xp33_ASAP7_75t_L     g08360(.A(\b[12] ), .B(new_n5240), .Y(new_n8617));
  AOI22xp33_ASAP7_75t_L     g08361(.A1(new_n5249), .A2(\b[13] ), .B1(new_n5247), .B2(new_n800), .Y(new_n8618));
  NAND4xp25_ASAP7_75t_L     g08362(.A(new_n8618), .B(\a[41] ), .C(new_n8616), .D(new_n8617), .Y(new_n8619));
  NAND3xp33_ASAP7_75t_L     g08363(.A(new_n8618), .B(new_n8617), .C(new_n8616), .Y(new_n8620));
  NAND2xp33_ASAP7_75t_L     g08364(.A(new_n5244), .B(new_n8620), .Y(new_n8621));
  A2O1A1O1Ixp25_ASAP7_75t_L g08365(.A1(new_n8024), .A2(new_n8034), .B(new_n8316), .C(new_n8365), .D(new_n8361), .Y(new_n8622));
  NOR3xp33_ASAP7_75t_L      g08366(.A(new_n8317), .B(new_n7995), .C(new_n7999), .Y(new_n8623));
  NAND2xp33_ASAP7_75t_L     g08367(.A(new_n8330), .B(new_n8329), .Y(new_n8624));
  MAJx2_ASAP7_75t_L         g08368(.A(new_n8624), .B(new_n8623), .C(new_n8322), .Y(new_n8625));
  NAND2xp33_ASAP7_75t_L     g08369(.A(\b[2] ), .B(new_n7993), .Y(new_n8626));
  NAND2xp33_ASAP7_75t_L     g08370(.A(\b[3] ), .B(new_n7649), .Y(new_n8627));
  AOI22xp33_ASAP7_75t_L     g08371(.A1(new_n7659), .A2(\b[4] ), .B1(new_n7656), .B2(new_n328), .Y(new_n8628));
  NAND4xp25_ASAP7_75t_L     g08372(.A(new_n8628), .B(\a[50] ), .C(new_n8626), .D(new_n8627), .Y(new_n8629));
  AOI31xp33_ASAP7_75t_L     g08373(.A1(new_n8628), .A2(new_n8627), .A3(new_n8626), .B(\a[50] ), .Y(new_n8630));
  INVx1_ASAP7_75t_L         g08374(.A(new_n8630), .Y(new_n8631));
  NAND2xp33_ASAP7_75t_L     g08375(.A(\a[53] ), .B(new_n8322), .Y(new_n8632));
  NAND2xp33_ASAP7_75t_L     g08376(.A(new_n8320), .B(new_n8319), .Y(new_n8633));
  XNOR2x2_ASAP7_75t_L       g08377(.A(\a[52] ), .B(\a[51] ), .Y(new_n8634));
  NOR2xp33_ASAP7_75t_L      g08378(.A(new_n8634), .B(new_n8633), .Y(new_n8635));
  NAND2xp33_ASAP7_75t_L     g08379(.A(\b[0] ), .B(new_n8635), .Y(new_n8636));
  INVx1_ASAP7_75t_L         g08380(.A(\a[52] ), .Y(new_n8637));
  NAND2xp33_ASAP7_75t_L     g08381(.A(\a[53] ), .B(new_n8637), .Y(new_n8638));
  INVx1_ASAP7_75t_L         g08382(.A(\a[53] ), .Y(new_n8639));
  NAND2xp33_ASAP7_75t_L     g08383(.A(\a[52] ), .B(new_n8639), .Y(new_n8640));
  AND2x2_ASAP7_75t_L        g08384(.A(new_n8638), .B(new_n8640), .Y(new_n8641));
  NOR2xp33_ASAP7_75t_L      g08385(.A(new_n8321), .B(new_n8641), .Y(new_n8642));
  NAND2xp33_ASAP7_75t_L     g08386(.A(new_n271), .B(new_n8642), .Y(new_n8643));
  NAND2xp33_ASAP7_75t_L     g08387(.A(new_n8640), .B(new_n8638), .Y(new_n8644));
  NOR2xp33_ASAP7_75t_L      g08388(.A(new_n8644), .B(new_n8321), .Y(new_n8645));
  NAND2xp33_ASAP7_75t_L     g08389(.A(\b[1] ), .B(new_n8645), .Y(new_n8646));
  NAND3xp33_ASAP7_75t_L     g08390(.A(new_n8643), .B(new_n8646), .C(new_n8636), .Y(new_n8647));
  XOR2x2_ASAP7_75t_L        g08391(.A(new_n8632), .B(new_n8647), .Y(new_n8648));
  NAND3xp33_ASAP7_75t_L     g08392(.A(new_n8631), .B(new_n8629), .C(new_n8648), .Y(new_n8649));
  INVx1_ASAP7_75t_L         g08393(.A(new_n8629), .Y(new_n8650));
  XNOR2x2_ASAP7_75t_L       g08394(.A(new_n8632), .B(new_n8647), .Y(new_n8651));
  OAI21xp33_ASAP7_75t_L     g08395(.A1(new_n8630), .A2(new_n8650), .B(new_n8651), .Y(new_n8652));
  NAND3xp33_ASAP7_75t_L     g08396(.A(new_n8625), .B(new_n8649), .C(new_n8652), .Y(new_n8653));
  MAJIxp5_ASAP7_75t_L       g08397(.A(new_n8624), .B(new_n8322), .C(new_n8623), .Y(new_n8654));
  NOR3xp33_ASAP7_75t_L      g08398(.A(new_n8650), .B(new_n8630), .C(new_n8651), .Y(new_n8655));
  AOI21xp33_ASAP7_75t_L     g08399(.A1(new_n8631), .A2(new_n8629), .B(new_n8648), .Y(new_n8656));
  OAI21xp33_ASAP7_75t_L     g08400(.A1(new_n8655), .A2(new_n8656), .B(new_n8654), .Y(new_n8657));
  AOI32xp33_ASAP7_75t_L     g08401(.A1(new_n424), .A2(new_n426), .A3(new_n6819), .B1(new_n6822), .B2(\b[7] ), .Y(new_n8658));
  OAI221xp5_ASAP7_75t_L     g08402(.A1(new_n7392), .A2(new_n382), .B1(new_n353), .B2(new_n7115), .C(new_n8658), .Y(new_n8659));
  NOR2xp33_ASAP7_75t_L      g08403(.A(new_n6816), .B(new_n8659), .Y(new_n8660));
  INVx1_ASAP7_75t_L         g08404(.A(new_n8660), .Y(new_n8661));
  NAND2xp33_ASAP7_75t_L     g08405(.A(new_n6816), .B(new_n8659), .Y(new_n8662));
  NAND4xp25_ASAP7_75t_L     g08406(.A(new_n8653), .B(new_n8661), .C(new_n8662), .D(new_n8657), .Y(new_n8663));
  NOR3xp33_ASAP7_75t_L      g08407(.A(new_n8654), .B(new_n8655), .C(new_n8656), .Y(new_n8664));
  AOI21xp33_ASAP7_75t_L     g08408(.A1(new_n8652), .A2(new_n8649), .B(new_n8625), .Y(new_n8665));
  INVx1_ASAP7_75t_L         g08409(.A(new_n8662), .Y(new_n8666));
  OAI22xp33_ASAP7_75t_L     g08410(.A1(new_n8665), .A2(new_n8664), .B1(new_n8666), .B2(new_n8660), .Y(new_n8667));
  NAND2xp33_ASAP7_75t_L     g08411(.A(new_n8663), .B(new_n8667), .Y(new_n8668));
  AND2x2_ASAP7_75t_L        g08412(.A(new_n8332), .B(new_n8331), .Y(new_n8669));
  NAND2xp33_ASAP7_75t_L     g08413(.A(new_n8336), .B(new_n8338), .Y(new_n8670));
  NAND2xp33_ASAP7_75t_L     g08414(.A(new_n8670), .B(new_n8669), .Y(new_n8671));
  A2O1A1Ixp33_ASAP7_75t_L   g08415(.A1(new_n8356), .A2(new_n8018), .B(new_n8341), .C(new_n8671), .Y(new_n8672));
  NOR2xp33_ASAP7_75t_L      g08416(.A(new_n8672), .B(new_n8668), .Y(new_n8673));
  AND3x1_ASAP7_75t_L        g08417(.A(new_n8670), .B(new_n8332), .C(new_n8331), .Y(new_n8674));
  O2A1O1Ixp33_ASAP7_75t_L   g08418(.A1(new_n8339), .A2(new_n8340), .B(new_n8357), .C(new_n8674), .Y(new_n8675));
  AOI21xp33_ASAP7_75t_L     g08419(.A1(new_n8667), .A2(new_n8663), .B(new_n8675), .Y(new_n8676));
  NAND2xp33_ASAP7_75t_L     g08420(.A(\b[8] ), .B(new_n6308), .Y(new_n8677));
  NAND2xp33_ASAP7_75t_L     g08421(.A(\b[9] ), .B(new_n5992), .Y(new_n8678));
  AOI22xp33_ASAP7_75t_L     g08422(.A1(new_n6002), .A2(\b[10] ), .B1(new_n5999), .B2(new_n852), .Y(new_n8679));
  NAND4xp25_ASAP7_75t_L     g08423(.A(new_n8679), .B(\a[44] ), .C(new_n8677), .D(new_n8678), .Y(new_n8680));
  NAND2xp33_ASAP7_75t_L     g08424(.A(new_n8678), .B(new_n8679), .Y(new_n8681));
  A2O1A1Ixp33_ASAP7_75t_L   g08425(.A1(\b[8] ), .A2(new_n6308), .B(new_n8681), .C(new_n5996), .Y(new_n8682));
  OAI211xp5_ASAP7_75t_L     g08426(.A1(new_n8676), .A2(new_n8673), .B(new_n8680), .C(new_n8682), .Y(new_n8683));
  NAND3xp33_ASAP7_75t_L     g08427(.A(new_n8675), .B(new_n8667), .C(new_n8663), .Y(new_n8684));
  A2O1A1Ixp33_ASAP7_75t_L   g08428(.A1(new_n8670), .A2(new_n8669), .B(new_n8359), .C(new_n8668), .Y(new_n8685));
  NAND2xp33_ASAP7_75t_L     g08429(.A(new_n8680), .B(new_n8682), .Y(new_n8686));
  NAND3xp33_ASAP7_75t_L     g08430(.A(new_n8686), .B(new_n8685), .C(new_n8684), .Y(new_n8687));
  NAND3xp33_ASAP7_75t_L     g08431(.A(new_n8622), .B(new_n8683), .C(new_n8687), .Y(new_n8688));
  AO21x2_ASAP7_75t_L        g08432(.A1(new_n8687), .A2(new_n8683), .B(new_n8622), .Y(new_n8689));
  NAND4xp25_ASAP7_75t_L     g08433(.A(new_n8689), .B(new_n8619), .C(new_n8621), .D(new_n8688), .Y(new_n8690));
  NAND2xp33_ASAP7_75t_L     g08434(.A(new_n8619), .B(new_n8621), .Y(new_n8691));
  AND3x1_ASAP7_75t_L        g08435(.A(new_n8622), .B(new_n8687), .C(new_n8683), .Y(new_n8692));
  AOI21xp33_ASAP7_75t_L     g08436(.A1(new_n8683), .A2(new_n8687), .B(new_n8622), .Y(new_n8693));
  OAI21xp33_ASAP7_75t_L     g08437(.A1(new_n8693), .A2(new_n8692), .B(new_n8691), .Y(new_n8694));
  NAND3xp33_ASAP7_75t_L     g08438(.A(new_n8614), .B(new_n8690), .C(new_n8694), .Y(new_n8695));
  O2A1O1Ixp33_ASAP7_75t_L   g08439(.A1(new_n8374), .A2(new_n8369), .B(new_n8308), .C(new_n8612), .Y(new_n8696));
  NAND2xp33_ASAP7_75t_L     g08440(.A(new_n8690), .B(new_n8694), .Y(new_n8697));
  NAND2xp33_ASAP7_75t_L     g08441(.A(new_n8697), .B(new_n8696), .Y(new_n8698));
  NAND2xp33_ASAP7_75t_L     g08442(.A(\b[14] ), .B(new_n4780), .Y(new_n8699));
  NAND2xp33_ASAP7_75t_L     g08443(.A(\b[15] ), .B(new_n4548), .Y(new_n8700));
  AOI22xp33_ASAP7_75t_L     g08444(.A1(new_n4544), .A2(\b[16] ), .B1(new_n4542), .B2(new_n1058), .Y(new_n8701));
  NAND4xp25_ASAP7_75t_L     g08445(.A(new_n8701), .B(\a[38] ), .C(new_n8699), .D(new_n8700), .Y(new_n8702));
  NAND2xp33_ASAP7_75t_L     g08446(.A(new_n8700), .B(new_n8701), .Y(new_n8703));
  A2O1A1Ixp33_ASAP7_75t_L   g08447(.A1(\b[14] ), .A2(new_n4780), .B(new_n8703), .C(new_n4539), .Y(new_n8704));
  AND2x2_ASAP7_75t_L        g08448(.A(new_n8702), .B(new_n8704), .Y(new_n8705));
  NAND3xp33_ASAP7_75t_L     g08449(.A(new_n8695), .B(new_n8698), .C(new_n8705), .Y(new_n8706));
  AO21x2_ASAP7_75t_L        g08450(.A1(new_n8698), .A2(new_n8695), .B(new_n8705), .Y(new_n8707));
  INVx1_ASAP7_75t_L         g08451(.A(new_n8390), .Y(new_n8708));
  NOR3xp33_ASAP7_75t_L      g08452(.A(new_n8386), .B(new_n8385), .C(new_n8384), .Y(new_n8709));
  A2O1A1O1Ixp25_ASAP7_75t_L g08453(.A1(new_n8059), .A2(new_n8058), .B(new_n8708), .C(new_n8387), .D(new_n8709), .Y(new_n8710));
  NAND3xp33_ASAP7_75t_L     g08454(.A(new_n8707), .B(new_n8710), .C(new_n8706), .Y(new_n8711));
  AO21x2_ASAP7_75t_L        g08455(.A1(new_n8706), .A2(new_n8707), .B(new_n8710), .Y(new_n8712));
  AOI22xp33_ASAP7_75t_L     g08456(.A1(new_n3884), .A2(\b[19] ), .B1(new_n3881), .B2(new_n1499), .Y(new_n8713));
  OAI221xp5_ASAP7_75t_L     g08457(.A1(new_n4312), .A2(new_n1356), .B1(new_n1244), .B2(new_n4986), .C(new_n8713), .Y(new_n8714));
  XNOR2x2_ASAP7_75t_L       g08458(.A(new_n3878), .B(new_n8714), .Y(new_n8715));
  AO21x2_ASAP7_75t_L        g08459(.A1(new_n8711), .A2(new_n8712), .B(new_n8715), .Y(new_n8716));
  NAND3xp33_ASAP7_75t_L     g08460(.A(new_n8712), .B(new_n8711), .C(new_n8715), .Y(new_n8717));
  NAND3xp33_ASAP7_75t_L     g08461(.A(new_n8611), .B(new_n8716), .C(new_n8717), .Y(new_n8718));
  INVx1_ASAP7_75t_L         g08462(.A(new_n8393), .Y(new_n8719));
  OAI21xp33_ASAP7_75t_L     g08463(.A1(new_n8397), .A2(new_n8400), .B(new_n8719), .Y(new_n8720));
  AOI21xp33_ASAP7_75t_L     g08464(.A1(new_n8712), .A2(new_n8711), .B(new_n8715), .Y(new_n8721));
  AND3x1_ASAP7_75t_L        g08465(.A(new_n8712), .B(new_n8715), .C(new_n8711), .Y(new_n8722));
  OAI21xp33_ASAP7_75t_L     g08466(.A1(new_n8721), .A2(new_n8722), .B(new_n8720), .Y(new_n8723));
  AOI21xp33_ASAP7_75t_L     g08467(.A1(new_n8723), .A2(new_n8718), .B(new_n8609), .Y(new_n8724));
  NAND2xp33_ASAP7_75t_L     g08468(.A(new_n8608), .B(new_n8607), .Y(new_n8725));
  AND3x1_ASAP7_75t_L        g08469(.A(new_n8611), .B(new_n8717), .C(new_n8716), .Y(new_n8726));
  AOI21xp33_ASAP7_75t_L     g08470(.A1(new_n8717), .A2(new_n8716), .B(new_n8611), .Y(new_n8727));
  NOR3xp33_ASAP7_75t_L      g08471(.A(new_n8726), .B(new_n8727), .C(new_n8725), .Y(new_n8728));
  OAI221xp5_ASAP7_75t_L     g08472(.A1(new_n8728), .A2(new_n8724), .B1(new_n8411), .B2(new_n8601), .C(new_n8603), .Y(new_n8729));
  MAJIxp5_ASAP7_75t_L       g08473(.A(new_n8411), .B(new_n8408), .C(new_n8602), .Y(new_n8730));
  NOR2xp33_ASAP7_75t_L      g08474(.A(new_n8724), .B(new_n8728), .Y(new_n8731));
  NAND2xp33_ASAP7_75t_L     g08475(.A(new_n8730), .B(new_n8731), .Y(new_n8732));
  NAND2xp33_ASAP7_75t_L     g08476(.A(\b[23] ), .B(new_n2931), .Y(new_n8733));
  NOR2xp33_ASAP7_75t_L      g08477(.A(new_n2180), .B(new_n2708), .Y(new_n8734));
  AOI221xp5_ASAP7_75t_L     g08478(.A1(new_n2706), .A2(\b[24] ), .B1(new_n2700), .B2(new_n2188), .C(new_n8734), .Y(new_n8735));
  AND3x1_ASAP7_75t_L        g08479(.A(new_n8735), .B(new_n8733), .C(\a[29] ), .Y(new_n8736));
  O2A1O1Ixp33_ASAP7_75t_L   g08480(.A1(new_n1995), .A2(new_n2932), .B(new_n8735), .C(\a[29] ), .Y(new_n8737));
  NOR2xp33_ASAP7_75t_L      g08481(.A(new_n8737), .B(new_n8736), .Y(new_n8738));
  NAND3xp33_ASAP7_75t_L     g08482(.A(new_n8732), .B(new_n8729), .C(new_n8738), .Y(new_n8739));
  NOR2xp33_ASAP7_75t_L      g08483(.A(new_n8730), .B(new_n8731), .Y(new_n8740));
  OAI21xp33_ASAP7_75t_L     g08484(.A1(new_n8727), .A2(new_n8726), .B(new_n8725), .Y(new_n8741));
  NAND3xp33_ASAP7_75t_L     g08485(.A(new_n8723), .B(new_n8718), .C(new_n8609), .Y(new_n8742));
  NAND2xp33_ASAP7_75t_L     g08486(.A(new_n8742), .B(new_n8741), .Y(new_n8743));
  O2A1O1Ixp33_ASAP7_75t_L   g08487(.A1(new_n8601), .A2(new_n8411), .B(new_n8603), .C(new_n8743), .Y(new_n8744));
  OR2x4_ASAP7_75t_L         g08488(.A(new_n8737), .B(new_n8736), .Y(new_n8745));
  OAI21xp33_ASAP7_75t_L     g08489(.A1(new_n8740), .A2(new_n8744), .B(new_n8745), .Y(new_n8746));
  AOI21xp33_ASAP7_75t_L     g08490(.A1(new_n8746), .A2(new_n8739), .B(new_n8600), .Y(new_n8747));
  A2O1A1Ixp33_ASAP7_75t_L   g08491(.A1(new_n8433), .A2(new_n7761), .B(new_n7962), .C(new_n8103), .Y(new_n8748));
  A2O1A1Ixp33_ASAP7_75t_L   g08492(.A1(new_n8748), .A2(new_n8104), .B(new_n8431), .C(new_n8428), .Y(new_n8749));
  NOR3xp33_ASAP7_75t_L      g08493(.A(new_n8744), .B(new_n8745), .C(new_n8740), .Y(new_n8750));
  AOI21xp33_ASAP7_75t_L     g08494(.A1(new_n8732), .A2(new_n8729), .B(new_n8738), .Y(new_n8751));
  NOR3xp33_ASAP7_75t_L      g08495(.A(new_n8749), .B(new_n8751), .C(new_n8750), .Y(new_n8752));
  NOR3xp33_ASAP7_75t_L      g08496(.A(new_n8599), .B(new_n8752), .C(new_n8747), .Y(new_n8753));
  NAND2xp33_ASAP7_75t_L     g08497(.A(new_n8596), .B(new_n8598), .Y(new_n8754));
  OAI21xp33_ASAP7_75t_L     g08498(.A1(new_n8750), .A2(new_n8751), .B(new_n8749), .Y(new_n8755));
  NAND3xp33_ASAP7_75t_L     g08499(.A(new_n8600), .B(new_n8739), .C(new_n8746), .Y(new_n8756));
  AOI21xp33_ASAP7_75t_L     g08500(.A1(new_n8756), .A2(new_n8755), .B(new_n8754), .Y(new_n8757));
  OAI221xp5_ASAP7_75t_L     g08501(.A1(new_n8458), .A2(new_n8293), .B1(new_n8753), .B2(new_n8757), .C(new_n8593), .Y(new_n8758));
  A2O1A1Ixp33_ASAP7_75t_L   g08502(.A1(new_n8444), .A2(new_n8447), .B(new_n8293), .C(new_n8593), .Y(new_n8759));
  NAND3xp33_ASAP7_75t_L     g08503(.A(new_n8756), .B(new_n8755), .C(new_n8754), .Y(new_n8760));
  OAI21xp33_ASAP7_75t_L     g08504(.A1(new_n8747), .A2(new_n8752), .B(new_n8599), .Y(new_n8761));
  NAND3xp33_ASAP7_75t_L     g08505(.A(new_n8759), .B(new_n8760), .C(new_n8761), .Y(new_n8762));
  AOI22xp33_ASAP7_75t_L     g08506(.A1(new_n1766), .A2(\b[31] ), .B1(new_n1764), .B2(new_n3426), .Y(new_n8763));
  OAI221xp5_ASAP7_75t_L     g08507(.A1(new_n1758), .A2(new_n3212), .B1(new_n2871), .B2(new_n1911), .C(new_n8763), .Y(new_n8764));
  XNOR2x2_ASAP7_75t_L       g08508(.A(\a[23] ), .B(new_n8764), .Y(new_n8765));
  AND3x1_ASAP7_75t_L        g08509(.A(new_n8762), .B(new_n8758), .C(new_n8765), .Y(new_n8766));
  AOI21xp33_ASAP7_75t_L     g08510(.A1(new_n8762), .A2(new_n8758), .B(new_n8765), .Y(new_n8767));
  NAND3xp33_ASAP7_75t_L     g08511(.A(new_n8455), .B(new_n8459), .C(new_n8454), .Y(new_n8768));
  OAI21xp33_ASAP7_75t_L     g08512(.A1(new_n8460), .A2(new_n8284), .B(new_n8768), .Y(new_n8769));
  NOR3xp33_ASAP7_75t_L      g08513(.A(new_n8769), .B(new_n8767), .C(new_n8766), .Y(new_n8770));
  NAND3xp33_ASAP7_75t_L     g08514(.A(new_n8762), .B(new_n8758), .C(new_n8765), .Y(new_n8771));
  AO21x2_ASAP7_75t_L        g08515(.A1(new_n8758), .A2(new_n8762), .B(new_n8765), .Y(new_n8772));
  OAI21xp33_ASAP7_75t_L     g08516(.A1(new_n8448), .A2(new_n8452), .B(new_n8290), .Y(new_n8773));
  A2O1A1O1Ixp25_ASAP7_75t_L g08517(.A1(new_n8117), .A2(new_n8128), .B(new_n8283), .C(new_n8773), .D(new_n8453), .Y(new_n8774));
  AOI21xp33_ASAP7_75t_L     g08518(.A1(new_n8772), .A2(new_n8771), .B(new_n8774), .Y(new_n8775));
  NAND2xp33_ASAP7_75t_L     g08519(.A(\b[32] ), .B(new_n1548), .Y(new_n8776));
  NAND2xp33_ASAP7_75t_L     g08520(.A(\b[33] ), .B(new_n1410), .Y(new_n8777));
  AOI22xp33_ASAP7_75t_L     g08521(.A1(new_n1406), .A2(\b[34] ), .B1(new_n1404), .B2(new_n3833), .Y(new_n8778));
  NAND4xp25_ASAP7_75t_L     g08522(.A(new_n8778), .B(\a[20] ), .C(new_n8776), .D(new_n8777), .Y(new_n8779));
  NAND2xp33_ASAP7_75t_L     g08523(.A(new_n8777), .B(new_n8778), .Y(new_n8780));
  A2O1A1Ixp33_ASAP7_75t_L   g08524(.A1(\b[32] ), .A2(new_n1548), .B(new_n8780), .C(new_n1401), .Y(new_n8781));
  NAND2xp33_ASAP7_75t_L     g08525(.A(new_n8779), .B(new_n8781), .Y(new_n8782));
  NOR3xp33_ASAP7_75t_L      g08526(.A(new_n8775), .B(new_n8770), .C(new_n8782), .Y(new_n8783));
  NAND3xp33_ASAP7_75t_L     g08527(.A(new_n8774), .B(new_n8772), .C(new_n8771), .Y(new_n8784));
  OAI21xp33_ASAP7_75t_L     g08528(.A1(new_n8767), .A2(new_n8766), .B(new_n8769), .Y(new_n8785));
  INVx1_ASAP7_75t_L         g08529(.A(new_n8782), .Y(new_n8786));
  AOI21xp33_ASAP7_75t_L     g08530(.A1(new_n8784), .A2(new_n8785), .B(new_n8786), .Y(new_n8787));
  NOR2xp33_ASAP7_75t_L      g08531(.A(new_n8787), .B(new_n8783), .Y(new_n8788));
  NOR2xp33_ASAP7_75t_L      g08532(.A(new_n8471), .B(new_n8472), .Y(new_n8789));
  MAJIxp5_ASAP7_75t_L       g08533(.A(new_n8479), .B(new_n8789), .C(new_n8473), .Y(new_n8790));
  NAND2xp33_ASAP7_75t_L     g08534(.A(new_n8790), .B(new_n8788), .Y(new_n8791));
  NAND2xp33_ASAP7_75t_L     g08535(.A(new_n8462), .B(new_n8461), .Y(new_n8792));
  MAJIxp5_ASAP7_75t_L       g08536(.A(new_n8282), .B(new_n8469), .C(new_n8792), .Y(new_n8793));
  OAI21xp33_ASAP7_75t_L     g08537(.A1(new_n8783), .A2(new_n8787), .B(new_n8793), .Y(new_n8794));
  NAND2xp33_ASAP7_75t_L     g08538(.A(\b[35] ), .B(new_n1194), .Y(new_n8795));
  NAND2xp33_ASAP7_75t_L     g08539(.A(\b[36] ), .B(new_n1103), .Y(new_n8796));
  AOI22xp33_ASAP7_75t_L     g08540(.A1(new_n1113), .A2(\b[37] ), .B1(new_n1110), .B2(new_n4709), .Y(new_n8797));
  NAND4xp25_ASAP7_75t_L     g08541(.A(new_n8797), .B(\a[17] ), .C(new_n8795), .D(new_n8796), .Y(new_n8798));
  INVx1_ASAP7_75t_L         g08542(.A(new_n8798), .Y(new_n8799));
  AOI31xp33_ASAP7_75t_L     g08543(.A1(new_n8797), .A2(new_n8796), .A3(new_n8795), .B(\a[17] ), .Y(new_n8800));
  NOR2xp33_ASAP7_75t_L      g08544(.A(new_n8800), .B(new_n8799), .Y(new_n8801));
  NAND3xp33_ASAP7_75t_L     g08545(.A(new_n8791), .B(new_n8794), .C(new_n8801), .Y(new_n8802));
  NOR3xp33_ASAP7_75t_L      g08546(.A(new_n8793), .B(new_n8787), .C(new_n8783), .Y(new_n8803));
  NAND3xp33_ASAP7_75t_L     g08547(.A(new_n8786), .B(new_n8784), .C(new_n8785), .Y(new_n8804));
  OAI21xp33_ASAP7_75t_L     g08548(.A1(new_n8770), .A2(new_n8775), .B(new_n8782), .Y(new_n8805));
  NAND2xp33_ASAP7_75t_L     g08549(.A(new_n8473), .B(new_n8789), .Y(new_n8806));
  AOI22xp33_ASAP7_75t_L     g08550(.A1(new_n8804), .A2(new_n8805), .B1(new_n8806), .B2(new_n8482), .Y(new_n8807));
  INVx1_ASAP7_75t_L         g08551(.A(new_n8800), .Y(new_n8808));
  NAND2xp33_ASAP7_75t_L     g08552(.A(new_n8798), .B(new_n8808), .Y(new_n8809));
  OAI21xp33_ASAP7_75t_L     g08553(.A1(new_n8803), .A2(new_n8807), .B(new_n8809), .Y(new_n8810));
  A2O1A1O1Ixp25_ASAP7_75t_L g08554(.A1(new_n8157), .A2(new_n8171), .B(new_n8274), .C(new_n8497), .D(new_n8477), .Y(new_n8811));
  NAND3xp33_ASAP7_75t_L     g08555(.A(new_n8811), .B(new_n8810), .C(new_n8802), .Y(new_n8812));
  NAND2xp33_ASAP7_75t_L     g08556(.A(new_n8802), .B(new_n8810), .Y(new_n8813));
  A2O1A1Ixp33_ASAP7_75t_L   g08557(.A1(new_n8487), .A2(new_n8486), .B(new_n8477), .C(new_n8813), .Y(new_n8814));
  NAND2xp33_ASAP7_75t_L     g08558(.A(\b[38] ), .B(new_n908), .Y(new_n8815));
  NAND2xp33_ASAP7_75t_L     g08559(.A(\b[39] ), .B(new_n817), .Y(new_n8816));
  AOI22xp33_ASAP7_75t_L     g08560(.A1(new_n826), .A2(\b[40] ), .B1(new_n823), .B2(new_n5194), .Y(new_n8817));
  NAND4xp25_ASAP7_75t_L     g08561(.A(new_n8817), .B(\a[14] ), .C(new_n8815), .D(new_n8816), .Y(new_n8818));
  NAND2xp33_ASAP7_75t_L     g08562(.A(new_n8816), .B(new_n8817), .Y(new_n8819));
  A2O1A1Ixp33_ASAP7_75t_L   g08563(.A1(\b[38] ), .A2(new_n908), .B(new_n8819), .C(new_n813), .Y(new_n8820));
  NAND2xp33_ASAP7_75t_L     g08564(.A(new_n8818), .B(new_n8820), .Y(new_n8821));
  INVx1_ASAP7_75t_L         g08565(.A(new_n8821), .Y(new_n8822));
  NAND3xp33_ASAP7_75t_L     g08566(.A(new_n8814), .B(new_n8822), .C(new_n8812), .Y(new_n8823));
  NOR3xp33_ASAP7_75t_L      g08567(.A(new_n8500), .B(new_n8813), .C(new_n8477), .Y(new_n8824));
  AOI21xp33_ASAP7_75t_L     g08568(.A1(new_n8810), .A2(new_n8802), .B(new_n8811), .Y(new_n8825));
  OAI21xp33_ASAP7_75t_L     g08569(.A1(new_n8825), .A2(new_n8824), .B(new_n8821), .Y(new_n8826));
  NAND2xp33_ASAP7_75t_L     g08570(.A(new_n8823), .B(new_n8826), .Y(new_n8827));
  NOR3xp33_ASAP7_75t_L      g08571(.A(new_n8500), .B(new_n8494), .C(new_n8498), .Y(new_n8828));
  INVx1_ASAP7_75t_L         g08572(.A(new_n8828), .Y(new_n8829));
  A2O1A1Ixp33_ASAP7_75t_L   g08573(.A1(new_n8502), .A2(new_n8495), .B(new_n8506), .C(new_n8829), .Y(new_n8830));
  NOR2xp33_ASAP7_75t_L      g08574(.A(new_n8830), .B(new_n8827), .Y(new_n8831));
  NOR3xp33_ASAP7_75t_L      g08575(.A(new_n8824), .B(new_n8825), .C(new_n8821), .Y(new_n8832));
  AOI21xp33_ASAP7_75t_L     g08576(.A1(new_n8814), .A2(new_n8812), .B(new_n8822), .Y(new_n8833));
  NOR2xp33_ASAP7_75t_L      g08577(.A(new_n8833), .B(new_n8832), .Y(new_n8834));
  NAND2xp33_ASAP7_75t_L     g08578(.A(new_n8175), .B(new_n8167), .Y(new_n8835));
  A2O1A1O1Ixp25_ASAP7_75t_L g08579(.A1(new_n8182), .A2(new_n8835), .B(new_n8518), .C(new_n8517), .D(new_n8828), .Y(new_n8836));
  NOR2xp33_ASAP7_75t_L      g08580(.A(new_n8834), .B(new_n8836), .Y(new_n8837));
  NAND2xp33_ASAP7_75t_L     g08581(.A(\b[42] ), .B(new_n590), .Y(new_n8838));
  AOI22xp33_ASAP7_75t_L     g08582(.A1(new_n600), .A2(\b[43] ), .B1(new_n597), .B2(new_n6202), .Y(new_n8839));
  NAND2xp33_ASAP7_75t_L     g08583(.A(new_n8838), .B(new_n8839), .Y(new_n8840));
  AOI211xp5_ASAP7_75t_L     g08584(.A1(\b[41] ), .A2(new_n674), .B(new_n594), .C(new_n8840), .Y(new_n8841));
  INVx1_ASAP7_75t_L         g08585(.A(new_n8840), .Y(new_n8842));
  O2A1O1Ixp33_ASAP7_75t_L   g08586(.A1(new_n5666), .A2(new_n1620), .B(new_n8842), .C(\a[11] ), .Y(new_n8843));
  NOR2xp33_ASAP7_75t_L      g08587(.A(new_n8841), .B(new_n8843), .Y(new_n8844));
  OAI21xp33_ASAP7_75t_L     g08588(.A1(new_n8831), .A2(new_n8837), .B(new_n8844), .Y(new_n8845));
  NAND2xp33_ASAP7_75t_L     g08589(.A(new_n8834), .B(new_n8836), .Y(new_n8846));
  INVx1_ASAP7_75t_L         g08590(.A(new_n8506), .Y(new_n8847));
  A2O1A1Ixp33_ASAP7_75t_L   g08591(.A1(new_n8517), .A2(new_n8847), .B(new_n8828), .C(new_n8827), .Y(new_n8848));
  OAI211xp5_ASAP7_75t_L     g08592(.A1(new_n8841), .A2(new_n8843), .B(new_n8848), .C(new_n8846), .Y(new_n8849));
  NAND3xp33_ASAP7_75t_L     g08593(.A(new_n8592), .B(new_n8849), .C(new_n8845), .Y(new_n8850));
  AO21x2_ASAP7_75t_L        g08594(.A1(new_n8849), .A2(new_n8845), .B(new_n8592), .Y(new_n8851));
  AOI21xp33_ASAP7_75t_L     g08595(.A1(new_n8851), .A2(new_n8850), .B(new_n8591), .Y(new_n8852));
  AND3x1_ASAP7_75t_L        g08596(.A(new_n8592), .B(new_n8849), .C(new_n8845), .Y(new_n8853));
  AOI21xp33_ASAP7_75t_L     g08597(.A1(new_n8849), .A2(new_n8845), .B(new_n8592), .Y(new_n8854));
  NOR3xp33_ASAP7_75t_L      g08598(.A(new_n8853), .B(new_n8854), .C(new_n8590), .Y(new_n8855));
  OAI221xp5_ASAP7_75t_L     g08599(.A1(new_n8545), .A2(new_n8546), .B1(new_n8852), .B2(new_n8855), .C(new_n8584), .Y(new_n8856));
  NAND2xp33_ASAP7_75t_L     g08600(.A(new_n8541), .B(new_n8540), .Y(new_n8857));
  MAJIxp5_ASAP7_75t_L       g08601(.A(new_n8546), .B(new_n8857), .C(new_n8537), .Y(new_n8858));
  OAI21xp33_ASAP7_75t_L     g08602(.A1(new_n8854), .A2(new_n8853), .B(new_n8590), .Y(new_n8859));
  NAND3xp33_ASAP7_75t_L     g08603(.A(new_n8851), .B(new_n8591), .C(new_n8850), .Y(new_n8860));
  NAND3xp33_ASAP7_75t_L     g08604(.A(new_n8858), .B(new_n8859), .C(new_n8860), .Y(new_n8861));
  NAND2xp33_ASAP7_75t_L     g08605(.A(\b[47] ), .B(new_n366), .Y(new_n8862));
  NAND2xp33_ASAP7_75t_L     g08606(.A(\b[48] ), .B(new_n334), .Y(new_n8863));
  AOI22xp33_ASAP7_75t_L     g08607(.A1(new_n345), .A2(\b[49] ), .B1(new_n342), .B2(new_n7914), .Y(new_n8864));
  AND4x1_ASAP7_75t_L        g08608(.A(new_n8864), .B(new_n8863), .C(new_n8862), .D(\a[5] ), .Y(new_n8865));
  AOI31xp33_ASAP7_75t_L     g08609(.A1(new_n8864), .A2(new_n8863), .A3(new_n8862), .B(\a[5] ), .Y(new_n8866));
  NOR2xp33_ASAP7_75t_L      g08610(.A(new_n8866), .B(new_n8865), .Y(new_n8867));
  NAND3xp33_ASAP7_75t_L     g08611(.A(new_n8861), .B(new_n8856), .C(new_n8867), .Y(new_n8868));
  AO21x2_ASAP7_75t_L        g08612(.A1(new_n8856), .A2(new_n8861), .B(new_n8867), .Y(new_n8869));
  AOI21xp33_ASAP7_75t_L     g08613(.A1(new_n8869), .A2(new_n8868), .B(new_n8583), .Y(new_n8870));
  OAI21xp33_ASAP7_75t_L     g08614(.A1(new_n8263), .A2(new_n8264), .B(new_n8225), .Y(new_n8871));
  INVx1_ASAP7_75t_L         g08615(.A(new_n8265), .Y(new_n8872));
  A2O1A1Ixp33_ASAP7_75t_L   g08616(.A1(new_n8871), .A2(new_n8872), .B(new_n8548), .C(new_n8559), .Y(new_n8873));
  NAND2xp33_ASAP7_75t_L     g08617(.A(new_n8868), .B(new_n8869), .Y(new_n8874));
  NOR2xp33_ASAP7_75t_L      g08618(.A(new_n8873), .B(new_n8874), .Y(new_n8875));
  NOR3xp33_ASAP7_75t_L      g08619(.A(new_n8875), .B(new_n8870), .C(new_n8582), .Y(new_n8876));
  INVx1_ASAP7_75t_L         g08620(.A(new_n8876), .Y(new_n8877));
  OAI21xp33_ASAP7_75t_L     g08621(.A1(new_n8870), .A2(new_n8875), .B(new_n8582), .Y(new_n8878));
  NAND2xp33_ASAP7_75t_L     g08622(.A(new_n8878), .B(new_n8877), .Y(new_n8879));
  XOR2x2_ASAP7_75t_L        g08623(.A(new_n8879), .B(new_n8567), .Y(\f[52] ));
  NOR2xp33_ASAP7_75t_L      g08624(.A(\b[52] ), .B(\b[53] ), .Y(new_n8881));
  INVx1_ASAP7_75t_L         g08625(.A(\b[53] ), .Y(new_n8882));
  NOR2xp33_ASAP7_75t_L      g08626(.A(new_n8569), .B(new_n8882), .Y(new_n8883));
  NOR2xp33_ASAP7_75t_L      g08627(.A(new_n8881), .B(new_n8883), .Y(new_n8884));
  A2O1A1Ixp33_ASAP7_75t_L   g08628(.A1(new_n8574), .A2(new_n8571), .B(new_n8570), .C(new_n8884), .Y(new_n8885));
  O2A1O1Ixp33_ASAP7_75t_L   g08629(.A1(new_n8250), .A2(new_n8253), .B(new_n8571), .C(new_n8570), .Y(new_n8886));
  OAI21xp33_ASAP7_75t_L     g08630(.A1(new_n8881), .A2(new_n8883), .B(new_n8886), .Y(new_n8887));
  NAND2xp33_ASAP7_75t_L     g08631(.A(new_n8887), .B(new_n8885), .Y(new_n8888));
  INVx1_ASAP7_75t_L         g08632(.A(new_n8888), .Y(new_n8889));
  AOI22xp33_ASAP7_75t_L     g08633(.A1(new_n272), .A2(\b[53] ), .B1(new_n269), .B2(new_n8889), .Y(new_n8890));
  OAI221xp5_ASAP7_75t_L     g08634(.A1(new_n261), .A2(new_n8569), .B1(new_n8249), .B2(new_n277), .C(new_n8890), .Y(new_n8891));
  XNOR2x2_ASAP7_75t_L       g08635(.A(\a[2] ), .B(new_n8891), .Y(new_n8892));
  OAI211xp5_ASAP7_75t_L     g08636(.A1(new_n8865), .A2(new_n8866), .B(new_n8861), .C(new_n8856), .Y(new_n8893));
  INVx1_ASAP7_75t_L         g08637(.A(new_n8893), .Y(new_n8894));
  A2O1A1O1Ixp25_ASAP7_75t_L g08638(.A1(new_n8558), .A2(new_n8557), .B(new_n8555), .C(new_n8874), .D(new_n8894), .Y(new_n8895));
  NOR2xp33_ASAP7_75t_L      g08639(.A(new_n6756), .B(new_n481), .Y(new_n8896));
  INVx1_ASAP7_75t_L         g08640(.A(new_n8896), .Y(new_n8897));
  NAND2xp33_ASAP7_75t_L     g08641(.A(\b[46] ), .B(new_n441), .Y(new_n8898));
  AOI22xp33_ASAP7_75t_L     g08642(.A1(new_n451), .A2(\b[47] ), .B1(new_n448), .B2(new_n7323), .Y(new_n8899));
  AND4x1_ASAP7_75t_L        g08643(.A(new_n8899), .B(new_n8898), .C(new_n8897), .D(\a[8] ), .Y(new_n8900));
  AOI31xp33_ASAP7_75t_L     g08644(.A1(new_n8899), .A2(new_n8898), .A3(new_n8897), .B(\a[8] ), .Y(new_n8901));
  NOR2xp33_ASAP7_75t_L      g08645(.A(new_n8901), .B(new_n8900), .Y(new_n8902));
  NAND2xp33_ASAP7_75t_L     g08646(.A(new_n8758), .B(new_n8762), .Y(new_n8903));
  MAJIxp5_ASAP7_75t_L       g08647(.A(new_n8774), .B(new_n8903), .C(new_n8765), .Y(new_n8904));
  NOR2xp33_ASAP7_75t_L      g08648(.A(new_n3212), .B(new_n1911), .Y(new_n8905));
  INVx1_ASAP7_75t_L         g08649(.A(new_n8905), .Y(new_n8906));
  NAND2xp33_ASAP7_75t_L     g08650(.A(\b[31] ), .B(new_n1770), .Y(new_n8907));
  AOI22xp33_ASAP7_75t_L     g08651(.A1(new_n1766), .A2(\b[32] ), .B1(new_n1764), .B2(new_n3450), .Y(new_n8908));
  AND4x1_ASAP7_75t_L        g08652(.A(new_n8908), .B(new_n8907), .C(new_n8906), .D(\a[23] ), .Y(new_n8909));
  AOI31xp33_ASAP7_75t_L     g08653(.A1(new_n8908), .A2(new_n8907), .A3(new_n8906), .B(\a[23] ), .Y(new_n8910));
  NOR2xp33_ASAP7_75t_L      g08654(.A(new_n8910), .B(new_n8909), .Y(new_n8911));
  NOR3xp33_ASAP7_75t_L      g08655(.A(new_n8446), .B(new_n8445), .C(new_n8443), .Y(new_n8912));
  A2O1A1O1Ixp25_ASAP7_75t_L g08656(.A1(new_n8450), .A2(new_n8451), .B(new_n8912), .C(new_n8761), .D(new_n8753), .Y(new_n8913));
  OAI22xp33_ASAP7_75t_L     g08657(.A1(new_n2881), .A2(new_n2233), .B1(new_n2871), .B2(new_n2234), .Y(new_n8914));
  AOI21xp33_ASAP7_75t_L     g08658(.A1(new_n2232), .A2(\b[28] ), .B(new_n8914), .Y(new_n8915));
  OA211x2_ASAP7_75t_L       g08659(.A1(new_n2387), .A2(new_n2650), .B(new_n8915), .C(\a[26] ), .Y(new_n8916));
  O2A1O1Ixp33_ASAP7_75t_L   g08660(.A1(new_n2650), .A2(new_n2387), .B(new_n8915), .C(\a[26] ), .Y(new_n8917));
  NOR2xp33_ASAP7_75t_L      g08661(.A(new_n8917), .B(new_n8916), .Y(new_n8918));
  INVx1_ASAP7_75t_L         g08662(.A(new_n8918), .Y(new_n8919));
  NAND2xp33_ASAP7_75t_L     g08663(.A(new_n8729), .B(new_n8732), .Y(new_n8920));
  MAJIxp5_ASAP7_75t_L       g08664(.A(new_n8600), .B(new_n8920), .C(new_n8738), .Y(new_n8921));
  OAI22xp33_ASAP7_75t_L     g08665(.A1(new_n2487), .A2(new_n2707), .B1(new_n2708), .B2(new_n2477), .Y(new_n8922));
  AOI221xp5_ASAP7_75t_L     g08666(.A1(\b[24] ), .A2(new_n2931), .B1(\b[25] ), .B2(new_n2706), .C(new_n8922), .Y(new_n8923));
  XNOR2x2_ASAP7_75t_L       g08667(.A(new_n2697), .B(new_n8923), .Y(new_n8924));
  NOR2xp33_ASAP7_75t_L      g08668(.A(new_n8408), .B(new_n8602), .Y(new_n8925));
  O2A1O1Ixp33_ASAP7_75t_L   g08669(.A1(new_n8424), .A2(new_n8425), .B(new_n8426), .C(new_n8925), .Y(new_n8926));
  AOI32xp33_ASAP7_75t_L     g08670(.A1(new_n1998), .A2(new_n2001), .A3(new_n3254), .B1(new_n3256), .B2(\b[23] ), .Y(new_n8927));
  OAI221xp5_ASAP7_75t_L     g08671(.A1(new_n3248), .A2(new_n1857), .B1(new_n1709), .B2(new_n3492), .C(new_n8927), .Y(new_n8928));
  XNOR2x2_ASAP7_75t_L       g08672(.A(\a[32] ), .B(new_n8928), .Y(new_n8929));
  XNOR2x2_ASAP7_75t_L       g08673(.A(new_n8697), .B(new_n8696), .Y(new_n8930));
  MAJIxp5_ASAP7_75t_L       g08674(.A(new_n8710), .B(new_n8705), .C(new_n8930), .Y(new_n8931));
  NAND2xp33_ASAP7_75t_L     g08675(.A(\b[16] ), .B(new_n4548), .Y(new_n8932));
  OAI221xp5_ASAP7_75t_L     g08676(.A1(new_n4550), .A2(new_n1244), .B1(new_n4549), .B2(new_n1251), .C(new_n8932), .Y(new_n8933));
  AOI21xp33_ASAP7_75t_L     g08677(.A1(new_n4780), .A2(\b[15] ), .B(new_n8933), .Y(new_n8934));
  NAND2xp33_ASAP7_75t_L     g08678(.A(\a[38] ), .B(new_n8934), .Y(new_n8935));
  A2O1A1Ixp33_ASAP7_75t_L   g08679(.A1(\b[15] ), .A2(new_n4780), .B(new_n8933), .C(new_n4539), .Y(new_n8936));
  NAND2xp33_ASAP7_75t_L     g08680(.A(new_n8936), .B(new_n8935), .Y(new_n8937));
  INVx1_ASAP7_75t_L         g08681(.A(new_n8694), .Y(new_n8938));
  O2A1O1Ixp33_ASAP7_75t_L   g08682(.A1(new_n8612), .A2(new_n8385), .B(new_n8690), .C(new_n8938), .Y(new_n8939));
  NOR2xp33_ASAP7_75t_L      g08683(.A(new_n559), .B(new_n6309), .Y(new_n8940));
  NAND2xp33_ASAP7_75t_L     g08684(.A(\b[10] ), .B(new_n5992), .Y(new_n8941));
  OAI221xp5_ASAP7_75t_L     g08685(.A1(new_n6312), .A2(new_n695), .B1(new_n6311), .B2(new_n701), .C(new_n8941), .Y(new_n8942));
  OR3x1_ASAP7_75t_L         g08686(.A(new_n8942), .B(new_n5996), .C(new_n8940), .Y(new_n8943));
  A2O1A1Ixp33_ASAP7_75t_L   g08687(.A1(\b[9] ), .A2(new_n6308), .B(new_n8942), .C(new_n5996), .Y(new_n8944));
  AND2x2_ASAP7_75t_L        g08688(.A(new_n8944), .B(new_n8943), .Y(new_n8945));
  OAI211xp5_ASAP7_75t_L     g08689(.A1(new_n8660), .A2(new_n8666), .B(new_n8653), .C(new_n8657), .Y(new_n8946));
  INVx1_ASAP7_75t_L         g08690(.A(new_n8946), .Y(new_n8947));
  O2A1O1Ixp33_ASAP7_75t_L   g08691(.A1(new_n8359), .A2(new_n8674), .B(new_n8668), .C(new_n8947), .Y(new_n8948));
  NAND2xp33_ASAP7_75t_L     g08692(.A(\b[7] ), .B(new_n6812), .Y(new_n8949));
  OAI221xp5_ASAP7_75t_L     g08693(.A1(new_n7118), .A2(new_n503), .B1(new_n7117), .B2(new_n509), .C(new_n8949), .Y(new_n8950));
  AOI21xp33_ASAP7_75t_L     g08694(.A1(new_n7124), .A2(\b[6] ), .B(new_n8950), .Y(new_n8951));
  NAND2xp33_ASAP7_75t_L     g08695(.A(\a[47] ), .B(new_n8951), .Y(new_n8952));
  A2O1A1Ixp33_ASAP7_75t_L   g08696(.A1(\b[6] ), .A2(new_n7124), .B(new_n8950), .C(new_n6816), .Y(new_n8953));
  AOI22xp33_ASAP7_75t_L     g08697(.A1(new_n8329), .A2(new_n8330), .B1(new_n8323), .B2(new_n8325), .Y(new_n8954));
  A2O1A1O1Ixp25_ASAP7_75t_L g08698(.A1(new_n8623), .A2(new_n8322), .B(new_n8954), .C(new_n8649), .D(new_n8656), .Y(new_n8955));
  NAND2xp33_ASAP7_75t_L     g08699(.A(\b[4] ), .B(new_n7649), .Y(new_n8956));
  OAI221xp5_ASAP7_75t_L     g08700(.A1(new_n7997), .A2(new_n353), .B1(new_n7996), .B2(new_n359), .C(new_n8956), .Y(new_n8957));
  AOI211xp5_ASAP7_75t_L     g08701(.A1(\b[3] ), .A2(new_n7993), .B(new_n7653), .C(new_n8957), .Y(new_n8958));
  NOR2xp33_ASAP7_75t_L      g08702(.A(new_n299), .B(new_n7994), .Y(new_n8959));
  OA21x2_ASAP7_75t_L        g08703(.A1(new_n8959), .A2(new_n8957), .B(new_n7653), .Y(new_n8960));
  NOR2xp33_ASAP7_75t_L      g08704(.A(new_n8958), .B(new_n8960), .Y(new_n8961));
  AND3x1_ASAP7_75t_L        g08705(.A(new_n8643), .B(new_n8646), .C(new_n8636), .Y(new_n8962));
  INVx1_ASAP7_75t_L         g08706(.A(new_n8634), .Y(new_n8963));
  NOR3xp33_ASAP7_75t_L      g08707(.A(new_n8641), .B(new_n8963), .C(new_n8633), .Y(new_n8964));
  INVx1_ASAP7_75t_L         g08708(.A(new_n8964), .Y(new_n8965));
  NOR2xp33_ASAP7_75t_L      g08709(.A(new_n258), .B(new_n8965), .Y(new_n8966));
  NAND2xp33_ASAP7_75t_L     g08710(.A(new_n8644), .B(new_n8633), .Y(new_n8967));
  NAND2xp33_ASAP7_75t_L     g08711(.A(new_n8633), .B(new_n8641), .Y(new_n8968));
  NAND2xp33_ASAP7_75t_L     g08712(.A(\b[1] ), .B(new_n8635), .Y(new_n8969));
  OAI221xp5_ASAP7_75t_L     g08713(.A1(new_n8967), .A2(new_n283), .B1(new_n278), .B2(new_n8968), .C(new_n8969), .Y(new_n8970));
  NOR2xp33_ASAP7_75t_L      g08714(.A(new_n8970), .B(new_n8966), .Y(new_n8971));
  A2O1A1Ixp33_ASAP7_75t_L   g08715(.A1(new_n8324), .A2(new_n8962), .B(new_n8639), .C(new_n8971), .Y(new_n8972));
  INVx1_ASAP7_75t_L         g08716(.A(new_n8972), .Y(new_n8973));
  A2O1A1Ixp33_ASAP7_75t_L   g08717(.A1(\b[0] ), .A2(new_n8633), .B(new_n8647), .C(\a[53] ), .Y(new_n8974));
  INVx1_ASAP7_75t_L         g08718(.A(new_n8970), .Y(new_n8975));
  O2A1O1Ixp33_ASAP7_75t_L   g08719(.A1(new_n8965), .A2(new_n258), .B(new_n8975), .C(new_n8974), .Y(new_n8976));
  OAI21xp33_ASAP7_75t_L     g08720(.A1(new_n8973), .A2(new_n8976), .B(new_n8961), .Y(new_n8977));
  O2A1O1Ixp33_ASAP7_75t_L   g08721(.A1(new_n258), .A2(new_n8321), .B(new_n8962), .C(new_n8639), .Y(new_n8978));
  A2O1A1Ixp33_ASAP7_75t_L   g08722(.A1(\b[0] ), .A2(new_n8964), .B(new_n8970), .C(new_n8978), .Y(new_n8979));
  OAI211xp5_ASAP7_75t_L     g08723(.A1(new_n8958), .A2(new_n8960), .B(new_n8979), .C(new_n8972), .Y(new_n8980));
  NAND3xp33_ASAP7_75t_L     g08724(.A(new_n8955), .B(new_n8980), .C(new_n8977), .Y(new_n8981));
  NAND2xp33_ASAP7_75t_L     g08725(.A(new_n8980), .B(new_n8977), .Y(new_n8982));
  A2O1A1Ixp33_ASAP7_75t_L   g08726(.A1(new_n8649), .A2(new_n8625), .B(new_n8656), .C(new_n8982), .Y(new_n8983));
  NAND4xp25_ASAP7_75t_L     g08727(.A(new_n8983), .B(new_n8952), .C(new_n8981), .D(new_n8953), .Y(new_n8984));
  AO22x1_ASAP7_75t_L        g08728(.A1(new_n8953), .A2(new_n8952), .B1(new_n8981), .B2(new_n8983), .Y(new_n8985));
  NAND2xp33_ASAP7_75t_L     g08729(.A(new_n8984), .B(new_n8985), .Y(new_n8986));
  NOR2xp33_ASAP7_75t_L      g08730(.A(new_n8986), .B(new_n8948), .Y(new_n8987));
  A2O1A1Ixp33_ASAP7_75t_L   g08731(.A1(new_n8667), .A2(new_n8663), .B(new_n8675), .C(new_n8946), .Y(new_n8988));
  AND4x1_ASAP7_75t_L        g08732(.A(new_n8952), .B(new_n8983), .C(new_n8981), .D(new_n8953), .Y(new_n8989));
  AOI22xp33_ASAP7_75t_L     g08733(.A1(new_n8952), .A2(new_n8953), .B1(new_n8981), .B2(new_n8983), .Y(new_n8990));
  NOR2xp33_ASAP7_75t_L      g08734(.A(new_n8990), .B(new_n8989), .Y(new_n8991));
  NOR2xp33_ASAP7_75t_L      g08735(.A(new_n8988), .B(new_n8991), .Y(new_n8992));
  OAI21xp33_ASAP7_75t_L     g08736(.A1(new_n8992), .A2(new_n8987), .B(new_n8945), .Y(new_n8993));
  NAND2xp33_ASAP7_75t_L     g08737(.A(new_n8944), .B(new_n8943), .Y(new_n8994));
  A2O1A1Ixp33_ASAP7_75t_L   g08738(.A1(new_n8672), .A2(new_n8668), .B(new_n8947), .C(new_n8991), .Y(new_n8995));
  NAND2xp33_ASAP7_75t_L     g08739(.A(new_n8986), .B(new_n8948), .Y(new_n8996));
  NAND3xp33_ASAP7_75t_L     g08740(.A(new_n8995), .B(new_n8996), .C(new_n8994), .Y(new_n8997));
  AOI21xp33_ASAP7_75t_L     g08741(.A1(new_n8685), .A2(new_n8684), .B(new_n8686), .Y(new_n8998));
  OAI21xp33_ASAP7_75t_L     g08742(.A1(new_n8998), .A2(new_n8622), .B(new_n8687), .Y(new_n8999));
  NAND3xp33_ASAP7_75t_L     g08743(.A(new_n8999), .B(new_n8997), .C(new_n8993), .Y(new_n9000));
  AOI21xp33_ASAP7_75t_L     g08744(.A1(new_n8995), .A2(new_n8996), .B(new_n8994), .Y(new_n9001));
  NOR3xp33_ASAP7_75t_L      g08745(.A(new_n8945), .B(new_n8987), .C(new_n8992), .Y(new_n9002));
  A2O1A1Ixp33_ASAP7_75t_L   g08746(.A1(new_n8372), .A2(new_n8365), .B(new_n8361), .C(new_n8683), .Y(new_n9003));
  OAI211xp5_ASAP7_75t_L     g08747(.A1(new_n9001), .A2(new_n9002), .B(new_n8687), .C(new_n9003), .Y(new_n9004));
  NAND2xp33_ASAP7_75t_L     g08748(.A(\b[12] ), .B(new_n5526), .Y(new_n9005));
  NAND2xp33_ASAP7_75t_L     g08749(.A(\b[13] ), .B(new_n5240), .Y(new_n9006));
  AOI32xp33_ASAP7_75t_L     g08750(.A1(new_n877), .A2(new_n874), .A3(new_n5247), .B1(\b[14] ), .B2(new_n5249), .Y(new_n9007));
  AND4x1_ASAP7_75t_L        g08751(.A(new_n9007), .B(new_n9006), .C(new_n9005), .D(\a[41] ), .Y(new_n9008));
  AOI31xp33_ASAP7_75t_L     g08752(.A1(new_n9007), .A2(new_n9006), .A3(new_n9005), .B(\a[41] ), .Y(new_n9009));
  NOR2xp33_ASAP7_75t_L      g08753(.A(new_n9009), .B(new_n9008), .Y(new_n9010));
  NAND3xp33_ASAP7_75t_L     g08754(.A(new_n9004), .B(new_n9000), .C(new_n9010), .Y(new_n9011));
  AND3x1_ASAP7_75t_L        g08755(.A(new_n8999), .B(new_n8997), .C(new_n8993), .Y(new_n9012));
  AOI21xp33_ASAP7_75t_L     g08756(.A1(new_n8997), .A2(new_n8993), .B(new_n8999), .Y(new_n9013));
  INVx1_ASAP7_75t_L         g08757(.A(new_n9010), .Y(new_n9014));
  OAI21xp33_ASAP7_75t_L     g08758(.A1(new_n9013), .A2(new_n9012), .B(new_n9014), .Y(new_n9015));
  AOI21xp33_ASAP7_75t_L     g08759(.A1(new_n9015), .A2(new_n9011), .B(new_n8939), .Y(new_n9016));
  A2O1A1Ixp33_ASAP7_75t_L   g08760(.A1(new_n8375), .A2(new_n8613), .B(new_n8697), .C(new_n8694), .Y(new_n9017));
  NAND2xp33_ASAP7_75t_L     g08761(.A(new_n9011), .B(new_n9015), .Y(new_n9018));
  NOR2xp33_ASAP7_75t_L      g08762(.A(new_n9018), .B(new_n9017), .Y(new_n9019));
  OAI21xp33_ASAP7_75t_L     g08763(.A1(new_n9019), .A2(new_n9016), .B(new_n8937), .Y(new_n9020));
  A2O1A1Ixp33_ASAP7_75t_L   g08764(.A1(new_n8690), .A2(new_n8614), .B(new_n8938), .C(new_n9018), .Y(new_n9021));
  NAND3xp33_ASAP7_75t_L     g08765(.A(new_n8939), .B(new_n9011), .C(new_n9015), .Y(new_n9022));
  NAND4xp25_ASAP7_75t_L     g08766(.A(new_n9022), .B(new_n9021), .C(new_n8935), .D(new_n8936), .Y(new_n9023));
  NAND3xp33_ASAP7_75t_L     g08767(.A(new_n8931), .B(new_n9023), .C(new_n9020), .Y(new_n9024));
  AO21x2_ASAP7_75t_L        g08768(.A1(new_n9023), .A2(new_n9020), .B(new_n8931), .Y(new_n9025));
  NOR2xp33_ASAP7_75t_L      g08769(.A(new_n1594), .B(new_n4115), .Y(new_n9026));
  AOI221xp5_ASAP7_75t_L     g08770(.A1(new_n3874), .A2(\b[19] ), .B1(new_n3881), .B2(new_n1600), .C(new_n9026), .Y(new_n9027));
  OA211x2_ASAP7_75t_L       g08771(.A1(new_n4986), .A2(new_n1356), .B(new_n9027), .C(\a[35] ), .Y(new_n9028));
  O2A1O1Ixp33_ASAP7_75t_L   g08772(.A1(new_n1356), .A2(new_n4986), .B(new_n9027), .C(\a[35] ), .Y(new_n9029));
  NOR2xp33_ASAP7_75t_L      g08773(.A(new_n9029), .B(new_n9028), .Y(new_n9030));
  AO21x2_ASAP7_75t_L        g08774(.A1(new_n9024), .A2(new_n9025), .B(new_n9030), .Y(new_n9031));
  NAND3xp33_ASAP7_75t_L     g08775(.A(new_n9025), .B(new_n9030), .C(new_n9024), .Y(new_n9032));
  OAI21xp33_ASAP7_75t_L     g08776(.A1(new_n8721), .A2(new_n8611), .B(new_n8717), .Y(new_n9033));
  NAND3xp33_ASAP7_75t_L     g08777(.A(new_n9033), .B(new_n9032), .C(new_n9031), .Y(new_n9034));
  AOI21xp33_ASAP7_75t_L     g08778(.A1(new_n9025), .A2(new_n9024), .B(new_n9030), .Y(new_n9035));
  AND3x1_ASAP7_75t_L        g08779(.A(new_n9025), .B(new_n9030), .C(new_n9024), .Y(new_n9036));
  NOR2xp33_ASAP7_75t_L      g08780(.A(new_n8070), .B(new_n8071), .Y(new_n9037));
  INVx1_ASAP7_75t_L         g08781(.A(new_n8295), .Y(new_n9038));
  A2O1A1Ixp33_ASAP7_75t_L   g08782(.A1(new_n7967), .A2(new_n7729), .B(new_n9037), .C(new_n9038), .Y(new_n9039));
  A2O1A1O1Ixp25_ASAP7_75t_L g08783(.A1(new_n8610), .A2(new_n9039), .B(new_n8393), .C(new_n8716), .D(new_n8722), .Y(new_n9040));
  OAI21xp33_ASAP7_75t_L     g08784(.A1(new_n9035), .A2(new_n9036), .B(new_n9040), .Y(new_n9041));
  AOI21xp33_ASAP7_75t_L     g08785(.A1(new_n9041), .A2(new_n9034), .B(new_n8929), .Y(new_n9042));
  AND3x1_ASAP7_75t_L        g08786(.A(new_n9041), .B(new_n9034), .C(new_n8929), .Y(new_n9043));
  NOR2xp33_ASAP7_75t_L      g08787(.A(new_n9042), .B(new_n9043), .Y(new_n9044));
  O2A1O1Ixp33_ASAP7_75t_L   g08788(.A1(new_n8926), .A2(new_n8728), .B(new_n8741), .C(new_n9044), .Y(new_n9045));
  AO21x2_ASAP7_75t_L        g08789(.A1(new_n8742), .A2(new_n8730), .B(new_n8724), .Y(new_n9046));
  AO21x2_ASAP7_75t_L        g08790(.A1(new_n9034), .A2(new_n9041), .B(new_n8929), .Y(new_n9047));
  NAND3xp33_ASAP7_75t_L     g08791(.A(new_n9041), .B(new_n9034), .C(new_n8929), .Y(new_n9048));
  NAND2xp33_ASAP7_75t_L     g08792(.A(new_n9048), .B(new_n9047), .Y(new_n9049));
  NOR2xp33_ASAP7_75t_L      g08793(.A(new_n9049), .B(new_n9046), .Y(new_n9050));
  OAI21xp33_ASAP7_75t_L     g08794(.A1(new_n9045), .A2(new_n9050), .B(new_n8924), .Y(new_n9051));
  INVx1_ASAP7_75t_L         g08795(.A(new_n8924), .Y(new_n9052));
  A2O1A1Ixp33_ASAP7_75t_L   g08796(.A1(new_n8742), .A2(new_n8730), .B(new_n8724), .C(new_n9049), .Y(new_n9053));
  O2A1O1Ixp33_ASAP7_75t_L   g08797(.A1(new_n8925), .A2(new_n8413), .B(new_n8742), .C(new_n8724), .Y(new_n9054));
  NAND2xp33_ASAP7_75t_L     g08798(.A(new_n9044), .B(new_n9054), .Y(new_n9055));
  NAND3xp33_ASAP7_75t_L     g08799(.A(new_n9052), .B(new_n9053), .C(new_n9055), .Y(new_n9056));
  NAND3xp33_ASAP7_75t_L     g08800(.A(new_n8921), .B(new_n9051), .C(new_n9056), .Y(new_n9057));
  AOI21xp33_ASAP7_75t_L     g08801(.A1(new_n9056), .A2(new_n9051), .B(new_n8921), .Y(new_n9058));
  INVx1_ASAP7_75t_L         g08802(.A(new_n9058), .Y(new_n9059));
  AOI21xp33_ASAP7_75t_L     g08803(.A1(new_n9059), .A2(new_n9057), .B(new_n8919), .Y(new_n9060));
  NOR2xp33_ASAP7_75t_L      g08804(.A(new_n8740), .B(new_n8744), .Y(new_n9061));
  MAJIxp5_ASAP7_75t_L       g08805(.A(new_n8749), .B(new_n8745), .C(new_n9061), .Y(new_n9062));
  AOI21xp33_ASAP7_75t_L     g08806(.A1(new_n9053), .A2(new_n9055), .B(new_n9052), .Y(new_n9063));
  NOR3xp33_ASAP7_75t_L      g08807(.A(new_n9050), .B(new_n9045), .C(new_n8924), .Y(new_n9064));
  NOR3xp33_ASAP7_75t_L      g08808(.A(new_n9062), .B(new_n9063), .C(new_n9064), .Y(new_n9065));
  NOR3xp33_ASAP7_75t_L      g08809(.A(new_n9065), .B(new_n9058), .C(new_n8918), .Y(new_n9066));
  NOR3xp33_ASAP7_75t_L      g08810(.A(new_n9060), .B(new_n9066), .C(new_n8913), .Y(new_n9067));
  AO21x2_ASAP7_75t_L        g08811(.A1(new_n8761), .A2(new_n8759), .B(new_n8753), .Y(new_n9068));
  OAI21xp33_ASAP7_75t_L     g08812(.A1(new_n9058), .A2(new_n9065), .B(new_n8918), .Y(new_n9069));
  INVx1_ASAP7_75t_L         g08813(.A(new_n9066), .Y(new_n9070));
  AOI21xp33_ASAP7_75t_L     g08814(.A1(new_n9070), .A2(new_n9069), .B(new_n9068), .Y(new_n9071));
  OAI21xp33_ASAP7_75t_L     g08815(.A1(new_n9067), .A2(new_n9071), .B(new_n8911), .Y(new_n9072));
  INVx1_ASAP7_75t_L         g08816(.A(new_n8911), .Y(new_n9073));
  NAND3xp33_ASAP7_75t_L     g08817(.A(new_n9068), .B(new_n9070), .C(new_n9069), .Y(new_n9074));
  OAI21xp33_ASAP7_75t_L     g08818(.A1(new_n9066), .A2(new_n9060), .B(new_n8913), .Y(new_n9075));
  NAND3xp33_ASAP7_75t_L     g08819(.A(new_n9074), .B(new_n9073), .C(new_n9075), .Y(new_n9076));
  NAND3xp33_ASAP7_75t_L     g08820(.A(new_n8904), .B(new_n9072), .C(new_n9076), .Y(new_n9077));
  NAND2xp33_ASAP7_75t_L     g08821(.A(new_n8760), .B(new_n8761), .Y(new_n9078));
  XNOR2x2_ASAP7_75t_L       g08822(.A(new_n8759), .B(new_n9078), .Y(new_n9079));
  INVx1_ASAP7_75t_L         g08823(.A(new_n8765), .Y(new_n9080));
  MAJIxp5_ASAP7_75t_L       g08824(.A(new_n8769), .B(new_n9080), .C(new_n9079), .Y(new_n9081));
  AOI21xp33_ASAP7_75t_L     g08825(.A1(new_n9074), .A2(new_n9075), .B(new_n9073), .Y(new_n9082));
  NOR3xp33_ASAP7_75t_L      g08826(.A(new_n9071), .B(new_n9067), .C(new_n8911), .Y(new_n9083));
  OAI21xp33_ASAP7_75t_L     g08827(.A1(new_n9083), .A2(new_n9082), .B(new_n9081), .Y(new_n9084));
  NOR2xp33_ASAP7_75t_L      g08828(.A(new_n3807), .B(new_n1549), .Y(new_n9085));
  INVx1_ASAP7_75t_L         g08829(.A(new_n9085), .Y(new_n9086));
  NAND2xp33_ASAP7_75t_L     g08830(.A(\b[34] ), .B(new_n1410), .Y(new_n9087));
  AOI22xp33_ASAP7_75t_L     g08831(.A1(new_n1406), .A2(\b[35] ), .B1(new_n1404), .B2(new_n5649), .Y(new_n9088));
  AND4x1_ASAP7_75t_L        g08832(.A(new_n9088), .B(new_n9087), .C(new_n9086), .D(\a[20] ), .Y(new_n9089));
  AOI31xp33_ASAP7_75t_L     g08833(.A1(new_n9088), .A2(new_n9087), .A3(new_n9086), .B(\a[20] ), .Y(new_n9090));
  NOR2xp33_ASAP7_75t_L      g08834(.A(new_n9090), .B(new_n9089), .Y(new_n9091));
  NAND3xp33_ASAP7_75t_L     g08835(.A(new_n9077), .B(new_n9084), .C(new_n9091), .Y(new_n9092));
  NOR3xp33_ASAP7_75t_L      g08836(.A(new_n9081), .B(new_n9082), .C(new_n9083), .Y(new_n9093));
  AOI21xp33_ASAP7_75t_L     g08837(.A1(new_n9076), .A2(new_n9072), .B(new_n8904), .Y(new_n9094));
  INVx1_ASAP7_75t_L         g08838(.A(new_n9091), .Y(new_n9095));
  OAI21xp33_ASAP7_75t_L     g08839(.A1(new_n9094), .A2(new_n9093), .B(new_n9095), .Y(new_n9096));
  NOR3xp33_ASAP7_75t_L      g08840(.A(new_n8786), .B(new_n8775), .C(new_n8770), .Y(new_n9097));
  O2A1O1Ixp33_ASAP7_75t_L   g08841(.A1(new_n8783), .A2(new_n8787), .B(new_n8793), .C(new_n9097), .Y(new_n9098));
  NAND3xp33_ASAP7_75t_L     g08842(.A(new_n9098), .B(new_n9096), .C(new_n9092), .Y(new_n9099));
  NAND2xp33_ASAP7_75t_L     g08843(.A(new_n9092), .B(new_n9096), .Y(new_n9100));
  INVx1_ASAP7_75t_L         g08844(.A(new_n9097), .Y(new_n9101));
  OAI21xp33_ASAP7_75t_L     g08845(.A1(new_n8790), .A2(new_n8788), .B(new_n9101), .Y(new_n9102));
  NAND2xp33_ASAP7_75t_L     g08846(.A(new_n9100), .B(new_n9102), .Y(new_n9103));
  NAND2xp33_ASAP7_75t_L     g08847(.A(\b[36] ), .B(new_n1194), .Y(new_n9104));
  NAND2xp33_ASAP7_75t_L     g08848(.A(\b[37] ), .B(new_n1103), .Y(new_n9105));
  AOI22xp33_ASAP7_75t_L     g08849(.A1(new_n1113), .A2(\b[38] ), .B1(new_n1110), .B2(new_n4923), .Y(new_n9106));
  AND4x1_ASAP7_75t_L        g08850(.A(new_n9106), .B(new_n9105), .C(new_n9104), .D(\a[17] ), .Y(new_n9107));
  AOI31xp33_ASAP7_75t_L     g08851(.A1(new_n9106), .A2(new_n9105), .A3(new_n9104), .B(\a[17] ), .Y(new_n9108));
  NOR2xp33_ASAP7_75t_L      g08852(.A(new_n9108), .B(new_n9107), .Y(new_n9109));
  NAND3xp33_ASAP7_75t_L     g08853(.A(new_n9103), .B(new_n9099), .C(new_n9109), .Y(new_n9110));
  AND4x1_ASAP7_75t_L        g08854(.A(new_n8794), .B(new_n9101), .C(new_n9092), .D(new_n9096), .Y(new_n9111));
  AOI21xp33_ASAP7_75t_L     g08855(.A1(new_n9096), .A2(new_n9092), .B(new_n9098), .Y(new_n9112));
  INVx1_ASAP7_75t_L         g08856(.A(new_n9109), .Y(new_n9113));
  OAI21xp33_ASAP7_75t_L     g08857(.A1(new_n9112), .A2(new_n9111), .B(new_n9113), .Y(new_n9114));
  NAND2xp33_ASAP7_75t_L     g08858(.A(new_n9114), .B(new_n9110), .Y(new_n9115));
  NAND3xp33_ASAP7_75t_L     g08859(.A(new_n8791), .B(new_n8794), .C(new_n8809), .Y(new_n9116));
  A2O1A1Ixp33_ASAP7_75t_L   g08860(.A1(new_n8810), .A2(new_n8802), .B(new_n8811), .C(new_n9116), .Y(new_n9117));
  NOR2xp33_ASAP7_75t_L      g08861(.A(new_n9117), .B(new_n9115), .Y(new_n9118));
  NOR3xp33_ASAP7_75t_L      g08862(.A(new_n9111), .B(new_n9112), .C(new_n9113), .Y(new_n9119));
  AOI21xp33_ASAP7_75t_L     g08863(.A1(new_n9103), .A2(new_n9099), .B(new_n9109), .Y(new_n9120));
  NOR2xp33_ASAP7_75t_L      g08864(.A(new_n9119), .B(new_n9120), .Y(new_n9121));
  AOI21xp33_ASAP7_75t_L     g08865(.A1(new_n8814), .A2(new_n9116), .B(new_n9121), .Y(new_n9122));
  NAND2xp33_ASAP7_75t_L     g08866(.A(\b[39] ), .B(new_n908), .Y(new_n9123));
  NAND2xp33_ASAP7_75t_L     g08867(.A(\b[40] ), .B(new_n817), .Y(new_n9124));
  AOI22xp33_ASAP7_75t_L     g08868(.A1(new_n826), .A2(\b[41] ), .B1(new_n823), .B2(new_n5669), .Y(new_n9125));
  AND4x1_ASAP7_75t_L        g08869(.A(new_n9125), .B(new_n9124), .C(new_n9123), .D(\a[14] ), .Y(new_n9126));
  AOI31xp33_ASAP7_75t_L     g08870(.A1(new_n9125), .A2(new_n9124), .A3(new_n9123), .B(\a[14] ), .Y(new_n9127));
  NOR2xp33_ASAP7_75t_L      g08871(.A(new_n9127), .B(new_n9126), .Y(new_n9128));
  INVx1_ASAP7_75t_L         g08872(.A(new_n9128), .Y(new_n9129));
  NOR3xp33_ASAP7_75t_L      g08873(.A(new_n9122), .B(new_n9129), .C(new_n9118), .Y(new_n9130));
  NAND4xp25_ASAP7_75t_L     g08874(.A(new_n8814), .B(new_n9116), .C(new_n9114), .D(new_n9110), .Y(new_n9131));
  NAND2xp33_ASAP7_75t_L     g08875(.A(new_n9117), .B(new_n9115), .Y(new_n9132));
  AOI21xp33_ASAP7_75t_L     g08876(.A1(new_n9131), .A2(new_n9132), .B(new_n9128), .Y(new_n9133));
  NOR2xp33_ASAP7_75t_L      g08877(.A(new_n9133), .B(new_n9130), .Y(new_n9134));
  NOR2xp33_ASAP7_75t_L      g08878(.A(new_n8825), .B(new_n8824), .Y(new_n9135));
  MAJIxp5_ASAP7_75t_L       g08879(.A(new_n8830), .B(new_n9135), .C(new_n8821), .Y(new_n9136));
  NAND2xp33_ASAP7_75t_L     g08880(.A(new_n9136), .B(new_n9134), .Y(new_n9137));
  NAND3xp33_ASAP7_75t_L     g08881(.A(new_n9131), .B(new_n9132), .C(new_n9128), .Y(new_n9138));
  OAI21xp33_ASAP7_75t_L     g08882(.A1(new_n9118), .A2(new_n9122), .B(new_n9129), .Y(new_n9139));
  NAND2xp33_ASAP7_75t_L     g08883(.A(new_n9138), .B(new_n9139), .Y(new_n9140));
  NAND2xp33_ASAP7_75t_L     g08884(.A(new_n8821), .B(new_n9135), .Y(new_n9141));
  INVx1_ASAP7_75t_L         g08885(.A(new_n9141), .Y(new_n9142));
  A2O1A1Ixp33_ASAP7_75t_L   g08886(.A1(new_n8827), .A2(new_n8830), .B(new_n9142), .C(new_n9140), .Y(new_n9143));
  NOR2xp33_ASAP7_75t_L      g08887(.A(new_n5680), .B(new_n1620), .Y(new_n9144));
  INVx1_ASAP7_75t_L         g08888(.A(new_n9144), .Y(new_n9145));
  NAND2xp33_ASAP7_75t_L     g08889(.A(\b[43] ), .B(new_n590), .Y(new_n9146));
  AOI22xp33_ASAP7_75t_L     g08890(.A1(new_n600), .A2(\b[44] ), .B1(new_n597), .B2(new_n7055), .Y(new_n9147));
  AND4x1_ASAP7_75t_L        g08891(.A(new_n9147), .B(new_n9146), .C(new_n9145), .D(\a[11] ), .Y(new_n9148));
  AOI31xp33_ASAP7_75t_L     g08892(.A1(new_n9147), .A2(new_n9146), .A3(new_n9145), .B(\a[11] ), .Y(new_n9149));
  NOR2xp33_ASAP7_75t_L      g08893(.A(new_n9149), .B(new_n9148), .Y(new_n9150));
  INVx1_ASAP7_75t_L         g08894(.A(new_n9150), .Y(new_n9151));
  NAND3xp33_ASAP7_75t_L     g08895(.A(new_n9143), .B(new_n9137), .C(new_n9151), .Y(new_n9152));
  OAI21xp33_ASAP7_75t_L     g08896(.A1(new_n8834), .A2(new_n8836), .B(new_n9141), .Y(new_n9153));
  NOR2xp33_ASAP7_75t_L      g08897(.A(new_n9140), .B(new_n9153), .Y(new_n9154));
  O2A1O1Ixp33_ASAP7_75t_L   g08898(.A1(new_n8836), .A2(new_n8834), .B(new_n9141), .C(new_n9134), .Y(new_n9155));
  OAI21xp33_ASAP7_75t_L     g08899(.A1(new_n9154), .A2(new_n9155), .B(new_n9150), .Y(new_n9156));
  NAND2xp33_ASAP7_75t_L     g08900(.A(new_n8846), .B(new_n8848), .Y(new_n9157));
  MAJIxp5_ASAP7_75t_L       g08901(.A(new_n8592), .B(new_n8844), .C(new_n9157), .Y(new_n9158));
  NAND3xp33_ASAP7_75t_L     g08902(.A(new_n9158), .B(new_n9156), .C(new_n9152), .Y(new_n9159));
  NOR3xp33_ASAP7_75t_L      g08903(.A(new_n9155), .B(new_n9154), .C(new_n9150), .Y(new_n9160));
  AOI21xp33_ASAP7_75t_L     g08904(.A1(new_n9143), .A2(new_n9137), .B(new_n9151), .Y(new_n9161));
  NOR3xp33_ASAP7_75t_L      g08905(.A(new_n8837), .B(new_n8844), .C(new_n8831), .Y(new_n9162));
  A2O1A1O1Ixp25_ASAP7_75t_L g08906(.A1(new_n8515), .A2(new_n8530), .B(new_n8528), .C(new_n8845), .D(new_n9162), .Y(new_n9163));
  OAI21xp33_ASAP7_75t_L     g08907(.A1(new_n9161), .A2(new_n9160), .B(new_n9163), .Y(new_n9164));
  NAND3xp33_ASAP7_75t_L     g08908(.A(new_n9159), .B(new_n8902), .C(new_n9164), .Y(new_n9165));
  NOR3xp33_ASAP7_75t_L      g08909(.A(new_n9163), .B(new_n9161), .C(new_n9160), .Y(new_n9166));
  AOI21xp33_ASAP7_75t_L     g08910(.A1(new_n9156), .A2(new_n9152), .B(new_n9158), .Y(new_n9167));
  OAI22xp33_ASAP7_75t_L     g08911(.A1(new_n9166), .A2(new_n9167), .B1(new_n8900), .B2(new_n8901), .Y(new_n9168));
  INVx1_ASAP7_75t_L         g08912(.A(new_n8584), .Y(new_n9169));
  A2O1A1O1Ixp25_ASAP7_75t_L g08913(.A1(new_n8543), .A2(new_n8553), .B(new_n9169), .C(new_n8860), .D(new_n8852), .Y(new_n9170));
  NAND3xp33_ASAP7_75t_L     g08914(.A(new_n9170), .B(new_n9168), .C(new_n9165), .Y(new_n9171));
  NAND2xp33_ASAP7_75t_L     g08915(.A(new_n9165), .B(new_n9168), .Y(new_n9172));
  A2O1A1Ixp33_ASAP7_75t_L   g08916(.A1(new_n8860), .A2(new_n8858), .B(new_n8852), .C(new_n9172), .Y(new_n9173));
  NOR2xp33_ASAP7_75t_L      g08917(.A(new_n7907), .B(new_n406), .Y(new_n9174));
  OAI22xp33_ASAP7_75t_L     g08918(.A1(new_n8234), .A2(new_n367), .B1(new_n8228), .B2(new_n368), .Y(new_n9175));
  NOR2xp33_ASAP7_75t_L      g08919(.A(new_n9174), .B(new_n9175), .Y(new_n9176));
  OAI21xp33_ASAP7_75t_L     g08920(.A1(new_n7333), .A2(new_n365), .B(new_n9176), .Y(new_n9177));
  NOR2xp33_ASAP7_75t_L      g08921(.A(new_n339), .B(new_n9177), .Y(new_n9178));
  O2A1O1Ixp33_ASAP7_75t_L   g08922(.A1(new_n7333), .A2(new_n365), .B(new_n9176), .C(\a[5] ), .Y(new_n9179));
  OAI211xp5_ASAP7_75t_L     g08923(.A1(new_n9178), .A2(new_n9179), .B(new_n9173), .C(new_n9171), .Y(new_n9180));
  A2O1A1Ixp33_ASAP7_75t_L   g08924(.A1(new_n8544), .A2(new_n8584), .B(new_n8855), .C(new_n8859), .Y(new_n9181));
  NOR2xp33_ASAP7_75t_L      g08925(.A(new_n9172), .B(new_n9181), .Y(new_n9182));
  AOI21xp33_ASAP7_75t_L     g08926(.A1(new_n9168), .A2(new_n9165), .B(new_n9170), .Y(new_n9183));
  NOR2xp33_ASAP7_75t_L      g08927(.A(new_n9179), .B(new_n9178), .Y(new_n9184));
  OAI21xp33_ASAP7_75t_L     g08928(.A1(new_n9183), .A2(new_n9182), .B(new_n9184), .Y(new_n9185));
  NAND2xp33_ASAP7_75t_L     g08929(.A(new_n9185), .B(new_n9180), .Y(new_n9186));
  NAND2xp33_ASAP7_75t_L     g08930(.A(new_n9186), .B(new_n8895), .Y(new_n9187));
  A2O1A1Ixp33_ASAP7_75t_L   g08931(.A1(new_n8868), .A2(new_n8869), .B(new_n8583), .C(new_n8893), .Y(new_n9188));
  NAND3xp33_ASAP7_75t_L     g08932(.A(new_n9188), .B(new_n9180), .C(new_n9185), .Y(new_n9189));
  NAND2xp33_ASAP7_75t_L     g08933(.A(new_n9189), .B(new_n9187), .Y(new_n9190));
  XNOR2x2_ASAP7_75t_L       g08934(.A(new_n8892), .B(new_n9190), .Y(new_n9191));
  O2A1O1Ixp33_ASAP7_75t_L   g08935(.A1(new_n8879), .A2(new_n8567), .B(new_n8877), .C(new_n9191), .Y(new_n9192));
  A2O1A1O1Ixp25_ASAP7_75t_L g08936(.A1(new_n8563), .A2(new_n8246), .B(new_n8561), .C(new_n8878), .D(new_n8876), .Y(new_n9193));
  AND2x2_ASAP7_75t_L        g08937(.A(new_n9193), .B(new_n9191), .Y(new_n9194));
  NOR2xp33_ASAP7_75t_L      g08938(.A(new_n9192), .B(new_n9194), .Y(\f[53] ));
  MAJIxp5_ASAP7_75t_L       g08939(.A(new_n9193), .B(new_n8892), .C(new_n9190), .Y(new_n9196));
  INVx1_ASAP7_75t_L         g08940(.A(new_n8883), .Y(new_n9197));
  NOR2xp33_ASAP7_75t_L      g08941(.A(\b[53] ), .B(\b[54] ), .Y(new_n9198));
  INVx1_ASAP7_75t_L         g08942(.A(\b[54] ), .Y(new_n9199));
  NOR2xp33_ASAP7_75t_L      g08943(.A(new_n8882), .B(new_n9199), .Y(new_n9200));
  NOR2xp33_ASAP7_75t_L      g08944(.A(new_n9198), .B(new_n9200), .Y(new_n9201));
  INVx1_ASAP7_75t_L         g08945(.A(new_n9201), .Y(new_n9202));
  O2A1O1Ixp33_ASAP7_75t_L   g08946(.A1(new_n8881), .A2(new_n8886), .B(new_n9197), .C(new_n9202), .Y(new_n9203));
  INVx1_ASAP7_75t_L         g08947(.A(new_n9203), .Y(new_n9204));
  A2O1A1O1Ixp25_ASAP7_75t_L g08948(.A1(new_n8571), .A2(new_n8574), .B(new_n8570), .C(new_n8884), .D(new_n8883), .Y(new_n9205));
  NAND2xp33_ASAP7_75t_L     g08949(.A(new_n9202), .B(new_n9205), .Y(new_n9206));
  NAND2xp33_ASAP7_75t_L     g08950(.A(new_n9204), .B(new_n9206), .Y(new_n9207));
  INVx1_ASAP7_75t_L         g08951(.A(new_n9207), .Y(new_n9208));
  NOR2xp33_ASAP7_75t_L      g08952(.A(new_n9199), .B(new_n632), .Y(new_n9209));
  AOI221xp5_ASAP7_75t_L     g08953(.A1(new_n380), .A2(\b[53] ), .B1(new_n269), .B2(new_n9208), .C(new_n9209), .Y(new_n9210));
  OA211x2_ASAP7_75t_L       g08954(.A1(new_n277), .A2(new_n8569), .B(new_n9210), .C(\a[2] ), .Y(new_n9211));
  O2A1O1Ixp33_ASAP7_75t_L   g08955(.A1(new_n8569), .A2(new_n277), .B(new_n9210), .C(\a[2] ), .Y(new_n9212));
  NOR2xp33_ASAP7_75t_L      g08956(.A(new_n9212), .B(new_n9211), .Y(new_n9213));
  NAND2xp33_ASAP7_75t_L     g08957(.A(\b[46] ), .B(new_n480), .Y(new_n9214));
  NAND2xp33_ASAP7_75t_L     g08958(.A(\b[47] ), .B(new_n441), .Y(new_n9215));
  AOI22xp33_ASAP7_75t_L     g08959(.A1(new_n451), .A2(\b[48] ), .B1(new_n448), .B2(new_n7341), .Y(new_n9216));
  AND4x1_ASAP7_75t_L        g08960(.A(new_n9216), .B(new_n9215), .C(new_n9214), .D(\a[8] ), .Y(new_n9217));
  AOI31xp33_ASAP7_75t_L     g08961(.A1(new_n9216), .A2(new_n9215), .A3(new_n9214), .B(\a[8] ), .Y(new_n9218));
  NOR2xp33_ASAP7_75t_L      g08962(.A(new_n9218), .B(new_n9217), .Y(new_n9219));
  NOR2xp33_ASAP7_75t_L      g08963(.A(new_n6195), .B(new_n1620), .Y(new_n9220));
  INVx1_ASAP7_75t_L         g08964(.A(new_n9220), .Y(new_n9221));
  NAND2xp33_ASAP7_75t_L     g08965(.A(\b[44] ), .B(new_n590), .Y(new_n9222));
  AOI22xp33_ASAP7_75t_L     g08966(.A1(new_n600), .A2(\b[45] ), .B1(new_n597), .B2(new_n6764), .Y(new_n9223));
  AND4x1_ASAP7_75t_L        g08967(.A(new_n9223), .B(new_n9222), .C(new_n9221), .D(\a[11] ), .Y(new_n9224));
  AOI31xp33_ASAP7_75t_L     g08968(.A1(new_n9223), .A2(new_n9222), .A3(new_n9221), .B(\a[11] ), .Y(new_n9225));
  NOR2xp33_ASAP7_75t_L      g08969(.A(new_n9225), .B(new_n9224), .Y(new_n9226));
  NAND2xp33_ASAP7_75t_L     g08970(.A(new_n9132), .B(new_n9131), .Y(new_n9227));
  MAJIxp5_ASAP7_75t_L       g08971(.A(new_n9136), .B(new_n9227), .C(new_n9128), .Y(new_n9228));
  NAND3xp33_ASAP7_75t_L     g08972(.A(new_n9077), .B(new_n9084), .C(new_n9095), .Y(new_n9229));
  INVx1_ASAP7_75t_L         g08973(.A(new_n9229), .Y(new_n9230));
  O2A1O1Ixp33_ASAP7_75t_L   g08974(.A1(new_n9097), .A2(new_n8807), .B(new_n9100), .C(new_n9230), .Y(new_n9231));
  NAND2xp33_ASAP7_75t_L     g08975(.A(\b[35] ), .B(new_n1410), .Y(new_n9232));
  AOI22xp33_ASAP7_75t_L     g08976(.A1(new_n1406), .A2(\b[36] ), .B1(new_n1404), .B2(new_n4473), .Y(new_n9233));
  NAND2xp33_ASAP7_75t_L     g08977(.A(new_n9232), .B(new_n9233), .Y(new_n9234));
  AOI21xp33_ASAP7_75t_L     g08978(.A1(new_n1548), .A2(\b[34] ), .B(new_n9234), .Y(new_n9235));
  NAND2xp33_ASAP7_75t_L     g08979(.A(\a[20] ), .B(new_n9235), .Y(new_n9236));
  A2O1A1Ixp33_ASAP7_75t_L   g08980(.A1(\b[34] ), .A2(new_n1548), .B(new_n9234), .C(new_n1401), .Y(new_n9237));
  NAND2xp33_ASAP7_75t_L     g08981(.A(new_n9237), .B(new_n9236), .Y(new_n9238));
  NAND2xp33_ASAP7_75t_L     g08982(.A(new_n9080), .B(new_n9079), .Y(new_n9239));
  A2O1A1Ixp33_ASAP7_75t_L   g08983(.A1(new_n8785), .A2(new_n9239), .B(new_n9082), .C(new_n9076), .Y(new_n9240));
  A2O1A1O1Ixp25_ASAP7_75t_L g08984(.A1(new_n8759), .A2(new_n8761), .B(new_n8753), .C(new_n9069), .D(new_n9066), .Y(new_n9241));
  NAND2xp33_ASAP7_75t_L     g08985(.A(new_n2226), .B(new_n3219), .Y(new_n9242));
  OAI221xp5_ASAP7_75t_L     g08986(.A1(new_n2234), .A2(new_n3212), .B1(new_n2871), .B2(new_n2220), .C(new_n9242), .Y(new_n9243));
  AOI21xp33_ASAP7_75t_L     g08987(.A1(new_n2386), .A2(\b[28] ), .B(new_n9243), .Y(new_n9244));
  NAND2xp33_ASAP7_75t_L     g08988(.A(\a[26] ), .B(new_n9244), .Y(new_n9245));
  A2O1A1Ixp33_ASAP7_75t_L   g08989(.A1(\b[28] ), .A2(new_n2386), .B(new_n9243), .C(new_n2223), .Y(new_n9246));
  AND2x2_ASAP7_75t_L        g08990(.A(new_n9246), .B(new_n9245), .Y(new_n9247));
  NAND2xp33_ASAP7_75t_L     g08991(.A(new_n8739), .B(new_n8746), .Y(new_n9248));
  NOR2xp33_ASAP7_75t_L      g08992(.A(new_n8738), .B(new_n8920), .Y(new_n9249));
  A2O1A1O1Ixp25_ASAP7_75t_L g08993(.A1(new_n8749), .A2(new_n9248), .B(new_n9249), .C(new_n9051), .D(new_n9064), .Y(new_n9250));
  NOR2xp33_ASAP7_75t_L      g08994(.A(new_n2180), .B(new_n2932), .Y(new_n9251));
  INVx1_ASAP7_75t_L         g08995(.A(new_n9251), .Y(new_n9252));
  NOR2xp33_ASAP7_75t_L      g08996(.A(new_n2477), .B(new_n2694), .Y(new_n9253));
  INVx1_ASAP7_75t_L         g08997(.A(new_n9253), .Y(new_n9254));
  AOI22xp33_ASAP7_75t_L     g08998(.A1(new_n2702), .A2(\b[27] ), .B1(new_n2700), .B2(new_n2657), .Y(new_n9255));
  AND4x1_ASAP7_75t_L        g08999(.A(new_n9255), .B(new_n9254), .C(new_n9252), .D(\a[29] ), .Y(new_n9256));
  AOI31xp33_ASAP7_75t_L     g09000(.A1(new_n9255), .A2(new_n9254), .A3(new_n9252), .B(\a[29] ), .Y(new_n9257));
  NOR2xp33_ASAP7_75t_L      g09001(.A(new_n9257), .B(new_n9256), .Y(new_n9258));
  INVx1_ASAP7_75t_L         g09002(.A(new_n8929), .Y(new_n9259));
  AND3x1_ASAP7_75t_L        g09003(.A(new_n9041), .B(new_n9034), .C(new_n9259), .Y(new_n9260));
  INVx1_ASAP7_75t_L         g09004(.A(new_n9260), .Y(new_n9261));
  NAND2xp33_ASAP7_75t_L     g09005(.A(\b[22] ), .B(new_n3491), .Y(new_n9262));
  NAND2xp33_ASAP7_75t_L     g09006(.A(\b[23] ), .B(new_n3260), .Y(new_n9263));
  AOI22xp33_ASAP7_75t_L     g09007(.A1(new_n3256), .A2(\b[24] ), .B1(new_n3254), .B2(new_n2027), .Y(new_n9264));
  NAND4xp25_ASAP7_75t_L     g09008(.A(new_n9264), .B(\a[32] ), .C(new_n9262), .D(new_n9263), .Y(new_n9265));
  NAND2xp33_ASAP7_75t_L     g09009(.A(new_n9263), .B(new_n9264), .Y(new_n9266));
  A2O1A1Ixp33_ASAP7_75t_L   g09010(.A1(\b[22] ), .A2(new_n3491), .B(new_n9266), .C(new_n3251), .Y(new_n9267));
  NAND2xp33_ASAP7_75t_L     g09011(.A(new_n9265), .B(new_n9267), .Y(new_n9268));
  A2O1A1Ixp33_ASAP7_75t_L   g09012(.A1(new_n9039), .A2(new_n8610), .B(new_n8393), .C(new_n8716), .Y(new_n9269));
  A2O1A1Ixp33_ASAP7_75t_L   g09013(.A1(new_n9269), .A2(new_n8717), .B(new_n9036), .C(new_n9031), .Y(new_n9270));
  NAND2xp33_ASAP7_75t_L     g09014(.A(\b[19] ), .B(new_n4111), .Y(new_n9271));
  NAND2xp33_ASAP7_75t_L     g09015(.A(\b[20] ), .B(new_n3874), .Y(new_n9272));
  AOI22xp33_ASAP7_75t_L     g09016(.A1(new_n3884), .A2(\b[21] ), .B1(new_n3881), .B2(new_n1715), .Y(new_n9273));
  NAND4xp25_ASAP7_75t_L     g09017(.A(new_n9273), .B(\a[35] ), .C(new_n9271), .D(new_n9272), .Y(new_n9274));
  NAND2xp33_ASAP7_75t_L     g09018(.A(new_n9272), .B(new_n9273), .Y(new_n9275));
  A2O1A1Ixp33_ASAP7_75t_L   g09019(.A1(\b[19] ), .A2(new_n4111), .B(new_n9275), .C(new_n3878), .Y(new_n9276));
  NAND2xp33_ASAP7_75t_L     g09020(.A(new_n9274), .B(new_n9276), .Y(new_n9277));
  NOR2xp33_ASAP7_75t_L      g09021(.A(new_n9019), .B(new_n9016), .Y(new_n9278));
  NAND2xp33_ASAP7_75t_L     g09022(.A(new_n8937), .B(new_n9278), .Y(new_n9279));
  AOI22xp33_ASAP7_75t_L     g09023(.A1(new_n8935), .A2(new_n8936), .B1(new_n9021), .B2(new_n9022), .Y(new_n9280));
  NOR3xp33_ASAP7_75t_L      g09024(.A(new_n9016), .B(new_n9019), .C(new_n8937), .Y(new_n9281));
  OAI21xp33_ASAP7_75t_L     g09025(.A1(new_n9280), .A2(new_n9281), .B(new_n8931), .Y(new_n9282));
  NOR2xp33_ASAP7_75t_L      g09026(.A(new_n1356), .B(new_n4550), .Y(new_n9283));
  AOI221xp5_ASAP7_75t_L     g09027(.A1(new_n4548), .A2(\b[17] ), .B1(new_n4542), .B2(new_n1363), .C(new_n9283), .Y(new_n9284));
  OAI21xp33_ASAP7_75t_L     g09028(.A1(new_n1051), .A2(new_n4781), .B(new_n9284), .Y(new_n9285));
  NOR2xp33_ASAP7_75t_L      g09029(.A(new_n4539), .B(new_n9285), .Y(new_n9286));
  O2A1O1Ixp33_ASAP7_75t_L   g09030(.A1(new_n1051), .A2(new_n4781), .B(new_n9284), .C(\a[38] ), .Y(new_n9287));
  OR2x4_ASAP7_75t_L         g09031(.A(new_n9287), .B(new_n9286), .Y(new_n9288));
  INVx1_ASAP7_75t_L         g09032(.A(new_n9018), .Y(new_n9289));
  NOR3xp33_ASAP7_75t_L      g09033(.A(new_n9012), .B(new_n9013), .C(new_n9010), .Y(new_n9290));
  INVx1_ASAP7_75t_L         g09034(.A(new_n9290), .Y(new_n9291));
  NOR2xp33_ASAP7_75t_L      g09035(.A(new_n793), .B(new_n5521), .Y(new_n9292));
  NAND2xp33_ASAP7_75t_L     g09036(.A(\b[14] ), .B(new_n5240), .Y(new_n9293));
  OAI221xp5_ASAP7_75t_L     g09037(.A1(new_n5253), .A2(new_n952), .B1(new_n5252), .B2(new_n2573), .C(new_n9293), .Y(new_n9294));
  OR3x1_ASAP7_75t_L         g09038(.A(new_n9294), .B(new_n5244), .C(new_n9292), .Y(new_n9295));
  A2O1A1Ixp33_ASAP7_75t_L   g09039(.A1(\b[13] ), .A2(new_n5526), .B(new_n9294), .C(new_n5244), .Y(new_n9296));
  NAND2xp33_ASAP7_75t_L     g09040(.A(new_n9296), .B(new_n9295), .Y(new_n9297));
  A2O1A1Ixp33_ASAP7_75t_L   g09041(.A1(new_n9003), .A2(new_n8687), .B(new_n9001), .C(new_n8997), .Y(new_n9298));
  NOR2xp33_ASAP7_75t_L      g09042(.A(new_n631), .B(new_n6309), .Y(new_n9299));
  NAND2xp33_ASAP7_75t_L     g09043(.A(\b[11] ), .B(new_n5992), .Y(new_n9300));
  OAI221xp5_ASAP7_75t_L     g09044(.A1(new_n6312), .A2(new_n763), .B1(new_n6311), .B2(new_n775), .C(new_n9300), .Y(new_n9301));
  OR3x1_ASAP7_75t_L         g09045(.A(new_n9301), .B(new_n5996), .C(new_n9299), .Y(new_n9302));
  A2O1A1Ixp33_ASAP7_75t_L   g09046(.A1(\b[10] ), .A2(new_n6308), .B(new_n9301), .C(new_n5996), .Y(new_n9303));
  NAND2xp33_ASAP7_75t_L     g09047(.A(new_n9303), .B(new_n9302), .Y(new_n9304));
  A2O1A1O1Ixp25_ASAP7_75t_L g09048(.A1(new_n8672), .A2(new_n8668), .B(new_n8947), .C(new_n8984), .D(new_n8990), .Y(new_n9305));
  NAND2xp33_ASAP7_75t_L     g09049(.A(\b[8] ), .B(new_n6812), .Y(new_n9306));
  OAI221xp5_ASAP7_75t_L     g09050(.A1(new_n7118), .A2(new_n559), .B1(new_n7117), .B2(new_n978), .C(new_n9306), .Y(new_n9307));
  AOI211xp5_ASAP7_75t_L     g09051(.A1(\b[7] ), .A2(new_n7124), .B(new_n6816), .C(new_n9307), .Y(new_n9308));
  NAND2xp33_ASAP7_75t_L     g09052(.A(\b[7] ), .B(new_n7124), .Y(new_n9309));
  AOI22xp33_ASAP7_75t_L     g09053(.A1(new_n6822), .A2(\b[9] ), .B1(new_n6819), .B2(new_n566), .Y(new_n9310));
  AOI31xp33_ASAP7_75t_L     g09054(.A1(new_n9310), .A2(new_n9306), .A3(new_n9309), .B(\a[47] ), .Y(new_n9311));
  NAND5xp2_ASAP7_75t_L      g09055(.A(new_n8646), .B(new_n8643), .C(new_n8636), .D(new_n8324), .E(\a[53] ), .Y(new_n9312));
  INVx1_ASAP7_75t_L         g09056(.A(\a[54] ), .Y(new_n9313));
  NAND2xp33_ASAP7_75t_L     g09057(.A(\a[53] ), .B(new_n9313), .Y(new_n9314));
  NAND2xp33_ASAP7_75t_L     g09058(.A(\a[54] ), .B(new_n8639), .Y(new_n9315));
  AND2x2_ASAP7_75t_L        g09059(.A(new_n9314), .B(new_n9315), .Y(new_n9316));
  NOR2xp33_ASAP7_75t_L      g09060(.A(new_n258), .B(new_n9316), .Y(new_n9317));
  OAI31xp33_ASAP7_75t_L     g09061(.A1(new_n9312), .A2(new_n8970), .A3(new_n8966), .B(new_n9317), .Y(new_n9318));
  INVx1_ASAP7_75t_L         g09062(.A(new_n9317), .Y(new_n9319));
  NAND5xp2_ASAP7_75t_L      g09063(.A(\a[53] ), .B(new_n8971), .C(new_n9319), .D(new_n8962), .E(new_n8324), .Y(new_n9320));
  NOR2xp33_ASAP7_75t_L      g09064(.A(new_n276), .B(new_n8965), .Y(new_n9321));
  NAND2xp33_ASAP7_75t_L     g09065(.A(new_n8963), .B(new_n8321), .Y(new_n9322));
  NAND2xp33_ASAP7_75t_L     g09066(.A(\b[3] ), .B(new_n8645), .Y(new_n9323));
  OAI221xp5_ASAP7_75t_L     g09067(.A1(new_n278), .A2(new_n9322), .B1(new_n8967), .B2(new_n303), .C(new_n9323), .Y(new_n9324));
  OR3x1_ASAP7_75t_L         g09068(.A(new_n9324), .B(new_n8639), .C(new_n9321), .Y(new_n9325));
  A2O1A1Ixp33_ASAP7_75t_L   g09069(.A1(\b[1] ), .A2(new_n8964), .B(new_n9324), .C(new_n8639), .Y(new_n9326));
  AOI22xp33_ASAP7_75t_L     g09070(.A1(new_n9325), .A2(new_n9326), .B1(new_n9318), .B2(new_n9320), .Y(new_n9327));
  INVx1_ASAP7_75t_L         g09071(.A(new_n9327), .Y(new_n9328));
  NAND4xp25_ASAP7_75t_L     g09072(.A(new_n9320), .B(new_n9318), .C(new_n9325), .D(new_n9326), .Y(new_n9329));
  NAND2xp33_ASAP7_75t_L     g09073(.A(\b[4] ), .B(new_n7993), .Y(new_n9330));
  NAND2xp33_ASAP7_75t_L     g09074(.A(\b[5] ), .B(new_n7649), .Y(new_n9331));
  AOI22xp33_ASAP7_75t_L     g09075(.A1(new_n7659), .A2(\b[6] ), .B1(new_n7656), .B2(new_n389), .Y(new_n9332));
  NAND4xp25_ASAP7_75t_L     g09076(.A(new_n9332), .B(\a[50] ), .C(new_n9330), .D(new_n9331), .Y(new_n9333));
  AOI31xp33_ASAP7_75t_L     g09077(.A1(new_n9332), .A2(new_n9331), .A3(new_n9330), .B(\a[50] ), .Y(new_n9334));
  INVx1_ASAP7_75t_L         g09078(.A(new_n9334), .Y(new_n9335));
  NAND4xp25_ASAP7_75t_L     g09079(.A(new_n9328), .B(new_n9335), .C(new_n9333), .D(new_n9329), .Y(new_n9336));
  AND4x1_ASAP7_75t_L        g09080(.A(new_n9320), .B(new_n9318), .C(new_n9326), .D(new_n9325), .Y(new_n9337));
  INVx1_ASAP7_75t_L         g09081(.A(new_n9333), .Y(new_n9338));
  OAI22xp33_ASAP7_75t_L     g09082(.A1(new_n9338), .A2(new_n9334), .B1(new_n9327), .B2(new_n9337), .Y(new_n9339));
  A2O1A1Ixp33_ASAP7_75t_L   g09083(.A1(new_n8625), .A2(new_n8649), .B(new_n8656), .C(new_n8977), .Y(new_n9340));
  AOI22xp33_ASAP7_75t_L     g09084(.A1(new_n9339), .A2(new_n9336), .B1(new_n8980), .B2(new_n9340), .Y(new_n9341));
  INVx1_ASAP7_75t_L         g09085(.A(new_n8980), .Y(new_n9342));
  NOR4xp25_ASAP7_75t_L      g09086(.A(new_n9338), .B(new_n9337), .C(new_n9334), .D(new_n9327), .Y(new_n9343));
  AOI22xp33_ASAP7_75t_L     g09087(.A1(new_n9333), .A2(new_n9335), .B1(new_n9329), .B2(new_n9328), .Y(new_n9344));
  AOI211xp5_ASAP7_75t_L     g09088(.A1(new_n8979), .A2(new_n8972), .B(new_n8958), .C(new_n8960), .Y(new_n9345));
  O2A1O1Ixp33_ASAP7_75t_L   g09089(.A1(new_n8654), .A2(new_n8655), .B(new_n8652), .C(new_n9345), .Y(new_n9346));
  NOR4xp25_ASAP7_75t_L      g09090(.A(new_n9344), .B(new_n9346), .C(new_n9342), .D(new_n9343), .Y(new_n9347));
  OAI22xp33_ASAP7_75t_L     g09091(.A1(new_n9341), .A2(new_n9347), .B1(new_n9308), .B2(new_n9311), .Y(new_n9348));
  NAND4xp25_ASAP7_75t_L     g09092(.A(new_n9310), .B(\a[47] ), .C(new_n9309), .D(new_n9306), .Y(new_n9349));
  A2O1A1Ixp33_ASAP7_75t_L   g09093(.A1(\b[7] ), .A2(new_n7124), .B(new_n9307), .C(new_n6816), .Y(new_n9350));
  OAI22xp33_ASAP7_75t_L     g09094(.A1(new_n9344), .A2(new_n9343), .B1(new_n9342), .B2(new_n9346), .Y(new_n9351));
  A2O1A1O1Ixp25_ASAP7_75t_L g09095(.A1(new_n8649), .A2(new_n8625), .B(new_n8656), .C(new_n8977), .D(new_n9342), .Y(new_n9352));
  NAND3xp33_ASAP7_75t_L     g09096(.A(new_n9352), .B(new_n9339), .C(new_n9336), .Y(new_n9353));
  NAND4xp25_ASAP7_75t_L     g09097(.A(new_n9353), .B(new_n9351), .C(new_n9349), .D(new_n9350), .Y(new_n9354));
  AOI21xp33_ASAP7_75t_L     g09098(.A1(new_n9354), .A2(new_n9348), .B(new_n9305), .Y(new_n9355));
  NAND2xp33_ASAP7_75t_L     g09099(.A(new_n9348), .B(new_n9354), .Y(new_n9356));
  AOI211xp5_ASAP7_75t_L     g09100(.A1(new_n8991), .A2(new_n8988), .B(new_n8990), .C(new_n9356), .Y(new_n9357));
  OAI21xp33_ASAP7_75t_L     g09101(.A1(new_n9355), .A2(new_n9357), .B(new_n9304), .Y(new_n9358));
  A2O1A1Ixp33_ASAP7_75t_L   g09102(.A1(new_n8991), .A2(new_n8988), .B(new_n8990), .C(new_n9356), .Y(new_n9359));
  NAND3xp33_ASAP7_75t_L     g09103(.A(new_n9305), .B(new_n9348), .C(new_n9354), .Y(new_n9360));
  NAND4xp25_ASAP7_75t_L     g09104(.A(new_n9359), .B(new_n9360), .C(new_n9302), .D(new_n9303), .Y(new_n9361));
  NAND2xp33_ASAP7_75t_L     g09105(.A(new_n9361), .B(new_n9358), .Y(new_n9362));
  NAND2xp33_ASAP7_75t_L     g09106(.A(new_n9298), .B(new_n9362), .Y(new_n9363));
  NOR2xp33_ASAP7_75t_L      g09107(.A(new_n8676), .B(new_n8673), .Y(new_n9364));
  O2A1O1Ixp33_ASAP7_75t_L   g09108(.A1(new_n8355), .A2(new_n8364), .B(new_n8366), .C(new_n8998), .Y(new_n9365));
  A2O1A1O1Ixp25_ASAP7_75t_L g09109(.A1(new_n9364), .A2(new_n8686), .B(new_n9365), .C(new_n8993), .D(new_n9002), .Y(new_n9366));
  NAND3xp33_ASAP7_75t_L     g09110(.A(new_n9366), .B(new_n9358), .C(new_n9361), .Y(new_n9367));
  NAND3xp33_ASAP7_75t_L     g09111(.A(new_n9367), .B(new_n9363), .C(new_n9297), .Y(new_n9368));
  AND2x2_ASAP7_75t_L        g09112(.A(new_n9296), .B(new_n9295), .Y(new_n9369));
  AOI21xp33_ASAP7_75t_L     g09113(.A1(new_n9361), .A2(new_n9358), .B(new_n9366), .Y(new_n9370));
  NOR2xp33_ASAP7_75t_L      g09114(.A(new_n9298), .B(new_n9362), .Y(new_n9371));
  OAI21xp33_ASAP7_75t_L     g09115(.A1(new_n9371), .A2(new_n9370), .B(new_n9369), .Y(new_n9372));
  NAND2xp33_ASAP7_75t_L     g09116(.A(new_n9368), .B(new_n9372), .Y(new_n9373));
  O2A1O1Ixp33_ASAP7_75t_L   g09117(.A1(new_n8939), .A2(new_n9289), .B(new_n9291), .C(new_n9373), .Y(new_n9374));
  AOI221xp5_ASAP7_75t_L     g09118(.A1(new_n9017), .A2(new_n9018), .B1(new_n9368), .B2(new_n9372), .C(new_n9290), .Y(new_n9375));
  OAI21xp33_ASAP7_75t_L     g09119(.A1(new_n9375), .A2(new_n9374), .B(new_n9288), .Y(new_n9376));
  NOR2xp33_ASAP7_75t_L      g09120(.A(new_n9287), .B(new_n9286), .Y(new_n9377));
  NOR3xp33_ASAP7_75t_L      g09121(.A(new_n9370), .B(new_n9371), .C(new_n9369), .Y(new_n9378));
  AOI21xp33_ASAP7_75t_L     g09122(.A1(new_n9367), .A2(new_n9363), .B(new_n9297), .Y(new_n9379));
  NOR2xp33_ASAP7_75t_L      g09123(.A(new_n9379), .B(new_n9378), .Y(new_n9380));
  A2O1A1Ixp33_ASAP7_75t_L   g09124(.A1(new_n9018), .A2(new_n9017), .B(new_n9290), .C(new_n9380), .Y(new_n9381));
  A2O1A1O1Ixp25_ASAP7_75t_L g09125(.A1(new_n8690), .A2(new_n8614), .B(new_n8938), .C(new_n9018), .D(new_n9290), .Y(new_n9382));
  NAND2xp33_ASAP7_75t_L     g09126(.A(new_n9373), .B(new_n9382), .Y(new_n9383));
  NAND3xp33_ASAP7_75t_L     g09127(.A(new_n9381), .B(new_n9383), .C(new_n9377), .Y(new_n9384));
  AO22x1_ASAP7_75t_L        g09128(.A1(new_n9384), .A2(new_n9376), .B1(new_n9279), .B2(new_n9282), .Y(new_n9385));
  AOI211xp5_ASAP7_75t_L     g09129(.A1(new_n8936), .A2(new_n8935), .B(new_n9019), .C(new_n9016), .Y(new_n9386));
  O2A1O1Ixp33_ASAP7_75t_L   g09130(.A1(new_n9280), .A2(new_n9281), .B(new_n8931), .C(new_n9386), .Y(new_n9387));
  NAND3xp33_ASAP7_75t_L     g09131(.A(new_n9387), .B(new_n9376), .C(new_n9384), .Y(new_n9388));
  NAND3xp33_ASAP7_75t_L     g09132(.A(new_n9385), .B(new_n9277), .C(new_n9388), .Y(new_n9389));
  AND2x2_ASAP7_75t_L        g09133(.A(new_n9274), .B(new_n9276), .Y(new_n9390));
  AOI21xp33_ASAP7_75t_L     g09134(.A1(new_n9384), .A2(new_n9376), .B(new_n9387), .Y(new_n9391));
  AND4x1_ASAP7_75t_L        g09135(.A(new_n9282), .B(new_n9279), .C(new_n9384), .D(new_n9376), .Y(new_n9392));
  OAI21xp33_ASAP7_75t_L     g09136(.A1(new_n9391), .A2(new_n9392), .B(new_n9390), .Y(new_n9393));
  NAND3xp33_ASAP7_75t_L     g09137(.A(new_n9270), .B(new_n9389), .C(new_n9393), .Y(new_n9394));
  A2O1A1O1Ixp25_ASAP7_75t_L g09138(.A1(new_n8716), .A2(new_n8720), .B(new_n8722), .C(new_n9032), .D(new_n9035), .Y(new_n9395));
  NOR3xp33_ASAP7_75t_L      g09139(.A(new_n9392), .B(new_n9391), .C(new_n9390), .Y(new_n9396));
  AOI21xp33_ASAP7_75t_L     g09140(.A1(new_n9385), .A2(new_n9388), .B(new_n9277), .Y(new_n9397));
  OAI21xp33_ASAP7_75t_L     g09141(.A1(new_n9396), .A2(new_n9397), .B(new_n9395), .Y(new_n9398));
  NAND3xp33_ASAP7_75t_L     g09142(.A(new_n9394), .B(new_n9268), .C(new_n9398), .Y(new_n9399));
  INVx1_ASAP7_75t_L         g09143(.A(new_n9268), .Y(new_n9400));
  NOR3xp33_ASAP7_75t_L      g09144(.A(new_n9395), .B(new_n9396), .C(new_n9397), .Y(new_n9401));
  AOI221xp5_ASAP7_75t_L     g09145(.A1(new_n9032), .A2(new_n9033), .B1(new_n9393), .B2(new_n9389), .C(new_n9035), .Y(new_n9402));
  OAI21xp33_ASAP7_75t_L     g09146(.A1(new_n9402), .A2(new_n9401), .B(new_n9400), .Y(new_n9403));
  NAND2xp33_ASAP7_75t_L     g09147(.A(new_n9403), .B(new_n9399), .Y(new_n9404));
  O2A1O1Ixp33_ASAP7_75t_L   g09148(.A1(new_n9054), .A2(new_n9044), .B(new_n9261), .C(new_n9404), .Y(new_n9405));
  AOI221xp5_ASAP7_75t_L     g09149(.A1(new_n9403), .A2(new_n9399), .B1(new_n9049), .B2(new_n9046), .C(new_n9260), .Y(new_n9406));
  NOR3xp33_ASAP7_75t_L      g09150(.A(new_n9405), .B(new_n9406), .C(new_n9258), .Y(new_n9407));
  INVx1_ASAP7_75t_L         g09151(.A(new_n9258), .Y(new_n9408));
  AND2x2_ASAP7_75t_L        g09152(.A(new_n9403), .B(new_n9399), .Y(new_n9409));
  A2O1A1Ixp33_ASAP7_75t_L   g09153(.A1(new_n9049), .A2(new_n9046), .B(new_n9260), .C(new_n9409), .Y(new_n9410));
  INVx1_ASAP7_75t_L         g09154(.A(new_n9406), .Y(new_n9411));
  AOI21xp33_ASAP7_75t_L     g09155(.A1(new_n9411), .A2(new_n9410), .B(new_n9408), .Y(new_n9412));
  NOR3xp33_ASAP7_75t_L      g09156(.A(new_n9250), .B(new_n9407), .C(new_n9412), .Y(new_n9413));
  NAND3xp33_ASAP7_75t_L     g09157(.A(new_n9411), .B(new_n9410), .C(new_n9408), .Y(new_n9414));
  OAI21xp33_ASAP7_75t_L     g09158(.A1(new_n9406), .A2(new_n9405), .B(new_n9258), .Y(new_n9415));
  AOI221xp5_ASAP7_75t_L     g09159(.A1(new_n8921), .A2(new_n9051), .B1(new_n9415), .B2(new_n9414), .C(new_n9064), .Y(new_n9416));
  NOR3xp33_ASAP7_75t_L      g09160(.A(new_n9416), .B(new_n9413), .C(new_n9247), .Y(new_n9417));
  OA21x2_ASAP7_75t_L        g09161(.A1(new_n9413), .A2(new_n9416), .B(new_n9247), .Y(new_n9418));
  NOR3xp33_ASAP7_75t_L      g09162(.A(new_n9418), .B(new_n9241), .C(new_n9417), .Y(new_n9419));
  OAI21xp33_ASAP7_75t_L     g09163(.A1(new_n8913), .A2(new_n9060), .B(new_n9070), .Y(new_n9420));
  OR3x1_ASAP7_75t_L         g09164(.A(new_n9416), .B(new_n9413), .C(new_n9247), .Y(new_n9421));
  OAI21xp33_ASAP7_75t_L     g09165(.A1(new_n9413), .A2(new_n9416), .B(new_n9247), .Y(new_n9422));
  AOI21xp33_ASAP7_75t_L     g09166(.A1(new_n9422), .A2(new_n9421), .B(new_n9420), .Y(new_n9423));
  NAND2xp33_ASAP7_75t_L     g09167(.A(\b[32] ), .B(new_n1770), .Y(new_n9424));
  AOI22xp33_ASAP7_75t_L     g09168(.A1(new_n1766), .A2(\b[33] ), .B1(new_n1764), .B2(new_n3813), .Y(new_n9425));
  NAND2xp33_ASAP7_75t_L     g09169(.A(new_n9424), .B(new_n9425), .Y(new_n9426));
  AOI211xp5_ASAP7_75t_L     g09170(.A1(\b[31] ), .A2(new_n1910), .B(new_n1761), .C(new_n9426), .Y(new_n9427));
  INVx1_ASAP7_75t_L         g09171(.A(new_n9426), .Y(new_n9428));
  O2A1O1Ixp33_ASAP7_75t_L   g09172(.A1(new_n3419), .A2(new_n1911), .B(new_n9428), .C(\a[23] ), .Y(new_n9429));
  NOR2xp33_ASAP7_75t_L      g09173(.A(new_n9427), .B(new_n9429), .Y(new_n9430));
  INVx1_ASAP7_75t_L         g09174(.A(new_n9430), .Y(new_n9431));
  NOR3xp33_ASAP7_75t_L      g09175(.A(new_n9431), .B(new_n9423), .C(new_n9419), .Y(new_n9432));
  NAND3xp33_ASAP7_75t_L     g09176(.A(new_n9420), .B(new_n9421), .C(new_n9422), .Y(new_n9433));
  OAI21xp33_ASAP7_75t_L     g09177(.A1(new_n9417), .A2(new_n9418), .B(new_n9241), .Y(new_n9434));
  AOI21xp33_ASAP7_75t_L     g09178(.A1(new_n9433), .A2(new_n9434), .B(new_n9430), .Y(new_n9435));
  OAI21xp33_ASAP7_75t_L     g09179(.A1(new_n9432), .A2(new_n9435), .B(new_n9240), .Y(new_n9436));
  NAND2xp33_ASAP7_75t_L     g09180(.A(new_n8771), .B(new_n8772), .Y(new_n9437));
  NOR2xp33_ASAP7_75t_L      g09181(.A(new_n8765), .B(new_n8903), .Y(new_n9438));
  A2O1A1O1Ixp25_ASAP7_75t_L g09182(.A1(new_n8769), .A2(new_n9437), .B(new_n9438), .C(new_n9072), .D(new_n9083), .Y(new_n9439));
  NAND3xp33_ASAP7_75t_L     g09183(.A(new_n9433), .B(new_n9434), .C(new_n9430), .Y(new_n9440));
  OAI21xp33_ASAP7_75t_L     g09184(.A1(new_n9419), .A2(new_n9423), .B(new_n9431), .Y(new_n9441));
  NAND3xp33_ASAP7_75t_L     g09185(.A(new_n9439), .B(new_n9440), .C(new_n9441), .Y(new_n9442));
  NAND3xp33_ASAP7_75t_L     g09186(.A(new_n9442), .B(new_n9436), .C(new_n9238), .Y(new_n9443));
  AND2x2_ASAP7_75t_L        g09187(.A(new_n9237), .B(new_n9236), .Y(new_n9444));
  AOI21xp33_ASAP7_75t_L     g09188(.A1(new_n9441), .A2(new_n9440), .B(new_n9439), .Y(new_n9445));
  NOR3xp33_ASAP7_75t_L      g09189(.A(new_n9240), .B(new_n9432), .C(new_n9435), .Y(new_n9446));
  OAI21xp33_ASAP7_75t_L     g09190(.A1(new_n9445), .A2(new_n9446), .B(new_n9444), .Y(new_n9447));
  NAND2xp33_ASAP7_75t_L     g09191(.A(new_n9443), .B(new_n9447), .Y(new_n9448));
  NAND2xp33_ASAP7_75t_L     g09192(.A(new_n9448), .B(new_n9231), .Y(new_n9449));
  A2O1A1Ixp33_ASAP7_75t_L   g09193(.A1(new_n9096), .A2(new_n9092), .B(new_n9098), .C(new_n9229), .Y(new_n9450));
  AND2x2_ASAP7_75t_L        g09194(.A(new_n9443), .B(new_n9447), .Y(new_n9451));
  NAND2xp33_ASAP7_75t_L     g09195(.A(new_n9450), .B(new_n9451), .Y(new_n9452));
  NAND2xp33_ASAP7_75t_L     g09196(.A(\b[37] ), .B(new_n1194), .Y(new_n9453));
  NAND2xp33_ASAP7_75t_L     g09197(.A(\b[38] ), .B(new_n1103), .Y(new_n9454));
  AOI22xp33_ASAP7_75t_L     g09198(.A1(new_n1113), .A2(\b[39] ), .B1(new_n1110), .B2(new_n5174), .Y(new_n9455));
  AND4x1_ASAP7_75t_L        g09199(.A(new_n9455), .B(new_n9454), .C(new_n9453), .D(\a[17] ), .Y(new_n9456));
  AOI31xp33_ASAP7_75t_L     g09200(.A1(new_n9455), .A2(new_n9454), .A3(new_n9453), .B(\a[17] ), .Y(new_n9457));
  NOR2xp33_ASAP7_75t_L      g09201(.A(new_n9457), .B(new_n9456), .Y(new_n9458));
  NAND3xp33_ASAP7_75t_L     g09202(.A(new_n9452), .B(new_n9449), .C(new_n9458), .Y(new_n9459));
  NOR2xp33_ASAP7_75t_L      g09203(.A(new_n9450), .B(new_n9451), .Y(new_n9460));
  A2O1A1O1Ixp25_ASAP7_75t_L g09204(.A1(new_n9096), .A2(new_n9092), .B(new_n9098), .C(new_n9229), .D(new_n9448), .Y(new_n9461));
  INVx1_ASAP7_75t_L         g09205(.A(new_n9458), .Y(new_n9462));
  OAI21xp33_ASAP7_75t_L     g09206(.A1(new_n9461), .A2(new_n9460), .B(new_n9462), .Y(new_n9463));
  NOR2xp33_ASAP7_75t_L      g09207(.A(new_n9112), .B(new_n9111), .Y(new_n9464));
  NAND2xp33_ASAP7_75t_L     g09208(.A(new_n9113), .B(new_n9464), .Y(new_n9465));
  AND4x1_ASAP7_75t_L        g09209(.A(new_n9132), .B(new_n9465), .C(new_n9459), .D(new_n9463), .Y(new_n9466));
  MAJIxp5_ASAP7_75t_L       g09210(.A(new_n9117), .B(new_n9464), .C(new_n9113), .Y(new_n9467));
  AOI21xp33_ASAP7_75t_L     g09211(.A1(new_n9463), .A2(new_n9459), .B(new_n9467), .Y(new_n9468));
  NAND2xp33_ASAP7_75t_L     g09212(.A(\b[40] ), .B(new_n908), .Y(new_n9469));
  NAND2xp33_ASAP7_75t_L     g09213(.A(\b[41] ), .B(new_n817), .Y(new_n9470));
  AOI22xp33_ASAP7_75t_L     g09214(.A1(new_n826), .A2(\b[42] ), .B1(new_n823), .B2(new_n5688), .Y(new_n9471));
  AND4x1_ASAP7_75t_L        g09215(.A(new_n9471), .B(new_n9470), .C(new_n9469), .D(\a[14] ), .Y(new_n9472));
  AOI31xp33_ASAP7_75t_L     g09216(.A1(new_n9471), .A2(new_n9470), .A3(new_n9469), .B(\a[14] ), .Y(new_n9473));
  NOR2xp33_ASAP7_75t_L      g09217(.A(new_n9473), .B(new_n9472), .Y(new_n9474));
  OAI21xp33_ASAP7_75t_L     g09218(.A1(new_n9468), .A2(new_n9466), .B(new_n9474), .Y(new_n9475));
  NAND3xp33_ASAP7_75t_L     g09219(.A(new_n9467), .B(new_n9463), .C(new_n9459), .Y(new_n9476));
  NAND2xp33_ASAP7_75t_L     g09220(.A(new_n9459), .B(new_n9463), .Y(new_n9477));
  A2O1A1Ixp33_ASAP7_75t_L   g09221(.A1(new_n8814), .A2(new_n9116), .B(new_n9121), .C(new_n9465), .Y(new_n9478));
  NAND2xp33_ASAP7_75t_L     g09222(.A(new_n9478), .B(new_n9477), .Y(new_n9479));
  INVx1_ASAP7_75t_L         g09223(.A(new_n9474), .Y(new_n9480));
  NAND3xp33_ASAP7_75t_L     g09224(.A(new_n9479), .B(new_n9480), .C(new_n9476), .Y(new_n9481));
  NAND3xp33_ASAP7_75t_L     g09225(.A(new_n9228), .B(new_n9475), .C(new_n9481), .Y(new_n9482));
  NOR2xp33_ASAP7_75t_L      g09226(.A(new_n9128), .B(new_n9227), .Y(new_n9483));
  INVx1_ASAP7_75t_L         g09227(.A(new_n9483), .Y(new_n9484));
  AOI21xp33_ASAP7_75t_L     g09228(.A1(new_n9479), .A2(new_n9476), .B(new_n9480), .Y(new_n9485));
  NOR3xp33_ASAP7_75t_L      g09229(.A(new_n9466), .B(new_n9474), .C(new_n9468), .Y(new_n9486));
  OAI221xp5_ASAP7_75t_L     g09230(.A1(new_n9136), .A2(new_n9134), .B1(new_n9485), .B2(new_n9486), .C(new_n9484), .Y(new_n9487));
  AOI21xp33_ASAP7_75t_L     g09231(.A1(new_n9482), .A2(new_n9487), .B(new_n9226), .Y(new_n9488));
  INVx1_ASAP7_75t_L         g09232(.A(new_n9226), .Y(new_n9489));
  NAND2xp33_ASAP7_75t_L     g09233(.A(new_n9481), .B(new_n9475), .Y(new_n9490));
  AOI21xp33_ASAP7_75t_L     g09234(.A1(new_n9143), .A2(new_n9484), .B(new_n9490), .Y(new_n9491));
  AOI21xp33_ASAP7_75t_L     g09235(.A1(new_n9481), .A2(new_n9475), .B(new_n9228), .Y(new_n9492));
  NOR3xp33_ASAP7_75t_L      g09236(.A(new_n9491), .B(new_n9492), .C(new_n9489), .Y(new_n9493));
  A2O1A1Ixp33_ASAP7_75t_L   g09237(.A1(new_n8530), .A2(new_n8515), .B(new_n8528), .C(new_n8845), .Y(new_n9494));
  A2O1A1Ixp33_ASAP7_75t_L   g09238(.A1(new_n9494), .A2(new_n8849), .B(new_n9161), .C(new_n9152), .Y(new_n9495));
  OAI21xp33_ASAP7_75t_L     g09239(.A1(new_n9488), .A2(new_n9493), .B(new_n9495), .Y(new_n9496));
  OAI21xp33_ASAP7_75t_L     g09240(.A1(new_n9492), .A2(new_n9491), .B(new_n9489), .Y(new_n9497));
  NAND3xp33_ASAP7_75t_L     g09241(.A(new_n9482), .B(new_n9226), .C(new_n9487), .Y(new_n9498));
  A2O1A1O1Ixp25_ASAP7_75t_L g09242(.A1(new_n7864), .A2(new_n7862), .B(new_n8196), .C(new_n8195), .D(new_n8524), .Y(new_n9499));
  OAI21xp33_ASAP7_75t_L     g09243(.A1(new_n8522), .A2(new_n9499), .B(new_n8521), .Y(new_n9500));
  A2O1A1O1Ixp25_ASAP7_75t_L g09244(.A1(new_n8845), .A2(new_n9500), .B(new_n9162), .C(new_n9156), .D(new_n9160), .Y(new_n9501));
  NAND3xp33_ASAP7_75t_L     g09245(.A(new_n9501), .B(new_n9498), .C(new_n9497), .Y(new_n9502));
  NAND3xp33_ASAP7_75t_L     g09246(.A(new_n9502), .B(new_n9496), .C(new_n9219), .Y(new_n9503));
  INVx1_ASAP7_75t_L         g09247(.A(new_n9219), .Y(new_n9504));
  AOI21xp33_ASAP7_75t_L     g09248(.A1(new_n9498), .A2(new_n9497), .B(new_n9501), .Y(new_n9505));
  NOR3xp33_ASAP7_75t_L      g09249(.A(new_n9495), .B(new_n9493), .C(new_n9488), .Y(new_n9506));
  OAI21xp33_ASAP7_75t_L     g09250(.A1(new_n9506), .A2(new_n9505), .B(new_n9504), .Y(new_n9507));
  NAND2xp33_ASAP7_75t_L     g09251(.A(new_n9503), .B(new_n9507), .Y(new_n9508));
  NAND2xp33_ASAP7_75t_L     g09252(.A(new_n9164), .B(new_n9159), .Y(new_n9509));
  MAJIxp5_ASAP7_75t_L       g09253(.A(new_n9170), .B(new_n8902), .C(new_n9509), .Y(new_n9510));
  NOR2xp33_ASAP7_75t_L      g09254(.A(new_n9510), .B(new_n9508), .Y(new_n9511));
  AND2x2_ASAP7_75t_L        g09255(.A(new_n9510), .B(new_n9508), .Y(new_n9512));
  NAND2xp33_ASAP7_75t_L     g09256(.A(\b[49] ), .B(new_n366), .Y(new_n9513));
  NAND2xp33_ASAP7_75t_L     g09257(.A(\b[50] ), .B(new_n334), .Y(new_n9514));
  AOI22xp33_ASAP7_75t_L     g09258(.A1(new_n345), .A2(\b[51] ), .B1(new_n342), .B2(new_n8257), .Y(new_n9515));
  NAND3xp33_ASAP7_75t_L     g09259(.A(new_n9515), .B(new_n9514), .C(new_n9513), .Y(new_n9516));
  XNOR2x2_ASAP7_75t_L       g09260(.A(\a[5] ), .B(new_n9516), .Y(new_n9517));
  OAI21xp33_ASAP7_75t_L     g09261(.A1(new_n9511), .A2(new_n9512), .B(new_n9517), .Y(new_n9518));
  OR3x1_ASAP7_75t_L         g09262(.A(new_n9512), .B(new_n9511), .C(new_n9517), .Y(new_n9519));
  NAND2xp33_ASAP7_75t_L     g09263(.A(new_n9518), .B(new_n9519), .Y(new_n9520));
  O2A1O1Ixp33_ASAP7_75t_L   g09264(.A1(new_n8895), .A2(new_n9186), .B(new_n9180), .C(new_n9520), .Y(new_n9521));
  OA21x2_ASAP7_75t_L        g09265(.A1(new_n9511), .A2(new_n9512), .B(new_n9517), .Y(new_n9522));
  NOR3xp33_ASAP7_75t_L      g09266(.A(new_n9512), .B(new_n9517), .C(new_n9511), .Y(new_n9523));
  NOR3xp33_ASAP7_75t_L      g09267(.A(new_n9182), .B(new_n9183), .C(new_n9184), .Y(new_n9524));
  A2O1A1O1Ixp25_ASAP7_75t_L g09268(.A1(new_n8873), .A2(new_n8874), .B(new_n8894), .C(new_n9185), .D(new_n9524), .Y(new_n9525));
  OA21x2_ASAP7_75t_L        g09269(.A1(new_n9523), .A2(new_n9522), .B(new_n9525), .Y(new_n9526));
  NOR3xp33_ASAP7_75t_L      g09270(.A(new_n9521), .B(new_n9526), .C(new_n9213), .Y(new_n9527));
  INVx1_ASAP7_75t_L         g09271(.A(new_n9527), .Y(new_n9528));
  OAI21xp33_ASAP7_75t_L     g09272(.A1(new_n9526), .A2(new_n9521), .B(new_n9213), .Y(new_n9529));
  NAND2xp33_ASAP7_75t_L     g09273(.A(new_n9529), .B(new_n9528), .Y(new_n9530));
  XNOR2x2_ASAP7_75t_L       g09274(.A(new_n9196), .B(new_n9530), .Y(\f[54] ));
  INVx1_ASAP7_75t_L         g09275(.A(new_n9196), .Y(new_n9532));
  NOR2xp33_ASAP7_75t_L      g09276(.A(\b[54] ), .B(\b[55] ), .Y(new_n9533));
  INVx1_ASAP7_75t_L         g09277(.A(\b[55] ), .Y(new_n9534));
  NOR2xp33_ASAP7_75t_L      g09278(.A(new_n9199), .B(new_n9534), .Y(new_n9535));
  NOR2xp33_ASAP7_75t_L      g09279(.A(new_n9533), .B(new_n9535), .Y(new_n9536));
  A2O1A1Ixp33_ASAP7_75t_L   g09280(.A1(\b[54] ), .A2(\b[53] ), .B(new_n9203), .C(new_n9536), .Y(new_n9537));
  INVx1_ASAP7_75t_L         g09281(.A(new_n9537), .Y(new_n9538));
  INVx1_ASAP7_75t_L         g09282(.A(new_n9200), .Y(new_n9539));
  A2O1A1Ixp33_ASAP7_75t_L   g09283(.A1(new_n8885), .A2(new_n9197), .B(new_n9198), .C(new_n9539), .Y(new_n9540));
  NOR2xp33_ASAP7_75t_L      g09284(.A(new_n9536), .B(new_n9540), .Y(new_n9541));
  NOR2xp33_ASAP7_75t_L      g09285(.A(new_n9538), .B(new_n9541), .Y(new_n9542));
  NOR2xp33_ASAP7_75t_L      g09286(.A(new_n9534), .B(new_n632), .Y(new_n9543));
  AOI221xp5_ASAP7_75t_L     g09287(.A1(new_n380), .A2(\b[54] ), .B1(new_n269), .B2(new_n9542), .C(new_n9543), .Y(new_n9544));
  OA211x2_ASAP7_75t_L       g09288(.A1(new_n277), .A2(new_n8882), .B(new_n9544), .C(\a[2] ), .Y(new_n9545));
  O2A1O1Ixp33_ASAP7_75t_L   g09289(.A1(new_n8882), .A2(new_n277), .B(new_n9544), .C(\a[2] ), .Y(new_n9546));
  NOR2xp33_ASAP7_75t_L      g09290(.A(new_n9546), .B(new_n9545), .Y(new_n9547));
  A2O1A1O1Ixp25_ASAP7_75t_L g09291(.A1(new_n9185), .A2(new_n9188), .B(new_n9524), .C(new_n9518), .D(new_n9523), .Y(new_n9548));
  NOR3xp33_ASAP7_75t_L      g09292(.A(new_n9505), .B(new_n9506), .C(new_n9219), .Y(new_n9549));
  NAND2xp33_ASAP7_75t_L     g09293(.A(new_n448), .B(new_n7914), .Y(new_n9550));
  OAI221xp5_ASAP7_75t_L     g09294(.A1(new_n667), .A2(new_n7907), .B1(new_n7333), .B2(new_n529), .C(new_n9550), .Y(new_n9551));
  AOI21xp33_ASAP7_75t_L     g09295(.A1(new_n480), .A2(\b[47] ), .B(new_n9551), .Y(new_n9552));
  NAND2xp33_ASAP7_75t_L     g09296(.A(\a[8] ), .B(new_n9552), .Y(new_n9553));
  A2O1A1Ixp33_ASAP7_75t_L   g09297(.A1(\b[47] ), .A2(new_n480), .B(new_n9551), .C(new_n445), .Y(new_n9554));
  NAND2xp33_ASAP7_75t_L     g09298(.A(new_n9554), .B(new_n9553), .Y(new_n9555));
  NAND2xp33_ASAP7_75t_L     g09299(.A(new_n9487), .B(new_n9482), .Y(new_n9556));
  MAJIxp5_ASAP7_75t_L       g09300(.A(new_n9501), .B(new_n9226), .C(new_n9556), .Y(new_n9557));
  NAND2xp33_ASAP7_75t_L     g09301(.A(\b[44] ), .B(new_n674), .Y(new_n9558));
  NAND2xp33_ASAP7_75t_L     g09302(.A(\b[45] ), .B(new_n590), .Y(new_n9559));
  AOI22xp33_ASAP7_75t_L     g09303(.A1(new_n600), .A2(\b[46] ), .B1(new_n597), .B2(new_n7041), .Y(new_n9560));
  AND4x1_ASAP7_75t_L        g09304(.A(new_n9560), .B(new_n9559), .C(new_n9558), .D(\a[11] ), .Y(new_n9561));
  AOI31xp33_ASAP7_75t_L     g09305(.A1(new_n9560), .A2(new_n9559), .A3(new_n9558), .B(\a[11] ), .Y(new_n9562));
  NOR2xp33_ASAP7_75t_L      g09306(.A(new_n9562), .B(new_n9561), .Y(new_n9563));
  A2O1A1O1Ixp25_ASAP7_75t_L g09307(.A1(new_n9140), .A2(new_n9153), .B(new_n9483), .C(new_n9475), .D(new_n9486), .Y(new_n9564));
  A2O1A1O1Ixp25_ASAP7_75t_L g09308(.A1(new_n9032), .A2(new_n9033), .B(new_n9035), .C(new_n9393), .D(new_n9396), .Y(new_n9565));
  NAND2xp33_ASAP7_75t_L     g09309(.A(\b[21] ), .B(new_n3874), .Y(new_n9566));
  OAI221xp5_ASAP7_75t_L     g09310(.A1(new_n4115), .A2(new_n1857), .B1(new_n4114), .B2(new_n1863), .C(new_n9566), .Y(new_n9567));
  AOI21xp33_ASAP7_75t_L     g09311(.A1(new_n4111), .A2(\b[20] ), .B(new_n9567), .Y(new_n9568));
  NAND2xp33_ASAP7_75t_L     g09312(.A(\a[35] ), .B(new_n9568), .Y(new_n9569));
  A2O1A1Ixp33_ASAP7_75t_L   g09313(.A1(\b[20] ), .A2(new_n4111), .B(new_n9567), .C(new_n3878), .Y(new_n9570));
  NAND2xp33_ASAP7_75t_L     g09314(.A(new_n9570), .B(new_n9569), .Y(new_n9571));
  INVx1_ASAP7_75t_L         g09315(.A(new_n9571), .Y(new_n9572));
  NOR3xp33_ASAP7_75t_L      g09316(.A(new_n9374), .B(new_n9375), .C(new_n9377), .Y(new_n9573));
  INVx1_ASAP7_75t_L         g09317(.A(new_n9573), .Y(new_n9574));
  NAND3xp33_ASAP7_75t_L     g09318(.A(new_n9304), .B(new_n9359), .C(new_n9360), .Y(new_n9575));
  A2O1A1Ixp33_ASAP7_75t_L   g09319(.A1(new_n9358), .A2(new_n9361), .B(new_n9366), .C(new_n9575), .Y(new_n9576));
  NOR2xp33_ASAP7_75t_L      g09320(.A(new_n695), .B(new_n6309), .Y(new_n9577));
  INVx1_ASAP7_75t_L         g09321(.A(new_n9577), .Y(new_n9578));
  NAND2xp33_ASAP7_75t_L     g09322(.A(\b[12] ), .B(new_n5992), .Y(new_n9579));
  AOI22xp33_ASAP7_75t_L     g09323(.A1(new_n6002), .A2(\b[13] ), .B1(new_n5999), .B2(new_n800), .Y(new_n9580));
  NAND4xp25_ASAP7_75t_L     g09324(.A(new_n9580), .B(\a[44] ), .C(new_n9578), .D(new_n9579), .Y(new_n9581));
  INVx1_ASAP7_75t_L         g09325(.A(new_n9581), .Y(new_n9582));
  AOI31xp33_ASAP7_75t_L     g09326(.A1(new_n9580), .A2(new_n9579), .A3(new_n9578), .B(\a[44] ), .Y(new_n9583));
  NOR2xp33_ASAP7_75t_L      g09327(.A(new_n9583), .B(new_n9582), .Y(new_n9584));
  AOI211xp5_ASAP7_75t_L     g09328(.A1(new_n9350), .A2(new_n9349), .B(new_n9347), .C(new_n9341), .Y(new_n9585));
  A2O1A1O1Ixp25_ASAP7_75t_L g09329(.A1(new_n8984), .A2(new_n8988), .B(new_n8990), .C(new_n9356), .D(new_n9585), .Y(new_n9586));
  NOR2xp33_ASAP7_75t_L      g09330(.A(new_n503), .B(new_n7115), .Y(new_n9587));
  INVx1_ASAP7_75t_L         g09331(.A(new_n9587), .Y(new_n9588));
  NAND2xp33_ASAP7_75t_L     g09332(.A(\b[9] ), .B(new_n6812), .Y(new_n9589));
  AOI22xp33_ASAP7_75t_L     g09333(.A1(new_n6822), .A2(\b[10] ), .B1(new_n6819), .B2(new_n852), .Y(new_n9590));
  AND4x1_ASAP7_75t_L        g09334(.A(new_n9590), .B(new_n9589), .C(new_n9588), .D(\a[47] ), .Y(new_n9591));
  AOI31xp33_ASAP7_75t_L     g09335(.A1(new_n9590), .A2(new_n9589), .A3(new_n9588), .B(\a[47] ), .Y(new_n9592));
  NOR2xp33_ASAP7_75t_L      g09336(.A(new_n9592), .B(new_n9591), .Y(new_n9593));
  OAI211xp5_ASAP7_75t_L     g09337(.A1(new_n9338), .A2(new_n9334), .B(new_n9328), .C(new_n9329), .Y(new_n9594));
  OAI22xp33_ASAP7_75t_L     g09338(.A1(new_n427), .A2(new_n7996), .B1(new_n7997), .B2(new_n421), .Y(new_n9595));
  AOI221xp5_ASAP7_75t_L     g09339(.A1(\b[5] ), .A2(new_n7993), .B1(\b[6] ), .B2(new_n7649), .C(new_n9595), .Y(new_n9596));
  NAND2xp33_ASAP7_75t_L     g09340(.A(\a[50] ), .B(new_n9596), .Y(new_n9597));
  INVx1_ASAP7_75t_L         g09341(.A(new_n9597), .Y(new_n9598));
  NOR2xp33_ASAP7_75t_L      g09342(.A(\a[50] ), .B(new_n9596), .Y(new_n9599));
  AND2x2_ASAP7_75t_L        g09343(.A(new_n9326), .B(new_n9325), .Y(new_n9600));
  NOR3xp33_ASAP7_75t_L      g09344(.A(new_n9312), .B(new_n8966), .C(new_n8970), .Y(new_n9601));
  NAND2xp33_ASAP7_75t_L     g09345(.A(new_n9317), .B(new_n9601), .Y(new_n9602));
  A2O1A1Ixp33_ASAP7_75t_L   g09346(.A1(new_n9320), .A2(new_n9318), .B(new_n9600), .C(new_n9602), .Y(new_n9603));
  NAND2xp33_ASAP7_75t_L     g09347(.A(\b[2] ), .B(new_n8964), .Y(new_n9604));
  NAND2xp33_ASAP7_75t_L     g09348(.A(\b[3] ), .B(new_n8635), .Y(new_n9605));
  AOI22xp33_ASAP7_75t_L     g09349(.A1(new_n8645), .A2(\b[4] ), .B1(new_n8642), .B2(new_n328), .Y(new_n9606));
  NAND4xp25_ASAP7_75t_L     g09350(.A(new_n9606), .B(\a[53] ), .C(new_n9604), .D(new_n9605), .Y(new_n9607));
  NAND2xp33_ASAP7_75t_L     g09351(.A(new_n9605), .B(new_n9606), .Y(new_n9608));
  A2O1A1Ixp33_ASAP7_75t_L   g09352(.A1(\b[2] ), .A2(new_n8964), .B(new_n9608), .C(new_n8639), .Y(new_n9609));
  INVx1_ASAP7_75t_L         g09353(.A(\a[56] ), .Y(new_n9610));
  NOR2xp33_ASAP7_75t_L      g09354(.A(new_n9610), .B(new_n9319), .Y(new_n9611));
  NAND2xp33_ASAP7_75t_L     g09355(.A(new_n9315), .B(new_n9314), .Y(new_n9612));
  XNOR2x2_ASAP7_75t_L       g09356(.A(\a[55] ), .B(\a[54] ), .Y(new_n9613));
  NOR2xp33_ASAP7_75t_L      g09357(.A(new_n9613), .B(new_n9612), .Y(new_n9614));
  NAND2xp33_ASAP7_75t_L     g09358(.A(\b[0] ), .B(new_n9614), .Y(new_n9615));
  INVx1_ASAP7_75t_L         g09359(.A(\a[55] ), .Y(new_n9616));
  NAND2xp33_ASAP7_75t_L     g09360(.A(\a[56] ), .B(new_n9616), .Y(new_n9617));
  NAND2xp33_ASAP7_75t_L     g09361(.A(\a[55] ), .B(new_n9610), .Y(new_n9618));
  AND2x2_ASAP7_75t_L        g09362(.A(new_n9617), .B(new_n9618), .Y(new_n9619));
  NOR2xp33_ASAP7_75t_L      g09363(.A(new_n9316), .B(new_n9619), .Y(new_n9620));
  NAND2xp33_ASAP7_75t_L     g09364(.A(new_n271), .B(new_n9620), .Y(new_n9621));
  NAND2xp33_ASAP7_75t_L     g09365(.A(new_n9618), .B(new_n9617), .Y(new_n9622));
  NOR2xp33_ASAP7_75t_L      g09366(.A(new_n9622), .B(new_n9316), .Y(new_n9623));
  NAND2xp33_ASAP7_75t_L     g09367(.A(\b[1] ), .B(new_n9623), .Y(new_n9624));
  NAND3xp33_ASAP7_75t_L     g09368(.A(new_n9621), .B(new_n9624), .C(new_n9615), .Y(new_n9625));
  XNOR2x2_ASAP7_75t_L       g09369(.A(new_n9611), .B(new_n9625), .Y(new_n9626));
  NAND3xp33_ASAP7_75t_L     g09370(.A(new_n9609), .B(new_n9607), .C(new_n9626), .Y(new_n9627));
  AOI21xp33_ASAP7_75t_L     g09371(.A1(new_n9609), .A2(new_n9607), .B(new_n9626), .Y(new_n9628));
  INVx1_ASAP7_75t_L         g09372(.A(new_n9628), .Y(new_n9629));
  NAND3xp33_ASAP7_75t_L     g09373(.A(new_n9629), .B(new_n9627), .C(new_n9603), .Y(new_n9630));
  AOI21xp33_ASAP7_75t_L     g09374(.A1(new_n9601), .A2(new_n9317), .B(new_n9327), .Y(new_n9631));
  INVx1_ASAP7_75t_L         g09375(.A(new_n9627), .Y(new_n9632));
  OAI21xp33_ASAP7_75t_L     g09376(.A1(new_n9628), .A2(new_n9632), .B(new_n9631), .Y(new_n9633));
  AOI211xp5_ASAP7_75t_L     g09377(.A1(new_n9630), .A2(new_n9633), .B(new_n9599), .C(new_n9598), .Y(new_n9634));
  AO21x2_ASAP7_75t_L        g09378(.A1(\b[6] ), .A2(new_n7649), .B(new_n9595), .Y(new_n9635));
  A2O1A1Ixp33_ASAP7_75t_L   g09379(.A1(\b[5] ), .A2(new_n7993), .B(new_n9635), .C(new_n7653), .Y(new_n9636));
  NOR3xp33_ASAP7_75t_L      g09380(.A(new_n9631), .B(new_n9632), .C(new_n9628), .Y(new_n9637));
  AOI21xp33_ASAP7_75t_L     g09381(.A1(new_n9629), .A2(new_n9627), .B(new_n9603), .Y(new_n9638));
  AOI211xp5_ASAP7_75t_L     g09382(.A1(new_n9636), .A2(new_n9597), .B(new_n9638), .C(new_n9637), .Y(new_n9639));
  AOI211xp5_ASAP7_75t_L     g09383(.A1(new_n9594), .A2(new_n9351), .B(new_n9639), .C(new_n9634), .Y(new_n9640));
  A2O1A1Ixp33_ASAP7_75t_L   g09384(.A1(new_n9339), .A2(new_n9336), .B(new_n9352), .C(new_n9594), .Y(new_n9641));
  OAI211xp5_ASAP7_75t_L     g09385(.A1(new_n9638), .A2(new_n9637), .B(new_n9636), .C(new_n9597), .Y(new_n9642));
  OAI211xp5_ASAP7_75t_L     g09386(.A1(new_n9599), .A2(new_n9598), .B(new_n9630), .C(new_n9633), .Y(new_n9643));
  AOI21xp33_ASAP7_75t_L     g09387(.A1(new_n9643), .A2(new_n9642), .B(new_n9641), .Y(new_n9644));
  OAI21xp33_ASAP7_75t_L     g09388(.A1(new_n9644), .A2(new_n9640), .B(new_n9593), .Y(new_n9645));
  NAND3xp33_ASAP7_75t_L     g09389(.A(new_n9641), .B(new_n9643), .C(new_n9642), .Y(new_n9646));
  OAI211xp5_ASAP7_75t_L     g09390(.A1(new_n9639), .A2(new_n9634), .B(new_n9594), .C(new_n9351), .Y(new_n9647));
  OAI211xp5_ASAP7_75t_L     g09391(.A1(new_n9591), .A2(new_n9592), .B(new_n9647), .C(new_n9646), .Y(new_n9648));
  NAND2xp33_ASAP7_75t_L     g09392(.A(new_n9645), .B(new_n9648), .Y(new_n9649));
  NOR2xp33_ASAP7_75t_L      g09393(.A(new_n9586), .B(new_n9649), .Y(new_n9650));
  INVx1_ASAP7_75t_L         g09394(.A(new_n9585), .Y(new_n9651));
  A2O1A1Ixp33_ASAP7_75t_L   g09395(.A1(new_n9348), .A2(new_n9354), .B(new_n9305), .C(new_n9651), .Y(new_n9652));
  AOI21xp33_ASAP7_75t_L     g09396(.A1(new_n9648), .A2(new_n9645), .B(new_n9652), .Y(new_n9653));
  OAI21xp33_ASAP7_75t_L     g09397(.A1(new_n9653), .A2(new_n9650), .B(new_n9584), .Y(new_n9654));
  INVx1_ASAP7_75t_L         g09398(.A(new_n9583), .Y(new_n9655));
  NAND2xp33_ASAP7_75t_L     g09399(.A(new_n9581), .B(new_n9655), .Y(new_n9656));
  NAND3xp33_ASAP7_75t_L     g09400(.A(new_n9652), .B(new_n9645), .C(new_n9648), .Y(new_n9657));
  NAND2xp33_ASAP7_75t_L     g09401(.A(new_n9586), .B(new_n9649), .Y(new_n9658));
  NAND3xp33_ASAP7_75t_L     g09402(.A(new_n9658), .B(new_n9657), .C(new_n9656), .Y(new_n9659));
  NAND3xp33_ASAP7_75t_L     g09403(.A(new_n9576), .B(new_n9654), .C(new_n9659), .Y(new_n9660));
  INVx1_ASAP7_75t_L         g09404(.A(new_n9575), .Y(new_n9661));
  A2O1A1O1Ixp25_ASAP7_75t_L g09405(.A1(new_n8993), .A2(new_n8999), .B(new_n9002), .C(new_n9362), .D(new_n9661), .Y(new_n9662));
  NAND2xp33_ASAP7_75t_L     g09406(.A(new_n9659), .B(new_n9654), .Y(new_n9663));
  NAND2xp33_ASAP7_75t_L     g09407(.A(new_n9663), .B(new_n9662), .Y(new_n9664));
  NAND2xp33_ASAP7_75t_L     g09408(.A(\b[14] ), .B(new_n5526), .Y(new_n9665));
  NAND2xp33_ASAP7_75t_L     g09409(.A(\b[15] ), .B(new_n5240), .Y(new_n9666));
  AOI22xp33_ASAP7_75t_L     g09410(.A1(new_n5249), .A2(\b[16] ), .B1(new_n5247), .B2(new_n1058), .Y(new_n9667));
  NAND4xp25_ASAP7_75t_L     g09411(.A(new_n9667), .B(\a[41] ), .C(new_n9665), .D(new_n9666), .Y(new_n9668));
  NAND2xp33_ASAP7_75t_L     g09412(.A(new_n9666), .B(new_n9667), .Y(new_n9669));
  A2O1A1Ixp33_ASAP7_75t_L   g09413(.A1(\b[14] ), .A2(new_n5526), .B(new_n9669), .C(new_n5244), .Y(new_n9670));
  AND2x2_ASAP7_75t_L        g09414(.A(new_n9668), .B(new_n9670), .Y(new_n9671));
  NAND3xp33_ASAP7_75t_L     g09415(.A(new_n9664), .B(new_n9660), .C(new_n9671), .Y(new_n9672));
  AO21x2_ASAP7_75t_L        g09416(.A1(new_n9660), .A2(new_n9664), .B(new_n9671), .Y(new_n9673));
  A2O1A1O1Ixp25_ASAP7_75t_L g09417(.A1(new_n9018), .A2(new_n9017), .B(new_n9290), .C(new_n9372), .D(new_n9378), .Y(new_n9674));
  AND3x1_ASAP7_75t_L        g09418(.A(new_n9674), .B(new_n9673), .C(new_n9672), .Y(new_n9675));
  AOI21xp33_ASAP7_75t_L     g09419(.A1(new_n9673), .A2(new_n9672), .B(new_n9674), .Y(new_n9676));
  NAND2xp33_ASAP7_75t_L     g09420(.A(\b[17] ), .B(new_n4780), .Y(new_n9677));
  NAND2xp33_ASAP7_75t_L     g09421(.A(\b[18] ), .B(new_n4548), .Y(new_n9678));
  AOI22xp33_ASAP7_75t_L     g09422(.A1(new_n4544), .A2(\b[19] ), .B1(new_n4542), .B2(new_n1499), .Y(new_n9679));
  NAND4xp25_ASAP7_75t_L     g09423(.A(new_n9679), .B(\a[38] ), .C(new_n9677), .D(new_n9678), .Y(new_n9680));
  NAND2xp33_ASAP7_75t_L     g09424(.A(new_n9678), .B(new_n9679), .Y(new_n9681));
  A2O1A1Ixp33_ASAP7_75t_L   g09425(.A1(\b[17] ), .A2(new_n4780), .B(new_n9681), .C(new_n4539), .Y(new_n9682));
  AND2x2_ASAP7_75t_L        g09426(.A(new_n9680), .B(new_n9682), .Y(new_n9683));
  OAI21xp33_ASAP7_75t_L     g09427(.A1(new_n9676), .A2(new_n9675), .B(new_n9683), .Y(new_n9684));
  NAND3xp33_ASAP7_75t_L     g09428(.A(new_n9674), .B(new_n9673), .C(new_n9672), .Y(new_n9685));
  AO21x2_ASAP7_75t_L        g09429(.A1(new_n9672), .A2(new_n9673), .B(new_n9674), .Y(new_n9686));
  NAND2xp33_ASAP7_75t_L     g09430(.A(new_n9680), .B(new_n9682), .Y(new_n9687));
  NAND3xp33_ASAP7_75t_L     g09431(.A(new_n9686), .B(new_n9685), .C(new_n9687), .Y(new_n9688));
  NAND4xp25_ASAP7_75t_L     g09432(.A(new_n9385), .B(new_n9688), .C(new_n9684), .D(new_n9574), .Y(new_n9689));
  MAJx2_ASAP7_75t_L         g09433(.A(new_n8931), .B(new_n8937), .C(new_n9278), .Y(new_n9690));
  NAND2xp33_ASAP7_75t_L     g09434(.A(new_n9376), .B(new_n9384), .Y(new_n9691));
  NAND2xp33_ASAP7_75t_L     g09435(.A(new_n9688), .B(new_n9684), .Y(new_n9692));
  A2O1A1Ixp33_ASAP7_75t_L   g09436(.A1(new_n9691), .A2(new_n9690), .B(new_n9573), .C(new_n9692), .Y(new_n9693));
  AOI21xp33_ASAP7_75t_L     g09437(.A1(new_n9689), .A2(new_n9693), .B(new_n9572), .Y(new_n9694));
  A2O1A1Ixp33_ASAP7_75t_L   g09438(.A1(new_n9376), .A2(new_n9384), .B(new_n9387), .C(new_n9574), .Y(new_n9695));
  NOR2xp33_ASAP7_75t_L      g09439(.A(new_n9692), .B(new_n9695), .Y(new_n9696));
  AOI22xp33_ASAP7_75t_L     g09440(.A1(new_n9684), .A2(new_n9688), .B1(new_n9574), .B2(new_n9385), .Y(new_n9697));
  NOR3xp33_ASAP7_75t_L      g09441(.A(new_n9697), .B(new_n9696), .C(new_n9571), .Y(new_n9698));
  OAI21xp33_ASAP7_75t_L     g09442(.A1(new_n9694), .A2(new_n9698), .B(new_n9565), .Y(new_n9699));
  OAI21xp33_ASAP7_75t_L     g09443(.A1(new_n9397), .A2(new_n9395), .B(new_n9389), .Y(new_n9700));
  OAI21xp33_ASAP7_75t_L     g09444(.A1(new_n9696), .A2(new_n9697), .B(new_n9571), .Y(new_n9701));
  NAND3xp33_ASAP7_75t_L     g09445(.A(new_n9572), .B(new_n9689), .C(new_n9693), .Y(new_n9702));
  NAND3xp33_ASAP7_75t_L     g09446(.A(new_n9700), .B(new_n9701), .C(new_n9702), .Y(new_n9703));
  NOR2xp33_ASAP7_75t_L      g09447(.A(new_n1995), .B(new_n3492), .Y(new_n9704));
  INVx1_ASAP7_75t_L         g09448(.A(new_n9704), .Y(new_n9705));
  NOR2xp33_ASAP7_75t_L      g09449(.A(new_n2180), .B(new_n3262), .Y(new_n9706));
  AOI221xp5_ASAP7_75t_L     g09450(.A1(new_n3260), .A2(\b[24] ), .B1(new_n3254), .B2(new_n2188), .C(new_n9706), .Y(new_n9707));
  AND3x1_ASAP7_75t_L        g09451(.A(new_n9707), .B(new_n9705), .C(\a[32] ), .Y(new_n9708));
  O2A1O1Ixp33_ASAP7_75t_L   g09452(.A1(new_n1995), .A2(new_n3492), .B(new_n9707), .C(\a[32] ), .Y(new_n9709));
  NOR2xp33_ASAP7_75t_L      g09453(.A(new_n9709), .B(new_n9708), .Y(new_n9710));
  NAND3xp33_ASAP7_75t_L     g09454(.A(new_n9703), .B(new_n9699), .C(new_n9710), .Y(new_n9711));
  AOI21xp33_ASAP7_75t_L     g09455(.A1(new_n9702), .A2(new_n9701), .B(new_n9700), .Y(new_n9712));
  NOR3xp33_ASAP7_75t_L      g09456(.A(new_n9698), .B(new_n9565), .C(new_n9694), .Y(new_n9713));
  NAND3xp33_ASAP7_75t_L     g09457(.A(new_n9707), .B(new_n9705), .C(\a[32] ), .Y(new_n9714));
  AO21x2_ASAP7_75t_L        g09458(.A1(new_n9705), .A2(new_n9707), .B(\a[32] ), .Y(new_n9715));
  NAND2xp33_ASAP7_75t_L     g09459(.A(new_n9714), .B(new_n9715), .Y(new_n9716));
  OAI21xp33_ASAP7_75t_L     g09460(.A1(new_n9712), .A2(new_n9713), .B(new_n9716), .Y(new_n9717));
  INVx1_ASAP7_75t_L         g09461(.A(new_n9399), .Y(new_n9718));
  A2O1A1O1Ixp25_ASAP7_75t_L g09462(.A1(new_n9049), .A2(new_n9046), .B(new_n9260), .C(new_n9403), .D(new_n9718), .Y(new_n9719));
  NAND3xp33_ASAP7_75t_L     g09463(.A(new_n9719), .B(new_n9717), .C(new_n9711), .Y(new_n9720));
  A2O1A1Ixp33_ASAP7_75t_L   g09464(.A1(new_n8732), .A2(new_n8741), .B(new_n9044), .C(new_n9261), .Y(new_n9721));
  NAND2xp33_ASAP7_75t_L     g09465(.A(new_n9711), .B(new_n9717), .Y(new_n9722));
  A2O1A1Ixp33_ASAP7_75t_L   g09466(.A1(new_n9409), .A2(new_n9721), .B(new_n9718), .C(new_n9722), .Y(new_n9723));
  AOI22xp33_ASAP7_75t_L     g09467(.A1(new_n2702), .A2(\b[28] ), .B1(new_n2700), .B2(new_n2858), .Y(new_n9724));
  OAI221xp5_ASAP7_75t_L     g09468(.A1(new_n2694), .A2(new_n2650), .B1(new_n2477), .B2(new_n2932), .C(new_n9724), .Y(new_n9725));
  XNOR2x2_ASAP7_75t_L       g09469(.A(\a[29] ), .B(new_n9725), .Y(new_n9726));
  NAND3xp33_ASAP7_75t_L     g09470(.A(new_n9720), .B(new_n9726), .C(new_n9723), .Y(new_n9727));
  AO21x2_ASAP7_75t_L        g09471(.A1(new_n9723), .A2(new_n9720), .B(new_n9726), .Y(new_n9728));
  A2O1A1O1Ixp25_ASAP7_75t_L g09472(.A1(new_n9051), .A2(new_n8921), .B(new_n9064), .C(new_n9415), .D(new_n9407), .Y(new_n9729));
  AND3x1_ASAP7_75t_L        g09473(.A(new_n9729), .B(new_n9728), .C(new_n9727), .Y(new_n9730));
  AOI21xp33_ASAP7_75t_L     g09474(.A1(new_n9728), .A2(new_n9727), .B(new_n9729), .Y(new_n9731));
  AOI22xp33_ASAP7_75t_L     g09475(.A1(new_n2228), .A2(\b[31] ), .B1(new_n2226), .B2(new_n3426), .Y(new_n9732));
  OAI221xp5_ASAP7_75t_L     g09476(.A1(new_n2220), .A2(new_n3212), .B1(new_n2871), .B2(new_n2387), .C(new_n9732), .Y(new_n9733));
  XNOR2x2_ASAP7_75t_L       g09477(.A(new_n2223), .B(new_n9733), .Y(new_n9734));
  NOR3xp33_ASAP7_75t_L      g09478(.A(new_n9730), .B(new_n9731), .C(new_n9734), .Y(new_n9735));
  NAND3xp33_ASAP7_75t_L     g09479(.A(new_n9729), .B(new_n9728), .C(new_n9727), .Y(new_n9736));
  AO21x2_ASAP7_75t_L        g09480(.A1(new_n9727), .A2(new_n9728), .B(new_n9729), .Y(new_n9737));
  XNOR2x2_ASAP7_75t_L       g09481(.A(\a[26] ), .B(new_n9733), .Y(new_n9738));
  AOI21xp33_ASAP7_75t_L     g09482(.A1(new_n9737), .A2(new_n9736), .B(new_n9738), .Y(new_n9739));
  NOR2xp33_ASAP7_75t_L      g09483(.A(new_n9739), .B(new_n9735), .Y(new_n9740));
  A2O1A1O1Ixp25_ASAP7_75t_L g09484(.A1(new_n9069), .A2(new_n9068), .B(new_n9066), .C(new_n9422), .D(new_n9417), .Y(new_n9741));
  NAND2xp33_ASAP7_75t_L     g09485(.A(new_n9741), .B(new_n9740), .Y(new_n9742));
  NAND3xp33_ASAP7_75t_L     g09486(.A(new_n9737), .B(new_n9736), .C(new_n9738), .Y(new_n9743));
  OAI21xp33_ASAP7_75t_L     g09487(.A1(new_n9731), .A2(new_n9730), .B(new_n9734), .Y(new_n9744));
  NAND2xp33_ASAP7_75t_L     g09488(.A(new_n9743), .B(new_n9744), .Y(new_n9745));
  A2O1A1Ixp33_ASAP7_75t_L   g09489(.A1(new_n9422), .A2(new_n9420), .B(new_n9417), .C(new_n9745), .Y(new_n9746));
  NAND2xp33_ASAP7_75t_L     g09490(.A(\b[33] ), .B(new_n1770), .Y(new_n9747));
  AOI22xp33_ASAP7_75t_L     g09491(.A1(new_n1766), .A2(\b[34] ), .B1(new_n1764), .B2(new_n3833), .Y(new_n9748));
  NAND2xp33_ASAP7_75t_L     g09492(.A(new_n9747), .B(new_n9748), .Y(new_n9749));
  AOI21xp33_ASAP7_75t_L     g09493(.A1(new_n1910), .A2(\b[32] ), .B(new_n9749), .Y(new_n9750));
  NAND2xp33_ASAP7_75t_L     g09494(.A(\a[23] ), .B(new_n9750), .Y(new_n9751));
  A2O1A1Ixp33_ASAP7_75t_L   g09495(.A1(\b[32] ), .A2(new_n1910), .B(new_n9749), .C(new_n1761), .Y(new_n9752));
  AND2x2_ASAP7_75t_L        g09496(.A(new_n9752), .B(new_n9751), .Y(new_n9753));
  NAND3xp33_ASAP7_75t_L     g09497(.A(new_n9746), .B(new_n9742), .C(new_n9753), .Y(new_n9754));
  OAI21xp33_ASAP7_75t_L     g09498(.A1(new_n9241), .A2(new_n9418), .B(new_n9421), .Y(new_n9755));
  NOR2xp33_ASAP7_75t_L      g09499(.A(new_n9755), .B(new_n9745), .Y(new_n9756));
  O2A1O1Ixp33_ASAP7_75t_L   g09500(.A1(new_n9241), .A2(new_n9418), .B(new_n9421), .C(new_n9740), .Y(new_n9757));
  NAND2xp33_ASAP7_75t_L     g09501(.A(new_n9752), .B(new_n9751), .Y(new_n9758));
  OAI21xp33_ASAP7_75t_L     g09502(.A1(new_n9756), .A2(new_n9757), .B(new_n9758), .Y(new_n9759));
  NOR2xp33_ASAP7_75t_L      g09503(.A(new_n9419), .B(new_n9423), .Y(new_n9760));
  NAND2xp33_ASAP7_75t_L     g09504(.A(new_n9431), .B(new_n9760), .Y(new_n9761));
  NAND4xp25_ASAP7_75t_L     g09505(.A(new_n9436), .B(new_n9761), .C(new_n9759), .D(new_n9754), .Y(new_n9762));
  NOR3xp33_ASAP7_75t_L      g09506(.A(new_n9757), .B(new_n9756), .C(new_n9758), .Y(new_n9763));
  AOI21xp33_ASAP7_75t_L     g09507(.A1(new_n9746), .A2(new_n9742), .B(new_n9753), .Y(new_n9764));
  NAND2xp33_ASAP7_75t_L     g09508(.A(new_n9434), .B(new_n9433), .Y(new_n9765));
  MAJIxp5_ASAP7_75t_L       g09509(.A(new_n9439), .B(new_n9765), .C(new_n9430), .Y(new_n9766));
  OAI21xp33_ASAP7_75t_L     g09510(.A1(new_n9763), .A2(new_n9764), .B(new_n9766), .Y(new_n9767));
  NAND2xp33_ASAP7_75t_L     g09511(.A(\b[36] ), .B(new_n1410), .Y(new_n9768));
  AOI22xp33_ASAP7_75t_L     g09512(.A1(new_n1406), .A2(\b[37] ), .B1(new_n1404), .B2(new_n4709), .Y(new_n9769));
  NAND2xp33_ASAP7_75t_L     g09513(.A(new_n9768), .B(new_n9769), .Y(new_n9770));
  AOI211xp5_ASAP7_75t_L     g09514(.A1(\b[35] ), .A2(new_n1548), .B(new_n1401), .C(new_n9770), .Y(new_n9771));
  AND2x2_ASAP7_75t_L        g09515(.A(new_n9768), .B(new_n9769), .Y(new_n9772));
  O2A1O1Ixp33_ASAP7_75t_L   g09516(.A1(new_n4053), .A2(new_n1549), .B(new_n9772), .C(\a[20] ), .Y(new_n9773));
  NOR2xp33_ASAP7_75t_L      g09517(.A(new_n9771), .B(new_n9773), .Y(new_n9774));
  NAND3xp33_ASAP7_75t_L     g09518(.A(new_n9767), .B(new_n9774), .C(new_n9762), .Y(new_n9775));
  AO21x2_ASAP7_75t_L        g09519(.A1(new_n9762), .A2(new_n9767), .B(new_n9774), .Y(new_n9776));
  NOR3xp33_ASAP7_75t_L      g09520(.A(new_n9446), .B(new_n9445), .C(new_n9444), .Y(new_n9777));
  A2O1A1O1Ixp25_ASAP7_75t_L g09521(.A1(new_n9100), .A2(new_n9102), .B(new_n9230), .C(new_n9447), .D(new_n9777), .Y(new_n9778));
  NAND3xp33_ASAP7_75t_L     g09522(.A(new_n9778), .B(new_n9776), .C(new_n9775), .Y(new_n9779));
  AO21x2_ASAP7_75t_L        g09523(.A1(new_n9775), .A2(new_n9776), .B(new_n9778), .Y(new_n9780));
  NAND2xp33_ASAP7_75t_L     g09524(.A(\b[38] ), .B(new_n1194), .Y(new_n9781));
  NAND2xp33_ASAP7_75t_L     g09525(.A(\b[39] ), .B(new_n1103), .Y(new_n9782));
  AOI22xp33_ASAP7_75t_L     g09526(.A1(new_n1113), .A2(\b[40] ), .B1(new_n1110), .B2(new_n5194), .Y(new_n9783));
  NAND4xp25_ASAP7_75t_L     g09527(.A(new_n9783), .B(\a[17] ), .C(new_n9781), .D(new_n9782), .Y(new_n9784));
  NAND2xp33_ASAP7_75t_L     g09528(.A(new_n9782), .B(new_n9783), .Y(new_n9785));
  A2O1A1Ixp33_ASAP7_75t_L   g09529(.A1(\b[38] ), .A2(new_n1194), .B(new_n9785), .C(new_n1107), .Y(new_n9786));
  AND2x2_ASAP7_75t_L        g09530(.A(new_n9784), .B(new_n9786), .Y(new_n9787));
  NAND3xp33_ASAP7_75t_L     g09531(.A(new_n9780), .B(new_n9779), .C(new_n9787), .Y(new_n9788));
  AND3x1_ASAP7_75t_L        g09532(.A(new_n9778), .B(new_n9776), .C(new_n9775), .Y(new_n9789));
  AOI21xp33_ASAP7_75t_L     g09533(.A1(new_n9776), .A2(new_n9775), .B(new_n9778), .Y(new_n9790));
  NAND2xp33_ASAP7_75t_L     g09534(.A(new_n9784), .B(new_n9786), .Y(new_n9791));
  OAI21xp33_ASAP7_75t_L     g09535(.A1(new_n9790), .A2(new_n9789), .B(new_n9791), .Y(new_n9792));
  NAND2xp33_ASAP7_75t_L     g09536(.A(new_n9788), .B(new_n9792), .Y(new_n9793));
  NAND2xp33_ASAP7_75t_L     g09537(.A(new_n9449), .B(new_n9452), .Y(new_n9794));
  MAJIxp5_ASAP7_75t_L       g09538(.A(new_n9467), .B(new_n9794), .C(new_n9458), .Y(new_n9795));
  NOR2xp33_ASAP7_75t_L      g09539(.A(new_n9793), .B(new_n9795), .Y(new_n9796));
  AND2x2_ASAP7_75t_L        g09540(.A(new_n9788), .B(new_n9792), .Y(new_n9797));
  O2A1O1Ixp33_ASAP7_75t_L   g09541(.A1(new_n9794), .A2(new_n9458), .B(new_n9479), .C(new_n9797), .Y(new_n9798));
  INVx1_ASAP7_75t_L         g09542(.A(new_n6202), .Y(new_n9799));
  NAND2xp33_ASAP7_75t_L     g09543(.A(\b[43] ), .B(new_n826), .Y(new_n9800));
  OAI221xp5_ASAP7_75t_L     g09544(.A1(new_n5680), .A2(new_n994), .B1(new_n911), .B2(new_n9799), .C(new_n9800), .Y(new_n9801));
  AOI21xp33_ASAP7_75t_L     g09545(.A1(new_n908), .A2(\b[41] ), .B(new_n9801), .Y(new_n9802));
  NAND2xp33_ASAP7_75t_L     g09546(.A(\a[14] ), .B(new_n9802), .Y(new_n9803));
  A2O1A1Ixp33_ASAP7_75t_L   g09547(.A1(\b[41] ), .A2(new_n908), .B(new_n9801), .C(new_n813), .Y(new_n9804));
  AND2x2_ASAP7_75t_L        g09548(.A(new_n9804), .B(new_n9803), .Y(new_n9805));
  OAI21xp33_ASAP7_75t_L     g09549(.A1(new_n9796), .A2(new_n9798), .B(new_n9805), .Y(new_n9806));
  OR3x1_ASAP7_75t_L         g09550(.A(new_n9798), .B(new_n9796), .C(new_n9805), .Y(new_n9807));
  NAND3xp33_ASAP7_75t_L     g09551(.A(new_n9807), .B(new_n9564), .C(new_n9806), .Y(new_n9808));
  A2O1A1Ixp33_ASAP7_75t_L   g09552(.A1(new_n9143), .A2(new_n9484), .B(new_n9485), .C(new_n9481), .Y(new_n9809));
  OA21x2_ASAP7_75t_L        g09553(.A1(new_n9796), .A2(new_n9798), .B(new_n9805), .Y(new_n9810));
  NOR3xp33_ASAP7_75t_L      g09554(.A(new_n9798), .B(new_n9805), .C(new_n9796), .Y(new_n9811));
  OAI21xp33_ASAP7_75t_L     g09555(.A1(new_n9810), .A2(new_n9811), .B(new_n9809), .Y(new_n9812));
  NAND3xp33_ASAP7_75t_L     g09556(.A(new_n9812), .B(new_n9563), .C(new_n9808), .Y(new_n9813));
  INVx1_ASAP7_75t_L         g09557(.A(new_n9563), .Y(new_n9814));
  AND3x1_ASAP7_75t_L        g09558(.A(new_n9807), .B(new_n9806), .C(new_n9564), .Y(new_n9815));
  AOI21xp33_ASAP7_75t_L     g09559(.A1(new_n9807), .A2(new_n9806), .B(new_n9564), .Y(new_n9816));
  OAI21xp33_ASAP7_75t_L     g09560(.A1(new_n9816), .A2(new_n9815), .B(new_n9814), .Y(new_n9817));
  NAND3xp33_ASAP7_75t_L     g09561(.A(new_n9557), .B(new_n9813), .C(new_n9817), .Y(new_n9818));
  NOR2xp33_ASAP7_75t_L      g09562(.A(new_n9492), .B(new_n9491), .Y(new_n9819));
  MAJIxp5_ASAP7_75t_L       g09563(.A(new_n9495), .B(new_n9489), .C(new_n9819), .Y(new_n9820));
  NOR3xp33_ASAP7_75t_L      g09564(.A(new_n9815), .B(new_n9816), .C(new_n9814), .Y(new_n9821));
  AOI21xp33_ASAP7_75t_L     g09565(.A1(new_n9812), .A2(new_n9808), .B(new_n9563), .Y(new_n9822));
  OAI21xp33_ASAP7_75t_L     g09566(.A1(new_n9821), .A2(new_n9822), .B(new_n9820), .Y(new_n9823));
  AOI21xp33_ASAP7_75t_L     g09567(.A1(new_n9818), .A2(new_n9823), .B(new_n9555), .Y(new_n9824));
  INVx1_ASAP7_75t_L         g09568(.A(new_n9555), .Y(new_n9825));
  NOR3xp33_ASAP7_75t_L      g09569(.A(new_n9820), .B(new_n9821), .C(new_n9822), .Y(new_n9826));
  NAND2xp33_ASAP7_75t_L     g09570(.A(new_n9498), .B(new_n9497), .Y(new_n9827));
  NOR2xp33_ASAP7_75t_L      g09571(.A(new_n9226), .B(new_n9556), .Y(new_n9828));
  AOI221xp5_ASAP7_75t_L     g09572(.A1(new_n9827), .A2(new_n9495), .B1(new_n9817), .B2(new_n9813), .C(new_n9828), .Y(new_n9829));
  NOR3xp33_ASAP7_75t_L      g09573(.A(new_n9826), .B(new_n9829), .C(new_n9825), .Y(new_n9830));
  NOR2xp33_ASAP7_75t_L      g09574(.A(new_n9830), .B(new_n9824), .Y(new_n9831));
  A2O1A1Ixp33_ASAP7_75t_L   g09575(.A1(new_n9510), .A2(new_n9508), .B(new_n9549), .C(new_n9831), .Y(new_n9832));
  NOR2xp33_ASAP7_75t_L      g09576(.A(new_n8902), .B(new_n9509), .Y(new_n9833));
  O2A1O1Ixp33_ASAP7_75t_L   g09577(.A1(new_n9833), .A2(new_n9183), .B(new_n9508), .C(new_n9549), .Y(new_n9834));
  OAI21xp33_ASAP7_75t_L     g09578(.A1(new_n9829), .A2(new_n9826), .B(new_n9825), .Y(new_n9835));
  NAND3xp33_ASAP7_75t_L     g09579(.A(new_n9818), .B(new_n9555), .C(new_n9823), .Y(new_n9836));
  NAND2xp33_ASAP7_75t_L     g09580(.A(new_n9835), .B(new_n9836), .Y(new_n9837));
  NAND2xp33_ASAP7_75t_L     g09581(.A(new_n9837), .B(new_n9834), .Y(new_n9838));
  NAND2xp33_ASAP7_75t_L     g09582(.A(\b[50] ), .B(new_n366), .Y(new_n9839));
  NAND2xp33_ASAP7_75t_L     g09583(.A(\b[51] ), .B(new_n334), .Y(new_n9840));
  AOI22xp33_ASAP7_75t_L     g09584(.A1(new_n345), .A2(\b[52] ), .B1(new_n342), .B2(new_n8577), .Y(new_n9841));
  AND4x1_ASAP7_75t_L        g09585(.A(new_n9841), .B(new_n9840), .C(new_n9839), .D(\a[5] ), .Y(new_n9842));
  AOI31xp33_ASAP7_75t_L     g09586(.A1(new_n9841), .A2(new_n9840), .A3(new_n9839), .B(\a[5] ), .Y(new_n9843));
  NOR2xp33_ASAP7_75t_L      g09587(.A(new_n9843), .B(new_n9842), .Y(new_n9844));
  NAND3xp33_ASAP7_75t_L     g09588(.A(new_n9832), .B(new_n9838), .C(new_n9844), .Y(new_n9845));
  NOR2xp33_ASAP7_75t_L      g09589(.A(new_n9837), .B(new_n9834), .Y(new_n9846));
  AOI221xp5_ASAP7_75t_L     g09590(.A1(new_n9508), .A2(new_n9510), .B1(new_n9835), .B2(new_n9836), .C(new_n9549), .Y(new_n9847));
  INVx1_ASAP7_75t_L         g09591(.A(new_n9844), .Y(new_n9848));
  OAI21xp33_ASAP7_75t_L     g09592(.A1(new_n9847), .A2(new_n9846), .B(new_n9848), .Y(new_n9849));
  AOI21xp33_ASAP7_75t_L     g09593(.A1(new_n9849), .A2(new_n9845), .B(new_n9548), .Y(new_n9850));
  OAI21xp33_ASAP7_75t_L     g09594(.A1(new_n9522), .A2(new_n9525), .B(new_n9519), .Y(new_n9851));
  NOR3xp33_ASAP7_75t_L      g09595(.A(new_n9846), .B(new_n9847), .C(new_n9848), .Y(new_n9852));
  AOI21xp33_ASAP7_75t_L     g09596(.A1(new_n9832), .A2(new_n9838), .B(new_n9844), .Y(new_n9853));
  NOR3xp33_ASAP7_75t_L      g09597(.A(new_n9851), .B(new_n9852), .C(new_n9853), .Y(new_n9854));
  NOR3xp33_ASAP7_75t_L      g09598(.A(new_n9854), .B(new_n9850), .C(new_n9547), .Y(new_n9855));
  INVx1_ASAP7_75t_L         g09599(.A(new_n9855), .Y(new_n9856));
  OAI21xp33_ASAP7_75t_L     g09600(.A1(new_n9850), .A2(new_n9854), .B(new_n9547), .Y(new_n9857));
  NAND2xp33_ASAP7_75t_L     g09601(.A(new_n9857), .B(new_n9856), .Y(new_n9858));
  O2A1O1Ixp33_ASAP7_75t_L   g09602(.A1(new_n9532), .A2(new_n9530), .B(new_n9528), .C(new_n9858), .Y(new_n9859));
  AOI221xp5_ASAP7_75t_L     g09603(.A1(new_n9529), .A2(new_n9196), .B1(new_n9857), .B2(new_n9856), .C(new_n9527), .Y(new_n9860));
  NOR2xp33_ASAP7_75t_L      g09604(.A(new_n9860), .B(new_n9859), .Y(\f[55] ));
  NOR3xp33_ASAP7_75t_L      g09605(.A(new_n9846), .B(new_n9847), .C(new_n9844), .Y(new_n9862));
  INVx1_ASAP7_75t_L         g09606(.A(new_n9862), .Y(new_n9863));
  A2O1A1Ixp33_ASAP7_75t_L   g09607(.A1(new_n9845), .A2(new_n9849), .B(new_n9548), .C(new_n9863), .Y(new_n9864));
  NAND2xp33_ASAP7_75t_L     g09608(.A(\b[51] ), .B(new_n366), .Y(new_n9865));
  NAND2xp33_ASAP7_75t_L     g09609(.A(\b[52] ), .B(new_n334), .Y(new_n9866));
  AOI22xp33_ASAP7_75t_L     g09610(.A1(new_n345), .A2(\b[53] ), .B1(new_n342), .B2(new_n8889), .Y(new_n9867));
  AND4x1_ASAP7_75t_L        g09611(.A(new_n9867), .B(new_n9866), .C(new_n9865), .D(\a[5] ), .Y(new_n9868));
  AOI31xp33_ASAP7_75t_L     g09612(.A1(new_n9867), .A2(new_n9866), .A3(new_n9865), .B(\a[5] ), .Y(new_n9869));
  NOR2xp33_ASAP7_75t_L      g09613(.A(new_n9869), .B(new_n9868), .Y(new_n9870));
  A2O1A1O1Ixp25_ASAP7_75t_L g09614(.A1(new_n9510), .A2(new_n9508), .B(new_n9549), .C(new_n9835), .D(new_n9830), .Y(new_n9871));
  NAND2xp33_ASAP7_75t_L     g09615(.A(\b[49] ), .B(new_n441), .Y(new_n9872));
  AOI22xp33_ASAP7_75t_L     g09616(.A1(new_n451), .A2(\b[50] ), .B1(new_n448), .B2(new_n8235), .Y(new_n9873));
  NAND2xp33_ASAP7_75t_L     g09617(.A(new_n9872), .B(new_n9873), .Y(new_n9874));
  AOI21xp33_ASAP7_75t_L     g09618(.A1(new_n480), .A2(\b[48] ), .B(new_n9874), .Y(new_n9875));
  NAND2xp33_ASAP7_75t_L     g09619(.A(\a[8] ), .B(new_n9875), .Y(new_n9876));
  A2O1A1Ixp33_ASAP7_75t_L   g09620(.A1(\b[48] ), .A2(new_n480), .B(new_n9874), .C(new_n445), .Y(new_n9877));
  AND2x2_ASAP7_75t_L        g09621(.A(new_n9877), .B(new_n9876), .Y(new_n9878));
  NAND2xp33_ASAP7_75t_L     g09622(.A(new_n9489), .B(new_n9819), .Y(new_n9879));
  A2O1A1Ixp33_ASAP7_75t_L   g09623(.A1(new_n9496), .A2(new_n9879), .B(new_n9821), .C(new_n9817), .Y(new_n9880));
  NOR2xp33_ASAP7_75t_L      g09624(.A(new_n6756), .B(new_n1620), .Y(new_n9881));
  INVx1_ASAP7_75t_L         g09625(.A(new_n9881), .Y(new_n9882));
  NOR2xp33_ASAP7_75t_L      g09626(.A(new_n7033), .B(new_n721), .Y(new_n9883));
  INVx1_ASAP7_75t_L         g09627(.A(new_n9883), .Y(new_n9884));
  AOI22xp33_ASAP7_75t_L     g09628(.A1(new_n600), .A2(\b[47] ), .B1(new_n597), .B2(new_n7323), .Y(new_n9885));
  AND4x1_ASAP7_75t_L        g09629(.A(new_n9885), .B(new_n9884), .C(new_n9882), .D(\a[11] ), .Y(new_n9886));
  AOI31xp33_ASAP7_75t_L     g09630(.A1(new_n9885), .A2(new_n9884), .A3(new_n9882), .B(\a[11] ), .Y(new_n9887));
  NOR2xp33_ASAP7_75t_L      g09631(.A(new_n9887), .B(new_n9886), .Y(new_n9888));
  NOR2xp33_ASAP7_75t_L      g09632(.A(new_n9458), .B(new_n9794), .Y(new_n9889));
  A2O1A1Ixp33_ASAP7_75t_L   g09633(.A1(new_n9477), .A2(new_n9478), .B(new_n9889), .C(new_n9793), .Y(new_n9890));
  NOR2xp33_ASAP7_75t_L      g09634(.A(new_n9731), .B(new_n9730), .Y(new_n9891));
  MAJIxp5_ASAP7_75t_L       g09635(.A(new_n9755), .B(new_n9891), .C(new_n9734), .Y(new_n9892));
  NAND2xp33_ASAP7_75t_L     g09636(.A(\b[30] ), .B(new_n2386), .Y(new_n9893));
  NAND2xp33_ASAP7_75t_L     g09637(.A(\b[31] ), .B(new_n2232), .Y(new_n9894));
  AOI22xp33_ASAP7_75t_L     g09638(.A1(new_n2228), .A2(\b[32] ), .B1(new_n2226), .B2(new_n3450), .Y(new_n9895));
  NAND4xp25_ASAP7_75t_L     g09639(.A(new_n9895), .B(\a[26] ), .C(new_n9893), .D(new_n9894), .Y(new_n9896));
  NAND2xp33_ASAP7_75t_L     g09640(.A(new_n9894), .B(new_n9895), .Y(new_n9897));
  A2O1A1Ixp33_ASAP7_75t_L   g09641(.A1(\b[30] ), .A2(new_n2386), .B(new_n9897), .C(new_n2223), .Y(new_n9898));
  NAND2xp33_ASAP7_75t_L     g09642(.A(new_n9896), .B(new_n9898), .Y(new_n9899));
  NAND2xp33_ASAP7_75t_L     g09643(.A(new_n9723), .B(new_n9720), .Y(new_n9900));
  MAJIxp5_ASAP7_75t_L       g09644(.A(new_n9729), .B(new_n9726), .C(new_n9900), .Y(new_n9901));
  OAI22xp33_ASAP7_75t_L     g09645(.A1(new_n2881), .A2(new_n2707), .B1(new_n2871), .B2(new_n2708), .Y(new_n9902));
  AOI221xp5_ASAP7_75t_L     g09646(.A1(\b[27] ), .A2(new_n2931), .B1(\b[28] ), .B2(new_n2706), .C(new_n9902), .Y(new_n9903));
  XNOR2x2_ASAP7_75t_L       g09647(.A(new_n2697), .B(new_n9903), .Y(new_n9904));
  NOR3xp33_ASAP7_75t_L      g09648(.A(new_n9713), .B(new_n9712), .C(new_n9710), .Y(new_n9905));
  A2O1A1O1Ixp25_ASAP7_75t_L g09649(.A1(new_n9721), .A2(new_n9409), .B(new_n9718), .C(new_n9722), .D(new_n9905), .Y(new_n9906));
  A2O1A1O1Ixp25_ASAP7_75t_L g09650(.A1(new_n9270), .A2(new_n9393), .B(new_n9396), .C(new_n9702), .D(new_n9694), .Y(new_n9907));
  NAND2xp33_ASAP7_75t_L     g09651(.A(\b[21] ), .B(new_n4111), .Y(new_n9908));
  NAND2xp33_ASAP7_75t_L     g09652(.A(\b[22] ), .B(new_n3874), .Y(new_n9909));
  AOI22xp33_ASAP7_75t_L     g09653(.A1(new_n3884), .A2(\b[23] ), .B1(new_n3881), .B2(new_n2002), .Y(new_n9910));
  NAND4xp25_ASAP7_75t_L     g09654(.A(new_n9910), .B(\a[35] ), .C(new_n9908), .D(new_n9909), .Y(new_n9911));
  AOI31xp33_ASAP7_75t_L     g09655(.A1(new_n9910), .A2(new_n9909), .A3(new_n9908), .B(\a[35] ), .Y(new_n9912));
  INVx1_ASAP7_75t_L         g09656(.A(new_n9912), .Y(new_n9913));
  AND2x2_ASAP7_75t_L        g09657(.A(new_n9911), .B(new_n9913), .Y(new_n9914));
  NAND2xp33_ASAP7_75t_L     g09658(.A(new_n9660), .B(new_n9664), .Y(new_n9915));
  MAJIxp5_ASAP7_75t_L       g09659(.A(new_n9674), .B(new_n9671), .C(new_n9915), .Y(new_n9916));
  NAND2xp33_ASAP7_75t_L     g09660(.A(\b[16] ), .B(new_n5240), .Y(new_n9917));
  OAI221xp5_ASAP7_75t_L     g09661(.A1(new_n5253), .A2(new_n1244), .B1(new_n5252), .B2(new_n1251), .C(new_n9917), .Y(new_n9918));
  AOI21xp33_ASAP7_75t_L     g09662(.A1(new_n5526), .A2(\b[15] ), .B(new_n9918), .Y(new_n9919));
  NAND2xp33_ASAP7_75t_L     g09663(.A(\a[41] ), .B(new_n9919), .Y(new_n9920));
  A2O1A1Ixp33_ASAP7_75t_L   g09664(.A1(\b[15] ), .A2(new_n5526), .B(new_n9918), .C(new_n5244), .Y(new_n9921));
  AND2x2_ASAP7_75t_L        g09665(.A(new_n9921), .B(new_n9920), .Y(new_n9922));
  NOR3xp33_ASAP7_75t_L      g09666(.A(new_n9650), .B(new_n9584), .C(new_n9653), .Y(new_n9923));
  A2O1A1O1Ixp25_ASAP7_75t_L g09667(.A1(new_n9298), .A2(new_n9362), .B(new_n9661), .C(new_n9654), .D(new_n9923), .Y(new_n9924));
  A2O1A1Ixp33_ASAP7_75t_L   g09668(.A1(new_n9359), .A2(new_n9651), .B(new_n9649), .C(new_n9648), .Y(new_n9925));
  NOR2xp33_ASAP7_75t_L      g09669(.A(new_n559), .B(new_n7115), .Y(new_n9926));
  INVx1_ASAP7_75t_L         g09670(.A(new_n9926), .Y(new_n9927));
  NAND2xp33_ASAP7_75t_L     g09671(.A(\b[10] ), .B(new_n6812), .Y(new_n9928));
  AOI32xp33_ASAP7_75t_L     g09672(.A1(new_n700), .A2(new_n698), .A3(new_n6819), .B1(\b[11] ), .B2(new_n6822), .Y(new_n9929));
  AND4x1_ASAP7_75t_L        g09673(.A(new_n9929), .B(new_n9928), .C(new_n9927), .D(\a[47] ), .Y(new_n9930));
  AOI31xp33_ASAP7_75t_L     g09674(.A1(new_n9929), .A2(new_n9928), .A3(new_n9927), .B(\a[47] ), .Y(new_n9931));
  NOR2xp33_ASAP7_75t_L      g09675(.A(new_n9931), .B(new_n9930), .Y(new_n9932));
  AOI21xp33_ASAP7_75t_L     g09676(.A1(new_n9641), .A2(new_n9642), .B(new_n9639), .Y(new_n9933));
  NAND2xp33_ASAP7_75t_L     g09677(.A(\b[7] ), .B(new_n7649), .Y(new_n9934));
  OAI221xp5_ASAP7_75t_L     g09678(.A1(new_n7997), .A2(new_n503), .B1(new_n7996), .B2(new_n509), .C(new_n9934), .Y(new_n9935));
  AOI21xp33_ASAP7_75t_L     g09679(.A1(new_n7993), .A2(\b[6] ), .B(new_n9935), .Y(new_n9936));
  NAND2xp33_ASAP7_75t_L     g09680(.A(\a[50] ), .B(new_n9936), .Y(new_n9937));
  A2O1A1Ixp33_ASAP7_75t_L   g09681(.A1(\b[6] ), .A2(new_n7993), .B(new_n9935), .C(new_n7653), .Y(new_n9938));
  A2O1A1O1Ixp25_ASAP7_75t_L g09682(.A1(new_n9601), .A2(new_n9317), .B(new_n9327), .C(new_n9627), .D(new_n9628), .Y(new_n9939));
  NAND2xp33_ASAP7_75t_L     g09683(.A(\b[3] ), .B(new_n8964), .Y(new_n9940));
  NAND2xp33_ASAP7_75t_L     g09684(.A(\b[4] ), .B(new_n8635), .Y(new_n9941));
  AOI22xp33_ASAP7_75t_L     g09685(.A1(new_n8645), .A2(\b[5] ), .B1(new_n8642), .B2(new_n360), .Y(new_n9942));
  NAND4xp25_ASAP7_75t_L     g09686(.A(new_n9942), .B(\a[53] ), .C(new_n9940), .D(new_n9941), .Y(new_n9943));
  AOI31xp33_ASAP7_75t_L     g09687(.A1(new_n9942), .A2(new_n9941), .A3(new_n9940), .B(\a[53] ), .Y(new_n9944));
  INVx1_ASAP7_75t_L         g09688(.A(new_n9944), .Y(new_n9945));
  AND3x1_ASAP7_75t_L        g09689(.A(new_n9621), .B(new_n9624), .C(new_n9615), .Y(new_n9946));
  INVx1_ASAP7_75t_L         g09690(.A(new_n9613), .Y(new_n9947));
  NOR3xp33_ASAP7_75t_L      g09691(.A(new_n9619), .B(new_n9947), .C(new_n9612), .Y(new_n9948));
  NAND2xp33_ASAP7_75t_L     g09692(.A(new_n9622), .B(new_n9612), .Y(new_n9949));
  NAND2xp33_ASAP7_75t_L     g09693(.A(new_n9612), .B(new_n9619), .Y(new_n9950));
  NAND2xp33_ASAP7_75t_L     g09694(.A(\b[1] ), .B(new_n9614), .Y(new_n9951));
  OAI221xp5_ASAP7_75t_L     g09695(.A1(new_n9949), .A2(new_n283), .B1(new_n278), .B2(new_n9950), .C(new_n9951), .Y(new_n9952));
  AOI21xp33_ASAP7_75t_L     g09696(.A1(new_n9948), .A2(\b[0] ), .B(new_n9952), .Y(new_n9953));
  A2O1A1Ixp33_ASAP7_75t_L   g09697(.A1(new_n9319), .A2(new_n9946), .B(new_n9610), .C(new_n9953), .Y(new_n9954));
  O2A1O1Ixp33_ASAP7_75t_L   g09698(.A1(new_n258), .A2(new_n9316), .B(new_n9946), .C(new_n9610), .Y(new_n9955));
  A2O1A1Ixp33_ASAP7_75t_L   g09699(.A1(\b[0] ), .A2(new_n9948), .B(new_n9952), .C(new_n9955), .Y(new_n9956));
  NAND2xp33_ASAP7_75t_L     g09700(.A(new_n9954), .B(new_n9956), .Y(new_n9957));
  NAND3xp33_ASAP7_75t_L     g09701(.A(new_n9957), .B(new_n9945), .C(new_n9943), .Y(new_n9958));
  INVx1_ASAP7_75t_L         g09702(.A(new_n9943), .Y(new_n9959));
  OAI211xp5_ASAP7_75t_L     g09703(.A1(new_n9944), .A2(new_n9959), .B(new_n9954), .C(new_n9956), .Y(new_n9960));
  NAND3xp33_ASAP7_75t_L     g09704(.A(new_n9939), .B(new_n9958), .C(new_n9960), .Y(new_n9961));
  A2O1A1Ixp33_ASAP7_75t_L   g09705(.A1(new_n9328), .A2(new_n9602), .B(new_n9632), .C(new_n9629), .Y(new_n9962));
  AOI211xp5_ASAP7_75t_L     g09706(.A1(new_n9954), .A2(new_n9956), .B(new_n9944), .C(new_n9959), .Y(new_n9963));
  AOI21xp33_ASAP7_75t_L     g09707(.A1(new_n9945), .A2(new_n9943), .B(new_n9957), .Y(new_n9964));
  OAI21xp33_ASAP7_75t_L     g09708(.A1(new_n9963), .A2(new_n9964), .B(new_n9962), .Y(new_n9965));
  AND4x1_ASAP7_75t_L        g09709(.A(new_n9965), .B(new_n9961), .C(new_n9938), .D(new_n9937), .Y(new_n9966));
  AOI22xp33_ASAP7_75t_L     g09710(.A1(new_n9937), .A2(new_n9938), .B1(new_n9961), .B2(new_n9965), .Y(new_n9967));
  NOR3xp33_ASAP7_75t_L      g09711(.A(new_n9933), .B(new_n9966), .C(new_n9967), .Y(new_n9968));
  A2O1A1Ixp33_ASAP7_75t_L   g09712(.A1(new_n9594), .A2(new_n9351), .B(new_n9634), .C(new_n9643), .Y(new_n9969));
  NAND4xp25_ASAP7_75t_L     g09713(.A(new_n9965), .B(new_n9961), .C(new_n9937), .D(new_n9938), .Y(new_n9970));
  AO22x1_ASAP7_75t_L        g09714(.A1(new_n9937), .A2(new_n9938), .B1(new_n9961), .B2(new_n9965), .Y(new_n9971));
  AOI21xp33_ASAP7_75t_L     g09715(.A1(new_n9971), .A2(new_n9970), .B(new_n9969), .Y(new_n9972));
  OAI21xp33_ASAP7_75t_L     g09716(.A1(new_n9972), .A2(new_n9968), .B(new_n9932), .Y(new_n9973));
  NAND3xp33_ASAP7_75t_L     g09717(.A(new_n9969), .B(new_n9971), .C(new_n9970), .Y(new_n9974));
  OAI21xp33_ASAP7_75t_L     g09718(.A1(new_n9966), .A2(new_n9967), .B(new_n9933), .Y(new_n9975));
  OAI211xp5_ASAP7_75t_L     g09719(.A1(new_n9931), .A2(new_n9930), .B(new_n9974), .C(new_n9975), .Y(new_n9976));
  AND2x2_ASAP7_75t_L        g09720(.A(new_n9976), .B(new_n9973), .Y(new_n9977));
  NAND2xp33_ASAP7_75t_L     g09721(.A(new_n9925), .B(new_n9977), .Y(new_n9978));
  INVx1_ASAP7_75t_L         g09722(.A(new_n9648), .Y(new_n9979));
  O2A1O1Ixp33_ASAP7_75t_L   g09723(.A1(new_n9585), .A2(new_n9355), .B(new_n9645), .C(new_n9979), .Y(new_n9980));
  NAND2xp33_ASAP7_75t_L     g09724(.A(new_n9976), .B(new_n9973), .Y(new_n9981));
  NAND2xp33_ASAP7_75t_L     g09725(.A(new_n9981), .B(new_n9980), .Y(new_n9982));
  NAND2xp33_ASAP7_75t_L     g09726(.A(\b[13] ), .B(new_n5992), .Y(new_n9983));
  OAI221xp5_ASAP7_75t_L     g09727(.A1(new_n6312), .A2(new_n871), .B1(new_n6311), .B2(new_n878), .C(new_n9983), .Y(new_n9984));
  AOI21xp33_ASAP7_75t_L     g09728(.A1(new_n6308), .A2(\b[12] ), .B(new_n9984), .Y(new_n9985));
  NAND2xp33_ASAP7_75t_L     g09729(.A(\a[44] ), .B(new_n9985), .Y(new_n9986));
  A2O1A1Ixp33_ASAP7_75t_L   g09730(.A1(\b[12] ), .A2(new_n6308), .B(new_n9984), .C(new_n5996), .Y(new_n9987));
  AND2x2_ASAP7_75t_L        g09731(.A(new_n9987), .B(new_n9986), .Y(new_n9988));
  NAND3xp33_ASAP7_75t_L     g09732(.A(new_n9978), .B(new_n9988), .C(new_n9982), .Y(new_n9989));
  O2A1O1Ixp33_ASAP7_75t_L   g09733(.A1(new_n9586), .A2(new_n9649), .B(new_n9648), .C(new_n9981), .Y(new_n9990));
  NOR2xp33_ASAP7_75t_L      g09734(.A(new_n9925), .B(new_n9977), .Y(new_n9991));
  NAND2xp33_ASAP7_75t_L     g09735(.A(new_n9987), .B(new_n9986), .Y(new_n9992));
  OAI21xp33_ASAP7_75t_L     g09736(.A1(new_n9990), .A2(new_n9991), .B(new_n9992), .Y(new_n9993));
  AO21x2_ASAP7_75t_L        g09737(.A1(new_n9989), .A2(new_n9993), .B(new_n9924), .Y(new_n9994));
  NAND3xp33_ASAP7_75t_L     g09738(.A(new_n9924), .B(new_n9993), .C(new_n9989), .Y(new_n9995));
  AOI21xp33_ASAP7_75t_L     g09739(.A1(new_n9994), .A2(new_n9995), .B(new_n9922), .Y(new_n9996));
  NAND2xp33_ASAP7_75t_L     g09740(.A(new_n9921), .B(new_n9920), .Y(new_n9997));
  AOI21xp33_ASAP7_75t_L     g09741(.A1(new_n9993), .A2(new_n9989), .B(new_n9924), .Y(new_n9998));
  AND3x1_ASAP7_75t_L        g09742(.A(new_n9924), .B(new_n9993), .C(new_n9989), .Y(new_n9999));
  NOR3xp33_ASAP7_75t_L      g09743(.A(new_n9999), .B(new_n9998), .C(new_n9997), .Y(new_n10000));
  NOR2xp33_ASAP7_75t_L      g09744(.A(new_n9996), .B(new_n10000), .Y(new_n10001));
  NAND2xp33_ASAP7_75t_L     g09745(.A(new_n9916), .B(new_n10001), .Y(new_n10002));
  AO21x2_ASAP7_75t_L        g09746(.A1(new_n9670), .A2(new_n9668), .B(new_n9915), .Y(new_n10003));
  OAI21xp33_ASAP7_75t_L     g09747(.A1(new_n9998), .A2(new_n9999), .B(new_n9997), .Y(new_n10004));
  NAND3xp33_ASAP7_75t_L     g09748(.A(new_n9922), .B(new_n9994), .C(new_n9995), .Y(new_n10005));
  NAND2xp33_ASAP7_75t_L     g09749(.A(new_n10004), .B(new_n10005), .Y(new_n10006));
  NAND3xp33_ASAP7_75t_L     g09750(.A(new_n9686), .B(new_n10006), .C(new_n10003), .Y(new_n10007));
  NOR2xp33_ASAP7_75t_L      g09751(.A(new_n1594), .B(new_n4550), .Y(new_n10008));
  AOI221xp5_ASAP7_75t_L     g09752(.A1(new_n4548), .A2(\b[19] ), .B1(new_n4542), .B2(new_n1600), .C(new_n10008), .Y(new_n10009));
  OAI211xp5_ASAP7_75t_L     g09753(.A1(new_n1356), .A2(new_n4781), .B(new_n10009), .C(\a[38] ), .Y(new_n10010));
  O2A1O1Ixp33_ASAP7_75t_L   g09754(.A1(new_n1356), .A2(new_n4781), .B(new_n10009), .C(\a[38] ), .Y(new_n10011));
  INVx1_ASAP7_75t_L         g09755(.A(new_n10011), .Y(new_n10012));
  AND2x2_ASAP7_75t_L        g09756(.A(new_n10010), .B(new_n10012), .Y(new_n10013));
  AOI21xp33_ASAP7_75t_L     g09757(.A1(new_n10007), .A2(new_n10002), .B(new_n10013), .Y(new_n10014));
  O2A1O1Ixp33_ASAP7_75t_L   g09758(.A1(new_n9915), .A2(new_n9671), .B(new_n9686), .C(new_n10006), .Y(new_n10015));
  NOR2xp33_ASAP7_75t_L      g09759(.A(new_n9916), .B(new_n10001), .Y(new_n10016));
  NAND2xp33_ASAP7_75t_L     g09760(.A(new_n10010), .B(new_n10012), .Y(new_n10017));
  NOR3xp33_ASAP7_75t_L      g09761(.A(new_n10015), .B(new_n10016), .C(new_n10017), .Y(new_n10018));
  NOR3xp33_ASAP7_75t_L      g09762(.A(new_n9683), .B(new_n9675), .C(new_n9676), .Y(new_n10019));
  A2O1A1O1Ixp25_ASAP7_75t_L g09763(.A1(new_n9691), .A2(new_n9690), .B(new_n9573), .C(new_n9684), .D(new_n10019), .Y(new_n10020));
  NOR3xp33_ASAP7_75t_L      g09764(.A(new_n10020), .B(new_n10018), .C(new_n10014), .Y(new_n10021));
  OAI21xp33_ASAP7_75t_L     g09765(.A1(new_n10016), .A2(new_n10015), .B(new_n10017), .Y(new_n10022));
  NAND3xp33_ASAP7_75t_L     g09766(.A(new_n10013), .B(new_n10007), .C(new_n10002), .Y(new_n10023));
  AOI21xp33_ASAP7_75t_L     g09767(.A1(new_n9686), .A2(new_n9685), .B(new_n9687), .Y(new_n10024));
  A2O1A1O1Ixp25_ASAP7_75t_L g09768(.A1(new_n9376), .A2(new_n9384), .B(new_n9387), .C(new_n9574), .D(new_n10024), .Y(new_n10025));
  AOI211xp5_ASAP7_75t_L     g09769(.A1(new_n10023), .A2(new_n10022), .B(new_n10025), .C(new_n10019), .Y(new_n10026));
  NOR3xp33_ASAP7_75t_L      g09770(.A(new_n9914), .B(new_n10021), .C(new_n10026), .Y(new_n10027));
  NAND2xp33_ASAP7_75t_L     g09771(.A(new_n9911), .B(new_n9913), .Y(new_n10028));
  OAI211xp5_ASAP7_75t_L     g09772(.A1(new_n10019), .A2(new_n10025), .B(new_n10022), .C(new_n10023), .Y(new_n10029));
  INVx1_ASAP7_75t_L         g09773(.A(new_n10026), .Y(new_n10030));
  AOI21xp33_ASAP7_75t_L     g09774(.A1(new_n10030), .A2(new_n10029), .B(new_n10028), .Y(new_n10031));
  OAI21xp33_ASAP7_75t_L     g09775(.A1(new_n10027), .A2(new_n10031), .B(new_n9907), .Y(new_n10032));
  OAI21xp33_ASAP7_75t_L     g09776(.A1(new_n9565), .A2(new_n9698), .B(new_n9701), .Y(new_n10033));
  NAND3xp33_ASAP7_75t_L     g09777(.A(new_n10030), .B(new_n10029), .C(new_n10028), .Y(new_n10034));
  OAI21xp33_ASAP7_75t_L     g09778(.A1(new_n10026), .A2(new_n10021), .B(new_n9914), .Y(new_n10035));
  NAND3xp33_ASAP7_75t_L     g09779(.A(new_n10033), .B(new_n10034), .C(new_n10035), .Y(new_n10036));
  AOI22xp33_ASAP7_75t_L     g09780(.A1(new_n3256), .A2(\b[26] ), .B1(new_n3254), .B2(new_n2888), .Y(new_n10037));
  OAI221xp5_ASAP7_75t_L     g09781(.A1(new_n3248), .A2(new_n2180), .B1(new_n2019), .B2(new_n3492), .C(new_n10037), .Y(new_n10038));
  XNOR2x2_ASAP7_75t_L       g09782(.A(new_n3251), .B(new_n10038), .Y(new_n10039));
  AOI21xp33_ASAP7_75t_L     g09783(.A1(new_n10032), .A2(new_n10036), .B(new_n10039), .Y(new_n10040));
  AOI21xp33_ASAP7_75t_L     g09784(.A1(new_n10034), .A2(new_n10035), .B(new_n10033), .Y(new_n10041));
  NOR3xp33_ASAP7_75t_L      g09785(.A(new_n10031), .B(new_n9907), .C(new_n10027), .Y(new_n10042));
  XNOR2x2_ASAP7_75t_L       g09786(.A(\a[32] ), .B(new_n10038), .Y(new_n10043));
  NOR3xp33_ASAP7_75t_L      g09787(.A(new_n10042), .B(new_n10041), .C(new_n10043), .Y(new_n10044));
  NOR2xp33_ASAP7_75t_L      g09788(.A(new_n10040), .B(new_n10044), .Y(new_n10045));
  NAND2xp33_ASAP7_75t_L     g09789(.A(new_n10045), .B(new_n9906), .Y(new_n10046));
  A2O1A1Ixp33_ASAP7_75t_L   g09790(.A1(new_n9053), .A2(new_n9261), .B(new_n9404), .C(new_n9399), .Y(new_n10047));
  OAI21xp33_ASAP7_75t_L     g09791(.A1(new_n10041), .A2(new_n10042), .B(new_n10043), .Y(new_n10048));
  NAND3xp33_ASAP7_75t_L     g09792(.A(new_n10032), .B(new_n10036), .C(new_n10039), .Y(new_n10049));
  NAND2xp33_ASAP7_75t_L     g09793(.A(new_n10049), .B(new_n10048), .Y(new_n10050));
  A2O1A1Ixp33_ASAP7_75t_L   g09794(.A1(new_n10047), .A2(new_n9722), .B(new_n9905), .C(new_n10050), .Y(new_n10051));
  NAND3xp33_ASAP7_75t_L     g09795(.A(new_n10051), .B(new_n10046), .C(new_n9904), .Y(new_n10052));
  INVx1_ASAP7_75t_L         g09796(.A(new_n9904), .Y(new_n10053));
  INVx1_ASAP7_75t_L         g09797(.A(new_n9905), .Y(new_n10054));
  A2O1A1Ixp33_ASAP7_75t_L   g09798(.A1(new_n9717), .A2(new_n9711), .B(new_n9719), .C(new_n10054), .Y(new_n10055));
  NOR2xp33_ASAP7_75t_L      g09799(.A(new_n10050), .B(new_n10055), .Y(new_n10056));
  NOR2xp33_ASAP7_75t_L      g09800(.A(new_n10045), .B(new_n9906), .Y(new_n10057));
  OAI21xp33_ASAP7_75t_L     g09801(.A1(new_n10057), .A2(new_n10056), .B(new_n10053), .Y(new_n10058));
  NAND3xp33_ASAP7_75t_L     g09802(.A(new_n9901), .B(new_n10052), .C(new_n10058), .Y(new_n10059));
  AND3x1_ASAP7_75t_L        g09803(.A(new_n9720), .B(new_n9726), .C(new_n9723), .Y(new_n10060));
  AOI21xp33_ASAP7_75t_L     g09804(.A1(new_n9720), .A2(new_n9723), .B(new_n9726), .Y(new_n10061));
  NOR2xp33_ASAP7_75t_L      g09805(.A(new_n10061), .B(new_n10060), .Y(new_n10062));
  NOR2xp33_ASAP7_75t_L      g09806(.A(new_n9726), .B(new_n9900), .Y(new_n10063));
  INVx1_ASAP7_75t_L         g09807(.A(new_n10063), .Y(new_n10064));
  NOR3xp33_ASAP7_75t_L      g09808(.A(new_n10056), .B(new_n10057), .C(new_n10053), .Y(new_n10065));
  AOI21xp33_ASAP7_75t_L     g09809(.A1(new_n10051), .A2(new_n10046), .B(new_n9904), .Y(new_n10066));
  OAI221xp5_ASAP7_75t_L     g09810(.A1(new_n10065), .A2(new_n10066), .B1(new_n9729), .B2(new_n10062), .C(new_n10064), .Y(new_n10067));
  AOI21xp33_ASAP7_75t_L     g09811(.A1(new_n10067), .A2(new_n10059), .B(new_n9899), .Y(new_n10068));
  AND3x1_ASAP7_75t_L        g09812(.A(new_n10067), .B(new_n10059), .C(new_n9899), .Y(new_n10069));
  NOR3xp33_ASAP7_75t_L      g09813(.A(new_n9892), .B(new_n10068), .C(new_n10069), .Y(new_n10070));
  NOR3xp33_ASAP7_75t_L      g09814(.A(new_n9730), .B(new_n9731), .C(new_n9738), .Y(new_n10071));
  INVx1_ASAP7_75t_L         g09815(.A(new_n10071), .Y(new_n10072));
  A2O1A1Ixp33_ASAP7_75t_L   g09816(.A1(new_n9744), .A2(new_n9743), .B(new_n9741), .C(new_n10072), .Y(new_n10073));
  AO21x2_ASAP7_75t_L        g09817(.A1(new_n10059), .A2(new_n10067), .B(new_n9899), .Y(new_n10074));
  NAND3xp33_ASAP7_75t_L     g09818(.A(new_n10067), .B(new_n10059), .C(new_n9899), .Y(new_n10075));
  AOI21xp33_ASAP7_75t_L     g09819(.A1(new_n10075), .A2(new_n10074), .B(new_n10073), .Y(new_n10076));
  NAND2xp33_ASAP7_75t_L     g09820(.A(\b[33] ), .B(new_n1910), .Y(new_n10077));
  NAND2xp33_ASAP7_75t_L     g09821(.A(\b[34] ), .B(new_n1770), .Y(new_n10078));
  AOI22xp33_ASAP7_75t_L     g09822(.A1(new_n1766), .A2(\b[35] ), .B1(new_n1764), .B2(new_n5649), .Y(new_n10079));
  AND4x1_ASAP7_75t_L        g09823(.A(new_n10079), .B(new_n10078), .C(new_n10077), .D(\a[23] ), .Y(new_n10080));
  AOI31xp33_ASAP7_75t_L     g09824(.A1(new_n10079), .A2(new_n10078), .A3(new_n10077), .B(\a[23] ), .Y(new_n10081));
  NOR2xp33_ASAP7_75t_L      g09825(.A(new_n10081), .B(new_n10080), .Y(new_n10082));
  INVx1_ASAP7_75t_L         g09826(.A(new_n10082), .Y(new_n10083));
  NOR3xp33_ASAP7_75t_L      g09827(.A(new_n10070), .B(new_n10076), .C(new_n10083), .Y(new_n10084));
  NAND3xp33_ASAP7_75t_L     g09828(.A(new_n10073), .B(new_n10074), .C(new_n10075), .Y(new_n10085));
  OAI21xp33_ASAP7_75t_L     g09829(.A1(new_n10068), .A2(new_n10069), .B(new_n9892), .Y(new_n10086));
  AOI21xp33_ASAP7_75t_L     g09830(.A1(new_n10085), .A2(new_n10086), .B(new_n10082), .Y(new_n10087));
  NOR2xp33_ASAP7_75t_L      g09831(.A(new_n10087), .B(new_n10084), .Y(new_n10088));
  NAND2xp33_ASAP7_75t_L     g09832(.A(new_n9742), .B(new_n9746), .Y(new_n10089));
  NOR2xp33_ASAP7_75t_L      g09833(.A(new_n9753), .B(new_n10089), .Y(new_n10090));
  O2A1O1Ixp33_ASAP7_75t_L   g09834(.A1(new_n9763), .A2(new_n9764), .B(new_n9766), .C(new_n10090), .Y(new_n10091));
  NAND2xp33_ASAP7_75t_L     g09835(.A(new_n10091), .B(new_n10088), .Y(new_n10092));
  NAND3xp33_ASAP7_75t_L     g09836(.A(new_n10085), .B(new_n10086), .C(new_n10082), .Y(new_n10093));
  OAI21xp33_ASAP7_75t_L     g09837(.A1(new_n10076), .A2(new_n10070), .B(new_n10083), .Y(new_n10094));
  NAND2xp33_ASAP7_75t_L     g09838(.A(new_n10093), .B(new_n10094), .Y(new_n10095));
  MAJIxp5_ASAP7_75t_L       g09839(.A(new_n9240), .B(new_n9431), .C(new_n9760), .Y(new_n10096));
  MAJIxp5_ASAP7_75t_L       g09840(.A(new_n10096), .B(new_n10089), .C(new_n9753), .Y(new_n10097));
  NAND2xp33_ASAP7_75t_L     g09841(.A(new_n10097), .B(new_n10095), .Y(new_n10098));
  AOI22xp33_ASAP7_75t_L     g09842(.A1(new_n1406), .A2(\b[38] ), .B1(new_n1404), .B2(new_n4923), .Y(new_n10099));
  OAI221xp5_ASAP7_75t_L     g09843(.A1(new_n1398), .A2(new_n4701), .B1(new_n4465), .B2(new_n1549), .C(new_n10099), .Y(new_n10100));
  XNOR2x2_ASAP7_75t_L       g09844(.A(new_n1401), .B(new_n10100), .Y(new_n10101));
  INVx1_ASAP7_75t_L         g09845(.A(new_n10101), .Y(new_n10102));
  NAND3xp33_ASAP7_75t_L     g09846(.A(new_n10102), .B(new_n10092), .C(new_n10098), .Y(new_n10103));
  NOR2xp33_ASAP7_75t_L      g09847(.A(new_n10097), .B(new_n10095), .Y(new_n10104));
  INVx1_ASAP7_75t_L         g09848(.A(new_n10090), .Y(new_n10105));
  AOI22xp33_ASAP7_75t_L     g09849(.A1(new_n10093), .A2(new_n10094), .B1(new_n10105), .B2(new_n9767), .Y(new_n10106));
  OAI21xp33_ASAP7_75t_L     g09850(.A1(new_n10106), .A2(new_n10104), .B(new_n10101), .Y(new_n10107));
  OAI211xp5_ASAP7_75t_L     g09851(.A1(new_n9771), .A2(new_n9773), .B(new_n9767), .C(new_n9762), .Y(new_n10108));
  NAND4xp25_ASAP7_75t_L     g09852(.A(new_n9780), .B(new_n10108), .C(new_n10107), .D(new_n10103), .Y(new_n10109));
  NOR3xp33_ASAP7_75t_L      g09853(.A(new_n10104), .B(new_n10106), .C(new_n10101), .Y(new_n10110));
  AOI21xp33_ASAP7_75t_L     g09854(.A1(new_n10092), .A2(new_n10098), .B(new_n10102), .Y(new_n10111));
  NAND2xp33_ASAP7_75t_L     g09855(.A(new_n9762), .B(new_n9767), .Y(new_n10112));
  MAJIxp5_ASAP7_75t_L       g09856(.A(new_n9778), .B(new_n10112), .C(new_n9774), .Y(new_n10113));
  OAI21xp33_ASAP7_75t_L     g09857(.A1(new_n10110), .A2(new_n10111), .B(new_n10113), .Y(new_n10114));
  NAND2xp33_ASAP7_75t_L     g09858(.A(\b[39] ), .B(new_n1194), .Y(new_n10115));
  NAND2xp33_ASAP7_75t_L     g09859(.A(\b[40] ), .B(new_n1103), .Y(new_n10116));
  AOI22xp33_ASAP7_75t_L     g09860(.A1(new_n1113), .A2(\b[41] ), .B1(new_n1110), .B2(new_n5669), .Y(new_n10117));
  AND4x1_ASAP7_75t_L        g09861(.A(new_n10117), .B(new_n10116), .C(new_n10115), .D(\a[17] ), .Y(new_n10118));
  AOI31xp33_ASAP7_75t_L     g09862(.A1(new_n10117), .A2(new_n10116), .A3(new_n10115), .B(\a[17] ), .Y(new_n10119));
  NOR2xp33_ASAP7_75t_L      g09863(.A(new_n10119), .B(new_n10118), .Y(new_n10120));
  NAND3xp33_ASAP7_75t_L     g09864(.A(new_n10109), .B(new_n10114), .C(new_n10120), .Y(new_n10121));
  NOR3xp33_ASAP7_75t_L      g09865(.A(new_n10113), .B(new_n10111), .C(new_n10110), .Y(new_n10122));
  OA21x2_ASAP7_75t_L        g09866(.A1(new_n10110), .A2(new_n10111), .B(new_n10113), .Y(new_n10123));
  INVx1_ASAP7_75t_L         g09867(.A(new_n10120), .Y(new_n10124));
  OAI21xp33_ASAP7_75t_L     g09868(.A1(new_n10122), .A2(new_n10123), .B(new_n10124), .Y(new_n10125));
  NAND2xp33_ASAP7_75t_L     g09869(.A(new_n9779), .B(new_n9780), .Y(new_n10126));
  NOR2xp33_ASAP7_75t_L      g09870(.A(new_n9787), .B(new_n10126), .Y(new_n10127));
  INVx1_ASAP7_75t_L         g09871(.A(new_n10127), .Y(new_n10128));
  NAND4xp25_ASAP7_75t_L     g09872(.A(new_n9890), .B(new_n10128), .C(new_n10125), .D(new_n10121), .Y(new_n10129));
  NAND2xp33_ASAP7_75t_L     g09873(.A(new_n10121), .B(new_n10125), .Y(new_n10130));
  A2O1A1Ixp33_ASAP7_75t_L   g09874(.A1(new_n9793), .A2(new_n9795), .B(new_n10127), .C(new_n10130), .Y(new_n10131));
  NOR2xp33_ASAP7_75t_L      g09875(.A(new_n5680), .B(new_n909), .Y(new_n10132));
  NAND2xp33_ASAP7_75t_L     g09876(.A(\b[43] ), .B(new_n817), .Y(new_n10133));
  AOI22xp33_ASAP7_75t_L     g09877(.A1(new_n826), .A2(\b[44] ), .B1(new_n823), .B2(new_n7055), .Y(new_n10134));
  NAND2xp33_ASAP7_75t_L     g09878(.A(new_n10133), .B(new_n10134), .Y(new_n10135));
  OR3x1_ASAP7_75t_L         g09879(.A(new_n10135), .B(new_n813), .C(new_n10132), .Y(new_n10136));
  A2O1A1Ixp33_ASAP7_75t_L   g09880(.A1(\b[42] ), .A2(new_n908), .B(new_n10135), .C(new_n813), .Y(new_n10137));
  NAND2xp33_ASAP7_75t_L     g09881(.A(new_n10137), .B(new_n10136), .Y(new_n10138));
  AOI21xp33_ASAP7_75t_L     g09882(.A1(new_n10131), .A2(new_n10129), .B(new_n10138), .Y(new_n10139));
  NAND3xp33_ASAP7_75t_L     g09883(.A(new_n9452), .B(new_n9462), .C(new_n9449), .Y(new_n10140));
  A2O1A1Ixp33_ASAP7_75t_L   g09884(.A1(new_n10140), .A2(new_n9479), .B(new_n9797), .C(new_n10128), .Y(new_n10141));
  NOR2xp33_ASAP7_75t_L      g09885(.A(new_n10130), .B(new_n10141), .Y(new_n10142));
  NOR3xp33_ASAP7_75t_L      g09886(.A(new_n10123), .B(new_n10124), .C(new_n10122), .Y(new_n10143));
  AOI21xp33_ASAP7_75t_L     g09887(.A1(new_n10109), .A2(new_n10114), .B(new_n10120), .Y(new_n10144));
  NOR2xp33_ASAP7_75t_L      g09888(.A(new_n10144), .B(new_n10143), .Y(new_n10145));
  O2A1O1Ixp33_ASAP7_75t_L   g09889(.A1(new_n9787), .A2(new_n10126), .B(new_n9890), .C(new_n10145), .Y(new_n10146));
  INVx1_ASAP7_75t_L         g09890(.A(new_n10138), .Y(new_n10147));
  NOR3xp33_ASAP7_75t_L      g09891(.A(new_n10142), .B(new_n10147), .C(new_n10146), .Y(new_n10148));
  A2O1A1O1Ixp25_ASAP7_75t_L g09892(.A1(new_n9475), .A2(new_n9228), .B(new_n9486), .C(new_n9806), .D(new_n9811), .Y(new_n10149));
  NOR3xp33_ASAP7_75t_L      g09893(.A(new_n10149), .B(new_n10148), .C(new_n10139), .Y(new_n10150));
  OAI21xp33_ASAP7_75t_L     g09894(.A1(new_n10146), .A2(new_n10142), .B(new_n10147), .Y(new_n10151));
  NAND3xp33_ASAP7_75t_L     g09895(.A(new_n10131), .B(new_n10129), .C(new_n10138), .Y(new_n10152));
  OAI21xp33_ASAP7_75t_L     g09896(.A1(new_n9810), .A2(new_n9564), .B(new_n9807), .Y(new_n10153));
  AOI21xp33_ASAP7_75t_L     g09897(.A1(new_n10152), .A2(new_n10151), .B(new_n10153), .Y(new_n10154));
  NOR3xp33_ASAP7_75t_L      g09898(.A(new_n10154), .B(new_n10150), .C(new_n9888), .Y(new_n10155));
  INVx1_ASAP7_75t_L         g09899(.A(new_n10155), .Y(new_n10156));
  OAI21xp33_ASAP7_75t_L     g09900(.A1(new_n10150), .A2(new_n10154), .B(new_n9888), .Y(new_n10157));
  NAND3xp33_ASAP7_75t_L     g09901(.A(new_n9880), .B(new_n10156), .C(new_n10157), .Y(new_n10158));
  A2O1A1O1Ixp25_ASAP7_75t_L g09902(.A1(new_n9495), .A2(new_n9827), .B(new_n9828), .C(new_n9813), .D(new_n9822), .Y(new_n10159));
  INVx1_ASAP7_75t_L         g09903(.A(new_n10157), .Y(new_n10160));
  OAI21xp33_ASAP7_75t_L     g09904(.A1(new_n10155), .A2(new_n10160), .B(new_n10159), .Y(new_n10161));
  AO21x2_ASAP7_75t_L        g09905(.A1(new_n10161), .A2(new_n10158), .B(new_n9878), .Y(new_n10162));
  NAND3xp33_ASAP7_75t_L     g09906(.A(new_n10158), .B(new_n9878), .C(new_n10161), .Y(new_n10163));
  AOI21xp33_ASAP7_75t_L     g09907(.A1(new_n10162), .A2(new_n10163), .B(new_n9871), .Y(new_n10164));
  NAND3xp33_ASAP7_75t_L     g09908(.A(new_n9871), .B(new_n10162), .C(new_n10163), .Y(new_n10165));
  INVx1_ASAP7_75t_L         g09909(.A(new_n10165), .Y(new_n10166));
  OAI21xp33_ASAP7_75t_L     g09910(.A1(new_n10164), .A2(new_n10166), .B(new_n9870), .Y(new_n10167));
  INVx1_ASAP7_75t_L         g09911(.A(new_n9870), .Y(new_n10168));
  INVx1_ASAP7_75t_L         g09912(.A(new_n10164), .Y(new_n10169));
  NAND3xp33_ASAP7_75t_L     g09913(.A(new_n10169), .B(new_n10168), .C(new_n10165), .Y(new_n10170));
  NAND3xp33_ASAP7_75t_L     g09914(.A(new_n9864), .B(new_n10167), .C(new_n10170), .Y(new_n10171));
  OAI21xp33_ASAP7_75t_L     g09915(.A1(new_n9852), .A2(new_n9853), .B(new_n9851), .Y(new_n10172));
  AOI21xp33_ASAP7_75t_L     g09916(.A1(new_n10169), .A2(new_n10165), .B(new_n10168), .Y(new_n10173));
  NOR3xp33_ASAP7_75t_L      g09917(.A(new_n10166), .B(new_n10164), .C(new_n9870), .Y(new_n10174));
  OAI211xp5_ASAP7_75t_L     g09918(.A1(new_n10173), .A2(new_n10174), .B(new_n10172), .C(new_n9863), .Y(new_n10175));
  NAND2xp33_ASAP7_75t_L     g09919(.A(new_n10175), .B(new_n10171), .Y(new_n10176));
  NOR2xp33_ASAP7_75t_L      g09920(.A(\b[55] ), .B(\b[56] ), .Y(new_n10177));
  INVx1_ASAP7_75t_L         g09921(.A(\b[56] ), .Y(new_n10178));
  NOR2xp33_ASAP7_75t_L      g09922(.A(new_n9534), .B(new_n10178), .Y(new_n10179));
  NOR2xp33_ASAP7_75t_L      g09923(.A(new_n10177), .B(new_n10179), .Y(new_n10180));
  A2O1A1Ixp33_ASAP7_75t_L   g09924(.A1(new_n9540), .A2(new_n9536), .B(new_n9535), .C(new_n10180), .Y(new_n10181));
  O2A1O1Ixp33_ASAP7_75t_L   g09925(.A1(new_n9200), .A2(new_n9203), .B(new_n9536), .C(new_n9535), .Y(new_n10182));
  OAI21xp33_ASAP7_75t_L     g09926(.A1(new_n10177), .A2(new_n10179), .B(new_n10182), .Y(new_n10183));
  NAND2xp33_ASAP7_75t_L     g09927(.A(new_n10181), .B(new_n10183), .Y(new_n10184));
  INVx1_ASAP7_75t_L         g09928(.A(new_n10184), .Y(new_n10185));
  AOI22xp33_ASAP7_75t_L     g09929(.A1(new_n272), .A2(\b[56] ), .B1(new_n269), .B2(new_n10185), .Y(new_n10186));
  OAI221xp5_ASAP7_75t_L     g09930(.A1(new_n261), .A2(new_n9534), .B1(new_n9199), .B2(new_n277), .C(new_n10186), .Y(new_n10187));
  XNOR2x2_ASAP7_75t_L       g09931(.A(\a[2] ), .B(new_n10187), .Y(new_n10188));
  XNOR2x2_ASAP7_75t_L       g09932(.A(new_n10188), .B(new_n10176), .Y(new_n10189));
  A2O1A1O1Ixp25_ASAP7_75t_L g09933(.A1(new_n9529), .A2(new_n9196), .B(new_n9527), .C(new_n9857), .D(new_n9855), .Y(new_n10190));
  XOR2x2_ASAP7_75t_L        g09934(.A(new_n10190), .B(new_n10189), .Y(\f[56] ));
  MAJIxp5_ASAP7_75t_L       g09935(.A(new_n10190), .B(new_n10188), .C(new_n10176), .Y(new_n10192));
  NOR2xp33_ASAP7_75t_L      g09936(.A(new_n8569), .B(new_n365), .Y(new_n10193));
  INVx1_ASAP7_75t_L         g09937(.A(new_n10193), .Y(new_n10194));
  NAND2xp33_ASAP7_75t_L     g09938(.A(\b[53] ), .B(new_n334), .Y(new_n10195));
  AOI22xp33_ASAP7_75t_L     g09939(.A1(new_n345), .A2(\b[54] ), .B1(new_n342), .B2(new_n9208), .Y(new_n10196));
  AND4x1_ASAP7_75t_L        g09940(.A(new_n10196), .B(new_n10195), .C(new_n10194), .D(\a[5] ), .Y(new_n10197));
  AOI31xp33_ASAP7_75t_L     g09941(.A1(new_n10196), .A2(new_n10195), .A3(new_n10194), .B(\a[5] ), .Y(new_n10198));
  NOR2xp33_ASAP7_75t_L      g09942(.A(new_n10198), .B(new_n10197), .Y(new_n10199));
  NAND2xp33_ASAP7_75t_L     g09943(.A(new_n10161), .B(new_n10158), .Y(new_n10200));
  MAJIxp5_ASAP7_75t_L       g09944(.A(new_n9871), .B(new_n9878), .C(new_n10200), .Y(new_n10201));
  NOR2xp33_ASAP7_75t_L      g09945(.A(new_n7907), .B(new_n481), .Y(new_n10202));
  INVx1_ASAP7_75t_L         g09946(.A(new_n10202), .Y(new_n10203));
  NAND2xp33_ASAP7_75t_L     g09947(.A(\b[50] ), .B(new_n441), .Y(new_n10204));
  AOI22xp33_ASAP7_75t_L     g09948(.A1(new_n451), .A2(\b[51] ), .B1(new_n448), .B2(new_n8257), .Y(new_n10205));
  AND4x1_ASAP7_75t_L        g09949(.A(new_n10205), .B(new_n10204), .C(new_n10203), .D(\a[8] ), .Y(new_n10206));
  AOI31xp33_ASAP7_75t_L     g09950(.A1(new_n10205), .A2(new_n10204), .A3(new_n10203), .B(\a[8] ), .Y(new_n10207));
  NOR2xp33_ASAP7_75t_L      g09951(.A(new_n10207), .B(new_n10206), .Y(new_n10208));
  INVx1_ASAP7_75t_L         g09952(.A(new_n10208), .Y(new_n10209));
  A2O1A1O1Ixp25_ASAP7_75t_L g09953(.A1(new_n9813), .A2(new_n9557), .B(new_n9822), .C(new_n10157), .D(new_n10155), .Y(new_n10210));
  NAND2xp33_ASAP7_75t_L     g09954(.A(\b[46] ), .B(new_n674), .Y(new_n10211));
  NAND2xp33_ASAP7_75t_L     g09955(.A(\b[47] ), .B(new_n590), .Y(new_n10212));
  AOI22xp33_ASAP7_75t_L     g09956(.A1(new_n600), .A2(\b[48] ), .B1(new_n597), .B2(new_n7341), .Y(new_n10213));
  AND4x1_ASAP7_75t_L        g09957(.A(new_n10213), .B(new_n10212), .C(new_n10211), .D(\a[11] ), .Y(new_n10214));
  AOI31xp33_ASAP7_75t_L     g09958(.A1(new_n10213), .A2(new_n10212), .A3(new_n10211), .B(\a[11] ), .Y(new_n10215));
  NOR2xp33_ASAP7_75t_L      g09959(.A(new_n10215), .B(new_n10214), .Y(new_n10216));
  INVx1_ASAP7_75t_L         g09960(.A(new_n10216), .Y(new_n10217));
  NAND2xp33_ASAP7_75t_L     g09961(.A(new_n823), .B(new_n6764), .Y(new_n10218));
  OAI221xp5_ASAP7_75t_L     g09962(.A1(new_n912), .A2(new_n6756), .B1(new_n6220), .B2(new_n994), .C(new_n10218), .Y(new_n10219));
  AOI21xp33_ASAP7_75t_L     g09963(.A1(new_n908), .A2(\b[43] ), .B(new_n10219), .Y(new_n10220));
  NAND2xp33_ASAP7_75t_L     g09964(.A(\a[14] ), .B(new_n10220), .Y(new_n10221));
  A2O1A1Ixp33_ASAP7_75t_L   g09965(.A1(\b[43] ), .A2(new_n908), .B(new_n10219), .C(new_n813), .Y(new_n10222));
  AND2x2_ASAP7_75t_L        g09966(.A(new_n10222), .B(new_n10221), .Y(new_n10223));
  NOR3xp33_ASAP7_75t_L      g09967(.A(new_n10123), .B(new_n10120), .C(new_n10122), .Y(new_n10224));
  INVx1_ASAP7_75t_L         g09968(.A(new_n10224), .Y(new_n10225));
  A2O1A1Ixp33_ASAP7_75t_L   g09969(.A1(new_n9890), .A2(new_n10128), .B(new_n10145), .C(new_n10225), .Y(new_n10226));
  NOR3xp33_ASAP7_75t_L      g09970(.A(new_n10070), .B(new_n10076), .C(new_n10082), .Y(new_n10227));
  O2A1O1Ixp33_ASAP7_75t_L   g09971(.A1(new_n10084), .A2(new_n10087), .B(new_n10097), .C(new_n10227), .Y(new_n10228));
  NAND2xp33_ASAP7_75t_L     g09972(.A(\b[35] ), .B(new_n1770), .Y(new_n10229));
  AOI22xp33_ASAP7_75t_L     g09973(.A1(new_n1766), .A2(\b[36] ), .B1(new_n1764), .B2(new_n4473), .Y(new_n10230));
  NAND2xp33_ASAP7_75t_L     g09974(.A(new_n10229), .B(new_n10230), .Y(new_n10231));
  AOI21xp33_ASAP7_75t_L     g09975(.A1(new_n1910), .A2(\b[34] ), .B(new_n10231), .Y(new_n10232));
  NAND2xp33_ASAP7_75t_L     g09976(.A(\a[23] ), .B(new_n10232), .Y(new_n10233));
  A2O1A1Ixp33_ASAP7_75t_L   g09977(.A1(\b[34] ), .A2(new_n1910), .B(new_n10231), .C(new_n1761), .Y(new_n10234));
  NAND2xp33_ASAP7_75t_L     g09978(.A(new_n10234), .B(new_n10233), .Y(new_n10235));
  A2O1A1O1Ixp25_ASAP7_75t_L g09979(.A1(new_n9755), .A2(new_n9745), .B(new_n10071), .C(new_n10074), .D(new_n10069), .Y(new_n10236));
  NAND2xp33_ASAP7_75t_L     g09980(.A(new_n2700), .B(new_n3219), .Y(new_n10237));
  OAI221xp5_ASAP7_75t_L     g09981(.A1(new_n2708), .A2(new_n3212), .B1(new_n2871), .B2(new_n2694), .C(new_n10237), .Y(new_n10238));
  AOI21xp33_ASAP7_75t_L     g09982(.A1(new_n2931), .A2(\b[28] ), .B(new_n10238), .Y(new_n10239));
  NAND2xp33_ASAP7_75t_L     g09983(.A(\a[29] ), .B(new_n10239), .Y(new_n10240));
  A2O1A1Ixp33_ASAP7_75t_L   g09984(.A1(\b[28] ), .A2(new_n2931), .B(new_n10238), .C(new_n2697), .Y(new_n10241));
  AND2x2_ASAP7_75t_L        g09985(.A(new_n10241), .B(new_n10240), .Y(new_n10242));
  A2O1A1Ixp33_ASAP7_75t_L   g09986(.A1(new_n9690), .A2(new_n9691), .B(new_n9573), .C(new_n9684), .Y(new_n10243));
  A2O1A1Ixp33_ASAP7_75t_L   g09987(.A1(new_n10243), .A2(new_n9688), .B(new_n10018), .C(new_n10022), .Y(new_n10244));
  AOI22xp33_ASAP7_75t_L     g09988(.A1(new_n4544), .A2(\b[21] ), .B1(new_n4542), .B2(new_n1715), .Y(new_n10245));
  OAI221xp5_ASAP7_75t_L     g09989(.A1(new_n4536), .A2(new_n1594), .B1(new_n1493), .B2(new_n4781), .C(new_n10245), .Y(new_n10246));
  XNOR2x2_ASAP7_75t_L       g09990(.A(\a[38] ), .B(new_n10246), .Y(new_n10247));
  INVx1_ASAP7_75t_L         g09991(.A(new_n10247), .Y(new_n10248));
  NOR3xp33_ASAP7_75t_L      g09992(.A(new_n9922), .B(new_n9999), .C(new_n9998), .Y(new_n10249));
  O2A1O1Ixp33_ASAP7_75t_L   g09993(.A1(new_n9996), .A2(new_n10000), .B(new_n9916), .C(new_n10249), .Y(new_n10250));
  AOI22xp33_ASAP7_75t_L     g09994(.A1(new_n5249), .A2(\b[18] ), .B1(new_n5247), .B2(new_n1363), .Y(new_n10251));
  OAI221xp5_ASAP7_75t_L     g09995(.A1(new_n5241), .A2(new_n1244), .B1(new_n1051), .B2(new_n5521), .C(new_n10251), .Y(new_n10252));
  XNOR2x2_ASAP7_75t_L       g09996(.A(\a[41] ), .B(new_n10252), .Y(new_n10253));
  NAND3xp33_ASAP7_75t_L     g09997(.A(new_n9978), .B(new_n9982), .C(new_n9992), .Y(new_n10254));
  A2O1A1Ixp33_ASAP7_75t_L   g09998(.A1(new_n9993), .A2(new_n9989), .B(new_n9924), .C(new_n10254), .Y(new_n10255));
  NAND2xp33_ASAP7_75t_L     g09999(.A(\b[13] ), .B(new_n6308), .Y(new_n10256));
  AOI22xp33_ASAP7_75t_L     g10000(.A1(new_n6002), .A2(\b[15] ), .B1(new_n5999), .B2(new_n959), .Y(new_n10257));
  OAI211xp5_ASAP7_75t_L     g10001(.A1(new_n871), .A2(new_n6544), .B(new_n10257), .C(new_n10256), .Y(new_n10258));
  XNOR2x2_ASAP7_75t_L       g10002(.A(\a[44] ), .B(new_n10258), .Y(new_n10259));
  NOR3xp33_ASAP7_75t_L      g10003(.A(new_n9968), .B(new_n9972), .C(new_n9932), .Y(new_n10260));
  A2O1A1O1Ixp25_ASAP7_75t_L g10004(.A1(new_n9645), .A2(new_n9652), .B(new_n9979), .C(new_n9973), .D(new_n10260), .Y(new_n10261));
  NAND2xp33_ASAP7_75t_L     g10005(.A(\b[10] ), .B(new_n7124), .Y(new_n10262));
  NAND2xp33_ASAP7_75t_L     g10006(.A(\b[11] ), .B(new_n6812), .Y(new_n10263));
  AOI22xp33_ASAP7_75t_L     g10007(.A1(new_n6822), .A2(\b[12] ), .B1(new_n6819), .B2(new_n970), .Y(new_n10264));
  NAND4xp25_ASAP7_75t_L     g10008(.A(new_n10264), .B(\a[47] ), .C(new_n10262), .D(new_n10263), .Y(new_n10265));
  NAND2xp33_ASAP7_75t_L     g10009(.A(new_n10263), .B(new_n10264), .Y(new_n10266));
  A2O1A1Ixp33_ASAP7_75t_L   g10010(.A1(\b[10] ), .A2(new_n7124), .B(new_n10266), .C(new_n6816), .Y(new_n10267));
  NAND2xp33_ASAP7_75t_L     g10011(.A(new_n10265), .B(new_n10267), .Y(new_n10268));
  A2O1A1Ixp33_ASAP7_75t_L   g10012(.A1(new_n9646), .A2(new_n9643), .B(new_n9966), .C(new_n9971), .Y(new_n10269));
  NAND3xp33_ASAP7_75t_L     g10013(.A(new_n9946), .B(new_n9319), .C(\a[56] ), .Y(new_n10270));
  AO21x2_ASAP7_75t_L        g10014(.A1(\b[0] ), .A2(new_n9948), .B(new_n9952), .Y(new_n10271));
  INVx1_ASAP7_75t_L         g10015(.A(\a[57] ), .Y(new_n10272));
  NAND2xp33_ASAP7_75t_L     g10016(.A(\a[56] ), .B(new_n10272), .Y(new_n10273));
  NAND2xp33_ASAP7_75t_L     g10017(.A(\a[57] ), .B(new_n9610), .Y(new_n10274));
  AND2x2_ASAP7_75t_L        g10018(.A(new_n10273), .B(new_n10274), .Y(new_n10275));
  NOR2xp33_ASAP7_75t_L      g10019(.A(new_n258), .B(new_n10275), .Y(new_n10276));
  OAI21xp33_ASAP7_75t_L     g10020(.A1(new_n10271), .A2(new_n10270), .B(new_n10276), .Y(new_n10277));
  INVx1_ASAP7_75t_L         g10021(.A(new_n10276), .Y(new_n10278));
  NAND5xp2_ASAP7_75t_L      g10022(.A(\a[56] ), .B(new_n9953), .C(new_n10278), .D(new_n9946), .E(new_n9319), .Y(new_n10279));
  INVx1_ASAP7_75t_L         g10023(.A(new_n9614), .Y(new_n10280));
  NAND2xp33_ASAP7_75t_L     g10024(.A(\b[3] ), .B(new_n9623), .Y(new_n10281));
  OAI221xp5_ASAP7_75t_L     g10025(.A1(new_n278), .A2(new_n10280), .B1(new_n9949), .B2(new_n303), .C(new_n10281), .Y(new_n10282));
  AOI21xp33_ASAP7_75t_L     g10026(.A1(new_n9948), .A2(\b[1] ), .B(new_n10282), .Y(new_n10283));
  NAND2xp33_ASAP7_75t_L     g10027(.A(\a[56] ), .B(new_n10283), .Y(new_n10284));
  A2O1A1Ixp33_ASAP7_75t_L   g10028(.A1(\b[1] ), .A2(new_n9948), .B(new_n10282), .C(new_n9610), .Y(new_n10285));
  AO22x1_ASAP7_75t_L        g10029(.A1(new_n10285), .A2(new_n10284), .B1(new_n10279), .B2(new_n10277), .Y(new_n10286));
  NAND4xp25_ASAP7_75t_L     g10030(.A(new_n10277), .B(new_n10285), .C(new_n10284), .D(new_n10279), .Y(new_n10287));
  NOR2xp33_ASAP7_75t_L      g10031(.A(new_n382), .B(new_n8968), .Y(new_n10288));
  AOI221xp5_ASAP7_75t_L     g10032(.A1(new_n8635), .A2(\b[5] ), .B1(new_n8642), .B2(new_n389), .C(new_n10288), .Y(new_n10289));
  OAI211xp5_ASAP7_75t_L     g10033(.A1(new_n323), .A2(new_n8965), .B(new_n10289), .C(\a[53] ), .Y(new_n10290));
  INVx1_ASAP7_75t_L         g10034(.A(new_n10289), .Y(new_n10291));
  A2O1A1Ixp33_ASAP7_75t_L   g10035(.A1(\b[4] ), .A2(new_n8964), .B(new_n10291), .C(new_n8639), .Y(new_n10292));
  AND4x1_ASAP7_75t_L        g10036(.A(new_n10286), .B(new_n10292), .C(new_n10287), .D(new_n10290), .Y(new_n10293));
  AOI22xp33_ASAP7_75t_L     g10037(.A1(new_n10286), .A2(new_n10287), .B1(new_n10290), .B2(new_n10292), .Y(new_n10294));
  NOR2xp33_ASAP7_75t_L      g10038(.A(new_n10294), .B(new_n10293), .Y(new_n10295));
  A2O1A1O1Ixp25_ASAP7_75t_L g10039(.A1(new_n9602), .A2(new_n9328), .B(new_n9632), .C(new_n9629), .D(new_n9963), .Y(new_n10296));
  OAI21xp33_ASAP7_75t_L     g10040(.A1(new_n10296), .A2(new_n9964), .B(new_n10295), .Y(new_n10297));
  A2O1A1O1Ixp25_ASAP7_75t_L g10041(.A1(new_n9627), .A2(new_n9603), .B(new_n9628), .C(new_n9958), .D(new_n9964), .Y(new_n10298));
  OAI21xp33_ASAP7_75t_L     g10042(.A1(new_n10293), .A2(new_n10294), .B(new_n10298), .Y(new_n10299));
  NAND2xp33_ASAP7_75t_L     g10043(.A(\b[7] ), .B(new_n7993), .Y(new_n10300));
  NAND2xp33_ASAP7_75t_L     g10044(.A(\b[8] ), .B(new_n7649), .Y(new_n10301));
  AOI22xp33_ASAP7_75t_L     g10045(.A1(new_n7659), .A2(\b[9] ), .B1(new_n7656), .B2(new_n566), .Y(new_n10302));
  NAND4xp25_ASAP7_75t_L     g10046(.A(new_n10302), .B(\a[50] ), .C(new_n10300), .D(new_n10301), .Y(new_n10303));
  NAND2xp33_ASAP7_75t_L     g10047(.A(new_n10301), .B(new_n10302), .Y(new_n10304));
  A2O1A1Ixp33_ASAP7_75t_L   g10048(.A1(\b[7] ), .A2(new_n7993), .B(new_n10304), .C(new_n7653), .Y(new_n10305));
  AO22x1_ASAP7_75t_L        g10049(.A1(new_n10305), .A2(new_n10303), .B1(new_n10299), .B2(new_n10297), .Y(new_n10306));
  NAND4xp25_ASAP7_75t_L     g10050(.A(new_n10297), .B(new_n10305), .C(new_n10303), .D(new_n10299), .Y(new_n10307));
  NAND3xp33_ASAP7_75t_L     g10051(.A(new_n10269), .B(new_n10306), .C(new_n10307), .Y(new_n10308));
  A2O1A1O1Ixp25_ASAP7_75t_L g10052(.A1(new_n9642), .A2(new_n9641), .B(new_n9639), .C(new_n9970), .D(new_n9967), .Y(new_n10309));
  AOI22xp33_ASAP7_75t_L     g10053(.A1(new_n10303), .A2(new_n10305), .B1(new_n10299), .B2(new_n10297), .Y(new_n10310));
  AND4x1_ASAP7_75t_L        g10054(.A(new_n10297), .B(new_n10305), .C(new_n10303), .D(new_n10299), .Y(new_n10311));
  OAI21xp33_ASAP7_75t_L     g10055(.A1(new_n10310), .A2(new_n10311), .B(new_n10309), .Y(new_n10312));
  AOI21xp33_ASAP7_75t_L     g10056(.A1(new_n10308), .A2(new_n10312), .B(new_n10268), .Y(new_n10313));
  NOR3xp33_ASAP7_75t_L      g10057(.A(new_n10309), .B(new_n10311), .C(new_n10310), .Y(new_n10314));
  INVx1_ASAP7_75t_L         g10058(.A(new_n10312), .Y(new_n10315));
  AOI211xp5_ASAP7_75t_L     g10059(.A1(new_n10265), .A2(new_n10267), .B(new_n10314), .C(new_n10315), .Y(new_n10316));
  NOR3xp33_ASAP7_75t_L      g10060(.A(new_n10316), .B(new_n10261), .C(new_n10313), .Y(new_n10317));
  OA21x2_ASAP7_75t_L        g10061(.A1(new_n10313), .A2(new_n10316), .B(new_n10261), .Y(new_n10318));
  OR3x1_ASAP7_75t_L         g10062(.A(new_n10259), .B(new_n10317), .C(new_n10318), .Y(new_n10319));
  OAI21xp33_ASAP7_75t_L     g10063(.A1(new_n10317), .A2(new_n10318), .B(new_n10259), .Y(new_n10320));
  NAND3xp33_ASAP7_75t_L     g10064(.A(new_n10255), .B(new_n10319), .C(new_n10320), .Y(new_n10321));
  NOR3xp33_ASAP7_75t_L      g10065(.A(new_n9991), .B(new_n9992), .C(new_n9990), .Y(new_n10322));
  AOI21xp33_ASAP7_75t_L     g10066(.A1(new_n9978), .A2(new_n9982), .B(new_n9988), .Y(new_n10323));
  NOR2xp33_ASAP7_75t_L      g10067(.A(new_n10323), .B(new_n10322), .Y(new_n10324));
  NOR3xp33_ASAP7_75t_L      g10068(.A(new_n10259), .B(new_n10318), .C(new_n10317), .Y(new_n10325));
  OA21x2_ASAP7_75t_L        g10069(.A1(new_n10317), .A2(new_n10318), .B(new_n10259), .Y(new_n10326));
  OAI221xp5_ASAP7_75t_L     g10070(.A1(new_n10326), .A2(new_n10325), .B1(new_n9924), .B2(new_n10324), .C(new_n10254), .Y(new_n10327));
  AO21x2_ASAP7_75t_L        g10071(.A1(new_n10321), .A2(new_n10327), .B(new_n10253), .Y(new_n10328));
  NAND3xp33_ASAP7_75t_L     g10072(.A(new_n10327), .B(new_n10321), .C(new_n10253), .Y(new_n10329));
  NAND2xp33_ASAP7_75t_L     g10073(.A(new_n10329), .B(new_n10328), .Y(new_n10330));
  XNOR2x2_ASAP7_75t_L       g10074(.A(new_n10250), .B(new_n10330), .Y(new_n10331));
  NAND2xp33_ASAP7_75t_L     g10075(.A(new_n10248), .B(new_n10331), .Y(new_n10332));
  INVx1_ASAP7_75t_L         g10076(.A(new_n10249), .Y(new_n10333));
  AOI21xp33_ASAP7_75t_L     g10077(.A1(new_n10327), .A2(new_n10321), .B(new_n10253), .Y(new_n10334));
  AND3x1_ASAP7_75t_L        g10078(.A(new_n10327), .B(new_n10321), .C(new_n10253), .Y(new_n10335));
  NOR2xp33_ASAP7_75t_L      g10079(.A(new_n10334), .B(new_n10335), .Y(new_n10336));
  A2O1A1O1Ixp25_ASAP7_75t_L g10080(.A1(new_n10003), .A2(new_n9686), .B(new_n10001), .C(new_n10333), .D(new_n10336), .Y(new_n10337));
  A2O1A1Ixp33_ASAP7_75t_L   g10081(.A1(new_n9686), .A2(new_n10003), .B(new_n10001), .C(new_n10333), .Y(new_n10338));
  NOR2xp33_ASAP7_75t_L      g10082(.A(new_n10330), .B(new_n10338), .Y(new_n10339));
  OAI21xp33_ASAP7_75t_L     g10083(.A1(new_n10339), .A2(new_n10337), .B(new_n10247), .Y(new_n10340));
  NAND3xp33_ASAP7_75t_L     g10084(.A(new_n10332), .B(new_n10244), .C(new_n10340), .Y(new_n10341));
  NOR3xp33_ASAP7_75t_L      g10085(.A(new_n10337), .B(new_n10339), .C(new_n10247), .Y(new_n10342));
  NOR2xp33_ASAP7_75t_L      g10086(.A(new_n10248), .B(new_n10331), .Y(new_n10343));
  OAI211xp5_ASAP7_75t_L     g10087(.A1(new_n10342), .A2(new_n10343), .B(new_n10029), .C(new_n10022), .Y(new_n10344));
  AOI22xp33_ASAP7_75t_L     g10088(.A1(new_n3884), .A2(\b[24] ), .B1(new_n3881), .B2(new_n2027), .Y(new_n10345));
  OAI221xp5_ASAP7_75t_L     g10089(.A1(new_n4312), .A2(new_n1995), .B1(new_n1857), .B2(new_n4986), .C(new_n10345), .Y(new_n10346));
  XNOR2x2_ASAP7_75t_L       g10090(.A(\a[35] ), .B(new_n10346), .Y(new_n10347));
  NAND3xp33_ASAP7_75t_L     g10091(.A(new_n10344), .B(new_n10347), .C(new_n10341), .Y(new_n10348));
  AOI211xp5_ASAP7_75t_L     g10092(.A1(new_n10022), .A2(new_n10029), .B(new_n10342), .C(new_n10343), .Y(new_n10349));
  AOI21xp33_ASAP7_75t_L     g10093(.A1(new_n10332), .A2(new_n10340), .B(new_n10244), .Y(new_n10350));
  INVx1_ASAP7_75t_L         g10094(.A(new_n10347), .Y(new_n10351));
  OAI21xp33_ASAP7_75t_L     g10095(.A1(new_n10350), .A2(new_n10349), .B(new_n10351), .Y(new_n10352));
  A2O1A1O1Ixp25_ASAP7_75t_L g10096(.A1(new_n9700), .A2(new_n9702), .B(new_n9694), .C(new_n10035), .D(new_n10027), .Y(new_n10353));
  AND3x1_ASAP7_75t_L        g10097(.A(new_n10353), .B(new_n10352), .C(new_n10348), .Y(new_n10354));
  AOI21xp33_ASAP7_75t_L     g10098(.A1(new_n10348), .A2(new_n10352), .B(new_n10353), .Y(new_n10355));
  NAND2xp33_ASAP7_75t_L     g10099(.A(new_n3254), .B(new_n2657), .Y(new_n10356));
  OAI221xp5_ASAP7_75t_L     g10100(.A1(new_n3262), .A2(new_n2650), .B1(new_n2477), .B2(new_n3248), .C(new_n10356), .Y(new_n10357));
  AOI21xp33_ASAP7_75t_L     g10101(.A1(new_n3491), .A2(\b[25] ), .B(new_n10357), .Y(new_n10358));
  NAND2xp33_ASAP7_75t_L     g10102(.A(\a[32] ), .B(new_n10358), .Y(new_n10359));
  A2O1A1Ixp33_ASAP7_75t_L   g10103(.A1(\b[25] ), .A2(new_n3491), .B(new_n10357), .C(new_n3251), .Y(new_n10360));
  AND2x2_ASAP7_75t_L        g10104(.A(new_n10360), .B(new_n10359), .Y(new_n10361));
  OAI21xp33_ASAP7_75t_L     g10105(.A1(new_n10355), .A2(new_n10354), .B(new_n10361), .Y(new_n10362));
  NAND3xp33_ASAP7_75t_L     g10106(.A(new_n10353), .B(new_n10348), .C(new_n10352), .Y(new_n10363));
  AO21x2_ASAP7_75t_L        g10107(.A1(new_n10348), .A2(new_n10352), .B(new_n10353), .Y(new_n10364));
  NAND2xp33_ASAP7_75t_L     g10108(.A(new_n10360), .B(new_n10359), .Y(new_n10365));
  NAND3xp33_ASAP7_75t_L     g10109(.A(new_n10364), .B(new_n10363), .C(new_n10365), .Y(new_n10366));
  NAND2xp33_ASAP7_75t_L     g10110(.A(new_n10366), .B(new_n10362), .Y(new_n10367));
  O2A1O1Ixp33_ASAP7_75t_L   g10111(.A1(new_n9906), .A2(new_n10040), .B(new_n10049), .C(new_n10367), .Y(new_n10368));
  A2O1A1O1Ixp25_ASAP7_75t_L g10112(.A1(new_n9717), .A2(new_n9711), .B(new_n9719), .C(new_n10054), .D(new_n10040), .Y(new_n10369));
  AOI211xp5_ASAP7_75t_L     g10113(.A1(new_n10362), .A2(new_n10366), .B(new_n10044), .C(new_n10369), .Y(new_n10370));
  NOR3xp33_ASAP7_75t_L      g10114(.A(new_n10368), .B(new_n10370), .C(new_n10242), .Y(new_n10371));
  NAND2xp33_ASAP7_75t_L     g10115(.A(new_n10241), .B(new_n10240), .Y(new_n10372));
  OAI211xp5_ASAP7_75t_L     g10116(.A1(new_n10044), .A2(new_n10369), .B(new_n10362), .C(new_n10366), .Y(new_n10373));
  A2O1A1O1Ixp25_ASAP7_75t_L g10117(.A1(new_n9722), .A2(new_n10047), .B(new_n9905), .C(new_n10048), .D(new_n10044), .Y(new_n10374));
  NAND2xp33_ASAP7_75t_L     g10118(.A(new_n10367), .B(new_n10374), .Y(new_n10375));
  AOI21xp33_ASAP7_75t_L     g10119(.A1(new_n10375), .A2(new_n10373), .B(new_n10372), .Y(new_n10376));
  NOR2xp33_ASAP7_75t_L      g10120(.A(new_n10376), .B(new_n10371), .Y(new_n10377));
  A2O1A1Ixp33_ASAP7_75t_L   g10121(.A1(new_n10052), .A2(new_n9901), .B(new_n10066), .C(new_n10377), .Y(new_n10378));
  O2A1O1Ixp33_ASAP7_75t_L   g10122(.A1(new_n10063), .A2(new_n9731), .B(new_n10052), .C(new_n10066), .Y(new_n10379));
  NAND3xp33_ASAP7_75t_L     g10123(.A(new_n10375), .B(new_n10373), .C(new_n10372), .Y(new_n10380));
  OAI21xp33_ASAP7_75t_L     g10124(.A1(new_n10370), .A2(new_n10368), .B(new_n10242), .Y(new_n10381));
  NAND2xp33_ASAP7_75t_L     g10125(.A(new_n10380), .B(new_n10381), .Y(new_n10382));
  NAND2xp33_ASAP7_75t_L     g10126(.A(new_n10379), .B(new_n10382), .Y(new_n10383));
  NAND2xp33_ASAP7_75t_L     g10127(.A(\b[31] ), .B(new_n2386), .Y(new_n10384));
  NAND2xp33_ASAP7_75t_L     g10128(.A(\b[32] ), .B(new_n2232), .Y(new_n10385));
  AOI22xp33_ASAP7_75t_L     g10129(.A1(new_n2228), .A2(\b[33] ), .B1(new_n2226), .B2(new_n3813), .Y(new_n10386));
  NAND4xp25_ASAP7_75t_L     g10130(.A(new_n10386), .B(\a[26] ), .C(new_n10384), .D(new_n10385), .Y(new_n10387));
  NAND2xp33_ASAP7_75t_L     g10131(.A(new_n10385), .B(new_n10386), .Y(new_n10388));
  A2O1A1Ixp33_ASAP7_75t_L   g10132(.A1(\b[31] ), .A2(new_n2386), .B(new_n10388), .C(new_n2223), .Y(new_n10389));
  NAND2xp33_ASAP7_75t_L     g10133(.A(new_n10387), .B(new_n10389), .Y(new_n10390));
  INVx1_ASAP7_75t_L         g10134(.A(new_n10390), .Y(new_n10391));
  NAND3xp33_ASAP7_75t_L     g10135(.A(new_n10378), .B(new_n10383), .C(new_n10391), .Y(new_n10392));
  INVx1_ASAP7_75t_L         g10136(.A(new_n9901), .Y(new_n10393));
  O2A1O1Ixp33_ASAP7_75t_L   g10137(.A1(new_n10393), .A2(new_n10065), .B(new_n10058), .C(new_n10382), .Y(new_n10394));
  A2O1A1Ixp33_ASAP7_75t_L   g10138(.A1(new_n9737), .A2(new_n10064), .B(new_n10065), .C(new_n10058), .Y(new_n10395));
  NOR2xp33_ASAP7_75t_L      g10139(.A(new_n10395), .B(new_n10377), .Y(new_n10396));
  OAI21xp33_ASAP7_75t_L     g10140(.A1(new_n10396), .A2(new_n10394), .B(new_n10390), .Y(new_n10397));
  AO21x2_ASAP7_75t_L        g10141(.A1(new_n10397), .A2(new_n10392), .B(new_n10236), .Y(new_n10398));
  NAND3xp33_ASAP7_75t_L     g10142(.A(new_n10236), .B(new_n10392), .C(new_n10397), .Y(new_n10399));
  NAND3xp33_ASAP7_75t_L     g10143(.A(new_n10398), .B(new_n10235), .C(new_n10399), .Y(new_n10400));
  INVx1_ASAP7_75t_L         g10144(.A(new_n10235), .Y(new_n10401));
  AOI21xp33_ASAP7_75t_L     g10145(.A1(new_n10397), .A2(new_n10392), .B(new_n10236), .Y(new_n10402));
  AND3x1_ASAP7_75t_L        g10146(.A(new_n10236), .B(new_n10397), .C(new_n10392), .Y(new_n10403));
  OAI21xp33_ASAP7_75t_L     g10147(.A1(new_n10402), .A2(new_n10403), .B(new_n10401), .Y(new_n10404));
  NAND2xp33_ASAP7_75t_L     g10148(.A(new_n10400), .B(new_n10404), .Y(new_n10405));
  NAND2xp33_ASAP7_75t_L     g10149(.A(new_n10405), .B(new_n10228), .Y(new_n10406));
  OAI211xp5_ASAP7_75t_L     g10150(.A1(new_n10227), .A2(new_n10106), .B(new_n10400), .C(new_n10404), .Y(new_n10407));
  NOR2xp33_ASAP7_75t_L      g10151(.A(new_n4701), .B(new_n1549), .Y(new_n10408));
  INVx1_ASAP7_75t_L         g10152(.A(new_n10408), .Y(new_n10409));
  NAND2xp33_ASAP7_75t_L     g10153(.A(\b[38] ), .B(new_n1410), .Y(new_n10410));
  AOI22xp33_ASAP7_75t_L     g10154(.A1(new_n1406), .A2(\b[39] ), .B1(new_n1404), .B2(new_n5174), .Y(new_n10411));
  AND4x1_ASAP7_75t_L        g10155(.A(new_n10411), .B(new_n10410), .C(new_n10409), .D(\a[20] ), .Y(new_n10412));
  AOI31xp33_ASAP7_75t_L     g10156(.A1(new_n10411), .A2(new_n10410), .A3(new_n10409), .B(\a[20] ), .Y(new_n10413));
  NOR2xp33_ASAP7_75t_L      g10157(.A(new_n10413), .B(new_n10412), .Y(new_n10414));
  NAND3xp33_ASAP7_75t_L     g10158(.A(new_n10407), .B(new_n10406), .C(new_n10414), .Y(new_n10415));
  AOI221xp5_ASAP7_75t_L     g10159(.A1(new_n10095), .A2(new_n10097), .B1(new_n10400), .B2(new_n10404), .C(new_n10227), .Y(new_n10416));
  NOR2xp33_ASAP7_75t_L      g10160(.A(new_n10405), .B(new_n10228), .Y(new_n10417));
  INVx1_ASAP7_75t_L         g10161(.A(new_n10414), .Y(new_n10418));
  OAI21xp33_ASAP7_75t_L     g10162(.A1(new_n10416), .A2(new_n10417), .B(new_n10418), .Y(new_n10419));
  NOR3xp33_ASAP7_75t_L      g10163(.A(new_n10104), .B(new_n10106), .C(new_n10102), .Y(new_n10420));
  O2A1O1Ixp33_ASAP7_75t_L   g10164(.A1(new_n10110), .A2(new_n10111), .B(new_n10113), .C(new_n10420), .Y(new_n10421));
  NAND3xp33_ASAP7_75t_L     g10165(.A(new_n10421), .B(new_n10419), .C(new_n10415), .Y(new_n10422));
  NOR2xp33_ASAP7_75t_L      g10166(.A(new_n10106), .B(new_n10104), .Y(new_n10423));
  NAND2xp33_ASAP7_75t_L     g10167(.A(new_n10101), .B(new_n10423), .Y(new_n10424));
  AO22x1_ASAP7_75t_L        g10168(.A1(new_n10415), .A2(new_n10419), .B1(new_n10424), .B2(new_n10114), .Y(new_n10425));
  NOR2xp33_ASAP7_75t_L      g10169(.A(new_n5186), .B(new_n1195), .Y(new_n10426));
  INVx1_ASAP7_75t_L         g10170(.A(new_n10426), .Y(new_n10427));
  NAND2xp33_ASAP7_75t_L     g10171(.A(\b[41] ), .B(new_n1103), .Y(new_n10428));
  AOI22xp33_ASAP7_75t_L     g10172(.A1(new_n1113), .A2(\b[42] ), .B1(new_n1110), .B2(new_n5688), .Y(new_n10429));
  AND4x1_ASAP7_75t_L        g10173(.A(new_n10429), .B(new_n10428), .C(new_n10427), .D(\a[17] ), .Y(new_n10430));
  AOI31xp33_ASAP7_75t_L     g10174(.A1(new_n10429), .A2(new_n10428), .A3(new_n10427), .B(\a[17] ), .Y(new_n10431));
  NOR2xp33_ASAP7_75t_L      g10175(.A(new_n10431), .B(new_n10430), .Y(new_n10432));
  INVx1_ASAP7_75t_L         g10176(.A(new_n10432), .Y(new_n10433));
  AOI21xp33_ASAP7_75t_L     g10177(.A1(new_n10425), .A2(new_n10422), .B(new_n10433), .Y(new_n10434));
  AND4x1_ASAP7_75t_L        g10178(.A(new_n10114), .B(new_n10424), .C(new_n10415), .D(new_n10419), .Y(new_n10435));
  AOI21xp33_ASAP7_75t_L     g10179(.A1(new_n10419), .A2(new_n10415), .B(new_n10421), .Y(new_n10436));
  NOR3xp33_ASAP7_75t_L      g10180(.A(new_n10435), .B(new_n10436), .C(new_n10432), .Y(new_n10437));
  NOR2xp33_ASAP7_75t_L      g10181(.A(new_n10437), .B(new_n10434), .Y(new_n10438));
  NAND2xp33_ASAP7_75t_L     g10182(.A(new_n10438), .B(new_n10226), .Y(new_n10439));
  A2O1A1O1Ixp25_ASAP7_75t_L g10183(.A1(new_n9795), .A2(new_n9793), .B(new_n10127), .C(new_n10130), .D(new_n10224), .Y(new_n10440));
  OAI21xp33_ASAP7_75t_L     g10184(.A1(new_n10436), .A2(new_n10435), .B(new_n10432), .Y(new_n10441));
  NAND3xp33_ASAP7_75t_L     g10185(.A(new_n10425), .B(new_n10422), .C(new_n10433), .Y(new_n10442));
  NAND2xp33_ASAP7_75t_L     g10186(.A(new_n10441), .B(new_n10442), .Y(new_n10443));
  NAND2xp33_ASAP7_75t_L     g10187(.A(new_n10443), .B(new_n10440), .Y(new_n10444));
  AOI21xp33_ASAP7_75t_L     g10188(.A1(new_n10439), .A2(new_n10444), .B(new_n10223), .Y(new_n10445));
  NAND2xp33_ASAP7_75t_L     g10189(.A(new_n10222), .B(new_n10221), .Y(new_n10446));
  A2O1A1O1Ixp25_ASAP7_75t_L g10190(.A1(new_n9478), .A2(new_n9477), .B(new_n9889), .C(new_n9793), .D(new_n10127), .Y(new_n10447));
  O2A1O1Ixp33_ASAP7_75t_L   g10191(.A1(new_n10145), .A2(new_n10447), .B(new_n10225), .C(new_n10443), .Y(new_n10448));
  AOI221xp5_ASAP7_75t_L     g10192(.A1(new_n10442), .A2(new_n10441), .B1(new_n10130), .B2(new_n10141), .C(new_n10224), .Y(new_n10449));
  NOR3xp33_ASAP7_75t_L      g10193(.A(new_n10448), .B(new_n10449), .C(new_n10446), .Y(new_n10450));
  O2A1O1Ixp33_ASAP7_75t_L   g10194(.A1(new_n9564), .A2(new_n9810), .B(new_n9807), .C(new_n10139), .Y(new_n10451));
  OA22x2_ASAP7_75t_L        g10195(.A1(new_n10445), .A2(new_n10450), .B1(new_n10148), .B2(new_n10451), .Y(new_n10452));
  NOR4xp25_ASAP7_75t_L      g10196(.A(new_n10451), .B(new_n10445), .C(new_n10450), .D(new_n10148), .Y(new_n10453));
  OAI21xp33_ASAP7_75t_L     g10197(.A1(new_n10453), .A2(new_n10452), .B(new_n10217), .Y(new_n10454));
  OAI22xp33_ASAP7_75t_L     g10198(.A1(new_n10450), .A2(new_n10445), .B1(new_n10148), .B2(new_n10451), .Y(new_n10455));
  OAI21xp33_ASAP7_75t_L     g10199(.A1(new_n10449), .A2(new_n10448), .B(new_n10446), .Y(new_n10456));
  NAND3xp33_ASAP7_75t_L     g10200(.A(new_n10439), .B(new_n10444), .C(new_n10223), .Y(new_n10457));
  A2O1A1Ixp33_ASAP7_75t_L   g10201(.A1(new_n9809), .A2(new_n9806), .B(new_n9811), .C(new_n10151), .Y(new_n10458));
  NAND4xp25_ASAP7_75t_L     g10202(.A(new_n10458), .B(new_n10152), .C(new_n10456), .D(new_n10457), .Y(new_n10459));
  NAND3xp33_ASAP7_75t_L     g10203(.A(new_n10459), .B(new_n10455), .C(new_n10216), .Y(new_n10460));
  AOI21xp33_ASAP7_75t_L     g10204(.A1(new_n10460), .A2(new_n10454), .B(new_n10210), .Y(new_n10461));
  OAI21xp33_ASAP7_75t_L     g10205(.A1(new_n10160), .A2(new_n10159), .B(new_n10156), .Y(new_n10462));
  NAND2xp33_ASAP7_75t_L     g10206(.A(new_n10460), .B(new_n10454), .Y(new_n10463));
  NOR2xp33_ASAP7_75t_L      g10207(.A(new_n10463), .B(new_n10462), .Y(new_n10464));
  OAI21xp33_ASAP7_75t_L     g10208(.A1(new_n10461), .A2(new_n10464), .B(new_n10209), .Y(new_n10465));
  NAND2xp33_ASAP7_75t_L     g10209(.A(new_n10463), .B(new_n10462), .Y(new_n10466));
  NAND3xp33_ASAP7_75t_L     g10210(.A(new_n10210), .B(new_n10454), .C(new_n10460), .Y(new_n10467));
  NAND3xp33_ASAP7_75t_L     g10211(.A(new_n10466), .B(new_n10208), .C(new_n10467), .Y(new_n10468));
  NAND2xp33_ASAP7_75t_L     g10212(.A(new_n10468), .B(new_n10465), .Y(new_n10469));
  NAND2xp33_ASAP7_75t_L     g10213(.A(new_n10201), .B(new_n10469), .Y(new_n10470));
  MAJx2_ASAP7_75t_L         g10214(.A(new_n9871), .B(new_n9878), .C(new_n10200), .Y(new_n10471));
  AOI21xp33_ASAP7_75t_L     g10215(.A1(new_n10466), .A2(new_n10467), .B(new_n10208), .Y(new_n10472));
  NOR3xp33_ASAP7_75t_L      g10216(.A(new_n10464), .B(new_n10209), .C(new_n10461), .Y(new_n10473));
  NOR2xp33_ASAP7_75t_L      g10217(.A(new_n10472), .B(new_n10473), .Y(new_n10474));
  NAND2xp33_ASAP7_75t_L     g10218(.A(new_n10474), .B(new_n10471), .Y(new_n10475));
  AOI21xp33_ASAP7_75t_L     g10219(.A1(new_n10475), .A2(new_n10470), .B(new_n10199), .Y(new_n10476));
  INVx1_ASAP7_75t_L         g10220(.A(new_n10199), .Y(new_n10477));
  OA21x2_ASAP7_75t_L        g10221(.A1(new_n10472), .A2(new_n10473), .B(new_n10201), .Y(new_n10478));
  NOR2xp33_ASAP7_75t_L      g10222(.A(new_n10201), .B(new_n10469), .Y(new_n10479));
  NOR3xp33_ASAP7_75t_L      g10223(.A(new_n10478), .B(new_n10479), .C(new_n10477), .Y(new_n10480));
  NOR2xp33_ASAP7_75t_L      g10224(.A(new_n10476), .B(new_n10480), .Y(new_n10481));
  A2O1A1Ixp33_ASAP7_75t_L   g10225(.A1(new_n10167), .A2(new_n9864), .B(new_n10174), .C(new_n10481), .Y(new_n10482));
  NAND2xp33_ASAP7_75t_L     g10226(.A(new_n9849), .B(new_n9845), .Y(new_n10483));
  A2O1A1O1Ixp25_ASAP7_75t_L g10227(.A1(new_n9851), .A2(new_n10483), .B(new_n9862), .C(new_n10167), .D(new_n10174), .Y(new_n10484));
  OAI21xp33_ASAP7_75t_L     g10228(.A1(new_n10476), .A2(new_n10480), .B(new_n10484), .Y(new_n10485));
  INVx1_ASAP7_75t_L         g10229(.A(new_n10179), .Y(new_n10486));
  NOR2xp33_ASAP7_75t_L      g10230(.A(\b[56] ), .B(\b[57] ), .Y(new_n10487));
  INVx1_ASAP7_75t_L         g10231(.A(\b[57] ), .Y(new_n10488));
  NOR2xp33_ASAP7_75t_L      g10232(.A(new_n10178), .B(new_n10488), .Y(new_n10489));
  NOR2xp33_ASAP7_75t_L      g10233(.A(new_n10487), .B(new_n10489), .Y(new_n10490));
  INVx1_ASAP7_75t_L         g10234(.A(new_n10490), .Y(new_n10491));
  O2A1O1Ixp33_ASAP7_75t_L   g10235(.A1(new_n10177), .A2(new_n10182), .B(new_n10486), .C(new_n10491), .Y(new_n10492));
  A2O1A1O1Ixp25_ASAP7_75t_L g10236(.A1(new_n9536), .A2(new_n9540), .B(new_n9535), .C(new_n10180), .D(new_n10179), .Y(new_n10493));
  AND2x2_ASAP7_75t_L        g10237(.A(new_n10491), .B(new_n10493), .Y(new_n10494));
  NOR2xp33_ASAP7_75t_L      g10238(.A(new_n10492), .B(new_n10494), .Y(new_n10495));
  NOR2xp33_ASAP7_75t_L      g10239(.A(new_n10488), .B(new_n632), .Y(new_n10496));
  AOI221xp5_ASAP7_75t_L     g10240(.A1(new_n380), .A2(\b[56] ), .B1(new_n269), .B2(new_n10495), .C(new_n10496), .Y(new_n10497));
  OA211x2_ASAP7_75t_L       g10241(.A1(new_n277), .A2(new_n9534), .B(new_n10497), .C(\a[2] ), .Y(new_n10498));
  O2A1O1Ixp33_ASAP7_75t_L   g10242(.A1(new_n9534), .A2(new_n277), .B(new_n10497), .C(\a[2] ), .Y(new_n10499));
  NOR2xp33_ASAP7_75t_L      g10243(.A(new_n10499), .B(new_n10498), .Y(new_n10500));
  AOI21xp33_ASAP7_75t_L     g10244(.A1(new_n10482), .A2(new_n10485), .B(new_n10500), .Y(new_n10501));
  INVx1_ASAP7_75t_L         g10245(.A(new_n10501), .Y(new_n10502));
  NAND3xp33_ASAP7_75t_L     g10246(.A(new_n10482), .B(new_n10500), .C(new_n10485), .Y(new_n10503));
  NAND2xp33_ASAP7_75t_L     g10247(.A(new_n10503), .B(new_n10502), .Y(new_n10504));
  XNOR2x2_ASAP7_75t_L       g10248(.A(new_n10192), .B(new_n10504), .Y(\f[57] ));
  OAI21xp33_ASAP7_75t_L     g10249(.A1(new_n10479), .A2(new_n10478), .B(new_n10477), .Y(new_n10506));
  NAND3xp33_ASAP7_75t_L     g10250(.A(new_n10475), .B(new_n10470), .C(new_n10199), .Y(new_n10507));
  NAND3xp33_ASAP7_75t_L     g10251(.A(new_n10475), .B(new_n10470), .C(new_n10477), .Y(new_n10508));
  A2O1A1Ixp33_ASAP7_75t_L   g10252(.A1(new_n10506), .A2(new_n10507), .B(new_n10484), .C(new_n10508), .Y(new_n10509));
  NAND2xp33_ASAP7_75t_L     g10253(.A(\b[54] ), .B(new_n334), .Y(new_n10510));
  AOI22xp33_ASAP7_75t_L     g10254(.A1(new_n345), .A2(\b[55] ), .B1(new_n342), .B2(new_n9542), .Y(new_n10511));
  NAND2xp33_ASAP7_75t_L     g10255(.A(new_n10510), .B(new_n10511), .Y(new_n10512));
  AOI211xp5_ASAP7_75t_L     g10256(.A1(\b[53] ), .A2(new_n366), .B(new_n339), .C(new_n10512), .Y(new_n10513));
  INVx1_ASAP7_75t_L         g10257(.A(new_n10512), .Y(new_n10514));
  O2A1O1Ixp33_ASAP7_75t_L   g10258(.A1(new_n8882), .A2(new_n365), .B(new_n10514), .C(\a[5] ), .Y(new_n10515));
  NOR2xp33_ASAP7_75t_L      g10259(.A(new_n10513), .B(new_n10515), .Y(new_n10516));
  NOR2xp33_ASAP7_75t_L      g10260(.A(new_n10461), .B(new_n10464), .Y(new_n10517));
  MAJIxp5_ASAP7_75t_L       g10261(.A(new_n10201), .B(new_n10209), .C(new_n10517), .Y(new_n10518));
  INVx1_ASAP7_75t_L         g10262(.A(new_n8577), .Y(new_n10519));
  NAND2xp33_ASAP7_75t_L     g10263(.A(\b[51] ), .B(new_n441), .Y(new_n10520));
  OAI221xp5_ASAP7_75t_L     g10264(.A1(new_n667), .A2(new_n8569), .B1(new_n482), .B2(new_n10519), .C(new_n10520), .Y(new_n10521));
  AOI21xp33_ASAP7_75t_L     g10265(.A1(new_n480), .A2(\b[50] ), .B(new_n10521), .Y(new_n10522));
  NAND2xp33_ASAP7_75t_L     g10266(.A(\a[8] ), .B(new_n10522), .Y(new_n10523));
  A2O1A1Ixp33_ASAP7_75t_L   g10267(.A1(\b[50] ), .A2(new_n480), .B(new_n10521), .C(new_n445), .Y(new_n10524));
  NAND2xp33_ASAP7_75t_L     g10268(.A(new_n10524), .B(new_n10523), .Y(new_n10525));
  NAND2xp33_ASAP7_75t_L     g10269(.A(new_n10455), .B(new_n10459), .Y(new_n10526));
  MAJIxp5_ASAP7_75t_L       g10270(.A(new_n10210), .B(new_n10216), .C(new_n10526), .Y(new_n10527));
  NAND2xp33_ASAP7_75t_L     g10271(.A(\b[47] ), .B(new_n674), .Y(new_n10528));
  NAND2xp33_ASAP7_75t_L     g10272(.A(\b[48] ), .B(new_n590), .Y(new_n10529));
  AOI22xp33_ASAP7_75t_L     g10273(.A1(new_n600), .A2(\b[49] ), .B1(new_n597), .B2(new_n7914), .Y(new_n10530));
  NAND4xp25_ASAP7_75t_L     g10274(.A(new_n10530), .B(\a[11] ), .C(new_n10528), .D(new_n10529), .Y(new_n10531));
  AOI31xp33_ASAP7_75t_L     g10275(.A1(new_n10530), .A2(new_n10529), .A3(new_n10528), .B(\a[11] ), .Y(new_n10532));
  INVx1_ASAP7_75t_L         g10276(.A(new_n10532), .Y(new_n10533));
  NAND2xp33_ASAP7_75t_L     g10277(.A(new_n10531), .B(new_n10533), .Y(new_n10534));
  INVx1_ASAP7_75t_L         g10278(.A(new_n10534), .Y(new_n10535));
  NOR3xp33_ASAP7_75t_L      g10279(.A(new_n10448), .B(new_n10223), .C(new_n10449), .Y(new_n10536));
  INVx1_ASAP7_75t_L         g10280(.A(new_n10536), .Y(new_n10537));
  NAND2xp33_ASAP7_75t_L     g10281(.A(\b[46] ), .B(new_n826), .Y(new_n10538));
  OAI221xp5_ASAP7_75t_L     g10282(.A1(new_n6756), .A2(new_n994), .B1(new_n911), .B2(new_n7887), .C(new_n10538), .Y(new_n10539));
  AOI21xp33_ASAP7_75t_L     g10283(.A1(new_n908), .A2(\b[44] ), .B(new_n10539), .Y(new_n10540));
  NAND2xp33_ASAP7_75t_L     g10284(.A(\a[14] ), .B(new_n10540), .Y(new_n10541));
  A2O1A1Ixp33_ASAP7_75t_L   g10285(.A1(\b[44] ), .A2(new_n908), .B(new_n10539), .C(new_n813), .Y(new_n10542));
  NAND2xp33_ASAP7_75t_L     g10286(.A(new_n10542), .B(new_n10541), .Y(new_n10543));
  A2O1A1Ixp33_ASAP7_75t_L   g10287(.A1(new_n10131), .A2(new_n10225), .B(new_n10434), .C(new_n10442), .Y(new_n10544));
  A2O1A1O1Ixp25_ASAP7_75t_L g10288(.A1(new_n10052), .A2(new_n9901), .B(new_n10066), .C(new_n10381), .D(new_n10371), .Y(new_n10545));
  A2O1A1Ixp33_ASAP7_75t_L   g10289(.A1(new_n10047), .A2(new_n9722), .B(new_n9905), .C(new_n10048), .Y(new_n10546));
  A2O1A1Ixp33_ASAP7_75t_L   g10290(.A1(new_n10049), .A2(new_n10546), .B(new_n10367), .C(new_n10366), .Y(new_n10547));
  O2A1O1Ixp33_ASAP7_75t_L   g10291(.A1(new_n10014), .A2(new_n10021), .B(new_n10340), .C(new_n10342), .Y(new_n10548));
  AOI22xp33_ASAP7_75t_L     g10292(.A1(new_n4544), .A2(\b[22] ), .B1(new_n4542), .B2(new_n1864), .Y(new_n10549));
  OAI221xp5_ASAP7_75t_L     g10293(.A1(new_n4536), .A2(new_n1709), .B1(new_n1594), .B2(new_n4781), .C(new_n10549), .Y(new_n10550));
  XNOR2x2_ASAP7_75t_L       g10294(.A(new_n4539), .B(new_n10550), .Y(new_n10551));
  INVx1_ASAP7_75t_L         g10295(.A(new_n10253), .Y(new_n10552));
  NAND3xp33_ASAP7_75t_L     g10296(.A(new_n10552), .B(new_n10321), .C(new_n10327), .Y(new_n10553));
  A2O1A1Ixp33_ASAP7_75t_L   g10297(.A1(new_n10328), .A2(new_n10329), .B(new_n10250), .C(new_n10553), .Y(new_n10554));
  A2O1A1Ixp33_ASAP7_75t_L   g10298(.A1(new_n9994), .A2(new_n10254), .B(new_n10326), .C(new_n10319), .Y(new_n10555));
  NAND2xp33_ASAP7_75t_L     g10299(.A(\b[14] ), .B(new_n6308), .Y(new_n10556));
  NAND2xp33_ASAP7_75t_L     g10300(.A(\b[15] ), .B(new_n5992), .Y(new_n10557));
  AOI22xp33_ASAP7_75t_L     g10301(.A1(new_n6002), .A2(\b[16] ), .B1(new_n5999), .B2(new_n1058), .Y(new_n10558));
  NAND4xp25_ASAP7_75t_L     g10302(.A(new_n10558), .B(\a[44] ), .C(new_n10556), .D(new_n10557), .Y(new_n10559));
  NAND2xp33_ASAP7_75t_L     g10303(.A(new_n10557), .B(new_n10558), .Y(new_n10560));
  A2O1A1Ixp33_ASAP7_75t_L   g10304(.A1(\b[14] ), .A2(new_n6308), .B(new_n10560), .C(new_n5996), .Y(new_n10561));
  AND2x2_ASAP7_75t_L        g10305(.A(new_n10559), .B(new_n10561), .Y(new_n10562));
  OAI211xp5_ASAP7_75t_L     g10306(.A1(new_n10314), .A2(new_n10315), .B(new_n10267), .C(new_n10265), .Y(new_n10563));
  A2O1A1O1Ixp25_ASAP7_75t_L g10307(.A1(new_n9973), .A2(new_n9925), .B(new_n10260), .C(new_n10563), .D(new_n10316), .Y(new_n10564));
  NAND2xp33_ASAP7_75t_L     g10308(.A(new_n10287), .B(new_n10286), .Y(new_n10565));
  AO21x2_ASAP7_75t_L        g10309(.A1(new_n10292), .A2(new_n10290), .B(new_n10565), .Y(new_n10566));
  OAI22xp33_ASAP7_75t_L     g10310(.A1(new_n10296), .A2(new_n9964), .B1(new_n10293), .B2(new_n10294), .Y(new_n10567));
  OAI22xp33_ASAP7_75t_L     g10311(.A1(new_n427), .A2(new_n8967), .B1(new_n8968), .B2(new_n421), .Y(new_n10568));
  AOI221xp5_ASAP7_75t_L     g10312(.A1(\b[5] ), .A2(new_n8964), .B1(\b[6] ), .B2(new_n8635), .C(new_n10568), .Y(new_n10569));
  NAND2xp33_ASAP7_75t_L     g10313(.A(\a[53] ), .B(new_n10569), .Y(new_n10570));
  INVx1_ASAP7_75t_L         g10314(.A(new_n10570), .Y(new_n10571));
  NOR2xp33_ASAP7_75t_L      g10315(.A(\a[53] ), .B(new_n10569), .Y(new_n10572));
  AOI22xp33_ASAP7_75t_L     g10316(.A1(new_n10284), .A2(new_n10285), .B1(new_n10279), .B2(new_n10277), .Y(new_n10573));
  NOR3xp33_ASAP7_75t_L      g10317(.A(new_n10270), .B(new_n10271), .C(new_n10278), .Y(new_n10574));
  NAND2xp33_ASAP7_75t_L     g10318(.A(\b[2] ), .B(new_n9948), .Y(new_n10575));
  NAND2xp33_ASAP7_75t_L     g10319(.A(\b[3] ), .B(new_n9614), .Y(new_n10576));
  AOI22xp33_ASAP7_75t_L     g10320(.A1(new_n9623), .A2(\b[4] ), .B1(new_n9620), .B2(new_n328), .Y(new_n10577));
  NAND4xp25_ASAP7_75t_L     g10321(.A(new_n10577), .B(\a[56] ), .C(new_n10575), .D(new_n10576), .Y(new_n10578));
  NAND2xp33_ASAP7_75t_L     g10322(.A(new_n10576), .B(new_n10577), .Y(new_n10579));
  A2O1A1Ixp33_ASAP7_75t_L   g10323(.A1(\b[2] ), .A2(new_n9948), .B(new_n10579), .C(new_n9610), .Y(new_n10580));
  NAND2xp33_ASAP7_75t_L     g10324(.A(\a[59] ), .B(new_n10276), .Y(new_n10581));
  NAND2xp33_ASAP7_75t_L     g10325(.A(new_n10274), .B(new_n10273), .Y(new_n10582));
  XNOR2x2_ASAP7_75t_L       g10326(.A(\a[58] ), .B(\a[57] ), .Y(new_n10583));
  NOR2xp33_ASAP7_75t_L      g10327(.A(new_n10583), .B(new_n10582), .Y(new_n10584));
  NAND2xp33_ASAP7_75t_L     g10328(.A(\b[0] ), .B(new_n10584), .Y(new_n10585));
  INVx1_ASAP7_75t_L         g10329(.A(\a[58] ), .Y(new_n10586));
  NAND2xp33_ASAP7_75t_L     g10330(.A(\a[59] ), .B(new_n10586), .Y(new_n10587));
  INVx1_ASAP7_75t_L         g10331(.A(\a[59] ), .Y(new_n10588));
  NAND2xp33_ASAP7_75t_L     g10332(.A(\a[58] ), .B(new_n10588), .Y(new_n10589));
  AND2x2_ASAP7_75t_L        g10333(.A(new_n10587), .B(new_n10589), .Y(new_n10590));
  NOR2xp33_ASAP7_75t_L      g10334(.A(new_n10275), .B(new_n10590), .Y(new_n10591));
  NAND2xp33_ASAP7_75t_L     g10335(.A(new_n271), .B(new_n10591), .Y(new_n10592));
  NAND2xp33_ASAP7_75t_L     g10336(.A(new_n10589), .B(new_n10587), .Y(new_n10593));
  NOR2xp33_ASAP7_75t_L      g10337(.A(new_n10593), .B(new_n10275), .Y(new_n10594));
  NAND2xp33_ASAP7_75t_L     g10338(.A(\b[1] ), .B(new_n10594), .Y(new_n10595));
  AND3x1_ASAP7_75t_L        g10339(.A(new_n10592), .B(new_n10595), .C(new_n10585), .Y(new_n10596));
  XNOR2x2_ASAP7_75t_L       g10340(.A(new_n10581), .B(new_n10596), .Y(new_n10597));
  NAND3xp33_ASAP7_75t_L     g10341(.A(new_n10580), .B(new_n10578), .C(new_n10597), .Y(new_n10598));
  AO21x2_ASAP7_75t_L        g10342(.A1(new_n10578), .A2(new_n10580), .B(new_n10597), .Y(new_n10599));
  OAI211xp5_ASAP7_75t_L     g10343(.A1(new_n10574), .A2(new_n10573), .B(new_n10598), .C(new_n10599), .Y(new_n10600));
  INVx1_ASAP7_75t_L         g10344(.A(new_n10574), .Y(new_n10601));
  INVx1_ASAP7_75t_L         g10345(.A(new_n10598), .Y(new_n10602));
  AOI21xp33_ASAP7_75t_L     g10346(.A1(new_n10580), .A2(new_n10578), .B(new_n10597), .Y(new_n10603));
  OAI211xp5_ASAP7_75t_L     g10347(.A1(new_n10603), .A2(new_n10602), .B(new_n10601), .C(new_n10286), .Y(new_n10604));
  AOI211xp5_ASAP7_75t_L     g10348(.A1(new_n10604), .A2(new_n10600), .B(new_n10571), .C(new_n10572), .Y(new_n10605));
  INVx1_ASAP7_75t_L         g10349(.A(new_n10572), .Y(new_n10606));
  INVx1_ASAP7_75t_L         g10350(.A(new_n10600), .Y(new_n10607));
  AOI211xp5_ASAP7_75t_L     g10351(.A1(new_n10599), .A2(new_n10598), .B(new_n10573), .C(new_n10574), .Y(new_n10608));
  AOI211xp5_ASAP7_75t_L     g10352(.A1(new_n10606), .A2(new_n10570), .B(new_n10607), .C(new_n10608), .Y(new_n10609));
  AOI211xp5_ASAP7_75t_L     g10353(.A1(new_n10567), .A2(new_n10566), .B(new_n10605), .C(new_n10609), .Y(new_n10610));
  AND2x2_ASAP7_75t_L        g10354(.A(new_n10290), .B(new_n10292), .Y(new_n10611));
  MAJIxp5_ASAP7_75t_L       g10355(.A(new_n10298), .B(new_n10565), .C(new_n10611), .Y(new_n10612));
  OAI211xp5_ASAP7_75t_L     g10356(.A1(new_n10608), .A2(new_n10607), .B(new_n10606), .C(new_n10570), .Y(new_n10613));
  OAI211xp5_ASAP7_75t_L     g10357(.A1(new_n10572), .A2(new_n10571), .B(new_n10600), .C(new_n10604), .Y(new_n10614));
  AOI21xp33_ASAP7_75t_L     g10358(.A1(new_n10613), .A2(new_n10614), .B(new_n10612), .Y(new_n10615));
  NAND2xp33_ASAP7_75t_L     g10359(.A(\b[8] ), .B(new_n7993), .Y(new_n10616));
  NAND2xp33_ASAP7_75t_L     g10360(.A(\b[9] ), .B(new_n7649), .Y(new_n10617));
  AOI22xp33_ASAP7_75t_L     g10361(.A1(new_n7659), .A2(\b[10] ), .B1(new_n7656), .B2(new_n852), .Y(new_n10618));
  NAND4xp25_ASAP7_75t_L     g10362(.A(new_n10618), .B(\a[50] ), .C(new_n10616), .D(new_n10617), .Y(new_n10619));
  NAND2xp33_ASAP7_75t_L     g10363(.A(new_n10617), .B(new_n10618), .Y(new_n10620));
  A2O1A1Ixp33_ASAP7_75t_L   g10364(.A1(\b[8] ), .A2(new_n7993), .B(new_n10620), .C(new_n7653), .Y(new_n10621));
  NAND2xp33_ASAP7_75t_L     g10365(.A(new_n10619), .B(new_n10621), .Y(new_n10622));
  NOR3xp33_ASAP7_75t_L      g10366(.A(new_n10622), .B(new_n10610), .C(new_n10615), .Y(new_n10623));
  NAND3xp33_ASAP7_75t_L     g10367(.A(new_n10613), .B(new_n10612), .C(new_n10614), .Y(new_n10624));
  OAI211xp5_ASAP7_75t_L     g10368(.A1(new_n10605), .A2(new_n10609), .B(new_n10567), .C(new_n10566), .Y(new_n10625));
  AND2x2_ASAP7_75t_L        g10369(.A(new_n10619), .B(new_n10621), .Y(new_n10626));
  AOI21xp33_ASAP7_75t_L     g10370(.A1(new_n10625), .A2(new_n10624), .B(new_n10626), .Y(new_n10627));
  OAI21xp33_ASAP7_75t_L     g10371(.A1(new_n10311), .A2(new_n10309), .B(new_n10306), .Y(new_n10628));
  NOR3xp33_ASAP7_75t_L      g10372(.A(new_n10628), .B(new_n10627), .C(new_n10623), .Y(new_n10629));
  NAND4xp25_ASAP7_75t_L     g10373(.A(new_n10625), .B(new_n10624), .C(new_n10619), .D(new_n10621), .Y(new_n10630));
  OAI21xp33_ASAP7_75t_L     g10374(.A1(new_n10615), .A2(new_n10610), .B(new_n10622), .Y(new_n10631));
  A2O1A1O1Ixp25_ASAP7_75t_L g10375(.A1(new_n9970), .A2(new_n9969), .B(new_n9967), .C(new_n10307), .D(new_n10310), .Y(new_n10632));
  AOI21xp33_ASAP7_75t_L     g10376(.A1(new_n10631), .A2(new_n10630), .B(new_n10632), .Y(new_n10633));
  NAND2xp33_ASAP7_75t_L     g10377(.A(\b[12] ), .B(new_n6812), .Y(new_n10634));
  NOR2xp33_ASAP7_75t_L      g10378(.A(new_n793), .B(new_n7118), .Y(new_n10635));
  AOI21xp33_ASAP7_75t_L     g10379(.A1(new_n800), .A2(new_n6819), .B(new_n10635), .Y(new_n10636));
  NAND2xp33_ASAP7_75t_L     g10380(.A(new_n10634), .B(new_n10636), .Y(new_n10637));
  AOI211xp5_ASAP7_75t_L     g10381(.A1(\b[11] ), .A2(new_n7124), .B(new_n6816), .C(new_n10637), .Y(new_n10638));
  AND2x2_ASAP7_75t_L        g10382(.A(new_n10634), .B(new_n10636), .Y(new_n10639));
  O2A1O1Ixp33_ASAP7_75t_L   g10383(.A1(new_n695), .A2(new_n7115), .B(new_n10639), .C(\a[47] ), .Y(new_n10640));
  NOR2xp33_ASAP7_75t_L      g10384(.A(new_n10638), .B(new_n10640), .Y(new_n10641));
  OAI21xp33_ASAP7_75t_L     g10385(.A1(new_n10629), .A2(new_n10633), .B(new_n10641), .Y(new_n10642));
  NAND3xp33_ASAP7_75t_L     g10386(.A(new_n10632), .B(new_n10631), .C(new_n10630), .Y(new_n10643));
  OAI21xp33_ASAP7_75t_L     g10387(.A1(new_n10623), .A2(new_n10627), .B(new_n10628), .Y(new_n10644));
  NAND2xp33_ASAP7_75t_L     g10388(.A(\b[11] ), .B(new_n7124), .Y(new_n10645));
  NAND3xp33_ASAP7_75t_L     g10389(.A(new_n10639), .B(new_n10645), .C(\a[47] ), .Y(new_n10646));
  A2O1A1Ixp33_ASAP7_75t_L   g10390(.A1(\b[11] ), .A2(new_n7124), .B(new_n10637), .C(new_n6816), .Y(new_n10647));
  NAND2xp33_ASAP7_75t_L     g10391(.A(new_n10647), .B(new_n10646), .Y(new_n10648));
  NAND3xp33_ASAP7_75t_L     g10392(.A(new_n10648), .B(new_n10643), .C(new_n10644), .Y(new_n10649));
  NAND3xp33_ASAP7_75t_L     g10393(.A(new_n10564), .B(new_n10642), .C(new_n10649), .Y(new_n10650));
  NAND3xp33_ASAP7_75t_L     g10394(.A(new_n10268), .B(new_n10308), .C(new_n10312), .Y(new_n10651));
  OAI21xp33_ASAP7_75t_L     g10395(.A1(new_n10313), .A2(new_n10261), .B(new_n10651), .Y(new_n10652));
  NAND2xp33_ASAP7_75t_L     g10396(.A(new_n10649), .B(new_n10642), .Y(new_n10653));
  NAND2xp33_ASAP7_75t_L     g10397(.A(new_n10652), .B(new_n10653), .Y(new_n10654));
  AOI21xp33_ASAP7_75t_L     g10398(.A1(new_n10654), .A2(new_n10650), .B(new_n10562), .Y(new_n10655));
  NAND2xp33_ASAP7_75t_L     g10399(.A(new_n10559), .B(new_n10561), .Y(new_n10656));
  NOR2xp33_ASAP7_75t_L      g10400(.A(new_n10652), .B(new_n10653), .Y(new_n10657));
  AOI21xp33_ASAP7_75t_L     g10401(.A1(new_n10649), .A2(new_n10642), .B(new_n10564), .Y(new_n10658));
  NOR3xp33_ASAP7_75t_L      g10402(.A(new_n10657), .B(new_n10658), .C(new_n10656), .Y(new_n10659));
  NOR2xp33_ASAP7_75t_L      g10403(.A(new_n10655), .B(new_n10659), .Y(new_n10660));
  NOR2xp33_ASAP7_75t_L      g10404(.A(new_n10660), .B(new_n10555), .Y(new_n10661));
  NOR2xp33_ASAP7_75t_L      g10405(.A(new_n9990), .B(new_n9991), .Y(new_n10662));
  A2O1A1O1Ixp25_ASAP7_75t_L g10406(.A1(new_n9992), .A2(new_n10662), .B(new_n9998), .C(new_n10320), .D(new_n10325), .Y(new_n10663));
  OAI21xp33_ASAP7_75t_L     g10407(.A1(new_n10658), .A2(new_n10657), .B(new_n10656), .Y(new_n10664));
  NAND3xp33_ASAP7_75t_L     g10408(.A(new_n10654), .B(new_n10650), .C(new_n10562), .Y(new_n10665));
  NAND2xp33_ASAP7_75t_L     g10409(.A(new_n10665), .B(new_n10664), .Y(new_n10666));
  NOR2xp33_ASAP7_75t_L      g10410(.A(new_n10663), .B(new_n10666), .Y(new_n10667));
  AOI22xp33_ASAP7_75t_L     g10411(.A1(new_n5249), .A2(\b[19] ), .B1(new_n5247), .B2(new_n1499), .Y(new_n10668));
  OAI221xp5_ASAP7_75t_L     g10412(.A1(new_n5241), .A2(new_n1356), .B1(new_n1244), .B2(new_n5521), .C(new_n10668), .Y(new_n10669));
  XNOR2x2_ASAP7_75t_L       g10413(.A(\a[41] ), .B(new_n10669), .Y(new_n10670));
  OAI21xp33_ASAP7_75t_L     g10414(.A1(new_n10667), .A2(new_n10661), .B(new_n10670), .Y(new_n10671));
  NAND2xp33_ASAP7_75t_L     g10415(.A(new_n10663), .B(new_n10666), .Y(new_n10672));
  A2O1A1Ixp33_ASAP7_75t_L   g10416(.A1(new_n10320), .A2(new_n10255), .B(new_n10325), .C(new_n10660), .Y(new_n10673));
  XNOR2x2_ASAP7_75t_L       g10417(.A(new_n5244), .B(new_n10669), .Y(new_n10674));
  NAND3xp33_ASAP7_75t_L     g10418(.A(new_n10673), .B(new_n10674), .C(new_n10672), .Y(new_n10675));
  NAND2xp33_ASAP7_75t_L     g10419(.A(new_n10671), .B(new_n10675), .Y(new_n10676));
  NOR2xp33_ASAP7_75t_L      g10420(.A(new_n10554), .B(new_n10676), .Y(new_n10677));
  AOI21xp33_ASAP7_75t_L     g10421(.A1(new_n10673), .A2(new_n10672), .B(new_n10674), .Y(new_n10678));
  NOR3xp33_ASAP7_75t_L      g10422(.A(new_n10661), .B(new_n10667), .C(new_n10670), .Y(new_n10679));
  NOR2xp33_ASAP7_75t_L      g10423(.A(new_n10679), .B(new_n10678), .Y(new_n10680));
  O2A1O1Ixp33_ASAP7_75t_L   g10424(.A1(new_n10250), .A2(new_n10336), .B(new_n10553), .C(new_n10680), .Y(new_n10681));
  OAI21xp33_ASAP7_75t_L     g10425(.A1(new_n10677), .A2(new_n10681), .B(new_n10551), .Y(new_n10682));
  XNOR2x2_ASAP7_75t_L       g10426(.A(\a[38] ), .B(new_n10550), .Y(new_n10683));
  INVx1_ASAP7_75t_L         g10427(.A(new_n10553), .Y(new_n10684));
  O2A1O1Ixp33_ASAP7_75t_L   g10428(.A1(new_n10334), .A2(new_n10335), .B(new_n10338), .C(new_n10684), .Y(new_n10685));
  NAND2xp33_ASAP7_75t_L     g10429(.A(new_n10680), .B(new_n10685), .Y(new_n10686));
  A2O1A1Ixp33_ASAP7_75t_L   g10430(.A1(new_n10330), .A2(new_n10338), .B(new_n10684), .C(new_n10676), .Y(new_n10687));
  NAND3xp33_ASAP7_75t_L     g10431(.A(new_n10686), .B(new_n10687), .C(new_n10683), .Y(new_n10688));
  NAND2xp33_ASAP7_75t_L     g10432(.A(new_n10688), .B(new_n10682), .Y(new_n10689));
  NAND2xp33_ASAP7_75t_L     g10433(.A(new_n10548), .B(new_n10689), .Y(new_n10690));
  AOI21xp33_ASAP7_75t_L     g10434(.A1(new_n10686), .A2(new_n10687), .B(new_n10683), .Y(new_n10691));
  NOR3xp33_ASAP7_75t_L      g10435(.A(new_n10681), .B(new_n10677), .C(new_n10551), .Y(new_n10692));
  NOR2xp33_ASAP7_75t_L      g10436(.A(new_n10691), .B(new_n10692), .Y(new_n10693));
  A2O1A1Ixp33_ASAP7_75t_L   g10437(.A1(new_n10340), .A2(new_n10244), .B(new_n10342), .C(new_n10693), .Y(new_n10694));
  AOI22xp33_ASAP7_75t_L     g10438(.A1(new_n3884), .A2(\b[25] ), .B1(new_n3881), .B2(new_n2188), .Y(new_n10695));
  OAI221xp5_ASAP7_75t_L     g10439(.A1(new_n4312), .A2(new_n2019), .B1(new_n1995), .B2(new_n4986), .C(new_n10695), .Y(new_n10696));
  XNOR2x2_ASAP7_75t_L       g10440(.A(\a[35] ), .B(new_n10696), .Y(new_n10697));
  NAND3xp33_ASAP7_75t_L     g10441(.A(new_n10694), .B(new_n10690), .C(new_n10697), .Y(new_n10698));
  A2O1A1Ixp33_ASAP7_75t_L   g10442(.A1(new_n10022), .A2(new_n10029), .B(new_n10343), .C(new_n10332), .Y(new_n10699));
  NOR2xp33_ASAP7_75t_L      g10443(.A(new_n10699), .B(new_n10693), .Y(new_n10700));
  INVx1_ASAP7_75t_L         g10444(.A(new_n10244), .Y(new_n10701));
  O2A1O1Ixp33_ASAP7_75t_L   g10445(.A1(new_n10701), .A2(new_n10343), .B(new_n10332), .C(new_n10689), .Y(new_n10702));
  XNOR2x2_ASAP7_75t_L       g10446(.A(new_n3878), .B(new_n10696), .Y(new_n10703));
  OAI21xp33_ASAP7_75t_L     g10447(.A1(new_n10700), .A2(new_n10702), .B(new_n10703), .Y(new_n10704));
  NAND3xp33_ASAP7_75t_L     g10448(.A(new_n10344), .B(new_n10341), .C(new_n10351), .Y(new_n10705));
  NAND4xp25_ASAP7_75t_L     g10449(.A(new_n10364), .B(new_n10698), .C(new_n10704), .D(new_n10705), .Y(new_n10706));
  NOR3xp33_ASAP7_75t_L      g10450(.A(new_n10702), .B(new_n10700), .C(new_n10703), .Y(new_n10707));
  AOI21xp33_ASAP7_75t_L     g10451(.A1(new_n10694), .A2(new_n10690), .B(new_n10697), .Y(new_n10708));
  A2O1A1Ixp33_ASAP7_75t_L   g10452(.A1(new_n10348), .A2(new_n10352), .B(new_n10353), .C(new_n10705), .Y(new_n10709));
  OAI21xp33_ASAP7_75t_L     g10453(.A1(new_n10707), .A2(new_n10708), .B(new_n10709), .Y(new_n10710));
  NAND2xp33_ASAP7_75t_L     g10454(.A(\b[26] ), .B(new_n3491), .Y(new_n10711));
  NAND2xp33_ASAP7_75t_L     g10455(.A(\b[27] ), .B(new_n3260), .Y(new_n10712));
  AOI22xp33_ASAP7_75t_L     g10456(.A1(new_n3256), .A2(\b[28] ), .B1(new_n3254), .B2(new_n2858), .Y(new_n10713));
  NAND4xp25_ASAP7_75t_L     g10457(.A(new_n10713), .B(\a[32] ), .C(new_n10711), .D(new_n10712), .Y(new_n10714));
  NAND2xp33_ASAP7_75t_L     g10458(.A(new_n10712), .B(new_n10713), .Y(new_n10715));
  A2O1A1Ixp33_ASAP7_75t_L   g10459(.A1(\b[26] ), .A2(new_n3491), .B(new_n10715), .C(new_n3251), .Y(new_n10716));
  AND2x2_ASAP7_75t_L        g10460(.A(new_n10714), .B(new_n10716), .Y(new_n10717));
  NAND3xp33_ASAP7_75t_L     g10461(.A(new_n10706), .B(new_n10710), .C(new_n10717), .Y(new_n10718));
  NOR3xp33_ASAP7_75t_L      g10462(.A(new_n10709), .B(new_n10708), .C(new_n10707), .Y(new_n10719));
  AOI22xp33_ASAP7_75t_L     g10463(.A1(new_n10698), .A2(new_n10704), .B1(new_n10705), .B2(new_n10364), .Y(new_n10720));
  NAND2xp33_ASAP7_75t_L     g10464(.A(new_n10714), .B(new_n10716), .Y(new_n10721));
  OAI21xp33_ASAP7_75t_L     g10465(.A1(new_n10719), .A2(new_n10720), .B(new_n10721), .Y(new_n10722));
  NAND3xp33_ASAP7_75t_L     g10466(.A(new_n10547), .B(new_n10718), .C(new_n10722), .Y(new_n10723));
  INVx1_ASAP7_75t_L         g10467(.A(new_n10366), .Y(new_n10724));
  O2A1O1Ixp33_ASAP7_75t_L   g10468(.A1(new_n10044), .A2(new_n10369), .B(new_n10362), .C(new_n10724), .Y(new_n10725));
  NAND2xp33_ASAP7_75t_L     g10469(.A(new_n10718), .B(new_n10722), .Y(new_n10726));
  NAND2xp33_ASAP7_75t_L     g10470(.A(new_n10725), .B(new_n10726), .Y(new_n10727));
  NAND2xp33_ASAP7_75t_L     g10471(.A(\b[31] ), .B(new_n2702), .Y(new_n10728));
  OAI221xp5_ASAP7_75t_L     g10472(.A1(new_n3212), .A2(new_n2694), .B1(new_n2707), .B2(new_n4030), .C(new_n10728), .Y(new_n10729));
  AOI21xp33_ASAP7_75t_L     g10473(.A1(new_n2931), .A2(\b[29] ), .B(new_n10729), .Y(new_n10730));
  NAND2xp33_ASAP7_75t_L     g10474(.A(\a[29] ), .B(new_n10730), .Y(new_n10731));
  A2O1A1Ixp33_ASAP7_75t_L   g10475(.A1(\b[29] ), .A2(new_n2931), .B(new_n10729), .C(new_n2697), .Y(new_n10732));
  AND2x2_ASAP7_75t_L        g10476(.A(new_n10732), .B(new_n10731), .Y(new_n10733));
  AOI21xp33_ASAP7_75t_L     g10477(.A1(new_n10723), .A2(new_n10727), .B(new_n10733), .Y(new_n10734));
  O2A1O1Ixp33_ASAP7_75t_L   g10478(.A1(new_n10367), .A2(new_n10374), .B(new_n10366), .C(new_n10726), .Y(new_n10735));
  AOI21xp33_ASAP7_75t_L     g10479(.A1(new_n10722), .A2(new_n10718), .B(new_n10547), .Y(new_n10736));
  INVx1_ASAP7_75t_L         g10480(.A(new_n10733), .Y(new_n10737));
  NOR3xp33_ASAP7_75t_L      g10481(.A(new_n10735), .B(new_n10736), .C(new_n10737), .Y(new_n10738));
  OAI21xp33_ASAP7_75t_L     g10482(.A1(new_n10734), .A2(new_n10738), .B(new_n10545), .Y(new_n10739));
  A2O1A1Ixp33_ASAP7_75t_L   g10483(.A1(new_n10059), .A2(new_n10058), .B(new_n10376), .C(new_n10380), .Y(new_n10740));
  OAI21xp33_ASAP7_75t_L     g10484(.A1(new_n10736), .A2(new_n10735), .B(new_n10737), .Y(new_n10741));
  NAND3xp33_ASAP7_75t_L     g10485(.A(new_n10723), .B(new_n10727), .C(new_n10733), .Y(new_n10742));
  NAND3xp33_ASAP7_75t_L     g10486(.A(new_n10740), .B(new_n10741), .C(new_n10742), .Y(new_n10743));
  NAND2xp33_ASAP7_75t_L     g10487(.A(\b[33] ), .B(new_n2232), .Y(new_n10744));
  AOI22xp33_ASAP7_75t_L     g10488(.A1(new_n2228), .A2(\b[34] ), .B1(new_n2226), .B2(new_n3833), .Y(new_n10745));
  NAND2xp33_ASAP7_75t_L     g10489(.A(new_n10744), .B(new_n10745), .Y(new_n10746));
  AOI21xp33_ASAP7_75t_L     g10490(.A1(new_n2386), .A2(\b[32] ), .B(new_n10746), .Y(new_n10747));
  NAND2xp33_ASAP7_75t_L     g10491(.A(\a[26] ), .B(new_n10747), .Y(new_n10748));
  A2O1A1Ixp33_ASAP7_75t_L   g10492(.A1(\b[32] ), .A2(new_n2386), .B(new_n10746), .C(new_n2223), .Y(new_n10749));
  NAND4xp25_ASAP7_75t_L     g10493(.A(new_n10743), .B(new_n10748), .C(new_n10749), .D(new_n10739), .Y(new_n10750));
  AOI21xp33_ASAP7_75t_L     g10494(.A1(new_n10742), .A2(new_n10741), .B(new_n10740), .Y(new_n10751));
  NOR3xp33_ASAP7_75t_L      g10495(.A(new_n10545), .B(new_n10738), .C(new_n10734), .Y(new_n10752));
  NAND2xp33_ASAP7_75t_L     g10496(.A(new_n10749), .B(new_n10748), .Y(new_n10753));
  OAI21xp33_ASAP7_75t_L     g10497(.A1(new_n10752), .A2(new_n10751), .B(new_n10753), .Y(new_n10754));
  NAND3xp33_ASAP7_75t_L     g10498(.A(new_n10378), .B(new_n10383), .C(new_n10390), .Y(new_n10755));
  NAND4xp25_ASAP7_75t_L     g10499(.A(new_n10398), .B(new_n10755), .C(new_n10754), .D(new_n10750), .Y(new_n10756));
  NAND2xp33_ASAP7_75t_L     g10500(.A(new_n10754), .B(new_n10750), .Y(new_n10757));
  A2O1A1Ixp33_ASAP7_75t_L   g10501(.A1(new_n10392), .A2(new_n10397), .B(new_n10236), .C(new_n10755), .Y(new_n10758));
  NAND2xp33_ASAP7_75t_L     g10502(.A(new_n10758), .B(new_n10757), .Y(new_n10759));
  AOI22xp33_ASAP7_75t_L     g10503(.A1(new_n1766), .A2(\b[37] ), .B1(new_n1764), .B2(new_n4709), .Y(new_n10760));
  OAI221xp5_ASAP7_75t_L     g10504(.A1(new_n1758), .A2(new_n4465), .B1(new_n4053), .B2(new_n1911), .C(new_n10760), .Y(new_n10761));
  XNOR2x2_ASAP7_75t_L       g10505(.A(\a[23] ), .B(new_n10761), .Y(new_n10762));
  NAND3xp33_ASAP7_75t_L     g10506(.A(new_n10759), .B(new_n10756), .C(new_n10762), .Y(new_n10763));
  AO21x2_ASAP7_75t_L        g10507(.A1(new_n10756), .A2(new_n10759), .B(new_n10762), .Y(new_n10764));
  NOR3xp33_ASAP7_75t_L      g10508(.A(new_n10403), .B(new_n10401), .C(new_n10402), .Y(new_n10765));
  A2O1A1O1Ixp25_ASAP7_75t_L g10509(.A1(new_n10097), .A2(new_n10095), .B(new_n10227), .C(new_n10404), .D(new_n10765), .Y(new_n10766));
  NAND3xp33_ASAP7_75t_L     g10510(.A(new_n10766), .B(new_n10764), .C(new_n10763), .Y(new_n10767));
  AO21x2_ASAP7_75t_L        g10511(.A1(new_n10764), .A2(new_n10763), .B(new_n10766), .Y(new_n10768));
  NAND2xp33_ASAP7_75t_L     g10512(.A(\b[38] ), .B(new_n1548), .Y(new_n10769));
  NAND2xp33_ASAP7_75t_L     g10513(.A(\b[39] ), .B(new_n1410), .Y(new_n10770));
  AOI22xp33_ASAP7_75t_L     g10514(.A1(new_n1406), .A2(\b[40] ), .B1(new_n1404), .B2(new_n5194), .Y(new_n10771));
  AND4x1_ASAP7_75t_L        g10515(.A(new_n10771), .B(new_n10770), .C(new_n10769), .D(\a[20] ), .Y(new_n10772));
  AOI31xp33_ASAP7_75t_L     g10516(.A1(new_n10771), .A2(new_n10770), .A3(new_n10769), .B(\a[20] ), .Y(new_n10773));
  NOR2xp33_ASAP7_75t_L      g10517(.A(new_n10773), .B(new_n10772), .Y(new_n10774));
  NAND3xp33_ASAP7_75t_L     g10518(.A(new_n10768), .B(new_n10774), .C(new_n10767), .Y(new_n10775));
  AND3x1_ASAP7_75t_L        g10519(.A(new_n10766), .B(new_n10764), .C(new_n10763), .Y(new_n10776));
  AOI21xp33_ASAP7_75t_L     g10520(.A1(new_n10763), .A2(new_n10764), .B(new_n10766), .Y(new_n10777));
  INVx1_ASAP7_75t_L         g10521(.A(new_n10774), .Y(new_n10778));
  OAI21xp33_ASAP7_75t_L     g10522(.A1(new_n10777), .A2(new_n10776), .B(new_n10778), .Y(new_n10779));
  NAND2xp33_ASAP7_75t_L     g10523(.A(new_n10775), .B(new_n10779), .Y(new_n10780));
  NOR2xp33_ASAP7_75t_L      g10524(.A(new_n10416), .B(new_n10417), .Y(new_n10781));
  NAND2xp33_ASAP7_75t_L     g10525(.A(new_n10418), .B(new_n10781), .Y(new_n10782));
  A2O1A1Ixp33_ASAP7_75t_L   g10526(.A1(new_n10419), .A2(new_n10415), .B(new_n10421), .C(new_n10782), .Y(new_n10783));
  NOR2xp33_ASAP7_75t_L      g10527(.A(new_n10780), .B(new_n10783), .Y(new_n10784));
  NOR3xp33_ASAP7_75t_L      g10528(.A(new_n10776), .B(new_n10777), .C(new_n10778), .Y(new_n10785));
  AOI21xp33_ASAP7_75t_L     g10529(.A1(new_n10768), .A2(new_n10767), .B(new_n10774), .Y(new_n10786));
  NOR2xp33_ASAP7_75t_L      g10530(.A(new_n10786), .B(new_n10785), .Y(new_n10787));
  A2O1A1O1Ixp25_ASAP7_75t_L g10531(.A1(new_n10419), .A2(new_n10415), .B(new_n10421), .C(new_n10782), .D(new_n10787), .Y(new_n10788));
  NAND2xp33_ASAP7_75t_L     g10532(.A(\b[43] ), .B(new_n1113), .Y(new_n10789));
  OAI221xp5_ASAP7_75t_L     g10533(.A1(new_n5680), .A2(new_n1298), .B1(new_n1197), .B2(new_n9799), .C(new_n10789), .Y(new_n10790));
  AOI21xp33_ASAP7_75t_L     g10534(.A1(new_n1194), .A2(\b[41] ), .B(new_n10790), .Y(new_n10791));
  NAND2xp33_ASAP7_75t_L     g10535(.A(\a[17] ), .B(new_n10791), .Y(new_n10792));
  A2O1A1Ixp33_ASAP7_75t_L   g10536(.A1(\b[41] ), .A2(new_n1194), .B(new_n10790), .C(new_n1107), .Y(new_n10793));
  NAND2xp33_ASAP7_75t_L     g10537(.A(new_n10793), .B(new_n10792), .Y(new_n10794));
  INVx1_ASAP7_75t_L         g10538(.A(new_n10794), .Y(new_n10795));
  OAI21xp33_ASAP7_75t_L     g10539(.A1(new_n10784), .A2(new_n10788), .B(new_n10795), .Y(new_n10796));
  NAND3xp33_ASAP7_75t_L     g10540(.A(new_n10787), .B(new_n10425), .C(new_n10782), .Y(new_n10797));
  A2O1A1Ixp33_ASAP7_75t_L   g10541(.A1(new_n10418), .A2(new_n10781), .B(new_n10436), .C(new_n10780), .Y(new_n10798));
  NAND3xp33_ASAP7_75t_L     g10542(.A(new_n10797), .B(new_n10798), .C(new_n10794), .Y(new_n10799));
  NAND2xp33_ASAP7_75t_L     g10543(.A(new_n10799), .B(new_n10796), .Y(new_n10800));
  NOR2xp33_ASAP7_75t_L      g10544(.A(new_n10544), .B(new_n10800), .Y(new_n10801));
  A2O1A1O1Ixp25_ASAP7_75t_L g10545(.A1(new_n10130), .A2(new_n10141), .B(new_n10224), .C(new_n10441), .D(new_n10437), .Y(new_n10802));
  AOI21xp33_ASAP7_75t_L     g10546(.A1(new_n10799), .A2(new_n10796), .B(new_n10802), .Y(new_n10803));
  NOR3xp33_ASAP7_75t_L      g10547(.A(new_n10801), .B(new_n10803), .C(new_n10543), .Y(new_n10804));
  INVx1_ASAP7_75t_L         g10548(.A(new_n10543), .Y(new_n10805));
  NAND3xp33_ASAP7_75t_L     g10549(.A(new_n10802), .B(new_n10796), .C(new_n10799), .Y(new_n10806));
  A2O1A1Ixp33_ASAP7_75t_L   g10550(.A1(new_n10441), .A2(new_n10226), .B(new_n10437), .C(new_n10800), .Y(new_n10807));
  AOI21xp33_ASAP7_75t_L     g10551(.A1(new_n10807), .A2(new_n10806), .B(new_n10805), .Y(new_n10808));
  AOI211xp5_ASAP7_75t_L     g10552(.A1(new_n10455), .A2(new_n10537), .B(new_n10804), .C(new_n10808), .Y(new_n10809));
  NAND3xp33_ASAP7_75t_L     g10553(.A(new_n10807), .B(new_n10806), .C(new_n10805), .Y(new_n10810));
  OAI21xp33_ASAP7_75t_L     g10554(.A1(new_n10803), .A2(new_n10801), .B(new_n10543), .Y(new_n10811));
  AOI211xp5_ASAP7_75t_L     g10555(.A1(new_n10810), .A2(new_n10811), .B(new_n10536), .C(new_n10452), .Y(new_n10812));
  OAI21xp33_ASAP7_75t_L     g10556(.A1(new_n10809), .A2(new_n10812), .B(new_n10535), .Y(new_n10813));
  A2O1A1O1Ixp25_ASAP7_75t_L g10557(.A1(new_n9806), .A2(new_n9809), .B(new_n9811), .C(new_n10151), .D(new_n10148), .Y(new_n10814));
  A2O1A1Ixp33_ASAP7_75t_L   g10558(.A1(new_n10457), .A2(new_n10456), .B(new_n10814), .C(new_n10537), .Y(new_n10815));
  NAND3xp33_ASAP7_75t_L     g10559(.A(new_n10815), .B(new_n10810), .C(new_n10811), .Y(new_n10816));
  OAI211xp5_ASAP7_75t_L     g10560(.A1(new_n10804), .A2(new_n10808), .B(new_n10537), .C(new_n10455), .Y(new_n10817));
  NAND3xp33_ASAP7_75t_L     g10561(.A(new_n10816), .B(new_n10534), .C(new_n10817), .Y(new_n10818));
  NAND3xp33_ASAP7_75t_L     g10562(.A(new_n10527), .B(new_n10813), .C(new_n10818), .Y(new_n10819));
  AOI21xp33_ASAP7_75t_L     g10563(.A1(new_n10459), .A2(new_n10455), .B(new_n10216), .Y(new_n10820));
  NOR3xp33_ASAP7_75t_L      g10564(.A(new_n10452), .B(new_n10453), .C(new_n10217), .Y(new_n10821));
  NOR2xp33_ASAP7_75t_L      g10565(.A(new_n10820), .B(new_n10821), .Y(new_n10822));
  NOR2xp33_ASAP7_75t_L      g10566(.A(new_n10216), .B(new_n10526), .Y(new_n10823));
  INVx1_ASAP7_75t_L         g10567(.A(new_n10823), .Y(new_n10824));
  AOI21xp33_ASAP7_75t_L     g10568(.A1(new_n10816), .A2(new_n10817), .B(new_n10534), .Y(new_n10825));
  NOR3xp33_ASAP7_75t_L      g10569(.A(new_n10812), .B(new_n10809), .C(new_n10535), .Y(new_n10826));
  OAI221xp5_ASAP7_75t_L     g10570(.A1(new_n10822), .A2(new_n10210), .B1(new_n10826), .B2(new_n10825), .C(new_n10824), .Y(new_n10827));
  AOI21xp33_ASAP7_75t_L     g10571(.A1(new_n10819), .A2(new_n10827), .B(new_n10525), .Y(new_n10828));
  AND3x1_ASAP7_75t_L        g10572(.A(new_n10819), .B(new_n10827), .C(new_n10525), .Y(new_n10829));
  NOR3xp33_ASAP7_75t_L      g10573(.A(new_n10518), .B(new_n10828), .C(new_n10829), .Y(new_n10830));
  NOR3xp33_ASAP7_75t_L      g10574(.A(new_n10464), .B(new_n10461), .C(new_n10208), .Y(new_n10831));
  AO21x2_ASAP7_75t_L        g10575(.A1(new_n10827), .A2(new_n10819), .B(new_n10525), .Y(new_n10832));
  NAND3xp33_ASAP7_75t_L     g10576(.A(new_n10819), .B(new_n10827), .C(new_n10525), .Y(new_n10833));
  AOI221xp5_ASAP7_75t_L     g10577(.A1(new_n10201), .A2(new_n10469), .B1(new_n10833), .B2(new_n10832), .C(new_n10831), .Y(new_n10834));
  OAI21xp33_ASAP7_75t_L     g10578(.A1(new_n10834), .A2(new_n10830), .B(new_n10516), .Y(new_n10835));
  INVx1_ASAP7_75t_L         g10579(.A(new_n10516), .Y(new_n10836));
  NOR2xp33_ASAP7_75t_L      g10580(.A(new_n10828), .B(new_n10829), .Y(new_n10837));
  OAI21xp33_ASAP7_75t_L     g10581(.A1(new_n10831), .A2(new_n10478), .B(new_n10837), .Y(new_n10838));
  OAI21xp33_ASAP7_75t_L     g10582(.A1(new_n10828), .A2(new_n10829), .B(new_n10518), .Y(new_n10839));
  NAND3xp33_ASAP7_75t_L     g10583(.A(new_n10838), .B(new_n10836), .C(new_n10839), .Y(new_n10840));
  NAND3xp33_ASAP7_75t_L     g10584(.A(new_n10509), .B(new_n10835), .C(new_n10840), .Y(new_n10841));
  AOI21xp33_ASAP7_75t_L     g10585(.A1(new_n10838), .A2(new_n10839), .B(new_n10836), .Y(new_n10842));
  NOR3xp33_ASAP7_75t_L      g10586(.A(new_n10830), .B(new_n10834), .C(new_n10516), .Y(new_n10843));
  OAI221xp5_ASAP7_75t_L     g10587(.A1(new_n10842), .A2(new_n10843), .B1(new_n10481), .B2(new_n10484), .C(new_n10508), .Y(new_n10844));
  NAND2xp33_ASAP7_75t_L     g10588(.A(\b[56] ), .B(new_n291), .Y(new_n10845));
  NAND2xp33_ASAP7_75t_L     g10589(.A(\b[57] ), .B(new_n380), .Y(new_n10846));
  NOR2xp33_ASAP7_75t_L      g10590(.A(\b[57] ), .B(\b[58] ), .Y(new_n10847));
  INVx1_ASAP7_75t_L         g10591(.A(\b[58] ), .Y(new_n10848));
  NOR2xp33_ASAP7_75t_L      g10592(.A(new_n10488), .B(new_n10848), .Y(new_n10849));
  NOR2xp33_ASAP7_75t_L      g10593(.A(new_n10847), .B(new_n10849), .Y(new_n10850));
  A2O1A1Ixp33_ASAP7_75t_L   g10594(.A1(\b[57] ), .A2(\b[56] ), .B(new_n10492), .C(new_n10850), .Y(new_n10851));
  INVx1_ASAP7_75t_L         g10595(.A(new_n10489), .Y(new_n10852));
  A2O1A1Ixp33_ASAP7_75t_L   g10596(.A1(new_n10181), .A2(new_n10486), .B(new_n10487), .C(new_n10852), .Y(new_n10853));
  NOR2xp33_ASAP7_75t_L      g10597(.A(new_n10850), .B(new_n10853), .Y(new_n10854));
  INVx1_ASAP7_75t_L         g10598(.A(new_n10854), .Y(new_n10855));
  NAND2xp33_ASAP7_75t_L     g10599(.A(new_n10851), .B(new_n10855), .Y(new_n10856));
  INVx1_ASAP7_75t_L         g10600(.A(new_n10856), .Y(new_n10857));
  AOI22xp33_ASAP7_75t_L     g10601(.A1(new_n272), .A2(\b[58] ), .B1(new_n269), .B2(new_n10857), .Y(new_n10858));
  NAND4xp25_ASAP7_75t_L     g10602(.A(new_n10858), .B(\a[2] ), .C(new_n10845), .D(new_n10846), .Y(new_n10859));
  NAND2xp33_ASAP7_75t_L     g10603(.A(new_n10846), .B(new_n10858), .Y(new_n10860));
  A2O1A1Ixp33_ASAP7_75t_L   g10604(.A1(\b[56] ), .A2(new_n291), .B(new_n10860), .C(new_n265), .Y(new_n10861));
  NAND2xp33_ASAP7_75t_L     g10605(.A(new_n10859), .B(new_n10861), .Y(new_n10862));
  INVx1_ASAP7_75t_L         g10606(.A(new_n10862), .Y(new_n10863));
  NAND3xp33_ASAP7_75t_L     g10607(.A(new_n10841), .B(new_n10863), .C(new_n10844), .Y(new_n10864));
  A2O1A1Ixp33_ASAP7_75t_L   g10608(.A1(new_n10172), .A2(new_n9863), .B(new_n10173), .C(new_n10170), .Y(new_n10865));
  OAI21xp33_ASAP7_75t_L     g10609(.A1(new_n10476), .A2(new_n10480), .B(new_n10865), .Y(new_n10866));
  NAND2xp33_ASAP7_75t_L     g10610(.A(new_n10835), .B(new_n10840), .Y(new_n10867));
  AOI21xp33_ASAP7_75t_L     g10611(.A1(new_n10866), .A2(new_n10508), .B(new_n10867), .Y(new_n10868));
  AOI21xp33_ASAP7_75t_L     g10612(.A1(new_n10840), .A2(new_n10835), .B(new_n10509), .Y(new_n10869));
  OAI21xp33_ASAP7_75t_L     g10613(.A1(new_n10869), .A2(new_n10868), .B(new_n10862), .Y(new_n10870));
  NAND2xp33_ASAP7_75t_L     g10614(.A(new_n10864), .B(new_n10870), .Y(new_n10871));
  A2O1A1Ixp33_ASAP7_75t_L   g10615(.A1(new_n10503), .A2(new_n10192), .B(new_n10501), .C(new_n10871), .Y(new_n10872));
  INVx1_ASAP7_75t_L         g10616(.A(new_n10872), .Y(new_n10873));
  AO21x2_ASAP7_75t_L        g10617(.A1(new_n10503), .A2(new_n10192), .B(new_n10501), .Y(new_n10874));
  NOR2xp33_ASAP7_75t_L      g10618(.A(new_n10874), .B(new_n10871), .Y(new_n10875));
  NOR2xp33_ASAP7_75t_L      g10619(.A(new_n10875), .B(new_n10873), .Y(\f[58] ));
  NAND2xp33_ASAP7_75t_L     g10620(.A(new_n10844), .B(new_n10841), .Y(new_n10877));
  A2O1A1Ixp33_ASAP7_75t_L   g10621(.A1(new_n10859), .A2(new_n10861), .B(new_n10877), .C(new_n10872), .Y(new_n10878));
  A2O1A1Ixp33_ASAP7_75t_L   g10622(.A1(new_n10866), .A2(new_n10508), .B(new_n10842), .C(new_n10840), .Y(new_n10879));
  NOR2xp33_ASAP7_75t_L      g10623(.A(\b[58] ), .B(\b[59] ), .Y(new_n10880));
  INVx1_ASAP7_75t_L         g10624(.A(\b[59] ), .Y(new_n10881));
  NOR2xp33_ASAP7_75t_L      g10625(.A(new_n10848), .B(new_n10881), .Y(new_n10882));
  NOR2xp33_ASAP7_75t_L      g10626(.A(new_n10880), .B(new_n10882), .Y(new_n10883));
  A2O1A1Ixp33_ASAP7_75t_L   g10627(.A1(new_n10853), .A2(new_n10850), .B(new_n10849), .C(new_n10883), .Y(new_n10884));
  INVx1_ASAP7_75t_L         g10628(.A(new_n10884), .Y(new_n10885));
  AOI211xp5_ASAP7_75t_L     g10629(.A1(new_n10853), .A2(new_n10850), .B(new_n10883), .C(new_n10849), .Y(new_n10886));
  NOR2xp33_ASAP7_75t_L      g10630(.A(new_n10886), .B(new_n10885), .Y(new_n10887));
  INVx1_ASAP7_75t_L         g10631(.A(new_n10887), .Y(new_n10888));
  NOR2xp33_ASAP7_75t_L      g10632(.A(new_n10848), .B(new_n261), .Y(new_n10889));
  AOI221xp5_ASAP7_75t_L     g10633(.A1(\b[57] ), .A2(new_n291), .B1(\b[59] ), .B2(new_n272), .C(new_n10889), .Y(new_n10890));
  OA211x2_ASAP7_75t_L       g10634(.A1(new_n292), .A2(new_n10888), .B(new_n10890), .C(\a[2] ), .Y(new_n10891));
  O2A1O1Ixp33_ASAP7_75t_L   g10635(.A1(new_n292), .A2(new_n10888), .B(new_n10890), .C(\a[2] ), .Y(new_n10892));
  NOR2xp33_ASAP7_75t_L      g10636(.A(new_n10892), .B(new_n10891), .Y(new_n10893));
  A2O1A1O1Ixp25_ASAP7_75t_L g10637(.A1(new_n10201), .A2(new_n10469), .B(new_n10831), .C(new_n10832), .D(new_n10829), .Y(new_n10894));
  NAND2xp33_ASAP7_75t_L     g10638(.A(\b[53] ), .B(new_n451), .Y(new_n10895));
  OAI221xp5_ASAP7_75t_L     g10639(.A1(new_n8569), .A2(new_n529), .B1(new_n482), .B2(new_n8888), .C(new_n10895), .Y(new_n10896));
  AOI21xp33_ASAP7_75t_L     g10640(.A1(new_n480), .A2(\b[51] ), .B(new_n10896), .Y(new_n10897));
  NAND2xp33_ASAP7_75t_L     g10641(.A(\a[8] ), .B(new_n10897), .Y(new_n10898));
  A2O1A1Ixp33_ASAP7_75t_L   g10642(.A1(\b[51] ), .A2(new_n480), .B(new_n10896), .C(new_n445), .Y(new_n10899));
  NAND2xp33_ASAP7_75t_L     g10643(.A(new_n10899), .B(new_n10898), .Y(new_n10900));
  INVx1_ASAP7_75t_L         g10644(.A(new_n10900), .Y(new_n10901));
  A2O1A1O1Ixp25_ASAP7_75t_L g10645(.A1(new_n10463), .A2(new_n10462), .B(new_n10823), .C(new_n10813), .D(new_n10826), .Y(new_n10902));
  A2O1A1Ixp33_ASAP7_75t_L   g10646(.A1(new_n10455), .A2(new_n10537), .B(new_n10804), .C(new_n10811), .Y(new_n10903));
  NOR2xp33_ASAP7_75t_L      g10647(.A(new_n6756), .B(new_n909), .Y(new_n10904));
  INVx1_ASAP7_75t_L         g10648(.A(new_n10904), .Y(new_n10905));
  NAND2xp33_ASAP7_75t_L     g10649(.A(\b[46] ), .B(new_n817), .Y(new_n10906));
  AOI22xp33_ASAP7_75t_L     g10650(.A1(new_n826), .A2(\b[47] ), .B1(new_n823), .B2(new_n7323), .Y(new_n10907));
  AND4x1_ASAP7_75t_L        g10651(.A(new_n10907), .B(new_n10906), .C(new_n10905), .D(\a[14] ), .Y(new_n10908));
  AOI31xp33_ASAP7_75t_L     g10652(.A1(new_n10907), .A2(new_n10906), .A3(new_n10905), .B(\a[14] ), .Y(new_n10909));
  NOR2xp33_ASAP7_75t_L      g10653(.A(new_n10909), .B(new_n10908), .Y(new_n10910));
  INVx1_ASAP7_75t_L         g10654(.A(new_n10910), .Y(new_n10911));
  NAND2xp33_ASAP7_75t_L     g10655(.A(\b[44] ), .B(new_n1113), .Y(new_n10912));
  OAI221xp5_ASAP7_75t_L     g10656(.A1(new_n6195), .A2(new_n1298), .B1(new_n1197), .B2(new_n6229), .C(new_n10912), .Y(new_n10913));
  AOI21xp33_ASAP7_75t_L     g10657(.A1(new_n1194), .A2(\b[42] ), .B(new_n10913), .Y(new_n10914));
  NAND2xp33_ASAP7_75t_L     g10658(.A(\a[17] ), .B(new_n10914), .Y(new_n10915));
  A2O1A1Ixp33_ASAP7_75t_L   g10659(.A1(\b[42] ), .A2(new_n1194), .B(new_n10913), .C(new_n1107), .Y(new_n10916));
  NAND2xp33_ASAP7_75t_L     g10660(.A(new_n10916), .B(new_n10915), .Y(new_n10917));
  NOR3xp33_ASAP7_75t_L      g10661(.A(new_n10776), .B(new_n10777), .C(new_n10774), .Y(new_n10918));
  INVx1_ASAP7_75t_L         g10662(.A(new_n10918), .Y(new_n10919));
  A2O1A1Ixp33_ASAP7_75t_L   g10663(.A1(new_n10782), .A2(new_n10425), .B(new_n10787), .C(new_n10919), .Y(new_n10920));
  OAI21xp33_ASAP7_75t_L     g10664(.A1(new_n10738), .A2(new_n10545), .B(new_n10741), .Y(new_n10921));
  NAND2xp33_ASAP7_75t_L     g10665(.A(new_n2700), .B(new_n3450), .Y(new_n10922));
  OAI221xp5_ASAP7_75t_L     g10666(.A1(new_n2708), .A2(new_n3443), .B1(new_n3419), .B2(new_n2694), .C(new_n10922), .Y(new_n10923));
  AOI21xp33_ASAP7_75t_L     g10667(.A1(new_n2931), .A2(\b[30] ), .B(new_n10923), .Y(new_n10924));
  NAND2xp33_ASAP7_75t_L     g10668(.A(\a[29] ), .B(new_n10924), .Y(new_n10925));
  A2O1A1Ixp33_ASAP7_75t_L   g10669(.A1(\b[30] ), .A2(new_n2931), .B(new_n10923), .C(new_n2697), .Y(new_n10926));
  AND2x2_ASAP7_75t_L        g10670(.A(new_n10926), .B(new_n10925), .Y(new_n10927));
  INVx1_ASAP7_75t_L         g10671(.A(new_n10374), .Y(new_n10928));
  NAND3xp33_ASAP7_75t_L     g10672(.A(new_n10706), .B(new_n10710), .C(new_n10721), .Y(new_n10929));
  INVx1_ASAP7_75t_L         g10673(.A(new_n10929), .Y(new_n10930));
  A2O1A1O1Ixp25_ASAP7_75t_L g10674(.A1(new_n10362), .A2(new_n10928), .B(new_n10724), .C(new_n10726), .D(new_n10930), .Y(new_n10931));
  A2O1A1O1Ixp25_ASAP7_75t_L g10675(.A1(new_n10244), .A2(new_n10340), .B(new_n10342), .C(new_n10688), .D(new_n10691), .Y(new_n10932));
  AOI32xp33_ASAP7_75t_L     g10676(.A1(new_n1998), .A2(new_n2001), .A3(new_n4542), .B1(new_n4544), .B2(\b[23] ), .Y(new_n10933));
  OAI221xp5_ASAP7_75t_L     g10677(.A1(new_n4536), .A2(new_n1857), .B1(new_n1709), .B2(new_n4781), .C(new_n10933), .Y(new_n10934));
  XNOR2x2_ASAP7_75t_L       g10678(.A(\a[38] ), .B(new_n10934), .Y(new_n10935));
  INVx1_ASAP7_75t_L         g10679(.A(new_n10935), .Y(new_n10936));
  NAND2xp33_ASAP7_75t_L     g10680(.A(\b[18] ), .B(new_n5526), .Y(new_n10937));
  NOR2xp33_ASAP7_75t_L      g10681(.A(new_n1594), .B(new_n5253), .Y(new_n10938));
  AOI221xp5_ASAP7_75t_L     g10682(.A1(new_n5240), .A2(\b[19] ), .B1(new_n5247), .B2(new_n1600), .C(new_n10938), .Y(new_n10939));
  NAND3xp33_ASAP7_75t_L     g10683(.A(new_n10939), .B(new_n10937), .C(\a[41] ), .Y(new_n10940));
  AO21x2_ASAP7_75t_L        g10684(.A1(new_n10937), .A2(new_n10939), .B(\a[41] ), .Y(new_n10941));
  NAND2xp33_ASAP7_75t_L     g10685(.A(new_n10940), .B(new_n10941), .Y(new_n10942));
  NOR2xp33_ASAP7_75t_L      g10686(.A(new_n952), .B(new_n6309), .Y(new_n10943));
  NAND2xp33_ASAP7_75t_L     g10687(.A(\b[17] ), .B(new_n6002), .Y(new_n10944));
  OAI221xp5_ASAP7_75t_L     g10688(.A1(new_n1051), .A2(new_n6544), .B1(new_n6311), .B2(new_n1251), .C(new_n10944), .Y(new_n10945));
  NOR3xp33_ASAP7_75t_L      g10689(.A(new_n10945), .B(new_n10943), .C(new_n5996), .Y(new_n10946));
  OA21x2_ASAP7_75t_L        g10690(.A1(new_n10943), .A2(new_n10945), .B(new_n5996), .Y(new_n10947));
  NOR2xp33_ASAP7_75t_L      g10691(.A(new_n10946), .B(new_n10947), .Y(new_n10948));
  INVx1_ASAP7_75t_L         g10692(.A(new_n10948), .Y(new_n10949));
  NAND2xp33_ASAP7_75t_L     g10693(.A(new_n10624), .B(new_n10625), .Y(new_n10950));
  MAJIxp5_ASAP7_75t_L       g10694(.A(new_n10632), .B(new_n10626), .C(new_n10950), .Y(new_n10951));
  NAND2xp33_ASAP7_75t_L     g10695(.A(\b[10] ), .B(new_n7649), .Y(new_n10952));
  OAI221xp5_ASAP7_75t_L     g10696(.A1(new_n7997), .A2(new_n695), .B1(new_n7996), .B2(new_n701), .C(new_n10952), .Y(new_n10953));
  AOI21xp33_ASAP7_75t_L     g10697(.A1(new_n7993), .A2(\b[9] ), .B(new_n10953), .Y(new_n10954));
  NAND2xp33_ASAP7_75t_L     g10698(.A(\a[50] ), .B(new_n10954), .Y(new_n10955));
  A2O1A1Ixp33_ASAP7_75t_L   g10699(.A1(\b[9] ), .A2(new_n7993), .B(new_n10953), .C(new_n7653), .Y(new_n10956));
  AOI21xp33_ASAP7_75t_L     g10700(.A1(new_n10613), .A2(new_n10612), .B(new_n10609), .Y(new_n10957));
  NAND2xp33_ASAP7_75t_L     g10701(.A(\b[6] ), .B(new_n8964), .Y(new_n10958));
  NAND2xp33_ASAP7_75t_L     g10702(.A(\b[7] ), .B(new_n8635), .Y(new_n10959));
  AOI22xp33_ASAP7_75t_L     g10703(.A1(new_n8645), .A2(\b[8] ), .B1(new_n8642), .B2(new_n510), .Y(new_n10960));
  NAND3xp33_ASAP7_75t_L     g10704(.A(new_n10960), .B(new_n10959), .C(new_n10958), .Y(new_n10961));
  NOR2xp33_ASAP7_75t_L      g10705(.A(new_n8639), .B(new_n10961), .Y(new_n10962));
  NAND2xp33_ASAP7_75t_L     g10706(.A(new_n8639), .B(new_n10961), .Y(new_n10963));
  INVx1_ASAP7_75t_L         g10707(.A(new_n10963), .Y(new_n10964));
  O2A1O1Ixp33_ASAP7_75t_L   g10708(.A1(new_n10574), .A2(new_n10573), .B(new_n10598), .C(new_n10603), .Y(new_n10965));
  NAND2xp33_ASAP7_75t_L     g10709(.A(\b[3] ), .B(new_n9948), .Y(new_n10966));
  NAND2xp33_ASAP7_75t_L     g10710(.A(\b[4] ), .B(new_n9614), .Y(new_n10967));
  AOI22xp33_ASAP7_75t_L     g10711(.A1(new_n9623), .A2(\b[5] ), .B1(new_n9620), .B2(new_n360), .Y(new_n10968));
  NAND4xp25_ASAP7_75t_L     g10712(.A(new_n10968), .B(\a[56] ), .C(new_n10966), .D(new_n10967), .Y(new_n10969));
  AOI31xp33_ASAP7_75t_L     g10713(.A1(new_n10968), .A2(new_n10967), .A3(new_n10966), .B(\a[56] ), .Y(new_n10970));
  INVx1_ASAP7_75t_L         g10714(.A(new_n10970), .Y(new_n10971));
  INVx1_ASAP7_75t_L         g10715(.A(new_n10583), .Y(new_n10972));
  NOR3xp33_ASAP7_75t_L      g10716(.A(new_n10590), .B(new_n10972), .C(new_n10582), .Y(new_n10973));
  NAND2xp33_ASAP7_75t_L     g10717(.A(new_n10593), .B(new_n10582), .Y(new_n10974));
  NAND2xp33_ASAP7_75t_L     g10718(.A(new_n10582), .B(new_n10590), .Y(new_n10975));
  NAND2xp33_ASAP7_75t_L     g10719(.A(\b[1] ), .B(new_n10584), .Y(new_n10976));
  OAI221xp5_ASAP7_75t_L     g10720(.A1(new_n10974), .A2(new_n283), .B1(new_n278), .B2(new_n10975), .C(new_n10976), .Y(new_n10977));
  AOI21xp33_ASAP7_75t_L     g10721(.A1(new_n10973), .A2(\b[0] ), .B(new_n10977), .Y(new_n10978));
  A2O1A1Ixp33_ASAP7_75t_L   g10722(.A1(new_n10278), .A2(new_n10596), .B(new_n10588), .C(new_n10978), .Y(new_n10979));
  O2A1O1Ixp33_ASAP7_75t_L   g10723(.A1(new_n258), .A2(new_n10275), .B(new_n10596), .C(new_n10588), .Y(new_n10980));
  A2O1A1Ixp33_ASAP7_75t_L   g10724(.A1(\b[0] ), .A2(new_n10973), .B(new_n10977), .C(new_n10980), .Y(new_n10981));
  NAND2xp33_ASAP7_75t_L     g10725(.A(new_n10979), .B(new_n10981), .Y(new_n10982));
  NAND3xp33_ASAP7_75t_L     g10726(.A(new_n10982), .B(new_n10971), .C(new_n10969), .Y(new_n10983));
  INVx1_ASAP7_75t_L         g10727(.A(new_n10969), .Y(new_n10984));
  AND2x2_ASAP7_75t_L        g10728(.A(new_n10979), .B(new_n10981), .Y(new_n10985));
  OAI21xp33_ASAP7_75t_L     g10729(.A1(new_n10970), .A2(new_n10984), .B(new_n10985), .Y(new_n10986));
  NAND3xp33_ASAP7_75t_L     g10730(.A(new_n10965), .B(new_n10983), .C(new_n10986), .Y(new_n10987));
  INVx1_ASAP7_75t_L         g10731(.A(new_n10987), .Y(new_n10988));
  AOI21xp33_ASAP7_75t_L     g10732(.A1(new_n10986), .A2(new_n10983), .B(new_n10965), .Y(new_n10989));
  NOR4xp25_ASAP7_75t_L      g10733(.A(new_n10964), .B(new_n10989), .C(new_n10962), .D(new_n10988), .Y(new_n10990));
  AND3x1_ASAP7_75t_L        g10734(.A(new_n10960), .B(new_n10959), .C(new_n10958), .Y(new_n10991));
  NAND2xp33_ASAP7_75t_L     g10735(.A(\a[53] ), .B(new_n10991), .Y(new_n10992));
  INVx1_ASAP7_75t_L         g10736(.A(new_n10989), .Y(new_n10993));
  AOI22xp33_ASAP7_75t_L     g10737(.A1(new_n10992), .A2(new_n10963), .B1(new_n10987), .B2(new_n10993), .Y(new_n10994));
  NOR3xp33_ASAP7_75t_L      g10738(.A(new_n10990), .B(new_n10994), .C(new_n10957), .Y(new_n10995));
  A2O1A1Ixp33_ASAP7_75t_L   g10739(.A1(new_n10567), .A2(new_n10566), .B(new_n10605), .C(new_n10614), .Y(new_n10996));
  NAND4xp25_ASAP7_75t_L     g10740(.A(new_n10993), .B(new_n10992), .C(new_n10963), .D(new_n10987), .Y(new_n10997));
  OAI22xp33_ASAP7_75t_L     g10741(.A1(new_n10964), .A2(new_n10962), .B1(new_n10989), .B2(new_n10988), .Y(new_n10998));
  AOI21xp33_ASAP7_75t_L     g10742(.A1(new_n10998), .A2(new_n10997), .B(new_n10996), .Y(new_n10999));
  OAI211xp5_ASAP7_75t_L     g10743(.A1(new_n10999), .A2(new_n10995), .B(new_n10956), .C(new_n10955), .Y(new_n11000));
  NAND2xp33_ASAP7_75t_L     g10744(.A(new_n10956), .B(new_n10955), .Y(new_n11001));
  NAND3xp33_ASAP7_75t_L     g10745(.A(new_n10998), .B(new_n10996), .C(new_n10997), .Y(new_n11002));
  OAI21xp33_ASAP7_75t_L     g10746(.A1(new_n10994), .A2(new_n10990), .B(new_n10957), .Y(new_n11003));
  NAND3xp33_ASAP7_75t_L     g10747(.A(new_n11003), .B(new_n11001), .C(new_n11002), .Y(new_n11004));
  NAND3xp33_ASAP7_75t_L     g10748(.A(new_n10951), .B(new_n11000), .C(new_n11004), .Y(new_n11005));
  NOR2xp33_ASAP7_75t_L      g10749(.A(new_n10615), .B(new_n10610), .Y(new_n11006));
  MAJIxp5_ASAP7_75t_L       g10750(.A(new_n10628), .B(new_n10622), .C(new_n11006), .Y(new_n11007));
  AOI21xp33_ASAP7_75t_L     g10751(.A1(new_n11003), .A2(new_n11002), .B(new_n11001), .Y(new_n11008));
  AOI211xp5_ASAP7_75t_L     g10752(.A1(new_n10956), .A2(new_n10955), .B(new_n10999), .C(new_n10995), .Y(new_n11009));
  OAI21xp33_ASAP7_75t_L     g10753(.A1(new_n11008), .A2(new_n11009), .B(new_n11007), .Y(new_n11010));
  NOR2xp33_ASAP7_75t_L      g10754(.A(new_n763), .B(new_n7115), .Y(new_n11011));
  NAND2xp33_ASAP7_75t_L     g10755(.A(\b[13] ), .B(new_n6812), .Y(new_n11012));
  OAI221xp5_ASAP7_75t_L     g10756(.A1(new_n7118), .A2(new_n871), .B1(new_n7117), .B2(new_n878), .C(new_n11012), .Y(new_n11013));
  OR3x1_ASAP7_75t_L         g10757(.A(new_n11013), .B(new_n6816), .C(new_n11011), .Y(new_n11014));
  A2O1A1Ixp33_ASAP7_75t_L   g10758(.A1(\b[12] ), .A2(new_n7124), .B(new_n11013), .C(new_n6816), .Y(new_n11015));
  AND2x2_ASAP7_75t_L        g10759(.A(new_n11015), .B(new_n11014), .Y(new_n11016));
  NAND3xp33_ASAP7_75t_L     g10760(.A(new_n11016), .B(new_n11005), .C(new_n11010), .Y(new_n11017));
  NOR3xp33_ASAP7_75t_L      g10761(.A(new_n11007), .B(new_n11008), .C(new_n11009), .Y(new_n11018));
  AOI21xp33_ASAP7_75t_L     g10762(.A1(new_n11000), .A2(new_n11004), .B(new_n10951), .Y(new_n11019));
  NAND2xp33_ASAP7_75t_L     g10763(.A(new_n11015), .B(new_n11014), .Y(new_n11020));
  OAI21xp33_ASAP7_75t_L     g10764(.A1(new_n11019), .A2(new_n11018), .B(new_n11020), .Y(new_n11021));
  NOR3xp33_ASAP7_75t_L      g10765(.A(new_n10641), .B(new_n10633), .C(new_n10629), .Y(new_n11022));
  AOI21xp33_ASAP7_75t_L     g10766(.A1(new_n10652), .A2(new_n10642), .B(new_n11022), .Y(new_n11023));
  AOI21xp33_ASAP7_75t_L     g10767(.A1(new_n11021), .A2(new_n11017), .B(new_n11023), .Y(new_n11024));
  NOR3xp33_ASAP7_75t_L      g10768(.A(new_n11018), .B(new_n11019), .C(new_n11020), .Y(new_n11025));
  AOI21xp33_ASAP7_75t_L     g10769(.A1(new_n11005), .A2(new_n11010), .B(new_n11016), .Y(new_n11026));
  AOI21xp33_ASAP7_75t_L     g10770(.A1(new_n10643), .A2(new_n10644), .B(new_n10648), .Y(new_n11027));
  O2A1O1Ixp33_ASAP7_75t_L   g10771(.A1(new_n10313), .A2(new_n10261), .B(new_n10651), .C(new_n11027), .Y(new_n11028));
  NOR4xp25_ASAP7_75t_L      g10772(.A(new_n11028), .B(new_n11025), .C(new_n11022), .D(new_n11026), .Y(new_n11029));
  OAI21xp33_ASAP7_75t_L     g10773(.A1(new_n11029), .A2(new_n11024), .B(new_n10949), .Y(new_n11030));
  OAI22xp33_ASAP7_75t_L     g10774(.A1(new_n11028), .A2(new_n11022), .B1(new_n11026), .B2(new_n11025), .Y(new_n11031));
  NAND3xp33_ASAP7_75t_L     g10775(.A(new_n11023), .B(new_n11021), .C(new_n11017), .Y(new_n11032));
  NAND3xp33_ASAP7_75t_L     g10776(.A(new_n11032), .B(new_n10948), .C(new_n11031), .Y(new_n11033));
  NAND2xp33_ASAP7_75t_L     g10777(.A(new_n11033), .B(new_n11030), .Y(new_n11034));
  A2O1A1Ixp33_ASAP7_75t_L   g10778(.A1(new_n10660), .A2(new_n10555), .B(new_n10655), .C(new_n11034), .Y(new_n11035));
  A2O1A1O1Ixp25_ASAP7_75t_L g10779(.A1(new_n10320), .A2(new_n10255), .B(new_n10325), .C(new_n10665), .D(new_n10655), .Y(new_n11036));
  NAND3xp33_ASAP7_75t_L     g10780(.A(new_n11036), .B(new_n11030), .C(new_n11033), .Y(new_n11037));
  NAND3xp33_ASAP7_75t_L     g10781(.A(new_n11035), .B(new_n10942), .C(new_n11037), .Y(new_n11038));
  AND2x2_ASAP7_75t_L        g10782(.A(new_n10940), .B(new_n10941), .Y(new_n11039));
  AOI21xp33_ASAP7_75t_L     g10783(.A1(new_n11033), .A2(new_n11030), .B(new_n11036), .Y(new_n11040));
  AND3x1_ASAP7_75t_L        g10784(.A(new_n11036), .B(new_n11033), .C(new_n11030), .Y(new_n11041));
  OAI21xp33_ASAP7_75t_L     g10785(.A1(new_n11040), .A2(new_n11041), .B(new_n11039), .Y(new_n11042));
  O2A1O1Ixp33_ASAP7_75t_L   g10786(.A1(new_n10250), .A2(new_n10336), .B(new_n10553), .C(new_n10678), .Y(new_n11043));
  OAI211xp5_ASAP7_75t_L     g10787(.A1(new_n10679), .A2(new_n11043), .B(new_n11038), .C(new_n11042), .Y(new_n11044));
  NAND2xp33_ASAP7_75t_L     g10788(.A(new_n11042), .B(new_n11038), .Y(new_n11045));
  A2O1A1O1Ixp25_ASAP7_75t_L g10789(.A1(new_n10330), .A2(new_n10338), .B(new_n10684), .C(new_n10671), .D(new_n10679), .Y(new_n11046));
  NAND2xp33_ASAP7_75t_L     g10790(.A(new_n11045), .B(new_n11046), .Y(new_n11047));
  NAND3xp33_ASAP7_75t_L     g10791(.A(new_n11044), .B(new_n10936), .C(new_n11047), .Y(new_n11048));
  O2A1O1Ixp33_ASAP7_75t_L   g10792(.A1(new_n10685), .A2(new_n10678), .B(new_n10675), .C(new_n11045), .Y(new_n11049));
  AOI211xp5_ASAP7_75t_L     g10793(.A1(new_n11038), .A2(new_n11042), .B(new_n10679), .C(new_n11043), .Y(new_n11050));
  OAI21xp33_ASAP7_75t_L     g10794(.A1(new_n11050), .A2(new_n11049), .B(new_n10935), .Y(new_n11051));
  NAND2xp33_ASAP7_75t_L     g10795(.A(new_n11048), .B(new_n11051), .Y(new_n11052));
  NAND2xp33_ASAP7_75t_L     g10796(.A(new_n10932), .B(new_n11052), .Y(new_n11053));
  NOR3xp33_ASAP7_75t_L      g10797(.A(new_n11049), .B(new_n11050), .C(new_n10935), .Y(new_n11054));
  AOI21xp33_ASAP7_75t_L     g10798(.A1(new_n11044), .A2(new_n11047), .B(new_n10936), .Y(new_n11055));
  NOR2xp33_ASAP7_75t_L      g10799(.A(new_n11055), .B(new_n11054), .Y(new_n11056));
  A2O1A1Ixp33_ASAP7_75t_L   g10800(.A1(new_n10688), .A2(new_n10699), .B(new_n10691), .C(new_n11056), .Y(new_n11057));
  OAI22xp33_ASAP7_75t_L     g10801(.A1(new_n2487), .A2(new_n4114), .B1(new_n4115), .B2(new_n2477), .Y(new_n11058));
  AOI221xp5_ASAP7_75t_L     g10802(.A1(\b[24] ), .A2(new_n4111), .B1(\b[25] ), .B2(new_n3874), .C(new_n11058), .Y(new_n11059));
  AND2x2_ASAP7_75t_L        g10803(.A(\a[35] ), .B(new_n11059), .Y(new_n11060));
  NOR2xp33_ASAP7_75t_L      g10804(.A(\a[35] ), .B(new_n11059), .Y(new_n11061));
  NOR2xp33_ASAP7_75t_L      g10805(.A(new_n11061), .B(new_n11060), .Y(new_n11062));
  NAND3xp33_ASAP7_75t_L     g10806(.A(new_n11057), .B(new_n11053), .C(new_n11062), .Y(new_n11063));
  AOI221xp5_ASAP7_75t_L     g10807(.A1(new_n11051), .A2(new_n11048), .B1(new_n10688), .B2(new_n10699), .C(new_n10691), .Y(new_n11064));
  O2A1O1Ixp33_ASAP7_75t_L   g10808(.A1(new_n10548), .A2(new_n10692), .B(new_n10682), .C(new_n11052), .Y(new_n11065));
  OR2x4_ASAP7_75t_L         g10809(.A(new_n11061), .B(new_n11060), .Y(new_n11066));
  OAI21xp33_ASAP7_75t_L     g10810(.A1(new_n11064), .A2(new_n11065), .B(new_n11066), .Y(new_n11067));
  XNOR2x2_ASAP7_75t_L       g10811(.A(new_n10699), .B(new_n10689), .Y(new_n11068));
  MAJIxp5_ASAP7_75t_L       g10812(.A(new_n10709), .B(new_n10703), .C(new_n11068), .Y(new_n11069));
  NAND3xp33_ASAP7_75t_L     g10813(.A(new_n11069), .B(new_n11067), .C(new_n11063), .Y(new_n11070));
  NAND2xp33_ASAP7_75t_L     g10814(.A(new_n11067), .B(new_n11063), .Y(new_n11071));
  A2O1A1Ixp33_ASAP7_75t_L   g10815(.A1(new_n10703), .A2(new_n11068), .B(new_n10720), .C(new_n11071), .Y(new_n11072));
  AOI22xp33_ASAP7_75t_L     g10816(.A1(new_n3256), .A2(\b[29] ), .B1(new_n3254), .B2(new_n5472), .Y(new_n11073));
  OAI221xp5_ASAP7_75t_L     g10817(.A1(new_n3248), .A2(new_n2852), .B1(new_n2650), .B2(new_n3492), .C(new_n11073), .Y(new_n11074));
  XNOR2x2_ASAP7_75t_L       g10818(.A(\a[32] ), .B(new_n11074), .Y(new_n11075));
  INVx1_ASAP7_75t_L         g10819(.A(new_n11075), .Y(new_n11076));
  AOI21xp33_ASAP7_75t_L     g10820(.A1(new_n11072), .A2(new_n11070), .B(new_n11076), .Y(new_n11077));
  NOR3xp33_ASAP7_75t_L      g10821(.A(new_n10702), .B(new_n10700), .C(new_n10697), .Y(new_n11078));
  NOR3xp33_ASAP7_75t_L      g10822(.A(new_n11071), .B(new_n10720), .C(new_n11078), .Y(new_n11079));
  AOI21xp33_ASAP7_75t_L     g10823(.A1(new_n11067), .A2(new_n11063), .B(new_n11069), .Y(new_n11080));
  NOR3xp33_ASAP7_75t_L      g10824(.A(new_n11079), .B(new_n11080), .C(new_n11075), .Y(new_n11081));
  NOR2xp33_ASAP7_75t_L      g10825(.A(new_n11077), .B(new_n11081), .Y(new_n11082));
  NAND2xp33_ASAP7_75t_L     g10826(.A(new_n10931), .B(new_n11082), .Y(new_n11083));
  OAI21xp33_ASAP7_75t_L     g10827(.A1(new_n11080), .A2(new_n11079), .B(new_n11075), .Y(new_n11084));
  NAND3xp33_ASAP7_75t_L     g10828(.A(new_n11072), .B(new_n11076), .C(new_n11070), .Y(new_n11085));
  NAND2xp33_ASAP7_75t_L     g10829(.A(new_n11085), .B(new_n11084), .Y(new_n11086));
  A2O1A1Ixp33_ASAP7_75t_L   g10830(.A1(new_n10726), .A2(new_n10547), .B(new_n10930), .C(new_n11086), .Y(new_n11087));
  NAND3xp33_ASAP7_75t_L     g10831(.A(new_n11087), .B(new_n11083), .C(new_n10927), .Y(new_n11088));
  NAND2xp33_ASAP7_75t_L     g10832(.A(new_n10926), .B(new_n10925), .Y(new_n11089));
  A2O1A1Ixp33_ASAP7_75t_L   g10833(.A1(new_n10718), .A2(new_n10722), .B(new_n10725), .C(new_n10929), .Y(new_n11090));
  NOR2xp33_ASAP7_75t_L      g10834(.A(new_n11090), .B(new_n11086), .Y(new_n11091));
  NOR2xp33_ASAP7_75t_L      g10835(.A(new_n10931), .B(new_n11082), .Y(new_n11092));
  OAI21xp33_ASAP7_75t_L     g10836(.A1(new_n11091), .A2(new_n11092), .B(new_n11089), .Y(new_n11093));
  NAND3xp33_ASAP7_75t_L     g10837(.A(new_n10921), .B(new_n11093), .C(new_n11088), .Y(new_n11094));
  AO21x2_ASAP7_75t_L        g10838(.A1(new_n11088), .A2(new_n11093), .B(new_n10921), .Y(new_n11095));
  NAND2xp33_ASAP7_75t_L     g10839(.A(\b[33] ), .B(new_n2386), .Y(new_n11096));
  NAND2xp33_ASAP7_75t_L     g10840(.A(\b[34] ), .B(new_n2232), .Y(new_n11097));
  AOI22xp33_ASAP7_75t_L     g10841(.A1(new_n2228), .A2(\b[35] ), .B1(new_n2226), .B2(new_n5649), .Y(new_n11098));
  NAND4xp25_ASAP7_75t_L     g10842(.A(new_n11098), .B(\a[26] ), .C(new_n11096), .D(new_n11097), .Y(new_n11099));
  NAND2xp33_ASAP7_75t_L     g10843(.A(new_n11097), .B(new_n11098), .Y(new_n11100));
  A2O1A1Ixp33_ASAP7_75t_L   g10844(.A1(\b[33] ), .A2(new_n2386), .B(new_n11100), .C(new_n2223), .Y(new_n11101));
  NAND2xp33_ASAP7_75t_L     g10845(.A(new_n11099), .B(new_n11101), .Y(new_n11102));
  INVx1_ASAP7_75t_L         g10846(.A(new_n11102), .Y(new_n11103));
  NAND3xp33_ASAP7_75t_L     g10847(.A(new_n11095), .B(new_n11103), .C(new_n11094), .Y(new_n11104));
  AND3x1_ASAP7_75t_L        g10848(.A(new_n10921), .B(new_n11093), .C(new_n11088), .Y(new_n11105));
  AOI21xp33_ASAP7_75t_L     g10849(.A1(new_n11093), .A2(new_n11088), .B(new_n10921), .Y(new_n11106));
  OAI21xp33_ASAP7_75t_L     g10850(.A1(new_n11106), .A2(new_n11105), .B(new_n11102), .Y(new_n11107));
  NAND2xp33_ASAP7_75t_L     g10851(.A(new_n11104), .B(new_n11107), .Y(new_n11108));
  NOR2xp33_ASAP7_75t_L      g10852(.A(new_n10752), .B(new_n10751), .Y(new_n11109));
  MAJx2_ASAP7_75t_L         g10853(.A(new_n10758), .B(new_n10753), .C(new_n11109), .Y(new_n11110));
  NOR2xp33_ASAP7_75t_L      g10854(.A(new_n11108), .B(new_n11110), .Y(new_n11111));
  MAJIxp5_ASAP7_75t_L       g10855(.A(new_n10758), .B(new_n10753), .C(new_n11109), .Y(new_n11112));
  AOI21xp33_ASAP7_75t_L     g10856(.A1(new_n11107), .A2(new_n11104), .B(new_n11112), .Y(new_n11113));
  NAND2xp33_ASAP7_75t_L     g10857(.A(\b[37] ), .B(new_n1770), .Y(new_n11114));
  AOI22xp33_ASAP7_75t_L     g10858(.A1(new_n1766), .A2(\b[38] ), .B1(new_n1764), .B2(new_n4923), .Y(new_n11115));
  NAND2xp33_ASAP7_75t_L     g10859(.A(new_n11114), .B(new_n11115), .Y(new_n11116));
  AOI21xp33_ASAP7_75t_L     g10860(.A1(new_n1910), .A2(\b[36] ), .B(new_n11116), .Y(new_n11117));
  NAND2xp33_ASAP7_75t_L     g10861(.A(\a[23] ), .B(new_n11117), .Y(new_n11118));
  A2O1A1Ixp33_ASAP7_75t_L   g10862(.A1(\b[36] ), .A2(new_n1910), .B(new_n11116), .C(new_n1761), .Y(new_n11119));
  NAND2xp33_ASAP7_75t_L     g10863(.A(new_n11119), .B(new_n11118), .Y(new_n11120));
  NOR3xp33_ASAP7_75t_L      g10864(.A(new_n11111), .B(new_n11113), .C(new_n11120), .Y(new_n11121));
  AND2x2_ASAP7_75t_L        g10865(.A(new_n11104), .B(new_n11107), .Y(new_n11122));
  NAND2xp33_ASAP7_75t_L     g10866(.A(new_n11112), .B(new_n11122), .Y(new_n11123));
  NAND2xp33_ASAP7_75t_L     g10867(.A(new_n11108), .B(new_n11110), .Y(new_n11124));
  AND2x2_ASAP7_75t_L        g10868(.A(new_n11119), .B(new_n11118), .Y(new_n11125));
  AOI21xp33_ASAP7_75t_L     g10869(.A1(new_n11123), .A2(new_n11124), .B(new_n11125), .Y(new_n11126));
  NAND2xp33_ASAP7_75t_L     g10870(.A(new_n10756), .B(new_n10759), .Y(new_n11127));
  MAJIxp5_ASAP7_75t_L       g10871(.A(new_n10766), .B(new_n10762), .C(new_n11127), .Y(new_n11128));
  NOR3xp33_ASAP7_75t_L      g10872(.A(new_n11128), .B(new_n11126), .C(new_n11121), .Y(new_n11129));
  OA21x2_ASAP7_75t_L        g10873(.A1(new_n11121), .A2(new_n11126), .B(new_n11128), .Y(new_n11130));
  NAND2xp33_ASAP7_75t_L     g10874(.A(\b[39] ), .B(new_n1548), .Y(new_n11131));
  NAND2xp33_ASAP7_75t_L     g10875(.A(\b[40] ), .B(new_n1410), .Y(new_n11132));
  AOI22xp33_ASAP7_75t_L     g10876(.A1(new_n1406), .A2(\b[41] ), .B1(new_n1404), .B2(new_n5669), .Y(new_n11133));
  NAND4xp25_ASAP7_75t_L     g10877(.A(new_n11133), .B(\a[20] ), .C(new_n11131), .D(new_n11132), .Y(new_n11134));
  NAND2xp33_ASAP7_75t_L     g10878(.A(new_n11132), .B(new_n11133), .Y(new_n11135));
  A2O1A1Ixp33_ASAP7_75t_L   g10879(.A1(\b[39] ), .A2(new_n1548), .B(new_n11135), .C(new_n1401), .Y(new_n11136));
  NAND2xp33_ASAP7_75t_L     g10880(.A(new_n11134), .B(new_n11136), .Y(new_n11137));
  INVx1_ASAP7_75t_L         g10881(.A(new_n11137), .Y(new_n11138));
  OAI21xp33_ASAP7_75t_L     g10882(.A1(new_n11129), .A2(new_n11130), .B(new_n11138), .Y(new_n11139));
  OR3x1_ASAP7_75t_L         g10883(.A(new_n11128), .B(new_n11121), .C(new_n11126), .Y(new_n11140));
  OAI21xp33_ASAP7_75t_L     g10884(.A1(new_n11121), .A2(new_n11126), .B(new_n11128), .Y(new_n11141));
  NAND3xp33_ASAP7_75t_L     g10885(.A(new_n11140), .B(new_n11141), .C(new_n11137), .Y(new_n11142));
  NAND2xp33_ASAP7_75t_L     g10886(.A(new_n11139), .B(new_n11142), .Y(new_n11143));
  NOR2xp33_ASAP7_75t_L      g10887(.A(new_n10920), .B(new_n11143), .Y(new_n11144));
  AOI21xp33_ASAP7_75t_L     g10888(.A1(new_n11140), .A2(new_n11141), .B(new_n11137), .Y(new_n11145));
  NOR3xp33_ASAP7_75t_L      g10889(.A(new_n11130), .B(new_n11138), .C(new_n11129), .Y(new_n11146));
  NOR2xp33_ASAP7_75t_L      g10890(.A(new_n11146), .B(new_n11145), .Y(new_n11147));
  A2O1A1O1Ixp25_ASAP7_75t_L g10891(.A1(new_n10425), .A2(new_n10782), .B(new_n10787), .C(new_n10919), .D(new_n11147), .Y(new_n11148));
  OAI21xp33_ASAP7_75t_L     g10892(.A1(new_n11144), .A2(new_n11148), .B(new_n10917), .Y(new_n11149));
  INVx1_ASAP7_75t_L         g10893(.A(new_n10917), .Y(new_n11150));
  O2A1O1Ixp33_ASAP7_75t_L   g10894(.A1(new_n10785), .A2(new_n10786), .B(new_n10783), .C(new_n10918), .Y(new_n11151));
  NAND2xp33_ASAP7_75t_L     g10895(.A(new_n11151), .B(new_n11147), .Y(new_n11152));
  A2O1A1Ixp33_ASAP7_75t_L   g10896(.A1(new_n10783), .A2(new_n10780), .B(new_n10918), .C(new_n11143), .Y(new_n11153));
  NAND3xp33_ASAP7_75t_L     g10897(.A(new_n11153), .B(new_n11152), .C(new_n11150), .Y(new_n11154));
  A2O1A1Ixp33_ASAP7_75t_L   g10898(.A1(new_n10438), .A2(new_n10226), .B(new_n10437), .C(new_n10796), .Y(new_n11155));
  NAND2xp33_ASAP7_75t_L     g10899(.A(new_n10799), .B(new_n11155), .Y(new_n11156));
  NAND3xp33_ASAP7_75t_L     g10900(.A(new_n11156), .B(new_n11154), .C(new_n11149), .Y(new_n11157));
  AOI21xp33_ASAP7_75t_L     g10901(.A1(new_n11153), .A2(new_n11152), .B(new_n11150), .Y(new_n11158));
  NOR3xp33_ASAP7_75t_L      g10902(.A(new_n11148), .B(new_n11144), .C(new_n10917), .Y(new_n11159));
  INVx1_ASAP7_75t_L         g10903(.A(new_n10799), .Y(new_n11160));
  A2O1A1O1Ixp25_ASAP7_75t_L g10904(.A1(new_n10226), .A2(new_n10438), .B(new_n10437), .C(new_n10796), .D(new_n11160), .Y(new_n11161));
  OAI21xp33_ASAP7_75t_L     g10905(.A1(new_n11158), .A2(new_n11159), .B(new_n11161), .Y(new_n11162));
  NAND3xp33_ASAP7_75t_L     g10906(.A(new_n11157), .B(new_n11162), .C(new_n10911), .Y(new_n11163));
  NOR3xp33_ASAP7_75t_L      g10907(.A(new_n11161), .B(new_n11159), .C(new_n11158), .Y(new_n11164));
  AOI21xp33_ASAP7_75t_L     g10908(.A1(new_n11154), .A2(new_n11149), .B(new_n11156), .Y(new_n11165));
  OAI21xp33_ASAP7_75t_L     g10909(.A1(new_n11164), .A2(new_n11165), .B(new_n10910), .Y(new_n11166));
  NAND3xp33_ASAP7_75t_L     g10910(.A(new_n10903), .B(new_n11166), .C(new_n11163), .Y(new_n11167));
  NAND2xp33_ASAP7_75t_L     g10911(.A(new_n10456), .B(new_n10457), .Y(new_n11168));
  A2O1A1Ixp33_ASAP7_75t_L   g10912(.A1(new_n9475), .A2(new_n9228), .B(new_n9486), .C(new_n9806), .Y(new_n11169));
  A2O1A1Ixp33_ASAP7_75t_L   g10913(.A1(new_n11169), .A2(new_n9807), .B(new_n10139), .C(new_n10152), .Y(new_n11170));
  A2O1A1O1Ixp25_ASAP7_75t_L g10914(.A1(new_n11170), .A2(new_n11168), .B(new_n10536), .C(new_n10810), .D(new_n10808), .Y(new_n11171));
  NOR3xp33_ASAP7_75t_L      g10915(.A(new_n11165), .B(new_n11164), .C(new_n10910), .Y(new_n11172));
  AOI21xp33_ASAP7_75t_L     g10916(.A1(new_n11157), .A2(new_n11162), .B(new_n10911), .Y(new_n11173));
  OAI21xp33_ASAP7_75t_L     g10917(.A1(new_n11173), .A2(new_n11172), .B(new_n11171), .Y(new_n11174));
  NAND2xp33_ASAP7_75t_L     g10918(.A(\b[49] ), .B(new_n590), .Y(new_n11175));
  AOI22xp33_ASAP7_75t_L     g10919(.A1(new_n600), .A2(\b[50] ), .B1(new_n597), .B2(new_n8235), .Y(new_n11176));
  NAND2xp33_ASAP7_75t_L     g10920(.A(new_n11175), .B(new_n11176), .Y(new_n11177));
  AOI21xp33_ASAP7_75t_L     g10921(.A1(new_n674), .A2(\b[48] ), .B(new_n11177), .Y(new_n11178));
  NAND2xp33_ASAP7_75t_L     g10922(.A(\a[11] ), .B(new_n11178), .Y(new_n11179));
  A2O1A1Ixp33_ASAP7_75t_L   g10923(.A1(\b[48] ), .A2(new_n674), .B(new_n11177), .C(new_n594), .Y(new_n11180));
  AND2x2_ASAP7_75t_L        g10924(.A(new_n11180), .B(new_n11179), .Y(new_n11181));
  NAND3xp33_ASAP7_75t_L     g10925(.A(new_n11174), .B(new_n11167), .C(new_n11181), .Y(new_n11182));
  AO21x2_ASAP7_75t_L        g10926(.A1(new_n11167), .A2(new_n11174), .B(new_n11181), .Y(new_n11183));
  AO21x2_ASAP7_75t_L        g10927(.A1(new_n11183), .A2(new_n11182), .B(new_n10902), .Y(new_n11184));
  NAND3xp33_ASAP7_75t_L     g10928(.A(new_n10902), .B(new_n11183), .C(new_n11182), .Y(new_n11185));
  AOI21xp33_ASAP7_75t_L     g10929(.A1(new_n11184), .A2(new_n11185), .B(new_n10901), .Y(new_n11186));
  AOI21xp33_ASAP7_75t_L     g10930(.A1(new_n11183), .A2(new_n11182), .B(new_n10902), .Y(new_n11187));
  AND3x1_ASAP7_75t_L        g10931(.A(new_n10902), .B(new_n11183), .C(new_n11182), .Y(new_n11188));
  NOR3xp33_ASAP7_75t_L      g10932(.A(new_n11188), .B(new_n11187), .C(new_n10900), .Y(new_n11189));
  NOR3xp33_ASAP7_75t_L      g10933(.A(new_n10894), .B(new_n11186), .C(new_n11189), .Y(new_n11190));
  INVx1_ASAP7_75t_L         g10934(.A(new_n10831), .Y(new_n11191));
  OAI21xp33_ASAP7_75t_L     g10935(.A1(new_n10474), .A2(new_n10471), .B(new_n11191), .Y(new_n11192));
  OAI21xp33_ASAP7_75t_L     g10936(.A1(new_n11187), .A2(new_n11188), .B(new_n10900), .Y(new_n11193));
  NAND3xp33_ASAP7_75t_L     g10937(.A(new_n11184), .B(new_n10901), .C(new_n11185), .Y(new_n11194));
  AOI221xp5_ASAP7_75t_L     g10938(.A1(new_n11194), .A2(new_n11193), .B1(new_n10837), .B2(new_n11192), .C(new_n10829), .Y(new_n11195));
  NAND2xp33_ASAP7_75t_L     g10939(.A(\b[56] ), .B(new_n345), .Y(new_n11196));
  OAI221xp5_ASAP7_75t_L     g10940(.A1(new_n9534), .A2(new_n406), .B1(new_n367), .B2(new_n10184), .C(new_n11196), .Y(new_n11197));
  AOI21xp33_ASAP7_75t_L     g10941(.A1(new_n366), .A2(\b[54] ), .B(new_n11197), .Y(new_n11198));
  NAND2xp33_ASAP7_75t_L     g10942(.A(\a[5] ), .B(new_n11198), .Y(new_n11199));
  A2O1A1Ixp33_ASAP7_75t_L   g10943(.A1(\b[54] ), .A2(new_n366), .B(new_n11197), .C(new_n339), .Y(new_n11200));
  NAND2xp33_ASAP7_75t_L     g10944(.A(new_n11200), .B(new_n11199), .Y(new_n11201));
  OAI21xp33_ASAP7_75t_L     g10945(.A1(new_n11195), .A2(new_n11190), .B(new_n11201), .Y(new_n11202));
  OAI21xp33_ASAP7_75t_L     g10946(.A1(new_n10828), .A2(new_n10518), .B(new_n10833), .Y(new_n11203));
  NOR2xp33_ASAP7_75t_L      g10947(.A(new_n11186), .B(new_n11189), .Y(new_n11204));
  NAND2xp33_ASAP7_75t_L     g10948(.A(new_n11203), .B(new_n11204), .Y(new_n11205));
  OAI21xp33_ASAP7_75t_L     g10949(.A1(new_n11186), .A2(new_n11189), .B(new_n10894), .Y(new_n11206));
  NAND4xp25_ASAP7_75t_L     g10950(.A(new_n11205), .B(new_n11200), .C(new_n11199), .D(new_n11206), .Y(new_n11207));
  NAND3xp33_ASAP7_75t_L     g10951(.A(new_n11207), .B(new_n11202), .C(new_n10893), .Y(new_n11208));
  INVx1_ASAP7_75t_L         g10952(.A(new_n10893), .Y(new_n11209));
  OA21x2_ASAP7_75t_L        g10953(.A1(new_n11195), .A2(new_n11190), .B(new_n11201), .Y(new_n11210));
  NOR3xp33_ASAP7_75t_L      g10954(.A(new_n11190), .B(new_n11195), .C(new_n11201), .Y(new_n11211));
  OAI21xp33_ASAP7_75t_L     g10955(.A1(new_n11211), .A2(new_n11210), .B(new_n11209), .Y(new_n11212));
  NAND3xp33_ASAP7_75t_L     g10956(.A(new_n10879), .B(new_n11212), .C(new_n11208), .Y(new_n11213));
  AOI21xp33_ASAP7_75t_L     g10957(.A1(new_n10509), .A2(new_n10835), .B(new_n10843), .Y(new_n11214));
  NOR3xp33_ASAP7_75t_L      g10958(.A(new_n11210), .B(new_n11211), .C(new_n11209), .Y(new_n11215));
  AOI21xp33_ASAP7_75t_L     g10959(.A1(new_n11207), .A2(new_n11202), .B(new_n10893), .Y(new_n11216));
  OAI21xp33_ASAP7_75t_L     g10960(.A1(new_n11216), .A2(new_n11215), .B(new_n11214), .Y(new_n11217));
  NAND2xp33_ASAP7_75t_L     g10961(.A(new_n11213), .B(new_n11217), .Y(new_n11218));
  XOR2x2_ASAP7_75t_L        g10962(.A(new_n11218), .B(new_n10878), .Y(\f[59] ));
  NOR2xp33_ASAP7_75t_L      g10963(.A(new_n11216), .B(new_n11215), .Y(new_n11220));
  NOR2xp33_ASAP7_75t_L      g10964(.A(new_n10863), .B(new_n10877), .Y(new_n11221));
  A2O1A1Ixp33_ASAP7_75t_L   g10965(.A1(new_n10871), .A2(new_n10874), .B(new_n11221), .C(new_n11218), .Y(new_n11222));
  O2A1O1Ixp33_ASAP7_75t_L   g10966(.A1(new_n10489), .A2(new_n10492), .B(new_n10850), .C(new_n10849), .Y(new_n11223));
  INVx1_ASAP7_75t_L         g10967(.A(new_n10882), .Y(new_n11224));
  NOR2xp33_ASAP7_75t_L      g10968(.A(\b[59] ), .B(\b[60] ), .Y(new_n11225));
  INVx1_ASAP7_75t_L         g10969(.A(\b[60] ), .Y(new_n11226));
  NOR2xp33_ASAP7_75t_L      g10970(.A(new_n10881), .B(new_n11226), .Y(new_n11227));
  NOR2xp33_ASAP7_75t_L      g10971(.A(new_n11225), .B(new_n11227), .Y(new_n11228));
  INVx1_ASAP7_75t_L         g10972(.A(new_n11228), .Y(new_n11229));
  O2A1O1Ixp33_ASAP7_75t_L   g10973(.A1(new_n10880), .A2(new_n11223), .B(new_n11224), .C(new_n11229), .Y(new_n11230));
  A2O1A1O1Ixp25_ASAP7_75t_L g10974(.A1(new_n10850), .A2(new_n10853), .B(new_n10849), .C(new_n10883), .D(new_n10882), .Y(new_n11231));
  NAND2xp33_ASAP7_75t_L     g10975(.A(new_n11229), .B(new_n11231), .Y(new_n11232));
  INVx1_ASAP7_75t_L         g10976(.A(new_n11232), .Y(new_n11233));
  NOR2xp33_ASAP7_75t_L      g10977(.A(new_n11230), .B(new_n11233), .Y(new_n11234));
  NOR2xp33_ASAP7_75t_L      g10978(.A(new_n10881), .B(new_n261), .Y(new_n11235));
  AOI221xp5_ASAP7_75t_L     g10979(.A1(\b[58] ), .A2(new_n291), .B1(\b[60] ), .B2(new_n272), .C(new_n11235), .Y(new_n11236));
  INVx1_ASAP7_75t_L         g10980(.A(new_n11236), .Y(new_n11237));
  AOI211xp5_ASAP7_75t_L     g10981(.A1(new_n11234), .A2(new_n269), .B(new_n11237), .C(new_n265), .Y(new_n11238));
  A2O1A1Ixp33_ASAP7_75t_L   g10982(.A1(new_n11234), .A2(new_n269), .B(new_n11237), .C(new_n265), .Y(new_n11239));
  INVx1_ASAP7_75t_L         g10983(.A(new_n11239), .Y(new_n11240));
  NOR2xp33_ASAP7_75t_L      g10984(.A(new_n11238), .B(new_n11240), .Y(new_n11241));
  INVx1_ASAP7_75t_L         g10985(.A(new_n11241), .Y(new_n11242));
  AOI22xp33_ASAP7_75t_L     g10986(.A1(new_n345), .A2(\b[57] ), .B1(new_n342), .B2(new_n10495), .Y(new_n11243));
  OAI221xp5_ASAP7_75t_L     g10987(.A1(new_n406), .A2(new_n10178), .B1(new_n9534), .B2(new_n365), .C(new_n11243), .Y(new_n11244));
  XNOR2x2_ASAP7_75t_L       g10988(.A(new_n339), .B(new_n11244), .Y(new_n11245));
  NAND3xp33_ASAP7_75t_L     g10989(.A(new_n11184), .B(new_n10900), .C(new_n11185), .Y(new_n11246));
  A2O1A1Ixp33_ASAP7_75t_L   g10990(.A1(new_n11193), .A2(new_n11194), .B(new_n10894), .C(new_n11246), .Y(new_n11247));
  NOR2xp33_ASAP7_75t_L      g10991(.A(new_n8569), .B(new_n481), .Y(new_n11248));
  INVx1_ASAP7_75t_L         g10992(.A(new_n11248), .Y(new_n11249));
  NAND2xp33_ASAP7_75t_L     g10993(.A(\b[53] ), .B(new_n441), .Y(new_n11250));
  AOI22xp33_ASAP7_75t_L     g10994(.A1(new_n451), .A2(\b[54] ), .B1(new_n448), .B2(new_n9208), .Y(new_n11251));
  AND4x1_ASAP7_75t_L        g10995(.A(new_n11251), .B(new_n11250), .C(new_n11249), .D(\a[8] ), .Y(new_n11252));
  AOI31xp33_ASAP7_75t_L     g10996(.A1(new_n11251), .A2(new_n11250), .A3(new_n11249), .B(\a[8] ), .Y(new_n11253));
  NOR2xp33_ASAP7_75t_L      g10997(.A(new_n11253), .B(new_n11252), .Y(new_n11254));
  INVx1_ASAP7_75t_L         g10998(.A(new_n11254), .Y(new_n11255));
  NAND2xp33_ASAP7_75t_L     g10999(.A(new_n11167), .B(new_n11174), .Y(new_n11256));
  MAJIxp5_ASAP7_75t_L       g11000(.A(new_n10902), .B(new_n11181), .C(new_n11256), .Y(new_n11257));
  NAND2xp33_ASAP7_75t_L     g11001(.A(\b[50] ), .B(new_n590), .Y(new_n11258));
  AOI22xp33_ASAP7_75t_L     g11002(.A1(new_n600), .A2(\b[51] ), .B1(new_n597), .B2(new_n8257), .Y(new_n11259));
  NAND2xp33_ASAP7_75t_L     g11003(.A(new_n11258), .B(new_n11259), .Y(new_n11260));
  AOI21xp33_ASAP7_75t_L     g11004(.A1(new_n674), .A2(\b[49] ), .B(new_n11260), .Y(new_n11261));
  NAND2xp33_ASAP7_75t_L     g11005(.A(\a[11] ), .B(new_n11261), .Y(new_n11262));
  A2O1A1Ixp33_ASAP7_75t_L   g11006(.A1(\b[49] ), .A2(new_n674), .B(new_n11260), .C(new_n594), .Y(new_n11263));
  NAND2xp33_ASAP7_75t_L     g11007(.A(new_n11263), .B(new_n11262), .Y(new_n11264));
  A2O1A1O1Ixp25_ASAP7_75t_L g11008(.A1(new_n10810), .A2(new_n10815), .B(new_n10808), .C(new_n11166), .D(new_n11172), .Y(new_n11265));
  NAND2xp33_ASAP7_75t_L     g11009(.A(\b[46] ), .B(new_n908), .Y(new_n11266));
  NAND2xp33_ASAP7_75t_L     g11010(.A(\b[47] ), .B(new_n817), .Y(new_n11267));
  AOI22xp33_ASAP7_75t_L     g11011(.A1(new_n826), .A2(\b[48] ), .B1(new_n823), .B2(new_n7341), .Y(new_n11268));
  AND4x1_ASAP7_75t_L        g11012(.A(new_n11268), .B(new_n11267), .C(new_n11266), .D(\a[14] ), .Y(new_n11269));
  AOI31xp33_ASAP7_75t_L     g11013(.A1(new_n11268), .A2(new_n11267), .A3(new_n11266), .B(\a[14] ), .Y(new_n11270));
  NOR2xp33_ASAP7_75t_L      g11014(.A(new_n11270), .B(new_n11269), .Y(new_n11271));
  INVx1_ASAP7_75t_L         g11015(.A(new_n11271), .Y(new_n11272));
  A2O1A1O1Ixp25_ASAP7_75t_L g11016(.A1(new_n10796), .A2(new_n10544), .B(new_n11160), .C(new_n11154), .D(new_n11158), .Y(new_n11273));
  NAND2xp33_ASAP7_75t_L     g11017(.A(new_n1110), .B(new_n6764), .Y(new_n11274));
  OAI221xp5_ASAP7_75t_L     g11018(.A1(new_n1198), .A2(new_n6756), .B1(new_n6220), .B2(new_n1298), .C(new_n11274), .Y(new_n11275));
  AOI21xp33_ASAP7_75t_L     g11019(.A1(new_n1194), .A2(\b[43] ), .B(new_n11275), .Y(new_n11276));
  NAND2xp33_ASAP7_75t_L     g11020(.A(\a[17] ), .B(new_n11276), .Y(new_n11277));
  A2O1A1Ixp33_ASAP7_75t_L   g11021(.A1(\b[43] ), .A2(new_n1194), .B(new_n11275), .C(new_n1107), .Y(new_n11278));
  AND2x2_ASAP7_75t_L        g11022(.A(new_n11278), .B(new_n11277), .Y(new_n11279));
  NOR3xp33_ASAP7_75t_L      g11023(.A(new_n11105), .B(new_n11106), .C(new_n11103), .Y(new_n11280));
  INVx1_ASAP7_75t_L         g11024(.A(new_n11280), .Y(new_n11281));
  NAND2xp33_ASAP7_75t_L     g11025(.A(\b[34] ), .B(new_n2386), .Y(new_n11282));
  NAND2xp33_ASAP7_75t_L     g11026(.A(\b[35] ), .B(new_n2232), .Y(new_n11283));
  AOI22xp33_ASAP7_75t_L     g11027(.A1(new_n2228), .A2(\b[36] ), .B1(new_n2226), .B2(new_n4473), .Y(new_n11284));
  AND4x1_ASAP7_75t_L        g11028(.A(new_n11284), .B(new_n11283), .C(new_n11282), .D(\a[26] ), .Y(new_n11285));
  AOI31xp33_ASAP7_75t_L     g11029(.A1(new_n11284), .A2(new_n11283), .A3(new_n11282), .B(\a[26] ), .Y(new_n11286));
  NOR2xp33_ASAP7_75t_L      g11030(.A(new_n11286), .B(new_n11285), .Y(new_n11287));
  AOI21xp33_ASAP7_75t_L     g11031(.A1(new_n11087), .A2(new_n11083), .B(new_n10927), .Y(new_n11288));
  A2O1A1O1Ixp25_ASAP7_75t_L g11032(.A1(new_n10740), .A2(new_n10742), .B(new_n10734), .C(new_n11088), .D(new_n11288), .Y(new_n11289));
  A2O1A1Ixp33_ASAP7_75t_L   g11033(.A1(new_n10338), .A2(new_n10330), .B(new_n10684), .C(new_n10671), .Y(new_n11290));
  A2O1A1Ixp33_ASAP7_75t_L   g11034(.A1(new_n10675), .A2(new_n11290), .B(new_n11045), .C(new_n11038), .Y(new_n11291));
  NAND2xp33_ASAP7_75t_L     g11035(.A(\b[19] ), .B(new_n5526), .Y(new_n11292));
  NAND2xp33_ASAP7_75t_L     g11036(.A(\b[20] ), .B(new_n5240), .Y(new_n11293));
  AOI22xp33_ASAP7_75t_L     g11037(.A1(new_n5249), .A2(\b[21] ), .B1(new_n5247), .B2(new_n1715), .Y(new_n11294));
  NAND4xp25_ASAP7_75t_L     g11038(.A(new_n11294), .B(\a[41] ), .C(new_n11292), .D(new_n11293), .Y(new_n11295));
  NAND2xp33_ASAP7_75t_L     g11039(.A(new_n11293), .B(new_n11294), .Y(new_n11296));
  A2O1A1Ixp33_ASAP7_75t_L   g11040(.A1(\b[19] ), .A2(new_n5526), .B(new_n11296), .C(new_n5244), .Y(new_n11297));
  NAND2xp33_ASAP7_75t_L     g11041(.A(new_n11295), .B(new_n11297), .Y(new_n11298));
  NOR3xp33_ASAP7_75t_L      g11042(.A(new_n11024), .B(new_n11029), .C(new_n10948), .Y(new_n11299));
  INVx1_ASAP7_75t_L         g11043(.A(new_n11299), .Y(new_n11300));
  A2O1A1Ixp33_ASAP7_75t_L   g11044(.A1(new_n11030), .A2(new_n11033), .B(new_n11036), .C(new_n11300), .Y(new_n11301));
  AOI22xp33_ASAP7_75t_L     g11045(.A1(new_n6002), .A2(\b[18] ), .B1(new_n5999), .B2(new_n1363), .Y(new_n11302));
  OAI221xp5_ASAP7_75t_L     g11046(.A1(new_n6544), .A2(new_n1244), .B1(new_n1051), .B2(new_n6309), .C(new_n11302), .Y(new_n11303));
  XNOR2x2_ASAP7_75t_L       g11047(.A(\a[44] ), .B(new_n11303), .Y(new_n11304));
  NOR3xp33_ASAP7_75t_L      g11048(.A(new_n11018), .B(new_n11016), .C(new_n11019), .Y(new_n11305));
  INVx1_ASAP7_75t_L         g11049(.A(new_n11305), .Y(new_n11306));
  A2O1A1Ixp33_ASAP7_75t_L   g11050(.A1(new_n11021), .A2(new_n11017), .B(new_n11023), .C(new_n11306), .Y(new_n11307));
  NAND2xp33_ASAP7_75t_L     g11051(.A(\b[13] ), .B(new_n7124), .Y(new_n11308));
  NAND2xp33_ASAP7_75t_L     g11052(.A(\b[14] ), .B(new_n6812), .Y(new_n11309));
  AOI22xp33_ASAP7_75t_L     g11053(.A1(new_n6822), .A2(\b[15] ), .B1(new_n6819), .B2(new_n959), .Y(new_n11310));
  NAND4xp25_ASAP7_75t_L     g11054(.A(new_n11310), .B(\a[47] ), .C(new_n11308), .D(new_n11309), .Y(new_n11311));
  NAND2xp33_ASAP7_75t_L     g11055(.A(new_n11309), .B(new_n11310), .Y(new_n11312));
  A2O1A1Ixp33_ASAP7_75t_L   g11056(.A1(\b[13] ), .A2(new_n7124), .B(new_n11312), .C(new_n6816), .Y(new_n11313));
  NAND2xp33_ASAP7_75t_L     g11057(.A(new_n11311), .B(new_n11313), .Y(new_n11314));
  NAND2xp33_ASAP7_75t_L     g11058(.A(new_n10622), .B(new_n11006), .Y(new_n11315));
  A2O1A1Ixp33_ASAP7_75t_L   g11059(.A1(new_n10644), .A2(new_n11315), .B(new_n11008), .C(new_n11004), .Y(new_n11316));
  AOI22xp33_ASAP7_75t_L     g11060(.A1(new_n7659), .A2(\b[12] ), .B1(new_n7656), .B2(new_n970), .Y(new_n11317));
  OAI221xp5_ASAP7_75t_L     g11061(.A1(new_n8326), .A2(new_n695), .B1(new_n631), .B2(new_n7994), .C(new_n11317), .Y(new_n11318));
  NOR2xp33_ASAP7_75t_L      g11062(.A(new_n7653), .B(new_n11318), .Y(new_n11319));
  INVx1_ASAP7_75t_L         g11063(.A(new_n11319), .Y(new_n11320));
  NAND2xp33_ASAP7_75t_L     g11064(.A(new_n7653), .B(new_n11318), .Y(new_n11321));
  A2O1A1O1Ixp25_ASAP7_75t_L g11065(.A1(new_n10613), .A2(new_n10612), .B(new_n10609), .C(new_n10997), .D(new_n10994), .Y(new_n11322));
  INVx1_ASAP7_75t_L         g11066(.A(\a[60] ), .Y(new_n11323));
  NAND2xp33_ASAP7_75t_L     g11067(.A(\a[59] ), .B(new_n11323), .Y(new_n11324));
  NAND2xp33_ASAP7_75t_L     g11068(.A(\a[60] ), .B(new_n10588), .Y(new_n11325));
  AND2x2_ASAP7_75t_L        g11069(.A(new_n11324), .B(new_n11325), .Y(new_n11326));
  NOR2xp33_ASAP7_75t_L      g11070(.A(new_n258), .B(new_n11326), .Y(new_n11327));
  INVx1_ASAP7_75t_L         g11071(.A(new_n11327), .Y(new_n11328));
  NAND3xp33_ASAP7_75t_L     g11072(.A(new_n10592), .B(new_n10595), .C(new_n10585), .Y(new_n11329));
  INVx1_ASAP7_75t_L         g11073(.A(new_n10973), .Y(new_n11330));
  NOR2xp33_ASAP7_75t_L      g11074(.A(new_n258), .B(new_n11330), .Y(new_n11331));
  NOR5xp2_ASAP7_75t_L       g11075(.A(new_n11329), .B(new_n11331), .C(new_n10977), .D(new_n10276), .E(new_n10588), .Y(new_n11332));
  NOR2xp33_ASAP7_75t_L      g11076(.A(new_n11328), .B(new_n11332), .Y(new_n11333));
  AND2x2_ASAP7_75t_L        g11077(.A(new_n11328), .B(new_n11332), .Y(new_n11334));
  INVx1_ASAP7_75t_L         g11078(.A(new_n10584), .Y(new_n11335));
  NAND2xp33_ASAP7_75t_L     g11079(.A(\b[3] ), .B(new_n10594), .Y(new_n11336));
  OAI221xp5_ASAP7_75t_L     g11080(.A1(new_n278), .A2(new_n11335), .B1(new_n10974), .B2(new_n303), .C(new_n11336), .Y(new_n11337));
  AOI21xp33_ASAP7_75t_L     g11081(.A1(new_n10973), .A2(\b[1] ), .B(new_n11337), .Y(new_n11338));
  NAND2xp33_ASAP7_75t_L     g11082(.A(\a[59] ), .B(new_n11338), .Y(new_n11339));
  A2O1A1Ixp33_ASAP7_75t_L   g11083(.A1(\b[1] ), .A2(new_n10973), .B(new_n11337), .C(new_n10588), .Y(new_n11340));
  NAND2xp33_ASAP7_75t_L     g11084(.A(new_n11340), .B(new_n11339), .Y(new_n11341));
  OAI21xp33_ASAP7_75t_L     g11085(.A1(new_n11333), .A2(new_n11334), .B(new_n11341), .Y(new_n11342));
  INVx1_ASAP7_75t_L         g11086(.A(new_n11333), .Y(new_n11343));
  A2O1A1Ixp33_ASAP7_75t_L   g11087(.A1(new_n11324), .A2(new_n11325), .B(new_n258), .C(new_n11332), .Y(new_n11344));
  AND2x2_ASAP7_75t_L        g11088(.A(new_n11340), .B(new_n11339), .Y(new_n11345));
  NAND3xp33_ASAP7_75t_L     g11089(.A(new_n11345), .B(new_n11343), .C(new_n11344), .Y(new_n11346));
  NAND2xp33_ASAP7_75t_L     g11090(.A(\b[4] ), .B(new_n9948), .Y(new_n11347));
  NAND2xp33_ASAP7_75t_L     g11091(.A(\b[5] ), .B(new_n9614), .Y(new_n11348));
  AOI22xp33_ASAP7_75t_L     g11092(.A1(new_n9623), .A2(\b[6] ), .B1(new_n9620), .B2(new_n389), .Y(new_n11349));
  NAND4xp25_ASAP7_75t_L     g11093(.A(new_n11349), .B(\a[56] ), .C(new_n11347), .D(new_n11348), .Y(new_n11350));
  NAND2xp33_ASAP7_75t_L     g11094(.A(new_n11348), .B(new_n11349), .Y(new_n11351));
  A2O1A1Ixp33_ASAP7_75t_L   g11095(.A1(\b[4] ), .A2(new_n9948), .B(new_n11351), .C(new_n9610), .Y(new_n11352));
  AND4x1_ASAP7_75t_L        g11096(.A(new_n11346), .B(new_n11342), .C(new_n11352), .D(new_n11350), .Y(new_n11353));
  AOI22xp33_ASAP7_75t_L     g11097(.A1(new_n11350), .A2(new_n11352), .B1(new_n11342), .B2(new_n11346), .Y(new_n11354));
  NOR2xp33_ASAP7_75t_L      g11098(.A(new_n11354), .B(new_n11353), .Y(new_n11355));
  NOR3xp33_ASAP7_75t_L      g11099(.A(new_n10985), .B(new_n10970), .C(new_n10984), .Y(new_n11356));
  A2O1A1Ixp33_ASAP7_75t_L   g11100(.A1(new_n10600), .A2(new_n10599), .B(new_n11356), .C(new_n10986), .Y(new_n11357));
  NAND2xp33_ASAP7_75t_L     g11101(.A(new_n11357), .B(new_n11355), .Y(new_n11358));
  OA21x2_ASAP7_75t_L        g11102(.A1(new_n11356), .A2(new_n10965), .B(new_n10986), .Y(new_n11359));
  OAI21xp33_ASAP7_75t_L     g11103(.A1(new_n11353), .A2(new_n11354), .B(new_n11359), .Y(new_n11360));
  NAND2xp33_ASAP7_75t_L     g11104(.A(\b[9] ), .B(new_n8645), .Y(new_n11361));
  OAI221xp5_ASAP7_75t_L     g11105(.A1(new_n503), .A2(new_n9322), .B1(new_n8967), .B2(new_n978), .C(new_n11361), .Y(new_n11362));
  AOI21xp33_ASAP7_75t_L     g11106(.A1(new_n8964), .A2(\b[7] ), .B(new_n11362), .Y(new_n11363));
  NAND2xp33_ASAP7_75t_L     g11107(.A(\a[53] ), .B(new_n11363), .Y(new_n11364));
  A2O1A1Ixp33_ASAP7_75t_L   g11108(.A1(\b[7] ), .A2(new_n8964), .B(new_n11362), .C(new_n8639), .Y(new_n11365));
  AOI22xp33_ASAP7_75t_L     g11109(.A1(new_n11364), .A2(new_n11365), .B1(new_n11360), .B2(new_n11358), .Y(new_n11366));
  AND4x1_ASAP7_75t_L        g11110(.A(new_n11358), .B(new_n11365), .C(new_n11364), .D(new_n11360), .Y(new_n11367));
  NOR3xp33_ASAP7_75t_L      g11111(.A(new_n11322), .B(new_n11366), .C(new_n11367), .Y(new_n11368));
  A2O1A1Ixp33_ASAP7_75t_L   g11112(.A1(new_n10624), .A2(new_n10614), .B(new_n10990), .C(new_n10998), .Y(new_n11369));
  AO22x1_ASAP7_75t_L        g11113(.A1(new_n11365), .A2(new_n11364), .B1(new_n11360), .B2(new_n11358), .Y(new_n11370));
  NAND4xp25_ASAP7_75t_L     g11114(.A(new_n11358), .B(new_n11364), .C(new_n11365), .D(new_n11360), .Y(new_n11371));
  AOI21xp33_ASAP7_75t_L     g11115(.A1(new_n11371), .A2(new_n11370), .B(new_n11369), .Y(new_n11372));
  OAI211xp5_ASAP7_75t_L     g11116(.A1(new_n11368), .A2(new_n11372), .B(new_n11321), .C(new_n11320), .Y(new_n11373));
  INVx1_ASAP7_75t_L         g11117(.A(new_n11321), .Y(new_n11374));
  NAND3xp33_ASAP7_75t_L     g11118(.A(new_n11369), .B(new_n11370), .C(new_n11371), .Y(new_n11375));
  OAI21xp33_ASAP7_75t_L     g11119(.A1(new_n11366), .A2(new_n11367), .B(new_n11322), .Y(new_n11376));
  OAI211xp5_ASAP7_75t_L     g11120(.A1(new_n11374), .A2(new_n11319), .B(new_n11375), .C(new_n11376), .Y(new_n11377));
  NAND3xp33_ASAP7_75t_L     g11121(.A(new_n11316), .B(new_n11377), .C(new_n11373), .Y(new_n11378));
  A2O1A1O1Ixp25_ASAP7_75t_L g11122(.A1(new_n10622), .A2(new_n11006), .B(new_n10633), .C(new_n11000), .D(new_n11009), .Y(new_n11379));
  AOI211xp5_ASAP7_75t_L     g11123(.A1(new_n11375), .A2(new_n11376), .B(new_n11374), .C(new_n11319), .Y(new_n11380));
  AOI211xp5_ASAP7_75t_L     g11124(.A1(new_n11320), .A2(new_n11321), .B(new_n11368), .C(new_n11372), .Y(new_n11381));
  OAI21xp33_ASAP7_75t_L     g11125(.A1(new_n11381), .A2(new_n11380), .B(new_n11379), .Y(new_n11382));
  NAND3xp33_ASAP7_75t_L     g11126(.A(new_n11378), .B(new_n11382), .C(new_n11314), .Y(new_n11383));
  AO21x2_ASAP7_75t_L        g11127(.A1(new_n11382), .A2(new_n11378), .B(new_n11314), .Y(new_n11384));
  NAND3xp33_ASAP7_75t_L     g11128(.A(new_n11307), .B(new_n11383), .C(new_n11384), .Y(new_n11385));
  NAND2xp33_ASAP7_75t_L     g11129(.A(new_n11017), .B(new_n11021), .Y(new_n11386));
  O2A1O1Ixp33_ASAP7_75t_L   g11130(.A1(new_n11022), .A2(new_n11028), .B(new_n11386), .C(new_n11305), .Y(new_n11387));
  NAND2xp33_ASAP7_75t_L     g11131(.A(new_n11383), .B(new_n11384), .Y(new_n11388));
  NAND2xp33_ASAP7_75t_L     g11132(.A(new_n11387), .B(new_n11388), .Y(new_n11389));
  AOI21xp33_ASAP7_75t_L     g11133(.A1(new_n11389), .A2(new_n11385), .B(new_n11304), .Y(new_n11390));
  AND3x1_ASAP7_75t_L        g11134(.A(new_n11389), .B(new_n11385), .C(new_n11304), .Y(new_n11391));
  OAI21xp33_ASAP7_75t_L     g11135(.A1(new_n11390), .A2(new_n11391), .B(new_n11301), .Y(new_n11392));
  A2O1A1O1Ixp25_ASAP7_75t_L g11136(.A1(new_n10555), .A2(new_n10660), .B(new_n10655), .C(new_n11034), .D(new_n11299), .Y(new_n11393));
  AO21x2_ASAP7_75t_L        g11137(.A1(new_n11385), .A2(new_n11389), .B(new_n11304), .Y(new_n11394));
  NAND3xp33_ASAP7_75t_L     g11138(.A(new_n11389), .B(new_n11385), .C(new_n11304), .Y(new_n11395));
  NAND3xp33_ASAP7_75t_L     g11139(.A(new_n11393), .B(new_n11394), .C(new_n11395), .Y(new_n11396));
  NAND3xp33_ASAP7_75t_L     g11140(.A(new_n11396), .B(new_n11392), .C(new_n11298), .Y(new_n11397));
  INVx1_ASAP7_75t_L         g11141(.A(new_n11298), .Y(new_n11398));
  AOI21xp33_ASAP7_75t_L     g11142(.A1(new_n11395), .A2(new_n11394), .B(new_n11393), .Y(new_n11399));
  NOR3xp33_ASAP7_75t_L      g11143(.A(new_n11301), .B(new_n11391), .C(new_n11390), .Y(new_n11400));
  OAI21xp33_ASAP7_75t_L     g11144(.A1(new_n11400), .A2(new_n11399), .B(new_n11398), .Y(new_n11401));
  NAND3xp33_ASAP7_75t_L     g11145(.A(new_n11291), .B(new_n11397), .C(new_n11401), .Y(new_n11402));
  INVx1_ASAP7_75t_L         g11146(.A(new_n11038), .Y(new_n11403));
  A2O1A1O1Ixp25_ASAP7_75t_L g11147(.A1(new_n10671), .A2(new_n10554), .B(new_n10679), .C(new_n11042), .D(new_n11403), .Y(new_n11404));
  NAND2xp33_ASAP7_75t_L     g11148(.A(new_n11397), .B(new_n11401), .Y(new_n11405));
  NAND2xp33_ASAP7_75t_L     g11149(.A(new_n11404), .B(new_n11405), .Y(new_n11406));
  NOR2xp33_ASAP7_75t_L      g11150(.A(new_n2019), .B(new_n4550), .Y(new_n11407));
  AOI221xp5_ASAP7_75t_L     g11151(.A1(new_n4548), .A2(\b[23] ), .B1(new_n4542), .B2(new_n2027), .C(new_n11407), .Y(new_n11408));
  OA211x2_ASAP7_75t_L       g11152(.A1(new_n4781), .A2(new_n1857), .B(new_n11408), .C(\a[38] ), .Y(new_n11409));
  O2A1O1Ixp33_ASAP7_75t_L   g11153(.A1(new_n1857), .A2(new_n4781), .B(new_n11408), .C(\a[38] ), .Y(new_n11410));
  NOR2xp33_ASAP7_75t_L      g11154(.A(new_n11410), .B(new_n11409), .Y(new_n11411));
  NAND3xp33_ASAP7_75t_L     g11155(.A(new_n11402), .B(new_n11406), .C(new_n11411), .Y(new_n11412));
  NOR2xp33_ASAP7_75t_L      g11156(.A(new_n11404), .B(new_n11405), .Y(new_n11413));
  AOI21xp33_ASAP7_75t_L     g11157(.A1(new_n11401), .A2(new_n11397), .B(new_n11291), .Y(new_n11414));
  INVx1_ASAP7_75t_L         g11158(.A(new_n11411), .Y(new_n11415));
  OAI21xp33_ASAP7_75t_L     g11159(.A1(new_n11414), .A2(new_n11413), .B(new_n11415), .Y(new_n11416));
  A2O1A1O1Ixp25_ASAP7_75t_L g11160(.A1(new_n10688), .A2(new_n10699), .B(new_n10691), .C(new_n11051), .D(new_n11054), .Y(new_n11417));
  NAND3xp33_ASAP7_75t_L     g11161(.A(new_n11417), .B(new_n11416), .C(new_n11412), .Y(new_n11418));
  NAND2xp33_ASAP7_75t_L     g11162(.A(new_n11412), .B(new_n11416), .Y(new_n11419));
  OAI21xp33_ASAP7_75t_L     g11163(.A1(new_n11055), .A2(new_n10932), .B(new_n11048), .Y(new_n11420));
  NAND2xp33_ASAP7_75t_L     g11164(.A(new_n11420), .B(new_n11419), .Y(new_n11421));
  NAND2xp33_ASAP7_75t_L     g11165(.A(\b[26] ), .B(new_n3874), .Y(new_n11422));
  AOI22xp33_ASAP7_75t_L     g11166(.A1(new_n3884), .A2(\b[27] ), .B1(new_n3881), .B2(new_n2657), .Y(new_n11423));
  NAND2xp33_ASAP7_75t_L     g11167(.A(new_n11422), .B(new_n11423), .Y(new_n11424));
  AOI211xp5_ASAP7_75t_L     g11168(.A1(\b[25] ), .A2(new_n4111), .B(new_n3878), .C(new_n11424), .Y(new_n11425));
  INVx1_ASAP7_75t_L         g11169(.A(new_n11424), .Y(new_n11426));
  O2A1O1Ixp33_ASAP7_75t_L   g11170(.A1(new_n2180), .A2(new_n4986), .B(new_n11426), .C(\a[35] ), .Y(new_n11427));
  NOR2xp33_ASAP7_75t_L      g11171(.A(new_n11425), .B(new_n11427), .Y(new_n11428));
  NAND3xp33_ASAP7_75t_L     g11172(.A(new_n11421), .B(new_n11428), .C(new_n11418), .Y(new_n11429));
  NOR2xp33_ASAP7_75t_L      g11173(.A(new_n11420), .B(new_n11419), .Y(new_n11430));
  AOI21xp33_ASAP7_75t_L     g11174(.A1(new_n11416), .A2(new_n11412), .B(new_n11417), .Y(new_n11431));
  OR2x4_ASAP7_75t_L         g11175(.A(new_n11425), .B(new_n11427), .Y(new_n11432));
  OAI21xp33_ASAP7_75t_L     g11176(.A1(new_n11431), .A2(new_n11430), .B(new_n11432), .Y(new_n11433));
  NAND2xp33_ASAP7_75t_L     g11177(.A(new_n11429), .B(new_n11433), .Y(new_n11434));
  NAND3xp33_ASAP7_75t_L     g11178(.A(new_n11066), .B(new_n11057), .C(new_n11053), .Y(new_n11435));
  A2O1A1Ixp33_ASAP7_75t_L   g11179(.A1(new_n11067), .A2(new_n11063), .B(new_n11069), .C(new_n11435), .Y(new_n11436));
  NOR2xp33_ASAP7_75t_L      g11180(.A(new_n11434), .B(new_n11436), .Y(new_n11437));
  NAND2xp33_ASAP7_75t_L     g11181(.A(new_n11053), .B(new_n11057), .Y(new_n11438));
  NOR3xp33_ASAP7_75t_L      g11182(.A(new_n11432), .B(new_n11430), .C(new_n11431), .Y(new_n11439));
  AOI21xp33_ASAP7_75t_L     g11183(.A1(new_n11421), .A2(new_n11418), .B(new_n11428), .Y(new_n11440));
  NOR2xp33_ASAP7_75t_L      g11184(.A(new_n11440), .B(new_n11439), .Y(new_n11441));
  O2A1O1Ixp33_ASAP7_75t_L   g11185(.A1(new_n11438), .A2(new_n11062), .B(new_n11072), .C(new_n11441), .Y(new_n11442));
  NAND2xp33_ASAP7_75t_L     g11186(.A(new_n3254), .B(new_n3219), .Y(new_n11443));
  OAI221xp5_ASAP7_75t_L     g11187(.A1(new_n3262), .A2(new_n3212), .B1(new_n2871), .B2(new_n3248), .C(new_n11443), .Y(new_n11444));
  AOI21xp33_ASAP7_75t_L     g11188(.A1(new_n3491), .A2(\b[28] ), .B(new_n11444), .Y(new_n11445));
  NAND2xp33_ASAP7_75t_L     g11189(.A(\a[32] ), .B(new_n11445), .Y(new_n11446));
  A2O1A1Ixp33_ASAP7_75t_L   g11190(.A1(\b[28] ), .A2(new_n3491), .B(new_n11444), .C(new_n3251), .Y(new_n11447));
  NAND2xp33_ASAP7_75t_L     g11191(.A(new_n11447), .B(new_n11446), .Y(new_n11448));
  INVx1_ASAP7_75t_L         g11192(.A(new_n11448), .Y(new_n11449));
  OAI21xp33_ASAP7_75t_L     g11193(.A1(new_n11437), .A2(new_n11442), .B(new_n11449), .Y(new_n11450));
  NAND3xp33_ASAP7_75t_L     g11194(.A(new_n11441), .B(new_n11072), .C(new_n11435), .Y(new_n11451));
  NAND2xp33_ASAP7_75t_L     g11195(.A(new_n11434), .B(new_n11436), .Y(new_n11452));
  NAND3xp33_ASAP7_75t_L     g11196(.A(new_n11451), .B(new_n11452), .C(new_n11448), .Y(new_n11453));
  A2O1A1O1Ixp25_ASAP7_75t_L g11197(.A1(new_n10718), .A2(new_n10722), .B(new_n10725), .C(new_n10929), .D(new_n11077), .Y(new_n11454));
  OAI211xp5_ASAP7_75t_L     g11198(.A1(new_n11081), .A2(new_n11454), .B(new_n11450), .C(new_n11453), .Y(new_n11455));
  AOI21xp33_ASAP7_75t_L     g11199(.A1(new_n11451), .A2(new_n11452), .B(new_n11448), .Y(new_n11456));
  NOR3xp33_ASAP7_75t_L      g11200(.A(new_n11442), .B(new_n11449), .C(new_n11437), .Y(new_n11457));
  A2O1A1O1Ixp25_ASAP7_75t_L g11201(.A1(new_n10547), .A2(new_n10726), .B(new_n10930), .C(new_n11084), .D(new_n11081), .Y(new_n11458));
  OAI21xp33_ASAP7_75t_L     g11202(.A1(new_n11456), .A2(new_n11457), .B(new_n11458), .Y(new_n11459));
  NAND2xp33_ASAP7_75t_L     g11203(.A(\b[32] ), .B(new_n2706), .Y(new_n11460));
  AOI22xp33_ASAP7_75t_L     g11204(.A1(new_n2702), .A2(\b[33] ), .B1(new_n2700), .B2(new_n3813), .Y(new_n11461));
  NAND2xp33_ASAP7_75t_L     g11205(.A(new_n11460), .B(new_n11461), .Y(new_n11462));
  AOI211xp5_ASAP7_75t_L     g11206(.A1(\b[31] ), .A2(new_n2931), .B(new_n2697), .C(new_n11462), .Y(new_n11463));
  INVx1_ASAP7_75t_L         g11207(.A(new_n11462), .Y(new_n11464));
  O2A1O1Ixp33_ASAP7_75t_L   g11208(.A1(new_n3419), .A2(new_n2932), .B(new_n11464), .C(\a[29] ), .Y(new_n11465));
  NOR2xp33_ASAP7_75t_L      g11209(.A(new_n11463), .B(new_n11465), .Y(new_n11466));
  NAND3xp33_ASAP7_75t_L     g11210(.A(new_n11455), .B(new_n11459), .C(new_n11466), .Y(new_n11467));
  NOR3xp33_ASAP7_75t_L      g11211(.A(new_n11458), .B(new_n11457), .C(new_n11456), .Y(new_n11468));
  AOI211xp5_ASAP7_75t_L     g11212(.A1(new_n11450), .A2(new_n11453), .B(new_n11081), .C(new_n11454), .Y(new_n11469));
  INVx1_ASAP7_75t_L         g11213(.A(new_n11466), .Y(new_n11470));
  OAI21xp33_ASAP7_75t_L     g11214(.A1(new_n11468), .A2(new_n11469), .B(new_n11470), .Y(new_n11471));
  AOI21xp33_ASAP7_75t_L     g11215(.A1(new_n11471), .A2(new_n11467), .B(new_n11289), .Y(new_n11472));
  AO21x2_ASAP7_75t_L        g11216(.A1(new_n11088), .A2(new_n10921), .B(new_n11288), .Y(new_n11473));
  NAND2xp33_ASAP7_75t_L     g11217(.A(new_n11467), .B(new_n11471), .Y(new_n11474));
  NOR2xp33_ASAP7_75t_L      g11218(.A(new_n11473), .B(new_n11474), .Y(new_n11475));
  NOR3xp33_ASAP7_75t_L      g11219(.A(new_n11475), .B(new_n11472), .C(new_n11287), .Y(new_n11476));
  INVx1_ASAP7_75t_L         g11220(.A(new_n11287), .Y(new_n11477));
  NAND2xp33_ASAP7_75t_L     g11221(.A(new_n11473), .B(new_n11474), .Y(new_n11478));
  NAND3xp33_ASAP7_75t_L     g11222(.A(new_n11289), .B(new_n11467), .C(new_n11471), .Y(new_n11479));
  AOI21xp33_ASAP7_75t_L     g11223(.A1(new_n11478), .A2(new_n11479), .B(new_n11477), .Y(new_n11480));
  OAI221xp5_ASAP7_75t_L     g11224(.A1(new_n11480), .A2(new_n11476), .B1(new_n11112), .B2(new_n11122), .C(new_n11281), .Y(new_n11481));
  A2O1A1Ixp33_ASAP7_75t_L   g11225(.A1(new_n11107), .A2(new_n11104), .B(new_n11112), .C(new_n11281), .Y(new_n11482));
  NOR2xp33_ASAP7_75t_L      g11226(.A(new_n11480), .B(new_n11476), .Y(new_n11483));
  NAND2xp33_ASAP7_75t_L     g11227(.A(new_n11482), .B(new_n11483), .Y(new_n11484));
  NAND2xp33_ASAP7_75t_L     g11228(.A(\b[38] ), .B(new_n1770), .Y(new_n11485));
  AOI22xp33_ASAP7_75t_L     g11229(.A1(new_n1766), .A2(\b[39] ), .B1(new_n1764), .B2(new_n5174), .Y(new_n11486));
  NAND2xp33_ASAP7_75t_L     g11230(.A(new_n11485), .B(new_n11486), .Y(new_n11487));
  AOI21xp33_ASAP7_75t_L     g11231(.A1(new_n1910), .A2(\b[37] ), .B(new_n11487), .Y(new_n11488));
  NAND2xp33_ASAP7_75t_L     g11232(.A(\a[23] ), .B(new_n11488), .Y(new_n11489));
  A2O1A1Ixp33_ASAP7_75t_L   g11233(.A1(\b[37] ), .A2(new_n1910), .B(new_n11487), .C(new_n1761), .Y(new_n11490));
  NAND2xp33_ASAP7_75t_L     g11234(.A(new_n11490), .B(new_n11489), .Y(new_n11491));
  INVx1_ASAP7_75t_L         g11235(.A(new_n11491), .Y(new_n11492));
  NAND3xp33_ASAP7_75t_L     g11236(.A(new_n11484), .B(new_n11492), .C(new_n11481), .Y(new_n11493));
  NOR2xp33_ASAP7_75t_L      g11237(.A(new_n11482), .B(new_n11483), .Y(new_n11494));
  NAND3xp33_ASAP7_75t_L     g11238(.A(new_n11478), .B(new_n11479), .C(new_n11477), .Y(new_n11495));
  OAI21xp33_ASAP7_75t_L     g11239(.A1(new_n11472), .A2(new_n11475), .B(new_n11287), .Y(new_n11496));
  NAND2xp33_ASAP7_75t_L     g11240(.A(new_n11495), .B(new_n11496), .Y(new_n11497));
  O2A1O1Ixp33_ASAP7_75t_L   g11241(.A1(new_n11122), .A2(new_n11112), .B(new_n11281), .C(new_n11497), .Y(new_n11498));
  OAI21xp33_ASAP7_75t_L     g11242(.A1(new_n11494), .A2(new_n11498), .B(new_n11491), .Y(new_n11499));
  NOR3xp33_ASAP7_75t_L      g11243(.A(new_n11125), .B(new_n11111), .C(new_n11113), .Y(new_n11500));
  O2A1O1Ixp33_ASAP7_75t_L   g11244(.A1(new_n11121), .A2(new_n11126), .B(new_n11128), .C(new_n11500), .Y(new_n11501));
  NAND3xp33_ASAP7_75t_L     g11245(.A(new_n11501), .B(new_n11499), .C(new_n11493), .Y(new_n11502));
  NAND2xp33_ASAP7_75t_L     g11246(.A(new_n11493), .B(new_n11499), .Y(new_n11503));
  OAI21xp33_ASAP7_75t_L     g11247(.A1(new_n11500), .A2(new_n11130), .B(new_n11503), .Y(new_n11504));
  NAND2xp33_ASAP7_75t_L     g11248(.A(\b[42] ), .B(new_n1406), .Y(new_n11505));
  OAI221xp5_ASAP7_75t_L     g11249(.A1(new_n5666), .A2(new_n1398), .B1(new_n1411), .B2(new_n5687), .C(new_n11505), .Y(new_n11506));
  AOI21xp33_ASAP7_75t_L     g11250(.A1(new_n1548), .A2(\b[40] ), .B(new_n11506), .Y(new_n11507));
  NAND2xp33_ASAP7_75t_L     g11251(.A(\a[20] ), .B(new_n11507), .Y(new_n11508));
  A2O1A1Ixp33_ASAP7_75t_L   g11252(.A1(\b[40] ), .A2(new_n1548), .B(new_n11506), .C(new_n1401), .Y(new_n11509));
  NAND2xp33_ASAP7_75t_L     g11253(.A(new_n11509), .B(new_n11508), .Y(new_n11510));
  AO21x2_ASAP7_75t_L        g11254(.A1(new_n11502), .A2(new_n11504), .B(new_n11510), .Y(new_n11511));
  NAND3xp33_ASAP7_75t_L     g11255(.A(new_n11504), .B(new_n11502), .C(new_n11510), .Y(new_n11512));
  A2O1A1O1Ixp25_ASAP7_75t_L g11256(.A1(new_n10425), .A2(new_n10782), .B(new_n10787), .C(new_n10919), .D(new_n11145), .Y(new_n11513));
  OAI211xp5_ASAP7_75t_L     g11257(.A1(new_n11146), .A2(new_n11513), .B(new_n11511), .C(new_n11512), .Y(new_n11514));
  AOI21xp33_ASAP7_75t_L     g11258(.A1(new_n11504), .A2(new_n11502), .B(new_n11510), .Y(new_n11515));
  AND3x1_ASAP7_75t_L        g11259(.A(new_n11504), .B(new_n11510), .C(new_n11502), .Y(new_n11516));
  A2O1A1O1Ixp25_ASAP7_75t_L g11260(.A1(new_n10780), .A2(new_n10783), .B(new_n10918), .C(new_n11139), .D(new_n11146), .Y(new_n11517));
  OAI21xp33_ASAP7_75t_L     g11261(.A1(new_n11515), .A2(new_n11516), .B(new_n11517), .Y(new_n11518));
  AOI21xp33_ASAP7_75t_L     g11262(.A1(new_n11514), .A2(new_n11518), .B(new_n11279), .Y(new_n11519));
  NAND2xp33_ASAP7_75t_L     g11263(.A(new_n11278), .B(new_n11277), .Y(new_n11520));
  NOR3xp33_ASAP7_75t_L      g11264(.A(new_n11516), .B(new_n11517), .C(new_n11515), .Y(new_n11521));
  AOI211xp5_ASAP7_75t_L     g11265(.A1(new_n11511), .A2(new_n11512), .B(new_n11513), .C(new_n11146), .Y(new_n11522));
  NOR3xp33_ASAP7_75t_L      g11266(.A(new_n11522), .B(new_n11521), .C(new_n11520), .Y(new_n11523));
  NOR2xp33_ASAP7_75t_L      g11267(.A(new_n11519), .B(new_n11523), .Y(new_n11524));
  NOR2xp33_ASAP7_75t_L      g11268(.A(new_n11273), .B(new_n11524), .Y(new_n11525));
  A2O1A1Ixp33_ASAP7_75t_L   g11269(.A1(new_n11155), .A2(new_n10799), .B(new_n11159), .C(new_n11149), .Y(new_n11526));
  OAI21xp33_ASAP7_75t_L     g11270(.A1(new_n11521), .A2(new_n11522), .B(new_n11520), .Y(new_n11527));
  NAND3xp33_ASAP7_75t_L     g11271(.A(new_n11514), .B(new_n11279), .C(new_n11518), .Y(new_n11528));
  NAND2xp33_ASAP7_75t_L     g11272(.A(new_n11528), .B(new_n11527), .Y(new_n11529));
  NOR2xp33_ASAP7_75t_L      g11273(.A(new_n11526), .B(new_n11529), .Y(new_n11530));
  OAI21xp33_ASAP7_75t_L     g11274(.A1(new_n11530), .A2(new_n11525), .B(new_n11272), .Y(new_n11531));
  NAND2xp33_ASAP7_75t_L     g11275(.A(new_n11526), .B(new_n11529), .Y(new_n11532));
  NAND2xp33_ASAP7_75t_L     g11276(.A(new_n11273), .B(new_n11524), .Y(new_n11533));
  NAND3xp33_ASAP7_75t_L     g11277(.A(new_n11533), .B(new_n11532), .C(new_n11271), .Y(new_n11534));
  AOI21xp33_ASAP7_75t_L     g11278(.A1(new_n11534), .A2(new_n11531), .B(new_n11265), .Y(new_n11535));
  OAI21xp33_ASAP7_75t_L     g11279(.A1(new_n11173), .A2(new_n11171), .B(new_n11163), .Y(new_n11536));
  NAND2xp33_ASAP7_75t_L     g11280(.A(new_n11534), .B(new_n11531), .Y(new_n11537));
  NOR2xp33_ASAP7_75t_L      g11281(.A(new_n11536), .B(new_n11537), .Y(new_n11538));
  OAI21xp33_ASAP7_75t_L     g11282(.A1(new_n11535), .A2(new_n11538), .B(new_n11264), .Y(new_n11539));
  INVx1_ASAP7_75t_L         g11283(.A(new_n11264), .Y(new_n11540));
  NAND2xp33_ASAP7_75t_L     g11284(.A(new_n11536), .B(new_n11537), .Y(new_n11541));
  NAND3xp33_ASAP7_75t_L     g11285(.A(new_n11265), .B(new_n11531), .C(new_n11534), .Y(new_n11542));
  NAND3xp33_ASAP7_75t_L     g11286(.A(new_n11541), .B(new_n11540), .C(new_n11542), .Y(new_n11543));
  NAND2xp33_ASAP7_75t_L     g11287(.A(new_n11543), .B(new_n11539), .Y(new_n11544));
  NAND2xp33_ASAP7_75t_L     g11288(.A(new_n11257), .B(new_n11544), .Y(new_n11545));
  MAJx2_ASAP7_75t_L         g11289(.A(new_n10902), .B(new_n11256), .C(new_n11181), .Y(new_n11546));
  AOI21xp33_ASAP7_75t_L     g11290(.A1(new_n11541), .A2(new_n11542), .B(new_n11540), .Y(new_n11547));
  NOR3xp33_ASAP7_75t_L      g11291(.A(new_n11538), .B(new_n11535), .C(new_n11264), .Y(new_n11548));
  NOR2xp33_ASAP7_75t_L      g11292(.A(new_n11547), .B(new_n11548), .Y(new_n11549));
  NAND2xp33_ASAP7_75t_L     g11293(.A(new_n11546), .B(new_n11549), .Y(new_n11550));
  NAND3xp33_ASAP7_75t_L     g11294(.A(new_n11550), .B(new_n11545), .C(new_n11255), .Y(new_n11551));
  NOR2xp33_ASAP7_75t_L      g11295(.A(new_n11546), .B(new_n11549), .Y(new_n11552));
  NOR2xp33_ASAP7_75t_L      g11296(.A(new_n11257), .B(new_n11544), .Y(new_n11553));
  OAI21xp33_ASAP7_75t_L     g11297(.A1(new_n11553), .A2(new_n11552), .B(new_n11254), .Y(new_n11554));
  NAND3xp33_ASAP7_75t_L     g11298(.A(new_n11247), .B(new_n11551), .C(new_n11554), .Y(new_n11555));
  NOR3xp33_ASAP7_75t_L      g11299(.A(new_n11552), .B(new_n11553), .C(new_n11254), .Y(new_n11556));
  AOI21xp33_ASAP7_75t_L     g11300(.A1(new_n11550), .A2(new_n11545), .B(new_n11255), .Y(new_n11557));
  OAI221xp5_ASAP7_75t_L     g11301(.A1(new_n11204), .A2(new_n10894), .B1(new_n11557), .B2(new_n11556), .C(new_n11246), .Y(new_n11558));
  NAND3xp33_ASAP7_75t_L     g11302(.A(new_n11558), .B(new_n11245), .C(new_n11555), .Y(new_n11559));
  AO21x2_ASAP7_75t_L        g11303(.A1(new_n11555), .A2(new_n11558), .B(new_n11245), .Y(new_n11560));
  NAND3xp33_ASAP7_75t_L     g11304(.A(new_n11560), .B(new_n11242), .C(new_n11559), .Y(new_n11561));
  AND3x1_ASAP7_75t_L        g11305(.A(new_n11558), .B(new_n11555), .C(new_n11245), .Y(new_n11562));
  AOI21xp33_ASAP7_75t_L     g11306(.A1(new_n11558), .A2(new_n11555), .B(new_n11245), .Y(new_n11563));
  OAI21xp33_ASAP7_75t_L     g11307(.A1(new_n11563), .A2(new_n11562), .B(new_n11241), .Y(new_n11564));
  NAND4xp25_ASAP7_75t_L     g11308(.A(new_n11564), .B(new_n11561), .C(new_n11207), .D(new_n11208), .Y(new_n11565));
  NOR3xp33_ASAP7_75t_L      g11309(.A(new_n11562), .B(new_n11563), .C(new_n11241), .Y(new_n11566));
  AOI21xp33_ASAP7_75t_L     g11310(.A1(new_n11560), .A2(new_n11559), .B(new_n11242), .Y(new_n11567));
  NAND2xp33_ASAP7_75t_L     g11311(.A(new_n11207), .B(new_n11208), .Y(new_n11568));
  OAI21xp33_ASAP7_75t_L     g11312(.A1(new_n11567), .A2(new_n11566), .B(new_n11568), .Y(new_n11569));
  NAND2xp33_ASAP7_75t_L     g11313(.A(new_n11565), .B(new_n11569), .Y(new_n11570));
  O2A1O1Ixp33_ASAP7_75t_L   g11314(.A1(new_n11214), .A2(new_n11220), .B(new_n11222), .C(new_n11570), .Y(new_n11571));
  A2O1A1O1Ixp25_ASAP7_75t_L g11315(.A1(new_n10866), .A2(new_n10508), .B(new_n10842), .C(new_n10840), .D(new_n11220), .Y(new_n11572));
  INVx1_ASAP7_75t_L         g11316(.A(new_n11572), .Y(new_n11573));
  AND3x1_ASAP7_75t_L        g11317(.A(new_n11570), .B(new_n11573), .C(new_n11222), .Y(new_n11574));
  NOR2xp33_ASAP7_75t_L      g11318(.A(new_n11571), .B(new_n11574), .Y(\f[60] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g11319(.A1(new_n10874), .A2(new_n10871), .B(new_n11221), .C(new_n11218), .D(new_n11572), .Y(new_n11576));
  NOR3xp33_ASAP7_75t_L      g11320(.A(new_n11538), .B(new_n11535), .C(new_n11540), .Y(new_n11577));
  NAND2xp33_ASAP7_75t_L     g11321(.A(\b[51] ), .B(new_n590), .Y(new_n11578));
  AOI22xp33_ASAP7_75t_L     g11322(.A1(new_n600), .A2(\b[52] ), .B1(new_n597), .B2(new_n8577), .Y(new_n11579));
  NAND2xp33_ASAP7_75t_L     g11323(.A(new_n11578), .B(new_n11579), .Y(new_n11580));
  AOI211xp5_ASAP7_75t_L     g11324(.A1(\b[50] ), .A2(new_n674), .B(new_n594), .C(new_n11580), .Y(new_n11581));
  INVx1_ASAP7_75t_L         g11325(.A(new_n11580), .Y(new_n11582));
  O2A1O1Ixp33_ASAP7_75t_L   g11326(.A1(new_n8228), .A2(new_n1620), .B(new_n11582), .C(\a[11] ), .Y(new_n11583));
  NOR2xp33_ASAP7_75t_L      g11327(.A(new_n11581), .B(new_n11583), .Y(new_n11584));
  INVx1_ASAP7_75t_L         g11328(.A(new_n11584), .Y(new_n11585));
  NOR3xp33_ASAP7_75t_L      g11329(.A(new_n11525), .B(new_n11530), .C(new_n11271), .Y(new_n11586));
  INVx1_ASAP7_75t_L         g11330(.A(new_n11586), .Y(new_n11587));
  A2O1A1Ixp33_ASAP7_75t_L   g11331(.A1(new_n11531), .A2(new_n11534), .B(new_n11265), .C(new_n11587), .Y(new_n11588));
  NAND2xp33_ASAP7_75t_L     g11332(.A(\b[47] ), .B(new_n908), .Y(new_n11589));
  NAND2xp33_ASAP7_75t_L     g11333(.A(\b[48] ), .B(new_n817), .Y(new_n11590));
  AOI22xp33_ASAP7_75t_L     g11334(.A1(new_n826), .A2(\b[49] ), .B1(new_n823), .B2(new_n7914), .Y(new_n11591));
  NAND4xp25_ASAP7_75t_L     g11335(.A(new_n11591), .B(\a[14] ), .C(new_n11589), .D(new_n11590), .Y(new_n11592));
  AOI31xp33_ASAP7_75t_L     g11336(.A1(new_n11591), .A2(new_n11590), .A3(new_n11589), .B(\a[14] ), .Y(new_n11593));
  INVx1_ASAP7_75t_L         g11337(.A(new_n11593), .Y(new_n11594));
  NAND2xp33_ASAP7_75t_L     g11338(.A(new_n11592), .B(new_n11594), .Y(new_n11595));
  INVx1_ASAP7_75t_L         g11339(.A(new_n11595), .Y(new_n11596));
  NOR3xp33_ASAP7_75t_L      g11340(.A(new_n11522), .B(new_n11279), .C(new_n11521), .Y(new_n11597));
  O2A1O1Ixp33_ASAP7_75t_L   g11341(.A1(new_n11519), .A2(new_n11523), .B(new_n11526), .C(new_n11597), .Y(new_n11598));
  NAND2xp33_ASAP7_75t_L     g11342(.A(\b[46] ), .B(new_n1113), .Y(new_n11599));
  OAI221xp5_ASAP7_75t_L     g11343(.A1(new_n6756), .A2(new_n1298), .B1(new_n1197), .B2(new_n7887), .C(new_n11599), .Y(new_n11600));
  AOI21xp33_ASAP7_75t_L     g11344(.A1(new_n1194), .A2(\b[44] ), .B(new_n11600), .Y(new_n11601));
  NAND2xp33_ASAP7_75t_L     g11345(.A(\a[17] ), .B(new_n11601), .Y(new_n11602));
  A2O1A1Ixp33_ASAP7_75t_L   g11346(.A1(\b[44] ), .A2(new_n1194), .B(new_n11600), .C(new_n1107), .Y(new_n11603));
  NAND2xp33_ASAP7_75t_L     g11347(.A(new_n11603), .B(new_n11602), .Y(new_n11604));
  A2O1A1Ixp33_ASAP7_75t_L   g11348(.A1(new_n10783), .A2(new_n10780), .B(new_n10918), .C(new_n11139), .Y(new_n11605));
  A2O1A1Ixp33_ASAP7_75t_L   g11349(.A1(new_n11605), .A2(new_n11142), .B(new_n11515), .C(new_n11512), .Y(new_n11606));
  NAND2xp33_ASAP7_75t_L     g11350(.A(new_n11459), .B(new_n11455), .Y(new_n11607));
  NOR2xp33_ASAP7_75t_L      g11351(.A(new_n11466), .B(new_n11607), .Y(new_n11608));
  A2O1A1O1Ixp25_ASAP7_75t_L g11352(.A1(new_n11084), .A2(new_n11090), .B(new_n11081), .C(new_n11450), .D(new_n11457), .Y(new_n11609));
  INVx1_ASAP7_75t_L         g11353(.A(new_n11397), .Y(new_n11610));
  O2A1O1Ixp33_ASAP7_75t_L   g11354(.A1(new_n11403), .A2(new_n11049), .B(new_n11401), .C(new_n11610), .Y(new_n11611));
  AOI22xp33_ASAP7_75t_L     g11355(.A1(new_n5249), .A2(\b[22] ), .B1(new_n5247), .B2(new_n1864), .Y(new_n11612));
  OAI221xp5_ASAP7_75t_L     g11356(.A1(new_n5241), .A2(new_n1709), .B1(new_n1594), .B2(new_n5521), .C(new_n11612), .Y(new_n11613));
  XNOR2x2_ASAP7_75t_L       g11357(.A(\a[41] ), .B(new_n11613), .Y(new_n11614));
  INVx1_ASAP7_75t_L         g11358(.A(new_n11304), .Y(new_n11615));
  NAND3xp33_ASAP7_75t_L     g11359(.A(new_n11389), .B(new_n11385), .C(new_n11615), .Y(new_n11616));
  INVx1_ASAP7_75t_L         g11360(.A(new_n11616), .Y(new_n11617));
  O2A1O1Ixp33_ASAP7_75t_L   g11361(.A1(new_n11390), .A2(new_n11391), .B(new_n11301), .C(new_n11617), .Y(new_n11618));
  AOI21xp33_ASAP7_75t_L     g11362(.A1(new_n11378), .A2(new_n11382), .B(new_n11314), .Y(new_n11619));
  A2O1A1Ixp33_ASAP7_75t_L   g11363(.A1(new_n11031), .A2(new_n11306), .B(new_n11619), .C(new_n11383), .Y(new_n11620));
  NOR2xp33_ASAP7_75t_L      g11364(.A(new_n1051), .B(new_n7118), .Y(new_n11621));
  AOI221xp5_ASAP7_75t_L     g11365(.A1(new_n6812), .A2(\b[15] ), .B1(new_n6819), .B2(new_n1058), .C(new_n11621), .Y(new_n11622));
  OA211x2_ASAP7_75t_L       g11366(.A1(new_n7115), .A2(new_n871), .B(new_n11622), .C(\a[47] ), .Y(new_n11623));
  O2A1O1Ixp33_ASAP7_75t_L   g11367(.A1(new_n871), .A2(new_n7115), .B(new_n11622), .C(\a[47] ), .Y(new_n11624));
  NOR2xp33_ASAP7_75t_L      g11368(.A(new_n11624), .B(new_n11623), .Y(new_n11625));
  A2O1A1O1Ixp25_ASAP7_75t_L g11369(.A1(new_n11000), .A2(new_n10951), .B(new_n11009), .C(new_n11373), .D(new_n11381), .Y(new_n11626));
  NAND2xp33_ASAP7_75t_L     g11370(.A(new_n11342), .B(new_n11346), .Y(new_n11627));
  AND2x2_ASAP7_75t_L        g11371(.A(new_n11350), .B(new_n11352), .Y(new_n11628));
  NOR2xp33_ASAP7_75t_L      g11372(.A(new_n11628), .B(new_n11627), .Y(new_n11629));
  O2A1O1Ixp33_ASAP7_75t_L   g11373(.A1(new_n11353), .A2(new_n11354), .B(new_n11357), .C(new_n11629), .Y(new_n11630));
  NAND2xp33_ASAP7_75t_L     g11374(.A(\b[7] ), .B(new_n9623), .Y(new_n11631));
  OAI221xp5_ASAP7_75t_L     g11375(.A1(new_n382), .A2(new_n10280), .B1(new_n9949), .B2(new_n427), .C(new_n11631), .Y(new_n11632));
  AOI21xp33_ASAP7_75t_L     g11376(.A1(new_n9948), .A2(\b[5] ), .B(new_n11632), .Y(new_n11633));
  NAND2xp33_ASAP7_75t_L     g11377(.A(\a[56] ), .B(new_n11633), .Y(new_n11634));
  INVx1_ASAP7_75t_L         g11378(.A(new_n11634), .Y(new_n11635));
  A2O1A1Ixp33_ASAP7_75t_L   g11379(.A1(\b[5] ), .A2(new_n9948), .B(new_n11632), .C(new_n9610), .Y(new_n11636));
  INVx1_ASAP7_75t_L         g11380(.A(new_n11636), .Y(new_n11637));
  NAND2xp33_ASAP7_75t_L     g11381(.A(new_n11327), .B(new_n11332), .Y(new_n11638));
  A2O1A1Ixp33_ASAP7_75t_L   g11382(.A1(new_n11343), .A2(new_n11344), .B(new_n11345), .C(new_n11638), .Y(new_n11639));
  AOI22xp33_ASAP7_75t_L     g11383(.A1(new_n10594), .A2(\b[4] ), .B1(new_n10591), .B2(new_n328), .Y(new_n11640));
  OAI221xp5_ASAP7_75t_L     g11384(.A1(new_n11335), .A2(new_n299), .B1(new_n278), .B2(new_n11330), .C(new_n11640), .Y(new_n11641));
  NOR2xp33_ASAP7_75t_L      g11385(.A(new_n10588), .B(new_n11641), .Y(new_n11642));
  AND2x2_ASAP7_75t_L        g11386(.A(new_n10588), .B(new_n11641), .Y(new_n11643));
  NAND2xp33_ASAP7_75t_L     g11387(.A(\a[62] ), .B(new_n11327), .Y(new_n11644));
  NAND2xp33_ASAP7_75t_L     g11388(.A(new_n11325), .B(new_n11324), .Y(new_n11645));
  XNOR2x2_ASAP7_75t_L       g11389(.A(\a[61] ), .B(\a[60] ), .Y(new_n11646));
  NOR2xp33_ASAP7_75t_L      g11390(.A(new_n11646), .B(new_n11645), .Y(new_n11647));
  NAND2xp33_ASAP7_75t_L     g11391(.A(\b[0] ), .B(new_n11647), .Y(new_n11648));
  INVx1_ASAP7_75t_L         g11392(.A(\a[61] ), .Y(new_n11649));
  NAND2xp33_ASAP7_75t_L     g11393(.A(\a[62] ), .B(new_n11649), .Y(new_n11650));
  INVx1_ASAP7_75t_L         g11394(.A(\a[62] ), .Y(new_n11651));
  NAND2xp33_ASAP7_75t_L     g11395(.A(\a[61] ), .B(new_n11651), .Y(new_n11652));
  AND2x2_ASAP7_75t_L        g11396(.A(new_n11650), .B(new_n11652), .Y(new_n11653));
  NOR2xp33_ASAP7_75t_L      g11397(.A(new_n11326), .B(new_n11653), .Y(new_n11654));
  NAND2xp33_ASAP7_75t_L     g11398(.A(new_n271), .B(new_n11654), .Y(new_n11655));
  AND3x1_ASAP7_75t_L        g11399(.A(new_n11645), .B(new_n11652), .C(new_n11650), .Y(new_n11656));
  NAND2xp33_ASAP7_75t_L     g11400(.A(\b[1] ), .B(new_n11656), .Y(new_n11657));
  NAND3xp33_ASAP7_75t_L     g11401(.A(new_n11655), .B(new_n11657), .C(new_n11648), .Y(new_n11658));
  XNOR2x2_ASAP7_75t_L       g11402(.A(new_n11644), .B(new_n11658), .Y(new_n11659));
  NOR3xp33_ASAP7_75t_L      g11403(.A(new_n11643), .B(new_n11642), .C(new_n11659), .Y(new_n11660));
  INVx1_ASAP7_75t_L         g11404(.A(new_n11660), .Y(new_n11661));
  OAI21xp33_ASAP7_75t_L     g11405(.A1(new_n11642), .A2(new_n11643), .B(new_n11659), .Y(new_n11662));
  NAND3xp33_ASAP7_75t_L     g11406(.A(new_n11661), .B(new_n11639), .C(new_n11662), .Y(new_n11663));
  AND2x2_ASAP7_75t_L        g11407(.A(new_n11327), .B(new_n11332), .Y(new_n11664));
  O2A1O1Ixp33_ASAP7_75t_L   g11408(.A1(new_n11333), .A2(new_n11334), .B(new_n11341), .C(new_n11664), .Y(new_n11665));
  INVx1_ASAP7_75t_L         g11409(.A(new_n11662), .Y(new_n11666));
  OAI21xp33_ASAP7_75t_L     g11410(.A1(new_n11660), .A2(new_n11666), .B(new_n11665), .Y(new_n11667));
  AOI211xp5_ASAP7_75t_L     g11411(.A1(new_n11667), .A2(new_n11663), .B(new_n11635), .C(new_n11637), .Y(new_n11668));
  OAI211xp5_ASAP7_75t_L     g11412(.A1(new_n11635), .A2(new_n11637), .B(new_n11667), .C(new_n11663), .Y(new_n11669));
  INVx1_ASAP7_75t_L         g11413(.A(new_n11669), .Y(new_n11670));
  NOR3xp33_ASAP7_75t_L      g11414(.A(new_n11670), .B(new_n11630), .C(new_n11668), .Y(new_n11671));
  MAJIxp5_ASAP7_75t_L       g11415(.A(new_n11359), .B(new_n11627), .C(new_n11628), .Y(new_n11672));
  NOR3xp33_ASAP7_75t_L      g11416(.A(new_n11666), .B(new_n11660), .C(new_n11665), .Y(new_n11673));
  AOI21xp33_ASAP7_75t_L     g11417(.A1(new_n11661), .A2(new_n11662), .B(new_n11639), .Y(new_n11674));
  OAI211xp5_ASAP7_75t_L     g11418(.A1(new_n11673), .A2(new_n11674), .B(new_n11636), .C(new_n11634), .Y(new_n11675));
  AOI21xp33_ASAP7_75t_L     g11419(.A1(new_n11669), .A2(new_n11675), .B(new_n11672), .Y(new_n11676));
  NAND2xp33_ASAP7_75t_L     g11420(.A(\b[8] ), .B(new_n8964), .Y(new_n11677));
  NAND2xp33_ASAP7_75t_L     g11421(.A(\b[9] ), .B(new_n8635), .Y(new_n11678));
  AOI22xp33_ASAP7_75t_L     g11422(.A1(new_n8645), .A2(\b[10] ), .B1(new_n8642), .B2(new_n852), .Y(new_n11679));
  NAND4xp25_ASAP7_75t_L     g11423(.A(new_n11679), .B(\a[53] ), .C(new_n11677), .D(new_n11678), .Y(new_n11680));
  NAND2xp33_ASAP7_75t_L     g11424(.A(new_n11678), .B(new_n11679), .Y(new_n11681));
  A2O1A1Ixp33_ASAP7_75t_L   g11425(.A1(\b[8] ), .A2(new_n8964), .B(new_n11681), .C(new_n8639), .Y(new_n11682));
  NAND2xp33_ASAP7_75t_L     g11426(.A(new_n11680), .B(new_n11682), .Y(new_n11683));
  NOR3xp33_ASAP7_75t_L      g11427(.A(new_n11671), .B(new_n11676), .C(new_n11683), .Y(new_n11684));
  NAND3xp33_ASAP7_75t_L     g11428(.A(new_n11672), .B(new_n11675), .C(new_n11669), .Y(new_n11685));
  OAI21xp33_ASAP7_75t_L     g11429(.A1(new_n11668), .A2(new_n11670), .B(new_n11630), .Y(new_n11686));
  INVx1_ASAP7_75t_L         g11430(.A(new_n11683), .Y(new_n11687));
  AOI21xp33_ASAP7_75t_L     g11431(.A1(new_n11686), .A2(new_n11685), .B(new_n11687), .Y(new_n11688));
  OAI21xp33_ASAP7_75t_L     g11432(.A1(new_n11367), .A2(new_n11322), .B(new_n11370), .Y(new_n11689));
  NOR3xp33_ASAP7_75t_L      g11433(.A(new_n11689), .B(new_n11688), .C(new_n11684), .Y(new_n11690));
  NAND3xp33_ASAP7_75t_L     g11434(.A(new_n11687), .B(new_n11686), .C(new_n11685), .Y(new_n11691));
  OAI21xp33_ASAP7_75t_L     g11435(.A1(new_n11676), .A2(new_n11671), .B(new_n11683), .Y(new_n11692));
  A2O1A1O1Ixp25_ASAP7_75t_L g11436(.A1(new_n10997), .A2(new_n10996), .B(new_n10994), .C(new_n11371), .D(new_n11366), .Y(new_n11693));
  AOI21xp33_ASAP7_75t_L     g11437(.A1(new_n11691), .A2(new_n11692), .B(new_n11693), .Y(new_n11694));
  NAND2xp33_ASAP7_75t_L     g11438(.A(new_n7656), .B(new_n800), .Y(new_n11695));
  OAI221xp5_ASAP7_75t_L     g11439(.A1(new_n7997), .A2(new_n793), .B1(new_n763), .B2(new_n8326), .C(new_n11695), .Y(new_n11696));
  AOI21xp33_ASAP7_75t_L     g11440(.A1(new_n7993), .A2(\b[11] ), .B(new_n11696), .Y(new_n11697));
  XNOR2x2_ASAP7_75t_L       g11441(.A(new_n7653), .B(new_n11697), .Y(new_n11698));
  OAI21xp33_ASAP7_75t_L     g11442(.A1(new_n11690), .A2(new_n11694), .B(new_n11698), .Y(new_n11699));
  NAND3xp33_ASAP7_75t_L     g11443(.A(new_n11691), .B(new_n11693), .C(new_n11692), .Y(new_n11700));
  OAI21xp33_ASAP7_75t_L     g11444(.A1(new_n11688), .A2(new_n11684), .B(new_n11689), .Y(new_n11701));
  NAND2xp33_ASAP7_75t_L     g11445(.A(\a[50] ), .B(new_n11697), .Y(new_n11702));
  A2O1A1Ixp33_ASAP7_75t_L   g11446(.A1(\b[11] ), .A2(new_n7993), .B(new_n11696), .C(new_n7653), .Y(new_n11703));
  NAND2xp33_ASAP7_75t_L     g11447(.A(new_n11703), .B(new_n11702), .Y(new_n11704));
  NAND3xp33_ASAP7_75t_L     g11448(.A(new_n11704), .B(new_n11701), .C(new_n11700), .Y(new_n11705));
  NAND3xp33_ASAP7_75t_L     g11449(.A(new_n11626), .B(new_n11699), .C(new_n11705), .Y(new_n11706));
  A2O1A1Ixp33_ASAP7_75t_L   g11450(.A1(new_n11005), .A2(new_n11004), .B(new_n11380), .C(new_n11377), .Y(new_n11707));
  AOI21xp33_ASAP7_75t_L     g11451(.A1(new_n11700), .A2(new_n11701), .B(new_n11704), .Y(new_n11708));
  NOR3xp33_ASAP7_75t_L      g11452(.A(new_n11698), .B(new_n11694), .C(new_n11690), .Y(new_n11709));
  OAI21xp33_ASAP7_75t_L     g11453(.A1(new_n11708), .A2(new_n11709), .B(new_n11707), .Y(new_n11710));
  AO21x2_ASAP7_75t_L        g11454(.A1(new_n11710), .A2(new_n11706), .B(new_n11625), .Y(new_n11711));
  NAND3xp33_ASAP7_75t_L     g11455(.A(new_n11706), .B(new_n11710), .C(new_n11625), .Y(new_n11712));
  AOI21xp33_ASAP7_75t_L     g11456(.A1(new_n11712), .A2(new_n11711), .B(new_n11620), .Y(new_n11713));
  INVx1_ASAP7_75t_L         g11457(.A(new_n11713), .Y(new_n11714));
  NAND3xp33_ASAP7_75t_L     g11458(.A(new_n11620), .B(new_n11711), .C(new_n11712), .Y(new_n11715));
  AOI22xp33_ASAP7_75t_L     g11459(.A1(new_n6002), .A2(\b[19] ), .B1(new_n5999), .B2(new_n1499), .Y(new_n11716));
  OAI221xp5_ASAP7_75t_L     g11460(.A1(new_n6544), .A2(new_n1356), .B1(new_n1244), .B2(new_n6309), .C(new_n11716), .Y(new_n11717));
  XNOR2x2_ASAP7_75t_L       g11461(.A(\a[44] ), .B(new_n11717), .Y(new_n11718));
  INVx1_ASAP7_75t_L         g11462(.A(new_n11718), .Y(new_n11719));
  AOI21xp33_ASAP7_75t_L     g11463(.A1(new_n11714), .A2(new_n11715), .B(new_n11719), .Y(new_n11720));
  INVx1_ASAP7_75t_L         g11464(.A(new_n11715), .Y(new_n11721));
  NOR3xp33_ASAP7_75t_L      g11465(.A(new_n11721), .B(new_n11718), .C(new_n11713), .Y(new_n11722));
  NOR2xp33_ASAP7_75t_L      g11466(.A(new_n11720), .B(new_n11722), .Y(new_n11723));
  NAND2xp33_ASAP7_75t_L     g11467(.A(new_n11618), .B(new_n11723), .Y(new_n11724));
  NAND2xp33_ASAP7_75t_L     g11468(.A(new_n11395), .B(new_n11394), .Y(new_n11725));
  OAI21xp33_ASAP7_75t_L     g11469(.A1(new_n11713), .A2(new_n11721), .B(new_n11718), .Y(new_n11726));
  NAND3xp33_ASAP7_75t_L     g11470(.A(new_n11719), .B(new_n11714), .C(new_n11715), .Y(new_n11727));
  NAND2xp33_ASAP7_75t_L     g11471(.A(new_n11726), .B(new_n11727), .Y(new_n11728));
  A2O1A1Ixp33_ASAP7_75t_L   g11472(.A1(new_n11725), .A2(new_n11301), .B(new_n11617), .C(new_n11728), .Y(new_n11729));
  AOI21xp33_ASAP7_75t_L     g11473(.A1(new_n11729), .A2(new_n11724), .B(new_n11614), .Y(new_n11730));
  NOR2xp33_ASAP7_75t_L      g11474(.A(new_n5244), .B(new_n11613), .Y(new_n11731));
  AND2x2_ASAP7_75t_L        g11475(.A(new_n5244), .B(new_n11613), .Y(new_n11732));
  A2O1A1Ixp33_ASAP7_75t_L   g11476(.A1(new_n11394), .A2(new_n11395), .B(new_n11393), .C(new_n11616), .Y(new_n11733));
  NOR2xp33_ASAP7_75t_L      g11477(.A(new_n11733), .B(new_n11728), .Y(new_n11734));
  NOR2xp33_ASAP7_75t_L      g11478(.A(new_n11618), .B(new_n11723), .Y(new_n11735));
  NOR4xp25_ASAP7_75t_L      g11479(.A(new_n11735), .B(new_n11734), .C(new_n11731), .D(new_n11732), .Y(new_n11736));
  OAI21xp33_ASAP7_75t_L     g11480(.A1(new_n11730), .A2(new_n11736), .B(new_n11611), .Y(new_n11737));
  A2O1A1Ixp33_ASAP7_75t_L   g11481(.A1(new_n11044), .A2(new_n11038), .B(new_n11405), .C(new_n11397), .Y(new_n11738));
  NOR2xp33_ASAP7_75t_L      g11482(.A(new_n11730), .B(new_n11736), .Y(new_n11739));
  NAND2xp33_ASAP7_75t_L     g11483(.A(new_n11738), .B(new_n11739), .Y(new_n11740));
  AOI22xp33_ASAP7_75t_L     g11484(.A1(new_n4544), .A2(\b[25] ), .B1(new_n4542), .B2(new_n2188), .Y(new_n11741));
  OAI221xp5_ASAP7_75t_L     g11485(.A1(new_n4536), .A2(new_n2019), .B1(new_n1995), .B2(new_n4781), .C(new_n11741), .Y(new_n11742));
  XNOR2x2_ASAP7_75t_L       g11486(.A(\a[38] ), .B(new_n11742), .Y(new_n11743));
  NAND3xp33_ASAP7_75t_L     g11487(.A(new_n11740), .B(new_n11737), .C(new_n11743), .Y(new_n11744));
  NOR2xp33_ASAP7_75t_L      g11488(.A(new_n11738), .B(new_n11739), .Y(new_n11745));
  NOR3xp33_ASAP7_75t_L      g11489(.A(new_n11611), .B(new_n11730), .C(new_n11736), .Y(new_n11746));
  INVx1_ASAP7_75t_L         g11490(.A(new_n11743), .Y(new_n11747));
  OAI21xp33_ASAP7_75t_L     g11491(.A1(new_n11746), .A2(new_n11745), .B(new_n11747), .Y(new_n11748));
  NAND3xp33_ASAP7_75t_L     g11492(.A(new_n11402), .B(new_n11406), .C(new_n11415), .Y(new_n11749));
  NAND4xp25_ASAP7_75t_L     g11493(.A(new_n11421), .B(new_n11749), .C(new_n11748), .D(new_n11744), .Y(new_n11750));
  NOR3xp33_ASAP7_75t_L      g11494(.A(new_n11745), .B(new_n11747), .C(new_n11746), .Y(new_n11751));
  AOI21xp33_ASAP7_75t_L     g11495(.A1(new_n11740), .A2(new_n11737), .B(new_n11743), .Y(new_n11752));
  A2O1A1Ixp33_ASAP7_75t_L   g11496(.A1(new_n11416), .A2(new_n11412), .B(new_n11417), .C(new_n11749), .Y(new_n11753));
  OAI21xp33_ASAP7_75t_L     g11497(.A1(new_n11752), .A2(new_n11751), .B(new_n11753), .Y(new_n11754));
  AOI22xp33_ASAP7_75t_L     g11498(.A1(new_n3884), .A2(\b[28] ), .B1(new_n3881), .B2(new_n2858), .Y(new_n11755));
  OAI221xp5_ASAP7_75t_L     g11499(.A1(new_n4312), .A2(new_n2650), .B1(new_n2477), .B2(new_n4986), .C(new_n11755), .Y(new_n11756));
  XNOR2x2_ASAP7_75t_L       g11500(.A(\a[35] ), .B(new_n11756), .Y(new_n11757));
  NAND3xp33_ASAP7_75t_L     g11501(.A(new_n11750), .B(new_n11754), .C(new_n11757), .Y(new_n11758));
  NOR3xp33_ASAP7_75t_L      g11502(.A(new_n11753), .B(new_n11751), .C(new_n11752), .Y(new_n11759));
  AOI22xp33_ASAP7_75t_L     g11503(.A1(new_n11744), .A2(new_n11748), .B1(new_n11749), .B2(new_n11421), .Y(new_n11760));
  INVx1_ASAP7_75t_L         g11504(.A(new_n11757), .Y(new_n11761));
  OAI21xp33_ASAP7_75t_L     g11505(.A1(new_n11759), .A2(new_n11760), .B(new_n11761), .Y(new_n11762));
  NAND2xp33_ASAP7_75t_L     g11506(.A(new_n11758), .B(new_n11762), .Y(new_n11763));
  NOR3xp33_ASAP7_75t_L      g11507(.A(new_n11430), .B(new_n11428), .C(new_n11431), .Y(new_n11764));
  INVx1_ASAP7_75t_L         g11508(.A(new_n11764), .Y(new_n11765));
  A2O1A1Ixp33_ASAP7_75t_L   g11509(.A1(new_n11072), .A2(new_n11435), .B(new_n11441), .C(new_n11765), .Y(new_n11766));
  NOR2xp33_ASAP7_75t_L      g11510(.A(new_n11763), .B(new_n11766), .Y(new_n11767));
  NOR3xp33_ASAP7_75t_L      g11511(.A(new_n11760), .B(new_n11759), .C(new_n11761), .Y(new_n11768));
  AOI21xp33_ASAP7_75t_L     g11512(.A1(new_n11750), .A2(new_n11754), .B(new_n11757), .Y(new_n11769));
  NOR2xp33_ASAP7_75t_L      g11513(.A(new_n11769), .B(new_n11768), .Y(new_n11770));
  O2A1O1Ixp33_ASAP7_75t_L   g11514(.A1(new_n11439), .A2(new_n11440), .B(new_n11436), .C(new_n11764), .Y(new_n11771));
  NOR2xp33_ASAP7_75t_L      g11515(.A(new_n11771), .B(new_n11770), .Y(new_n11772));
  NOR2xp33_ASAP7_75t_L      g11516(.A(new_n3419), .B(new_n3262), .Y(new_n11773));
  AOI221xp5_ASAP7_75t_L     g11517(.A1(new_n3260), .A2(\b[30] ), .B1(new_n3254), .B2(new_n3426), .C(new_n11773), .Y(new_n11774));
  OAI21xp33_ASAP7_75t_L     g11518(.A1(new_n2871), .A2(new_n3492), .B(new_n11774), .Y(new_n11775));
  NOR2xp33_ASAP7_75t_L      g11519(.A(new_n3251), .B(new_n11775), .Y(new_n11776));
  O2A1O1Ixp33_ASAP7_75t_L   g11520(.A1(new_n2871), .A2(new_n3492), .B(new_n11774), .C(\a[32] ), .Y(new_n11777));
  NOR2xp33_ASAP7_75t_L      g11521(.A(new_n11777), .B(new_n11776), .Y(new_n11778));
  INVx1_ASAP7_75t_L         g11522(.A(new_n11778), .Y(new_n11779));
  NOR3xp33_ASAP7_75t_L      g11523(.A(new_n11767), .B(new_n11772), .C(new_n11779), .Y(new_n11780));
  NAND2xp33_ASAP7_75t_L     g11524(.A(new_n11771), .B(new_n11770), .Y(new_n11781));
  A2O1A1Ixp33_ASAP7_75t_L   g11525(.A1(new_n11434), .A2(new_n11436), .B(new_n11764), .C(new_n11763), .Y(new_n11782));
  AOI21xp33_ASAP7_75t_L     g11526(.A1(new_n11782), .A2(new_n11781), .B(new_n11778), .Y(new_n11783));
  NOR3xp33_ASAP7_75t_L      g11527(.A(new_n11609), .B(new_n11780), .C(new_n11783), .Y(new_n11784));
  A2O1A1Ixp33_ASAP7_75t_L   g11528(.A1(new_n10547), .A2(new_n10726), .B(new_n10930), .C(new_n11084), .Y(new_n11785));
  A2O1A1Ixp33_ASAP7_75t_L   g11529(.A1(new_n11785), .A2(new_n11085), .B(new_n11456), .C(new_n11453), .Y(new_n11786));
  NAND3xp33_ASAP7_75t_L     g11530(.A(new_n11782), .B(new_n11781), .C(new_n11778), .Y(new_n11787));
  OAI21xp33_ASAP7_75t_L     g11531(.A1(new_n11772), .A2(new_n11767), .B(new_n11779), .Y(new_n11788));
  AOI21xp33_ASAP7_75t_L     g11532(.A1(new_n11788), .A2(new_n11787), .B(new_n11786), .Y(new_n11789));
  NAND2xp33_ASAP7_75t_L     g11533(.A(\b[33] ), .B(new_n2706), .Y(new_n11790));
  AOI22xp33_ASAP7_75t_L     g11534(.A1(new_n2702), .A2(\b[34] ), .B1(new_n2700), .B2(new_n3833), .Y(new_n11791));
  NAND2xp33_ASAP7_75t_L     g11535(.A(new_n11790), .B(new_n11791), .Y(new_n11792));
  AOI21xp33_ASAP7_75t_L     g11536(.A1(new_n2931), .A2(\b[32] ), .B(new_n11792), .Y(new_n11793));
  NAND2xp33_ASAP7_75t_L     g11537(.A(\a[29] ), .B(new_n11793), .Y(new_n11794));
  A2O1A1Ixp33_ASAP7_75t_L   g11538(.A1(\b[32] ), .A2(new_n2931), .B(new_n11792), .C(new_n2697), .Y(new_n11795));
  NAND2xp33_ASAP7_75t_L     g11539(.A(new_n11795), .B(new_n11794), .Y(new_n11796));
  OAI21xp33_ASAP7_75t_L     g11540(.A1(new_n11789), .A2(new_n11784), .B(new_n11796), .Y(new_n11797));
  NAND3xp33_ASAP7_75t_L     g11541(.A(new_n11786), .B(new_n11787), .C(new_n11788), .Y(new_n11798));
  OAI21xp33_ASAP7_75t_L     g11542(.A1(new_n11783), .A2(new_n11780), .B(new_n11609), .Y(new_n11799));
  AND2x2_ASAP7_75t_L        g11543(.A(new_n11795), .B(new_n11794), .Y(new_n11800));
  NAND3xp33_ASAP7_75t_L     g11544(.A(new_n11798), .B(new_n11799), .C(new_n11800), .Y(new_n11801));
  AO221x2_ASAP7_75t_L       g11545(.A1(new_n11474), .A2(new_n11473), .B1(new_n11797), .B2(new_n11801), .C(new_n11608), .Y(new_n11802));
  MAJIxp5_ASAP7_75t_L       g11546(.A(new_n11289), .B(new_n11607), .C(new_n11466), .Y(new_n11803));
  NAND3xp33_ASAP7_75t_L     g11547(.A(new_n11803), .B(new_n11797), .C(new_n11801), .Y(new_n11804));
  NAND2xp33_ASAP7_75t_L     g11548(.A(\b[36] ), .B(new_n2232), .Y(new_n11805));
  AOI22xp33_ASAP7_75t_L     g11549(.A1(new_n2228), .A2(\b[37] ), .B1(new_n2226), .B2(new_n4709), .Y(new_n11806));
  NAND2xp33_ASAP7_75t_L     g11550(.A(new_n11805), .B(new_n11806), .Y(new_n11807));
  AOI211xp5_ASAP7_75t_L     g11551(.A1(\b[35] ), .A2(new_n2386), .B(new_n2223), .C(new_n11807), .Y(new_n11808));
  AND2x2_ASAP7_75t_L        g11552(.A(new_n11805), .B(new_n11806), .Y(new_n11809));
  O2A1O1Ixp33_ASAP7_75t_L   g11553(.A1(new_n4053), .A2(new_n2387), .B(new_n11809), .C(\a[26] ), .Y(new_n11810));
  NOR2xp33_ASAP7_75t_L      g11554(.A(new_n11808), .B(new_n11810), .Y(new_n11811));
  NAND3xp33_ASAP7_75t_L     g11555(.A(new_n11804), .B(new_n11802), .C(new_n11811), .Y(new_n11812));
  AOI21xp33_ASAP7_75t_L     g11556(.A1(new_n11801), .A2(new_n11797), .B(new_n11803), .Y(new_n11813));
  INVx1_ASAP7_75t_L         g11557(.A(new_n11608), .Y(new_n11814));
  NAND2xp33_ASAP7_75t_L     g11558(.A(new_n11801), .B(new_n11797), .Y(new_n11815));
  AOI21xp33_ASAP7_75t_L     g11559(.A1(new_n11478), .A2(new_n11814), .B(new_n11815), .Y(new_n11816));
  INVx1_ASAP7_75t_L         g11560(.A(new_n11811), .Y(new_n11817));
  OAI21xp33_ASAP7_75t_L     g11561(.A1(new_n11813), .A2(new_n11816), .B(new_n11817), .Y(new_n11818));
  NAND2xp33_ASAP7_75t_L     g11562(.A(new_n11812), .B(new_n11818), .Y(new_n11819));
  NOR3xp33_ASAP7_75t_L      g11563(.A(new_n11498), .B(new_n11819), .C(new_n11476), .Y(new_n11820));
  A2O1A1O1Ixp25_ASAP7_75t_L g11564(.A1(new_n11108), .A2(new_n11110), .B(new_n11280), .C(new_n11496), .D(new_n11476), .Y(new_n11821));
  AOI21xp33_ASAP7_75t_L     g11565(.A1(new_n11818), .A2(new_n11812), .B(new_n11821), .Y(new_n11822));
  INVx1_ASAP7_75t_L         g11566(.A(new_n5194), .Y(new_n11823));
  NAND2xp33_ASAP7_75t_L     g11567(.A(\b[40] ), .B(new_n1766), .Y(new_n11824));
  OAI221xp5_ASAP7_75t_L     g11568(.A1(new_n5166), .A2(new_n1758), .B1(new_n1771), .B2(new_n11823), .C(new_n11824), .Y(new_n11825));
  AOI21xp33_ASAP7_75t_L     g11569(.A1(new_n1910), .A2(\b[38] ), .B(new_n11825), .Y(new_n11826));
  NAND2xp33_ASAP7_75t_L     g11570(.A(\a[23] ), .B(new_n11826), .Y(new_n11827));
  A2O1A1Ixp33_ASAP7_75t_L   g11571(.A1(\b[38] ), .A2(new_n1910), .B(new_n11825), .C(new_n1761), .Y(new_n11828));
  NAND2xp33_ASAP7_75t_L     g11572(.A(new_n11828), .B(new_n11827), .Y(new_n11829));
  NOR3xp33_ASAP7_75t_L      g11573(.A(new_n11820), .B(new_n11822), .C(new_n11829), .Y(new_n11830));
  NAND3xp33_ASAP7_75t_L     g11574(.A(new_n11821), .B(new_n11818), .C(new_n11812), .Y(new_n11831));
  A2O1A1Ixp33_ASAP7_75t_L   g11575(.A1(new_n11483), .A2(new_n11482), .B(new_n11476), .C(new_n11819), .Y(new_n11832));
  INVx1_ASAP7_75t_L         g11576(.A(new_n11829), .Y(new_n11833));
  AOI21xp33_ASAP7_75t_L     g11577(.A1(new_n11832), .A2(new_n11831), .B(new_n11833), .Y(new_n11834));
  NOR2xp33_ASAP7_75t_L      g11578(.A(new_n11834), .B(new_n11830), .Y(new_n11835));
  NOR3xp33_ASAP7_75t_L      g11579(.A(new_n11498), .B(new_n11494), .C(new_n11492), .Y(new_n11836));
  O2A1O1Ixp33_ASAP7_75t_L   g11580(.A1(new_n11130), .A2(new_n11500), .B(new_n11503), .C(new_n11836), .Y(new_n11837));
  NAND2xp33_ASAP7_75t_L     g11581(.A(new_n11837), .B(new_n11835), .Y(new_n11838));
  NAND3xp33_ASAP7_75t_L     g11582(.A(new_n11832), .B(new_n11833), .C(new_n11831), .Y(new_n11839));
  OAI21xp33_ASAP7_75t_L     g11583(.A1(new_n11822), .A2(new_n11820), .B(new_n11829), .Y(new_n11840));
  NAND2xp33_ASAP7_75t_L     g11584(.A(new_n11839), .B(new_n11840), .Y(new_n11841));
  INVx1_ASAP7_75t_L         g11585(.A(new_n11836), .Y(new_n11842));
  A2O1A1Ixp33_ASAP7_75t_L   g11586(.A1(new_n11499), .A2(new_n11493), .B(new_n11501), .C(new_n11842), .Y(new_n11843));
  NAND2xp33_ASAP7_75t_L     g11587(.A(new_n11843), .B(new_n11841), .Y(new_n11844));
  NAND2xp33_ASAP7_75t_L     g11588(.A(\b[41] ), .B(new_n1548), .Y(new_n11845));
  NAND2xp33_ASAP7_75t_L     g11589(.A(\b[42] ), .B(new_n1410), .Y(new_n11846));
  AOI22xp33_ASAP7_75t_L     g11590(.A1(new_n1406), .A2(\b[43] ), .B1(new_n1404), .B2(new_n6202), .Y(new_n11847));
  NAND4xp25_ASAP7_75t_L     g11591(.A(new_n11847), .B(\a[20] ), .C(new_n11845), .D(new_n11846), .Y(new_n11848));
  NAND2xp33_ASAP7_75t_L     g11592(.A(new_n11846), .B(new_n11847), .Y(new_n11849));
  A2O1A1Ixp33_ASAP7_75t_L   g11593(.A1(\b[41] ), .A2(new_n1548), .B(new_n11849), .C(new_n1401), .Y(new_n11850));
  NAND2xp33_ASAP7_75t_L     g11594(.A(new_n11848), .B(new_n11850), .Y(new_n11851));
  AOI21xp33_ASAP7_75t_L     g11595(.A1(new_n11838), .A2(new_n11844), .B(new_n11851), .Y(new_n11852));
  NOR2xp33_ASAP7_75t_L      g11596(.A(new_n11843), .B(new_n11841), .Y(new_n11853));
  NOR2xp33_ASAP7_75t_L      g11597(.A(new_n11837), .B(new_n11835), .Y(new_n11854));
  INVx1_ASAP7_75t_L         g11598(.A(new_n11851), .Y(new_n11855));
  NOR3xp33_ASAP7_75t_L      g11599(.A(new_n11854), .B(new_n11853), .C(new_n11855), .Y(new_n11856));
  NOR3xp33_ASAP7_75t_L      g11600(.A(new_n11856), .B(new_n11852), .C(new_n11606), .Y(new_n11857));
  OA21x2_ASAP7_75t_L        g11601(.A1(new_n11852), .A2(new_n11856), .B(new_n11606), .Y(new_n11858));
  NOR3xp33_ASAP7_75t_L      g11602(.A(new_n11858), .B(new_n11857), .C(new_n11604), .Y(new_n11859));
  INVx1_ASAP7_75t_L         g11603(.A(new_n11604), .Y(new_n11860));
  OR3x1_ASAP7_75t_L         g11604(.A(new_n11856), .B(new_n11852), .C(new_n11606), .Y(new_n11861));
  OAI21xp33_ASAP7_75t_L     g11605(.A1(new_n11852), .A2(new_n11856), .B(new_n11606), .Y(new_n11862));
  AOI21xp33_ASAP7_75t_L     g11606(.A1(new_n11861), .A2(new_n11862), .B(new_n11860), .Y(new_n11863));
  NOR3xp33_ASAP7_75t_L      g11607(.A(new_n11598), .B(new_n11859), .C(new_n11863), .Y(new_n11864));
  INVx1_ASAP7_75t_L         g11608(.A(new_n11597), .Y(new_n11865));
  A2O1A1Ixp33_ASAP7_75t_L   g11609(.A1(new_n11527), .A2(new_n11528), .B(new_n11273), .C(new_n11865), .Y(new_n11866));
  NAND3xp33_ASAP7_75t_L     g11610(.A(new_n11861), .B(new_n11860), .C(new_n11862), .Y(new_n11867));
  INVx1_ASAP7_75t_L         g11611(.A(new_n11863), .Y(new_n11868));
  AOI21xp33_ASAP7_75t_L     g11612(.A1(new_n11868), .A2(new_n11867), .B(new_n11866), .Y(new_n11869));
  OAI21xp33_ASAP7_75t_L     g11613(.A1(new_n11869), .A2(new_n11864), .B(new_n11596), .Y(new_n11870));
  NAND3xp33_ASAP7_75t_L     g11614(.A(new_n11866), .B(new_n11867), .C(new_n11868), .Y(new_n11871));
  OAI21xp33_ASAP7_75t_L     g11615(.A1(new_n11859), .A2(new_n11863), .B(new_n11598), .Y(new_n11872));
  NAND3xp33_ASAP7_75t_L     g11616(.A(new_n11871), .B(new_n11595), .C(new_n11872), .Y(new_n11873));
  NAND3xp33_ASAP7_75t_L     g11617(.A(new_n11588), .B(new_n11870), .C(new_n11873), .Y(new_n11874));
  AOI21xp33_ASAP7_75t_L     g11618(.A1(new_n11537), .A2(new_n11536), .B(new_n11586), .Y(new_n11875));
  NAND2xp33_ASAP7_75t_L     g11619(.A(new_n11873), .B(new_n11870), .Y(new_n11876));
  NAND2xp33_ASAP7_75t_L     g11620(.A(new_n11875), .B(new_n11876), .Y(new_n11877));
  AOI21xp33_ASAP7_75t_L     g11621(.A1(new_n11877), .A2(new_n11874), .B(new_n11585), .Y(new_n11878));
  NOR2xp33_ASAP7_75t_L      g11622(.A(new_n11875), .B(new_n11876), .Y(new_n11879));
  AOI21xp33_ASAP7_75t_L     g11623(.A1(new_n11873), .A2(new_n11870), .B(new_n11588), .Y(new_n11880));
  NOR3xp33_ASAP7_75t_L      g11624(.A(new_n11879), .B(new_n11880), .C(new_n11584), .Y(new_n11881));
  NOR2xp33_ASAP7_75t_L      g11625(.A(new_n11878), .B(new_n11881), .Y(new_n11882));
  A2O1A1Ixp33_ASAP7_75t_L   g11626(.A1(new_n11544), .A2(new_n11257), .B(new_n11577), .C(new_n11882), .Y(new_n11883));
  O2A1O1Ixp33_ASAP7_75t_L   g11627(.A1(new_n11547), .A2(new_n11548), .B(new_n11257), .C(new_n11577), .Y(new_n11884));
  OAI21xp33_ASAP7_75t_L     g11628(.A1(new_n11880), .A2(new_n11879), .B(new_n11584), .Y(new_n11885));
  NAND3xp33_ASAP7_75t_L     g11629(.A(new_n11877), .B(new_n11874), .C(new_n11585), .Y(new_n11886));
  NAND2xp33_ASAP7_75t_L     g11630(.A(new_n11886), .B(new_n11885), .Y(new_n11887));
  NAND2xp33_ASAP7_75t_L     g11631(.A(new_n11884), .B(new_n11887), .Y(new_n11888));
  AOI22xp33_ASAP7_75t_L     g11632(.A1(new_n451), .A2(\b[55] ), .B1(new_n448), .B2(new_n9542), .Y(new_n11889));
  OAI221xp5_ASAP7_75t_L     g11633(.A1(new_n529), .A2(new_n9199), .B1(new_n8882), .B2(new_n481), .C(new_n11889), .Y(new_n11890));
  XNOR2x2_ASAP7_75t_L       g11634(.A(\a[8] ), .B(new_n11890), .Y(new_n11891));
  NAND3xp33_ASAP7_75t_L     g11635(.A(new_n11883), .B(new_n11891), .C(new_n11888), .Y(new_n11892));
  INVx1_ASAP7_75t_L         g11636(.A(new_n11577), .Y(new_n11893));
  O2A1O1Ixp33_ASAP7_75t_L   g11637(.A1(new_n11546), .A2(new_n11549), .B(new_n11893), .C(new_n11887), .Y(new_n11894));
  A2O1A1Ixp33_ASAP7_75t_L   g11638(.A1(new_n11539), .A2(new_n11543), .B(new_n11546), .C(new_n11893), .Y(new_n11895));
  NOR2xp33_ASAP7_75t_L      g11639(.A(new_n11895), .B(new_n11882), .Y(new_n11896));
  INVx1_ASAP7_75t_L         g11640(.A(new_n11891), .Y(new_n11897));
  OAI21xp33_ASAP7_75t_L     g11641(.A1(new_n11896), .A2(new_n11894), .B(new_n11897), .Y(new_n11898));
  AOI21xp33_ASAP7_75t_L     g11642(.A1(new_n11247), .A2(new_n11554), .B(new_n11556), .Y(new_n11899));
  NAND3xp33_ASAP7_75t_L     g11643(.A(new_n11899), .B(new_n11892), .C(new_n11898), .Y(new_n11900));
  AO21x2_ASAP7_75t_L        g11644(.A1(new_n11892), .A2(new_n11898), .B(new_n11899), .Y(new_n11901));
  AOI22xp33_ASAP7_75t_L     g11645(.A1(new_n345), .A2(\b[58] ), .B1(new_n342), .B2(new_n10857), .Y(new_n11902));
  OAI221xp5_ASAP7_75t_L     g11646(.A1(new_n406), .A2(new_n10488), .B1(new_n10178), .B2(new_n365), .C(new_n11902), .Y(new_n11903));
  XNOR2x2_ASAP7_75t_L       g11647(.A(\a[5] ), .B(new_n11903), .Y(new_n11904));
  INVx1_ASAP7_75t_L         g11648(.A(new_n11904), .Y(new_n11905));
  AOI21xp33_ASAP7_75t_L     g11649(.A1(new_n11901), .A2(new_n11900), .B(new_n11905), .Y(new_n11906));
  AND3x1_ASAP7_75t_L        g11650(.A(new_n11899), .B(new_n11898), .C(new_n11892), .Y(new_n11907));
  AOI21xp33_ASAP7_75t_L     g11651(.A1(new_n11892), .A2(new_n11898), .B(new_n11899), .Y(new_n11908));
  NOR3xp33_ASAP7_75t_L      g11652(.A(new_n11907), .B(new_n11904), .C(new_n11908), .Y(new_n11909));
  NOR2xp33_ASAP7_75t_L      g11653(.A(\b[60] ), .B(\b[61] ), .Y(new_n11910));
  INVx1_ASAP7_75t_L         g11654(.A(\b[61] ), .Y(new_n11911));
  NOR2xp33_ASAP7_75t_L      g11655(.A(new_n11226), .B(new_n11911), .Y(new_n11912));
  NOR2xp33_ASAP7_75t_L      g11656(.A(new_n11910), .B(new_n11912), .Y(new_n11913));
  A2O1A1Ixp33_ASAP7_75t_L   g11657(.A1(\b[60] ), .A2(\b[59] ), .B(new_n11230), .C(new_n11913), .Y(new_n11914));
  INVx1_ASAP7_75t_L         g11658(.A(new_n11227), .Y(new_n11915));
  A2O1A1Ixp33_ASAP7_75t_L   g11659(.A1(new_n10884), .A2(new_n11224), .B(new_n11225), .C(new_n11915), .Y(new_n11916));
  NOR2xp33_ASAP7_75t_L      g11660(.A(new_n11913), .B(new_n11916), .Y(new_n11917));
  INVx1_ASAP7_75t_L         g11661(.A(new_n11917), .Y(new_n11918));
  AND2x2_ASAP7_75t_L        g11662(.A(new_n11914), .B(new_n11918), .Y(new_n11919));
  INVx1_ASAP7_75t_L         g11663(.A(new_n11919), .Y(new_n11920));
  NOR2xp33_ASAP7_75t_L      g11664(.A(new_n11226), .B(new_n261), .Y(new_n11921));
  AOI221xp5_ASAP7_75t_L     g11665(.A1(\b[59] ), .A2(new_n291), .B1(\b[61] ), .B2(new_n272), .C(new_n11921), .Y(new_n11922));
  OAI211xp5_ASAP7_75t_L     g11666(.A1(new_n292), .A2(new_n11920), .B(\a[2] ), .C(new_n11922), .Y(new_n11923));
  INVx1_ASAP7_75t_L         g11667(.A(new_n11922), .Y(new_n11924));
  A2O1A1Ixp33_ASAP7_75t_L   g11668(.A1(new_n11919), .A2(new_n269), .B(new_n11924), .C(new_n265), .Y(new_n11925));
  NAND2xp33_ASAP7_75t_L     g11669(.A(new_n11925), .B(new_n11923), .Y(new_n11926));
  NOR3xp33_ASAP7_75t_L      g11670(.A(new_n11909), .B(new_n11906), .C(new_n11926), .Y(new_n11927));
  OAI21xp33_ASAP7_75t_L     g11671(.A1(new_n11908), .A2(new_n11907), .B(new_n11904), .Y(new_n11928));
  NAND3xp33_ASAP7_75t_L     g11672(.A(new_n11901), .B(new_n11905), .C(new_n11900), .Y(new_n11929));
  INVx1_ASAP7_75t_L         g11673(.A(new_n11926), .Y(new_n11930));
  AOI21xp33_ASAP7_75t_L     g11674(.A1(new_n11928), .A2(new_n11929), .B(new_n11930), .Y(new_n11931));
  O2A1O1Ixp33_ASAP7_75t_L   g11675(.A1(new_n11240), .A2(new_n11238), .B(new_n11560), .C(new_n11562), .Y(new_n11932));
  INVx1_ASAP7_75t_L         g11676(.A(new_n11932), .Y(new_n11933));
  NOR3xp33_ASAP7_75t_L      g11677(.A(new_n11927), .B(new_n11931), .C(new_n11933), .Y(new_n11934));
  NAND3xp33_ASAP7_75t_L     g11678(.A(new_n11928), .B(new_n11929), .C(new_n11930), .Y(new_n11935));
  OAI21xp33_ASAP7_75t_L     g11679(.A1(new_n11906), .A2(new_n11909), .B(new_n11926), .Y(new_n11936));
  AOI21xp33_ASAP7_75t_L     g11680(.A1(new_n11936), .A2(new_n11935), .B(new_n11932), .Y(new_n11937));
  NOR2xp33_ASAP7_75t_L      g11681(.A(new_n11937), .B(new_n11934), .Y(new_n11938));
  INVx1_ASAP7_75t_L         g11682(.A(new_n11938), .Y(new_n11939));
  O2A1O1Ixp33_ASAP7_75t_L   g11683(.A1(new_n11576), .A2(new_n11570), .B(new_n11565), .C(new_n11939), .Y(new_n11940));
  A2O1A1Ixp33_ASAP7_75t_L   g11684(.A1(new_n11222), .A2(new_n11573), .B(new_n11570), .C(new_n11565), .Y(new_n11941));
  NOR2xp33_ASAP7_75t_L      g11685(.A(new_n11938), .B(new_n11941), .Y(new_n11942));
  NOR2xp33_ASAP7_75t_L      g11686(.A(new_n11942), .B(new_n11940), .Y(\f[61] ));
  NAND2xp33_ASAP7_75t_L     g11687(.A(new_n11938), .B(new_n11941), .Y(new_n11944));
  A2O1A1Ixp33_ASAP7_75t_L   g11688(.A1(new_n11936), .A2(new_n11935), .B(new_n11932), .C(new_n11944), .Y(new_n11945));
  A2O1A1O1Ixp25_ASAP7_75t_L g11689(.A1(new_n11257), .A2(new_n11544), .B(new_n11577), .C(new_n11885), .D(new_n11881), .Y(new_n11946));
  NAND2xp33_ASAP7_75t_L     g11690(.A(\b[52] ), .B(new_n590), .Y(new_n11947));
  AOI22xp33_ASAP7_75t_L     g11691(.A1(new_n600), .A2(\b[53] ), .B1(new_n597), .B2(new_n8889), .Y(new_n11948));
  NAND2xp33_ASAP7_75t_L     g11692(.A(new_n11947), .B(new_n11948), .Y(new_n11949));
  AOI211xp5_ASAP7_75t_L     g11693(.A1(\b[51] ), .A2(new_n674), .B(new_n594), .C(new_n11949), .Y(new_n11950));
  INVx1_ASAP7_75t_L         g11694(.A(new_n11949), .Y(new_n11951));
  O2A1O1Ixp33_ASAP7_75t_L   g11695(.A1(new_n8249), .A2(new_n1620), .B(new_n11951), .C(\a[11] ), .Y(new_n11952));
  NOR2xp33_ASAP7_75t_L      g11696(.A(new_n11950), .B(new_n11952), .Y(new_n11953));
  NOR3xp33_ASAP7_75t_L      g11697(.A(new_n11864), .B(new_n11869), .C(new_n11596), .Y(new_n11954));
  A2O1A1O1Ixp25_ASAP7_75t_L g11698(.A1(new_n11536), .A2(new_n11537), .B(new_n11586), .C(new_n11870), .D(new_n11954), .Y(new_n11955));
  NOR2xp33_ASAP7_75t_L      g11699(.A(new_n6756), .B(new_n1195), .Y(new_n11956));
  INVx1_ASAP7_75t_L         g11700(.A(new_n11956), .Y(new_n11957));
  NAND2xp33_ASAP7_75t_L     g11701(.A(\b[46] ), .B(new_n1103), .Y(new_n11958));
  AOI22xp33_ASAP7_75t_L     g11702(.A1(new_n1113), .A2(\b[47] ), .B1(new_n1110), .B2(new_n7323), .Y(new_n11959));
  AND4x1_ASAP7_75t_L        g11703(.A(new_n11959), .B(new_n11958), .C(new_n11957), .D(\a[17] ), .Y(new_n11960));
  AOI31xp33_ASAP7_75t_L     g11704(.A1(new_n11959), .A2(new_n11958), .A3(new_n11957), .B(\a[17] ), .Y(new_n11961));
  NOR2xp33_ASAP7_75t_L      g11705(.A(new_n11961), .B(new_n11960), .Y(new_n11962));
  NAND2xp33_ASAP7_75t_L     g11706(.A(\b[44] ), .B(new_n1406), .Y(new_n11963));
  OAI221xp5_ASAP7_75t_L     g11707(.A1(new_n6195), .A2(new_n1398), .B1(new_n1411), .B2(new_n6229), .C(new_n11963), .Y(new_n11964));
  AOI21xp33_ASAP7_75t_L     g11708(.A1(new_n1548), .A2(\b[42] ), .B(new_n11964), .Y(new_n11965));
  NAND2xp33_ASAP7_75t_L     g11709(.A(\a[20] ), .B(new_n11965), .Y(new_n11966));
  A2O1A1Ixp33_ASAP7_75t_L   g11710(.A1(\b[42] ), .A2(new_n1548), .B(new_n11964), .C(new_n1401), .Y(new_n11967));
  NAND2xp33_ASAP7_75t_L     g11711(.A(new_n11967), .B(new_n11966), .Y(new_n11968));
  INVx1_ASAP7_75t_L         g11712(.A(new_n11968), .Y(new_n11969));
  NOR3xp33_ASAP7_75t_L      g11713(.A(new_n11820), .B(new_n11822), .C(new_n11833), .Y(new_n11970));
  O2A1O1Ixp33_ASAP7_75t_L   g11714(.A1(new_n11830), .A2(new_n11834), .B(new_n11843), .C(new_n11970), .Y(new_n11971));
  AOI21xp33_ASAP7_75t_L     g11715(.A1(new_n11798), .A2(new_n11799), .B(new_n11800), .Y(new_n11972));
  A2O1A1O1Ixp25_ASAP7_75t_L g11716(.A1(new_n11473), .A2(new_n11474), .B(new_n11608), .C(new_n11801), .D(new_n11972), .Y(new_n11973));
  NAND2xp33_ASAP7_75t_L     g11717(.A(\b[35] ), .B(new_n2702), .Y(new_n11974));
  OAI221xp5_ASAP7_75t_L     g11718(.A1(new_n3827), .A2(new_n2694), .B1(new_n2707), .B2(new_n4060), .C(new_n11974), .Y(new_n11975));
  AOI21xp33_ASAP7_75t_L     g11719(.A1(new_n2931), .A2(\b[33] ), .B(new_n11975), .Y(new_n11976));
  NAND2xp33_ASAP7_75t_L     g11720(.A(\a[29] ), .B(new_n11976), .Y(new_n11977));
  A2O1A1Ixp33_ASAP7_75t_L   g11721(.A1(\b[33] ), .A2(new_n2931), .B(new_n11975), .C(new_n2697), .Y(new_n11978));
  NAND3xp33_ASAP7_75t_L     g11722(.A(new_n11782), .B(new_n11781), .C(new_n11779), .Y(new_n11979));
  OAI21xp33_ASAP7_75t_L     g11723(.A1(new_n11783), .A2(new_n11780), .B(new_n11786), .Y(new_n11980));
  NAND3xp33_ASAP7_75t_L     g11724(.A(new_n11729), .B(new_n11724), .C(new_n11614), .Y(new_n11981));
  NAND2xp33_ASAP7_75t_L     g11725(.A(\b[22] ), .B(new_n5240), .Y(new_n11982));
  OAI221xp5_ASAP7_75t_L     g11726(.A1(new_n5253), .A2(new_n1995), .B1(new_n5252), .B2(new_n4860), .C(new_n11982), .Y(new_n11983));
  AOI21xp33_ASAP7_75t_L     g11727(.A1(new_n5526), .A2(\b[21] ), .B(new_n11983), .Y(new_n11984));
  NAND2xp33_ASAP7_75t_L     g11728(.A(\a[41] ), .B(new_n11984), .Y(new_n11985));
  A2O1A1Ixp33_ASAP7_75t_L   g11729(.A1(\b[21] ), .A2(new_n5526), .B(new_n11983), .C(new_n5244), .Y(new_n11986));
  NAND2xp33_ASAP7_75t_L     g11730(.A(new_n11986), .B(new_n11985), .Y(new_n11987));
  NOR2xp33_ASAP7_75t_L      g11731(.A(new_n1356), .B(new_n6309), .Y(new_n11988));
  NAND2xp33_ASAP7_75t_L     g11732(.A(\b[19] ), .B(new_n5992), .Y(new_n11989));
  OAI221xp5_ASAP7_75t_L     g11733(.A1(new_n6312), .A2(new_n1594), .B1(new_n6311), .B2(new_n3001), .C(new_n11989), .Y(new_n11990));
  OR3x1_ASAP7_75t_L         g11734(.A(new_n11990), .B(new_n5996), .C(new_n11988), .Y(new_n11991));
  A2O1A1Ixp33_ASAP7_75t_L   g11735(.A1(\b[18] ), .A2(new_n6308), .B(new_n11990), .C(new_n5996), .Y(new_n11992));
  NAND2xp33_ASAP7_75t_L     g11736(.A(new_n11992), .B(new_n11991), .Y(new_n11993));
  AOI21xp33_ASAP7_75t_L     g11737(.A1(new_n11706), .A2(new_n11710), .B(new_n11625), .Y(new_n11994));
  NAND2xp33_ASAP7_75t_L     g11738(.A(\b[16] ), .B(new_n6812), .Y(new_n11995));
  OAI221xp5_ASAP7_75t_L     g11739(.A1(new_n7118), .A2(new_n1244), .B1(new_n7117), .B2(new_n1251), .C(new_n11995), .Y(new_n11996));
  AOI21xp33_ASAP7_75t_L     g11740(.A1(new_n7124), .A2(\b[15] ), .B(new_n11996), .Y(new_n11997));
  NAND2xp33_ASAP7_75t_L     g11741(.A(\a[47] ), .B(new_n11997), .Y(new_n11998));
  A2O1A1Ixp33_ASAP7_75t_L   g11742(.A1(\b[15] ), .A2(new_n7124), .B(new_n11996), .C(new_n6816), .Y(new_n11999));
  NAND2xp33_ASAP7_75t_L     g11743(.A(new_n11999), .B(new_n11998), .Y(new_n12000));
  NAND2xp33_ASAP7_75t_L     g11744(.A(new_n11685), .B(new_n11686), .Y(new_n12001));
  MAJIxp5_ASAP7_75t_L       g11745(.A(new_n11693), .B(new_n11687), .C(new_n12001), .Y(new_n12002));
  NAND2xp33_ASAP7_75t_L     g11746(.A(\b[10] ), .B(new_n8635), .Y(new_n12003));
  OAI221xp5_ASAP7_75t_L     g11747(.A1(new_n8968), .A2(new_n695), .B1(new_n8967), .B2(new_n701), .C(new_n12003), .Y(new_n12004));
  AOI21xp33_ASAP7_75t_L     g11748(.A1(new_n8964), .A2(\b[9] ), .B(new_n12004), .Y(new_n12005));
  NAND2xp33_ASAP7_75t_L     g11749(.A(\a[53] ), .B(new_n12005), .Y(new_n12006));
  A2O1A1Ixp33_ASAP7_75t_L   g11750(.A1(\b[9] ), .A2(new_n8964), .B(new_n12004), .C(new_n8639), .Y(new_n12007));
  NAND2xp33_ASAP7_75t_L     g11751(.A(new_n12007), .B(new_n12006), .Y(new_n12008));
  OAI21xp33_ASAP7_75t_L     g11752(.A1(new_n11668), .A2(new_n11630), .B(new_n11669), .Y(new_n12009));
  INVx1_ASAP7_75t_L         g11753(.A(new_n9948), .Y(new_n12010));
  AOI22xp33_ASAP7_75t_L     g11754(.A1(new_n9623), .A2(\b[8] ), .B1(new_n9620), .B2(new_n510), .Y(new_n12011));
  OAI221xp5_ASAP7_75t_L     g11755(.A1(new_n10280), .A2(new_n421), .B1(new_n382), .B2(new_n12010), .C(new_n12011), .Y(new_n12012));
  NOR2xp33_ASAP7_75t_L      g11756(.A(new_n9610), .B(new_n12012), .Y(new_n12013));
  INVx1_ASAP7_75t_L         g11757(.A(new_n12013), .Y(new_n12014));
  NAND2xp33_ASAP7_75t_L     g11758(.A(new_n9610), .B(new_n12012), .Y(new_n12015));
  AOI22xp33_ASAP7_75t_L     g11759(.A1(new_n10594), .A2(\b[5] ), .B1(new_n10591), .B2(new_n360), .Y(new_n12016));
  OAI221xp5_ASAP7_75t_L     g11760(.A1(new_n11335), .A2(new_n323), .B1(new_n299), .B2(new_n11330), .C(new_n12016), .Y(new_n12017));
  XNOR2x2_ASAP7_75t_L       g11761(.A(new_n10588), .B(new_n12017), .Y(new_n12018));
  INVx1_ASAP7_75t_L         g11762(.A(new_n11658), .Y(new_n12019));
  INVx1_ASAP7_75t_L         g11763(.A(new_n11646), .Y(new_n12020));
  NOR3xp33_ASAP7_75t_L      g11764(.A(new_n11653), .B(new_n12020), .C(new_n11645), .Y(new_n12021));
  INVx1_ASAP7_75t_L         g11765(.A(new_n11654), .Y(new_n12022));
  INVx1_ASAP7_75t_L         g11766(.A(new_n11656), .Y(new_n12023));
  NAND2xp33_ASAP7_75t_L     g11767(.A(\b[1] ), .B(new_n11647), .Y(new_n12024));
  OAI221xp5_ASAP7_75t_L     g11768(.A1(new_n12023), .A2(new_n278), .B1(new_n283), .B2(new_n12022), .C(new_n12024), .Y(new_n12025));
  AOI21xp33_ASAP7_75t_L     g11769(.A1(new_n12021), .A2(\b[0] ), .B(new_n12025), .Y(new_n12026));
  A2O1A1Ixp33_ASAP7_75t_L   g11770(.A1(new_n11328), .A2(new_n12019), .B(new_n11651), .C(new_n12026), .Y(new_n12027));
  O2A1O1Ixp33_ASAP7_75t_L   g11771(.A1(new_n258), .A2(new_n11326), .B(new_n12019), .C(new_n11651), .Y(new_n12028));
  A2O1A1Ixp33_ASAP7_75t_L   g11772(.A1(\b[0] ), .A2(new_n12021), .B(new_n12025), .C(new_n12028), .Y(new_n12029));
  AND2x2_ASAP7_75t_L        g11773(.A(new_n12027), .B(new_n12029), .Y(new_n12030));
  NOR2xp33_ASAP7_75t_L      g11774(.A(new_n12018), .B(new_n12030), .Y(new_n12031));
  XNOR2x2_ASAP7_75t_L       g11775(.A(\a[59] ), .B(new_n12017), .Y(new_n12032));
  NAND2xp33_ASAP7_75t_L     g11776(.A(new_n12027), .B(new_n12029), .Y(new_n12033));
  NOR2xp33_ASAP7_75t_L      g11777(.A(new_n12033), .B(new_n12032), .Y(new_n12034));
  NOR2xp33_ASAP7_75t_L      g11778(.A(new_n12034), .B(new_n12031), .Y(new_n12035));
  NAND3xp33_ASAP7_75t_L     g11779(.A(new_n12035), .B(new_n11663), .C(new_n11662), .Y(new_n12036));
  NAND2xp33_ASAP7_75t_L     g11780(.A(new_n12033), .B(new_n12032), .Y(new_n12037));
  NAND2xp33_ASAP7_75t_L     g11781(.A(new_n12018), .B(new_n12030), .Y(new_n12038));
  NAND2xp33_ASAP7_75t_L     g11782(.A(new_n12037), .B(new_n12038), .Y(new_n12039));
  A2O1A1Ixp33_ASAP7_75t_L   g11783(.A1(new_n11661), .A2(new_n11639), .B(new_n11666), .C(new_n12039), .Y(new_n12040));
  NAND4xp25_ASAP7_75t_L     g11784(.A(new_n12036), .B(new_n12014), .C(new_n12040), .D(new_n12015), .Y(new_n12041));
  INVx1_ASAP7_75t_L         g11785(.A(new_n12015), .Y(new_n12042));
  A2O1A1Ixp33_ASAP7_75t_L   g11786(.A1(new_n11342), .A2(new_n11638), .B(new_n11660), .C(new_n11662), .Y(new_n12043));
  NOR2xp33_ASAP7_75t_L      g11787(.A(new_n12043), .B(new_n12039), .Y(new_n12044));
  O2A1O1Ixp33_ASAP7_75t_L   g11788(.A1(new_n11665), .A2(new_n11660), .B(new_n11662), .C(new_n12035), .Y(new_n12045));
  OAI22xp33_ASAP7_75t_L     g11789(.A1(new_n12045), .A2(new_n12044), .B1(new_n12042), .B2(new_n12013), .Y(new_n12046));
  NAND3xp33_ASAP7_75t_L     g11790(.A(new_n12046), .B(new_n12009), .C(new_n12041), .Y(new_n12047));
  AO21x2_ASAP7_75t_L        g11791(.A1(new_n12041), .A2(new_n12046), .B(new_n12009), .Y(new_n12048));
  AO21x2_ASAP7_75t_L        g11792(.A1(new_n12047), .A2(new_n12048), .B(new_n12008), .Y(new_n12049));
  NAND3xp33_ASAP7_75t_L     g11793(.A(new_n12048), .B(new_n12047), .C(new_n12008), .Y(new_n12050));
  NAND3xp33_ASAP7_75t_L     g11794(.A(new_n12049), .B(new_n12002), .C(new_n12050), .Y(new_n12051));
  NOR2xp33_ASAP7_75t_L      g11795(.A(new_n11676), .B(new_n11671), .Y(new_n12052));
  MAJIxp5_ASAP7_75t_L       g11796(.A(new_n11689), .B(new_n11683), .C(new_n12052), .Y(new_n12053));
  AOI21xp33_ASAP7_75t_L     g11797(.A1(new_n12048), .A2(new_n12047), .B(new_n12008), .Y(new_n12054));
  AND3x1_ASAP7_75t_L        g11798(.A(new_n12048), .B(new_n12047), .C(new_n12008), .Y(new_n12055));
  OAI21xp33_ASAP7_75t_L     g11799(.A1(new_n12054), .A2(new_n12055), .B(new_n12053), .Y(new_n12056));
  NAND2xp33_ASAP7_75t_L     g11800(.A(\b[13] ), .B(new_n7649), .Y(new_n12057));
  OAI221xp5_ASAP7_75t_L     g11801(.A1(new_n7997), .A2(new_n871), .B1(new_n7996), .B2(new_n878), .C(new_n12057), .Y(new_n12058));
  AOI21xp33_ASAP7_75t_L     g11802(.A1(new_n7993), .A2(\b[12] ), .B(new_n12058), .Y(new_n12059));
  NAND2xp33_ASAP7_75t_L     g11803(.A(\a[50] ), .B(new_n12059), .Y(new_n12060));
  A2O1A1Ixp33_ASAP7_75t_L   g11804(.A1(\b[12] ), .A2(new_n7993), .B(new_n12058), .C(new_n7653), .Y(new_n12061));
  AND2x2_ASAP7_75t_L        g11805(.A(new_n12061), .B(new_n12060), .Y(new_n12062));
  NAND3xp33_ASAP7_75t_L     g11806(.A(new_n12062), .B(new_n12056), .C(new_n12051), .Y(new_n12063));
  AO21x2_ASAP7_75t_L        g11807(.A1(new_n12051), .A2(new_n12056), .B(new_n12062), .Y(new_n12064));
  A2O1A1Ixp33_ASAP7_75t_L   g11808(.A1(new_n11373), .A2(new_n11316), .B(new_n11381), .C(new_n11699), .Y(new_n12065));
  AOI22xp33_ASAP7_75t_L     g11809(.A1(new_n12064), .A2(new_n12063), .B1(new_n11705), .B2(new_n12065), .Y(new_n12066));
  AND3x1_ASAP7_75t_L        g11810(.A(new_n12062), .B(new_n12056), .C(new_n12051), .Y(new_n12067));
  AOI21xp33_ASAP7_75t_L     g11811(.A1(new_n12056), .A2(new_n12051), .B(new_n12062), .Y(new_n12068));
  O2A1O1Ixp33_ASAP7_75t_L   g11812(.A1(new_n11380), .A2(new_n11379), .B(new_n11377), .C(new_n11708), .Y(new_n12069));
  NOR4xp25_ASAP7_75t_L      g11813(.A(new_n12069), .B(new_n12067), .C(new_n11709), .D(new_n12068), .Y(new_n12070));
  OAI21xp33_ASAP7_75t_L     g11814(.A1(new_n12066), .A2(new_n12070), .B(new_n12000), .Y(new_n12071));
  AND2x2_ASAP7_75t_L        g11815(.A(new_n11999), .B(new_n11998), .Y(new_n12072));
  OAI22xp33_ASAP7_75t_L     g11816(.A1(new_n12069), .A2(new_n11709), .B1(new_n12067), .B2(new_n12068), .Y(new_n12073));
  NAND4xp25_ASAP7_75t_L     g11817(.A(new_n12065), .B(new_n12064), .C(new_n11705), .D(new_n12063), .Y(new_n12074));
  NAND3xp33_ASAP7_75t_L     g11818(.A(new_n12073), .B(new_n12072), .C(new_n12074), .Y(new_n12075));
  NAND2xp33_ASAP7_75t_L     g11819(.A(new_n12075), .B(new_n12071), .Y(new_n12076));
  A2O1A1Ixp33_ASAP7_75t_L   g11820(.A1(new_n11712), .A2(new_n11620), .B(new_n11994), .C(new_n12076), .Y(new_n12077));
  INVx1_ASAP7_75t_L         g11821(.A(new_n11383), .Y(new_n12078));
  A2O1A1O1Ixp25_ASAP7_75t_L g11822(.A1(new_n11384), .A2(new_n11307), .B(new_n12078), .C(new_n11712), .D(new_n11994), .Y(new_n12079));
  AOI21xp33_ASAP7_75t_L     g11823(.A1(new_n12073), .A2(new_n12074), .B(new_n12072), .Y(new_n12080));
  NOR3xp33_ASAP7_75t_L      g11824(.A(new_n12070), .B(new_n12066), .C(new_n12000), .Y(new_n12081));
  NOR2xp33_ASAP7_75t_L      g11825(.A(new_n12080), .B(new_n12081), .Y(new_n12082));
  NAND2xp33_ASAP7_75t_L     g11826(.A(new_n12079), .B(new_n12082), .Y(new_n12083));
  NAND3xp33_ASAP7_75t_L     g11827(.A(new_n12077), .B(new_n12083), .C(new_n11993), .Y(new_n12084));
  AND2x2_ASAP7_75t_L        g11828(.A(new_n11992), .B(new_n11991), .Y(new_n12085));
  NOR2xp33_ASAP7_75t_L      g11829(.A(new_n12079), .B(new_n12082), .Y(new_n12086));
  AO21x2_ASAP7_75t_L        g11830(.A1(new_n11712), .A2(new_n11620), .B(new_n11994), .Y(new_n12087));
  NOR2xp33_ASAP7_75t_L      g11831(.A(new_n12087), .B(new_n12076), .Y(new_n12088));
  OAI21xp33_ASAP7_75t_L     g11832(.A1(new_n12088), .A2(new_n12086), .B(new_n12085), .Y(new_n12089));
  A2O1A1Ixp33_ASAP7_75t_L   g11833(.A1(new_n11392), .A2(new_n11616), .B(new_n11720), .C(new_n11727), .Y(new_n12090));
  NAND3xp33_ASAP7_75t_L     g11834(.A(new_n12090), .B(new_n12089), .C(new_n12084), .Y(new_n12091));
  NAND2xp33_ASAP7_75t_L     g11835(.A(new_n12084), .B(new_n12089), .Y(new_n12092));
  A2O1A1O1Ixp25_ASAP7_75t_L g11836(.A1(new_n11301), .A2(new_n11725), .B(new_n11617), .C(new_n11726), .D(new_n11722), .Y(new_n12093));
  NAND2xp33_ASAP7_75t_L     g11837(.A(new_n12093), .B(new_n12092), .Y(new_n12094));
  NAND3xp33_ASAP7_75t_L     g11838(.A(new_n12094), .B(new_n12091), .C(new_n11987), .Y(new_n12095));
  AND2x2_ASAP7_75t_L        g11839(.A(new_n11986), .B(new_n11985), .Y(new_n12096));
  O2A1O1Ixp33_ASAP7_75t_L   g11840(.A1(new_n11618), .A2(new_n11720), .B(new_n11727), .C(new_n12092), .Y(new_n12097));
  AOI21xp33_ASAP7_75t_L     g11841(.A1(new_n12089), .A2(new_n12084), .B(new_n12090), .Y(new_n12098));
  OAI21xp33_ASAP7_75t_L     g11842(.A1(new_n12098), .A2(new_n12097), .B(new_n12096), .Y(new_n12099));
  AOI221xp5_ASAP7_75t_L     g11843(.A1(new_n11738), .A2(new_n11981), .B1(new_n12095), .B2(new_n12099), .C(new_n11730), .Y(new_n12100));
  INVx1_ASAP7_75t_L         g11844(.A(new_n11730), .Y(new_n12101));
  NAND2xp33_ASAP7_75t_L     g11845(.A(new_n12095), .B(new_n12099), .Y(new_n12102));
  O2A1O1Ixp33_ASAP7_75t_L   g11846(.A1(new_n11611), .A2(new_n11736), .B(new_n12101), .C(new_n12102), .Y(new_n12103));
  OAI22xp33_ASAP7_75t_L     g11847(.A1(new_n2487), .A2(new_n4549), .B1(new_n4550), .B2(new_n2477), .Y(new_n12104));
  AOI221xp5_ASAP7_75t_L     g11848(.A1(\b[24] ), .A2(new_n4780), .B1(\b[25] ), .B2(new_n4548), .C(new_n12104), .Y(new_n12105));
  XNOR2x2_ASAP7_75t_L       g11849(.A(new_n4539), .B(new_n12105), .Y(new_n12106));
  INVx1_ASAP7_75t_L         g11850(.A(new_n12106), .Y(new_n12107));
  NOR3xp33_ASAP7_75t_L      g11851(.A(new_n12103), .B(new_n12107), .C(new_n12100), .Y(new_n12108));
  A2O1A1O1Ixp25_ASAP7_75t_L g11852(.A1(new_n11291), .A2(new_n11401), .B(new_n11610), .C(new_n11981), .D(new_n11730), .Y(new_n12109));
  NAND2xp33_ASAP7_75t_L     g11853(.A(new_n12109), .B(new_n12102), .Y(new_n12110));
  NOR3xp33_ASAP7_75t_L      g11854(.A(new_n12097), .B(new_n12098), .C(new_n12096), .Y(new_n12111));
  AOI21xp33_ASAP7_75t_L     g11855(.A1(new_n12094), .A2(new_n12091), .B(new_n11987), .Y(new_n12112));
  NOR2xp33_ASAP7_75t_L      g11856(.A(new_n12112), .B(new_n12111), .Y(new_n12113));
  A2O1A1Ixp33_ASAP7_75t_L   g11857(.A1(new_n11739), .A2(new_n11738), .B(new_n11730), .C(new_n12113), .Y(new_n12114));
  AOI21xp33_ASAP7_75t_L     g11858(.A1(new_n12114), .A2(new_n12110), .B(new_n12106), .Y(new_n12115));
  NOR2xp33_ASAP7_75t_L      g11859(.A(new_n12108), .B(new_n12115), .Y(new_n12116));
  NOR3xp33_ASAP7_75t_L      g11860(.A(new_n11745), .B(new_n11746), .C(new_n11743), .Y(new_n12117));
  O2A1O1Ixp33_ASAP7_75t_L   g11861(.A1(new_n11752), .A2(new_n11751), .B(new_n11753), .C(new_n12117), .Y(new_n12118));
  NAND2xp33_ASAP7_75t_L     g11862(.A(new_n12118), .B(new_n12116), .Y(new_n12119));
  NOR2xp33_ASAP7_75t_L      g11863(.A(new_n11746), .B(new_n11745), .Y(new_n12120));
  NAND3xp33_ASAP7_75t_L     g11864(.A(new_n12114), .B(new_n12110), .C(new_n12106), .Y(new_n12121));
  OAI21xp33_ASAP7_75t_L     g11865(.A1(new_n12100), .A2(new_n12103), .B(new_n12107), .Y(new_n12122));
  NAND2xp33_ASAP7_75t_L     g11866(.A(new_n12122), .B(new_n12121), .Y(new_n12123));
  A2O1A1Ixp33_ASAP7_75t_L   g11867(.A1(new_n11747), .A2(new_n12120), .B(new_n11760), .C(new_n12123), .Y(new_n12124));
  AOI22xp33_ASAP7_75t_L     g11868(.A1(new_n3884), .A2(\b[29] ), .B1(new_n3881), .B2(new_n5472), .Y(new_n12125));
  OAI221xp5_ASAP7_75t_L     g11869(.A1(new_n4312), .A2(new_n2852), .B1(new_n2650), .B2(new_n4986), .C(new_n12125), .Y(new_n12126));
  XNOR2x2_ASAP7_75t_L       g11870(.A(\a[35] ), .B(new_n12126), .Y(new_n12127));
  NAND3xp33_ASAP7_75t_L     g11871(.A(new_n12124), .B(new_n12119), .C(new_n12127), .Y(new_n12128));
  NOR3xp33_ASAP7_75t_L      g11872(.A(new_n12123), .B(new_n12117), .C(new_n11760), .Y(new_n12129));
  NOR2xp33_ASAP7_75t_L      g11873(.A(new_n12118), .B(new_n12116), .Y(new_n12130));
  INVx1_ASAP7_75t_L         g11874(.A(new_n12127), .Y(new_n12131));
  OAI21xp33_ASAP7_75t_L     g11875(.A1(new_n12130), .A2(new_n12129), .B(new_n12131), .Y(new_n12132));
  NAND2xp33_ASAP7_75t_L     g11876(.A(new_n12128), .B(new_n12132), .Y(new_n12133));
  NOR2xp33_ASAP7_75t_L      g11877(.A(new_n11759), .B(new_n11760), .Y(new_n12134));
  NAND2xp33_ASAP7_75t_L     g11878(.A(new_n11761), .B(new_n12134), .Y(new_n12135));
  A2O1A1Ixp33_ASAP7_75t_L   g11879(.A1(new_n11762), .A2(new_n11758), .B(new_n11771), .C(new_n12135), .Y(new_n12136));
  NOR2xp33_ASAP7_75t_L      g11880(.A(new_n12136), .B(new_n12133), .Y(new_n12137));
  NOR3xp33_ASAP7_75t_L      g11881(.A(new_n12129), .B(new_n12130), .C(new_n12131), .Y(new_n12138));
  AOI21xp33_ASAP7_75t_L     g11882(.A1(new_n12124), .A2(new_n12119), .B(new_n12127), .Y(new_n12139));
  NOR2xp33_ASAP7_75t_L      g11883(.A(new_n12139), .B(new_n12138), .Y(new_n12140));
  O2A1O1Ixp33_ASAP7_75t_L   g11884(.A1(new_n11771), .A2(new_n11770), .B(new_n12135), .C(new_n12140), .Y(new_n12141));
  AOI22xp33_ASAP7_75t_L     g11885(.A1(new_n3256), .A2(\b[32] ), .B1(new_n3254), .B2(new_n3450), .Y(new_n12142));
  OAI221xp5_ASAP7_75t_L     g11886(.A1(new_n3248), .A2(new_n3419), .B1(new_n3212), .B2(new_n3492), .C(new_n12142), .Y(new_n12143));
  XNOR2x2_ASAP7_75t_L       g11887(.A(\a[32] ), .B(new_n12143), .Y(new_n12144));
  OAI21xp33_ASAP7_75t_L     g11888(.A1(new_n12137), .A2(new_n12141), .B(new_n12144), .Y(new_n12145));
  NAND3xp33_ASAP7_75t_L     g11889(.A(new_n12140), .B(new_n11782), .C(new_n12135), .Y(new_n12146));
  A2O1A1Ixp33_ASAP7_75t_L   g11890(.A1(new_n11761), .A2(new_n12134), .B(new_n11772), .C(new_n12133), .Y(new_n12147));
  INVx1_ASAP7_75t_L         g11891(.A(new_n12144), .Y(new_n12148));
  NAND3xp33_ASAP7_75t_L     g11892(.A(new_n12146), .B(new_n12147), .C(new_n12148), .Y(new_n12149));
  NAND4xp25_ASAP7_75t_L     g11893(.A(new_n12145), .B(new_n12149), .C(new_n11979), .D(new_n11980), .Y(new_n12150));
  A2O1A1Ixp33_ASAP7_75t_L   g11894(.A1(new_n11788), .A2(new_n11787), .B(new_n11609), .C(new_n11979), .Y(new_n12151));
  AOI21xp33_ASAP7_75t_L     g11895(.A1(new_n12146), .A2(new_n12147), .B(new_n12148), .Y(new_n12152));
  NOR3xp33_ASAP7_75t_L      g11896(.A(new_n12141), .B(new_n12144), .C(new_n12137), .Y(new_n12153));
  OAI21xp33_ASAP7_75t_L     g11897(.A1(new_n12152), .A2(new_n12153), .B(new_n12151), .Y(new_n12154));
  AOI22xp33_ASAP7_75t_L     g11898(.A1(new_n11977), .A2(new_n11978), .B1(new_n12150), .B2(new_n12154), .Y(new_n12155));
  AND4x1_ASAP7_75t_L        g11899(.A(new_n12154), .B(new_n12150), .C(new_n11978), .D(new_n11977), .Y(new_n12156));
  OA21x2_ASAP7_75t_L        g11900(.A1(new_n12155), .A2(new_n12156), .B(new_n11973), .Y(new_n12157));
  NOR3xp33_ASAP7_75t_L      g11901(.A(new_n11973), .B(new_n12156), .C(new_n12155), .Y(new_n12158));
  NAND2xp33_ASAP7_75t_L     g11902(.A(\b[36] ), .B(new_n2386), .Y(new_n12159));
  NAND2xp33_ASAP7_75t_L     g11903(.A(\b[37] ), .B(new_n2232), .Y(new_n12160));
  AOI22xp33_ASAP7_75t_L     g11904(.A1(new_n2228), .A2(\b[38] ), .B1(new_n2226), .B2(new_n4923), .Y(new_n12161));
  NAND4xp25_ASAP7_75t_L     g11905(.A(new_n12161), .B(\a[26] ), .C(new_n12159), .D(new_n12160), .Y(new_n12162));
  NAND2xp33_ASAP7_75t_L     g11906(.A(new_n12160), .B(new_n12161), .Y(new_n12163));
  A2O1A1Ixp33_ASAP7_75t_L   g11907(.A1(\b[36] ), .A2(new_n2386), .B(new_n12163), .C(new_n2223), .Y(new_n12164));
  NAND2xp33_ASAP7_75t_L     g11908(.A(new_n12162), .B(new_n12164), .Y(new_n12165));
  NOR3xp33_ASAP7_75t_L      g11909(.A(new_n12157), .B(new_n12165), .C(new_n12158), .Y(new_n12166));
  OA21x2_ASAP7_75t_L        g11910(.A1(new_n12158), .A2(new_n12157), .B(new_n12165), .Y(new_n12167));
  NOR2xp33_ASAP7_75t_L      g11911(.A(new_n12166), .B(new_n12167), .Y(new_n12168));
  NAND3xp33_ASAP7_75t_L     g11912(.A(new_n11817), .B(new_n11804), .C(new_n11802), .Y(new_n12169));
  INVx1_ASAP7_75t_L         g11913(.A(new_n12169), .Y(new_n12170));
  A2O1A1O1Ixp25_ASAP7_75t_L g11914(.A1(new_n11482), .A2(new_n11483), .B(new_n11476), .C(new_n11819), .D(new_n12170), .Y(new_n12171));
  NAND2xp33_ASAP7_75t_L     g11915(.A(new_n12168), .B(new_n12171), .Y(new_n12172));
  OR3x1_ASAP7_75t_L         g11916(.A(new_n12157), .B(new_n12158), .C(new_n12165), .Y(new_n12173));
  OAI21xp33_ASAP7_75t_L     g11917(.A1(new_n12158), .A2(new_n12157), .B(new_n12165), .Y(new_n12174));
  NAND2xp33_ASAP7_75t_L     g11918(.A(new_n12174), .B(new_n12173), .Y(new_n12175));
  A2O1A1Ixp33_ASAP7_75t_L   g11919(.A1(new_n11818), .A2(new_n11812), .B(new_n11821), .C(new_n12169), .Y(new_n12176));
  NAND2xp33_ASAP7_75t_L     g11920(.A(new_n12176), .B(new_n12175), .Y(new_n12177));
  AOI22xp33_ASAP7_75t_L     g11921(.A1(new_n1766), .A2(\b[41] ), .B1(new_n1764), .B2(new_n5669), .Y(new_n12178));
  OAI221xp5_ASAP7_75t_L     g11922(.A1(new_n1758), .A2(new_n5186), .B1(new_n5166), .B2(new_n1911), .C(new_n12178), .Y(new_n12179));
  XNOR2x2_ASAP7_75t_L       g11923(.A(\a[23] ), .B(new_n12179), .Y(new_n12180));
  INVx1_ASAP7_75t_L         g11924(.A(new_n12180), .Y(new_n12181));
  AOI21xp33_ASAP7_75t_L     g11925(.A1(new_n12177), .A2(new_n12172), .B(new_n12181), .Y(new_n12182));
  NOR2xp33_ASAP7_75t_L      g11926(.A(new_n12176), .B(new_n12175), .Y(new_n12183));
  A2O1A1O1Ixp25_ASAP7_75t_L g11927(.A1(new_n11818), .A2(new_n11812), .B(new_n11821), .C(new_n12169), .D(new_n12168), .Y(new_n12184));
  NOR3xp33_ASAP7_75t_L      g11928(.A(new_n12184), .B(new_n12183), .C(new_n12180), .Y(new_n12185));
  NOR2xp33_ASAP7_75t_L      g11929(.A(new_n12182), .B(new_n12185), .Y(new_n12186));
  NAND2xp33_ASAP7_75t_L     g11930(.A(new_n11971), .B(new_n12186), .Y(new_n12187));
  OAI21xp33_ASAP7_75t_L     g11931(.A1(new_n12183), .A2(new_n12184), .B(new_n12180), .Y(new_n12188));
  NAND3xp33_ASAP7_75t_L     g11932(.A(new_n12177), .B(new_n12172), .C(new_n12181), .Y(new_n12189));
  NAND2xp33_ASAP7_75t_L     g11933(.A(new_n12189), .B(new_n12188), .Y(new_n12190));
  A2O1A1Ixp33_ASAP7_75t_L   g11934(.A1(new_n11843), .A2(new_n11841), .B(new_n11970), .C(new_n12190), .Y(new_n12191));
  AOI21xp33_ASAP7_75t_L     g11935(.A1(new_n12191), .A2(new_n12187), .B(new_n11969), .Y(new_n12192));
  INVx1_ASAP7_75t_L         g11936(.A(new_n11970), .Y(new_n12193));
  A2O1A1Ixp33_ASAP7_75t_L   g11937(.A1(new_n11840), .A2(new_n11839), .B(new_n11837), .C(new_n12193), .Y(new_n12194));
  NOR2xp33_ASAP7_75t_L      g11938(.A(new_n12194), .B(new_n12190), .Y(new_n12195));
  NOR2xp33_ASAP7_75t_L      g11939(.A(new_n11971), .B(new_n12186), .Y(new_n12196));
  NOR3xp33_ASAP7_75t_L      g11940(.A(new_n12196), .B(new_n12195), .C(new_n11968), .Y(new_n12197));
  INVx1_ASAP7_75t_L         g11941(.A(new_n11517), .Y(new_n12198));
  OAI21xp33_ASAP7_75t_L     g11942(.A1(new_n11853), .A2(new_n11854), .B(new_n11855), .Y(new_n12199));
  A2O1A1O1Ixp25_ASAP7_75t_L g11943(.A1(new_n11511), .A2(new_n12198), .B(new_n11516), .C(new_n12199), .D(new_n11856), .Y(new_n12200));
  NOR3xp33_ASAP7_75t_L      g11944(.A(new_n12200), .B(new_n12192), .C(new_n12197), .Y(new_n12201));
  OAI21xp33_ASAP7_75t_L     g11945(.A1(new_n12195), .A2(new_n12196), .B(new_n11968), .Y(new_n12202));
  NAND3xp33_ASAP7_75t_L     g11946(.A(new_n12191), .B(new_n12187), .C(new_n11969), .Y(new_n12203));
  O2A1O1Ixp33_ASAP7_75t_L   g11947(.A1(new_n11515), .A2(new_n11517), .B(new_n11512), .C(new_n11852), .Y(new_n12204));
  AOI211xp5_ASAP7_75t_L     g11948(.A1(new_n12202), .A2(new_n12203), .B(new_n12204), .C(new_n11856), .Y(new_n12205));
  NOR3xp33_ASAP7_75t_L      g11949(.A(new_n12205), .B(new_n12201), .C(new_n11962), .Y(new_n12206));
  INVx1_ASAP7_75t_L         g11950(.A(new_n11962), .Y(new_n12207));
  OAI211xp5_ASAP7_75t_L     g11951(.A1(new_n11856), .A2(new_n12204), .B(new_n12202), .C(new_n12203), .Y(new_n12208));
  OAI21xp33_ASAP7_75t_L     g11952(.A1(new_n12197), .A2(new_n12192), .B(new_n12200), .Y(new_n12209));
  AOI21xp33_ASAP7_75t_L     g11953(.A1(new_n12209), .A2(new_n12208), .B(new_n12207), .Y(new_n12210));
  NOR2xp33_ASAP7_75t_L      g11954(.A(new_n12210), .B(new_n12206), .Y(new_n12211));
  A2O1A1Ixp33_ASAP7_75t_L   g11955(.A1(new_n11867), .A2(new_n11866), .B(new_n11863), .C(new_n12211), .Y(new_n12212));
  A2O1A1O1Ixp25_ASAP7_75t_L g11956(.A1(new_n11526), .A2(new_n11529), .B(new_n11597), .C(new_n11867), .D(new_n11863), .Y(new_n12213));
  NAND3xp33_ASAP7_75t_L     g11957(.A(new_n12209), .B(new_n12208), .C(new_n12207), .Y(new_n12214));
  OAI21xp33_ASAP7_75t_L     g11958(.A1(new_n12201), .A2(new_n12205), .B(new_n11962), .Y(new_n12215));
  NAND2xp33_ASAP7_75t_L     g11959(.A(new_n12214), .B(new_n12215), .Y(new_n12216));
  NAND2xp33_ASAP7_75t_L     g11960(.A(new_n12213), .B(new_n12216), .Y(new_n12217));
  NAND2xp33_ASAP7_75t_L     g11961(.A(\b[48] ), .B(new_n908), .Y(new_n12218));
  NAND2xp33_ASAP7_75t_L     g11962(.A(\b[49] ), .B(new_n817), .Y(new_n12219));
  AOI22xp33_ASAP7_75t_L     g11963(.A1(new_n826), .A2(\b[50] ), .B1(new_n823), .B2(new_n8235), .Y(new_n12220));
  AND4x1_ASAP7_75t_L        g11964(.A(new_n12220), .B(new_n12219), .C(new_n12218), .D(\a[14] ), .Y(new_n12221));
  AOI31xp33_ASAP7_75t_L     g11965(.A1(new_n12220), .A2(new_n12219), .A3(new_n12218), .B(\a[14] ), .Y(new_n12222));
  NOR2xp33_ASAP7_75t_L      g11966(.A(new_n12222), .B(new_n12221), .Y(new_n12223));
  NAND3xp33_ASAP7_75t_L     g11967(.A(new_n12212), .B(new_n12217), .C(new_n12223), .Y(new_n12224));
  O2A1O1Ixp33_ASAP7_75t_L   g11968(.A1(new_n11598), .A2(new_n11859), .B(new_n11868), .C(new_n12216), .Y(new_n12225));
  AOI221xp5_ASAP7_75t_L     g11969(.A1(new_n11866), .A2(new_n11867), .B1(new_n12214), .B2(new_n12215), .C(new_n11863), .Y(new_n12226));
  INVx1_ASAP7_75t_L         g11970(.A(new_n12223), .Y(new_n12227));
  OAI21xp33_ASAP7_75t_L     g11971(.A1(new_n12226), .A2(new_n12225), .B(new_n12227), .Y(new_n12228));
  AOI21xp33_ASAP7_75t_L     g11972(.A1(new_n12228), .A2(new_n12224), .B(new_n11955), .Y(new_n12229));
  AND3x1_ASAP7_75t_L        g11973(.A(new_n11955), .B(new_n12228), .C(new_n12224), .Y(new_n12230));
  NOR3xp33_ASAP7_75t_L      g11974(.A(new_n12230), .B(new_n12229), .C(new_n11953), .Y(new_n12231));
  INVx1_ASAP7_75t_L         g11975(.A(new_n11953), .Y(new_n12232));
  AO21x2_ASAP7_75t_L        g11976(.A1(new_n12228), .A2(new_n12224), .B(new_n11955), .Y(new_n12233));
  NAND3xp33_ASAP7_75t_L     g11977(.A(new_n11955), .B(new_n12224), .C(new_n12228), .Y(new_n12234));
  AOI21xp33_ASAP7_75t_L     g11978(.A1(new_n12233), .A2(new_n12234), .B(new_n12232), .Y(new_n12235));
  NOR3xp33_ASAP7_75t_L      g11979(.A(new_n11946), .B(new_n12231), .C(new_n12235), .Y(new_n12236));
  OAI21xp33_ASAP7_75t_L     g11980(.A1(new_n11878), .A2(new_n11884), .B(new_n11886), .Y(new_n12237));
  NAND3xp33_ASAP7_75t_L     g11981(.A(new_n12233), .B(new_n12232), .C(new_n12234), .Y(new_n12238));
  OAI21xp33_ASAP7_75t_L     g11982(.A1(new_n12229), .A2(new_n12230), .B(new_n11953), .Y(new_n12239));
  AOI21xp33_ASAP7_75t_L     g11983(.A1(new_n12239), .A2(new_n12238), .B(new_n12237), .Y(new_n12240));
  NAND2xp33_ASAP7_75t_L     g11984(.A(\b[55] ), .B(new_n441), .Y(new_n12241));
  AOI22xp33_ASAP7_75t_L     g11985(.A1(new_n451), .A2(\b[56] ), .B1(new_n448), .B2(new_n10185), .Y(new_n12242));
  NAND2xp33_ASAP7_75t_L     g11986(.A(new_n12241), .B(new_n12242), .Y(new_n12243));
  AOI211xp5_ASAP7_75t_L     g11987(.A1(\b[54] ), .A2(new_n480), .B(new_n445), .C(new_n12243), .Y(new_n12244));
  INVx1_ASAP7_75t_L         g11988(.A(new_n12243), .Y(new_n12245));
  O2A1O1Ixp33_ASAP7_75t_L   g11989(.A1(new_n9199), .A2(new_n481), .B(new_n12245), .C(\a[8] ), .Y(new_n12246));
  NOR2xp33_ASAP7_75t_L      g11990(.A(new_n12244), .B(new_n12246), .Y(new_n12247));
  OAI21xp33_ASAP7_75t_L     g11991(.A1(new_n12240), .A2(new_n12236), .B(new_n12247), .Y(new_n12248));
  NAND3xp33_ASAP7_75t_L     g11992(.A(new_n12237), .B(new_n12238), .C(new_n12239), .Y(new_n12249));
  OAI21xp33_ASAP7_75t_L     g11993(.A1(new_n12231), .A2(new_n12235), .B(new_n11946), .Y(new_n12250));
  INVx1_ASAP7_75t_L         g11994(.A(new_n12247), .Y(new_n12251));
  NAND3xp33_ASAP7_75t_L     g11995(.A(new_n12249), .B(new_n12250), .C(new_n12251), .Y(new_n12252));
  NAND2xp33_ASAP7_75t_L     g11996(.A(\b[59] ), .B(new_n345), .Y(new_n12253));
  OAI221xp5_ASAP7_75t_L     g11997(.A1(new_n10848), .A2(new_n406), .B1(new_n367), .B2(new_n10888), .C(new_n12253), .Y(new_n12254));
  AOI21xp33_ASAP7_75t_L     g11998(.A1(new_n366), .A2(\b[57] ), .B(new_n12254), .Y(new_n12255));
  NAND2xp33_ASAP7_75t_L     g11999(.A(\a[5] ), .B(new_n12255), .Y(new_n12256));
  A2O1A1Ixp33_ASAP7_75t_L   g12000(.A1(\b[57] ), .A2(new_n366), .B(new_n12254), .C(new_n339), .Y(new_n12257));
  AND2x2_ASAP7_75t_L        g12001(.A(new_n12257), .B(new_n12256), .Y(new_n12258));
  NAND3xp33_ASAP7_75t_L     g12002(.A(new_n12248), .B(new_n12252), .C(new_n12258), .Y(new_n12259));
  AOI21xp33_ASAP7_75t_L     g12003(.A1(new_n12249), .A2(new_n12250), .B(new_n12251), .Y(new_n12260));
  NOR3xp33_ASAP7_75t_L      g12004(.A(new_n12236), .B(new_n12240), .C(new_n12247), .Y(new_n12261));
  NAND2xp33_ASAP7_75t_L     g12005(.A(new_n12257), .B(new_n12256), .Y(new_n12262));
  OAI21xp33_ASAP7_75t_L     g12006(.A1(new_n12260), .A2(new_n12261), .B(new_n12262), .Y(new_n12263));
  NAND2xp33_ASAP7_75t_L     g12007(.A(new_n11888), .B(new_n11883), .Y(new_n12264));
  MAJx2_ASAP7_75t_L         g12008(.A(new_n11899), .B(new_n11891), .C(new_n12264), .Y(new_n12265));
  NAND3xp33_ASAP7_75t_L     g12009(.A(new_n12265), .B(new_n12263), .C(new_n12259), .Y(new_n12266));
  NOR3xp33_ASAP7_75t_L      g12010(.A(new_n12261), .B(new_n12260), .C(new_n12262), .Y(new_n12267));
  AOI21xp33_ASAP7_75t_L     g12011(.A1(new_n12248), .A2(new_n12252), .B(new_n12258), .Y(new_n12268));
  NAND3xp33_ASAP7_75t_L     g12012(.A(new_n11883), .B(new_n11888), .C(new_n11897), .Y(new_n12269));
  A2O1A1Ixp33_ASAP7_75t_L   g12013(.A1(new_n11892), .A2(new_n11898), .B(new_n11899), .C(new_n12269), .Y(new_n12270));
  OAI21xp33_ASAP7_75t_L     g12014(.A1(new_n12268), .A2(new_n12267), .B(new_n12270), .Y(new_n12271));
  NOR2xp33_ASAP7_75t_L      g12015(.A(\b[61] ), .B(\b[62] ), .Y(new_n12272));
  INVx1_ASAP7_75t_L         g12016(.A(\b[62] ), .Y(new_n12273));
  NOR2xp33_ASAP7_75t_L      g12017(.A(new_n11911), .B(new_n12273), .Y(new_n12274));
  NOR2xp33_ASAP7_75t_L      g12018(.A(new_n12272), .B(new_n12274), .Y(new_n12275));
  A2O1A1Ixp33_ASAP7_75t_L   g12019(.A1(new_n11916), .A2(new_n11913), .B(new_n11912), .C(new_n12275), .Y(new_n12276));
  INVx1_ASAP7_75t_L         g12020(.A(new_n12276), .Y(new_n12277));
  OAI21xp33_ASAP7_75t_L     g12021(.A1(new_n11226), .A2(new_n11911), .B(new_n11914), .Y(new_n12278));
  NOR2xp33_ASAP7_75t_L      g12022(.A(new_n12275), .B(new_n12278), .Y(new_n12279));
  NOR2xp33_ASAP7_75t_L      g12023(.A(new_n12277), .B(new_n12279), .Y(new_n12280));
  INVx1_ASAP7_75t_L         g12024(.A(new_n12280), .Y(new_n12281));
  NOR2xp33_ASAP7_75t_L      g12025(.A(new_n11911), .B(new_n261), .Y(new_n12282));
  AOI221xp5_ASAP7_75t_L     g12026(.A1(\b[60] ), .A2(new_n291), .B1(\b[62] ), .B2(new_n272), .C(new_n12282), .Y(new_n12283));
  OAI211xp5_ASAP7_75t_L     g12027(.A1(new_n292), .A2(new_n12281), .B(\a[2] ), .C(new_n12283), .Y(new_n12284));
  INVx1_ASAP7_75t_L         g12028(.A(new_n12283), .Y(new_n12285));
  A2O1A1Ixp33_ASAP7_75t_L   g12029(.A1(new_n12280), .A2(new_n269), .B(new_n12285), .C(new_n265), .Y(new_n12286));
  NAND2xp33_ASAP7_75t_L     g12030(.A(new_n12286), .B(new_n12284), .Y(new_n12287));
  AOI21xp33_ASAP7_75t_L     g12031(.A1(new_n12266), .A2(new_n12271), .B(new_n12287), .Y(new_n12288));
  NOR3xp33_ASAP7_75t_L      g12032(.A(new_n12267), .B(new_n12268), .C(new_n12270), .Y(new_n12289));
  AOI21xp33_ASAP7_75t_L     g12033(.A1(new_n12263), .A2(new_n12259), .B(new_n12265), .Y(new_n12290));
  INVx1_ASAP7_75t_L         g12034(.A(new_n12287), .Y(new_n12291));
  NOR3xp33_ASAP7_75t_L      g12035(.A(new_n12289), .B(new_n12290), .C(new_n12291), .Y(new_n12292));
  OAI21xp33_ASAP7_75t_L     g12036(.A1(new_n11926), .A2(new_n11909), .B(new_n11928), .Y(new_n12293));
  NOR3xp33_ASAP7_75t_L      g12037(.A(new_n12292), .B(new_n12288), .C(new_n12293), .Y(new_n12294));
  OAI21xp33_ASAP7_75t_L     g12038(.A1(new_n12290), .A2(new_n12289), .B(new_n12291), .Y(new_n12295));
  NAND3xp33_ASAP7_75t_L     g12039(.A(new_n12266), .B(new_n12271), .C(new_n12287), .Y(new_n12296));
  AOI22xp33_ASAP7_75t_L     g12040(.A1(new_n11935), .A2(new_n11928), .B1(new_n12296), .B2(new_n12295), .Y(new_n12297));
  NOR2xp33_ASAP7_75t_L      g12041(.A(new_n12297), .B(new_n12294), .Y(new_n12298));
  XOR2x2_ASAP7_75t_L        g12042(.A(new_n12298), .B(new_n11945), .Y(\f[62] ));
  NAND3xp33_ASAP7_75t_L     g12043(.A(new_n12212), .B(new_n12217), .C(new_n12227), .Y(new_n12300));
  NAND2xp33_ASAP7_75t_L     g12044(.A(new_n823), .B(new_n8257), .Y(new_n12301));
  OAI221xp5_ASAP7_75t_L     g12045(.A1(new_n912), .A2(new_n8249), .B1(new_n8228), .B2(new_n994), .C(new_n12301), .Y(new_n12302));
  AOI21xp33_ASAP7_75t_L     g12046(.A1(new_n908), .A2(\b[49] ), .B(new_n12302), .Y(new_n12303));
  NAND2xp33_ASAP7_75t_L     g12047(.A(\a[14] ), .B(new_n12303), .Y(new_n12304));
  A2O1A1Ixp33_ASAP7_75t_L   g12048(.A1(\b[49] ), .A2(new_n908), .B(new_n12302), .C(new_n813), .Y(new_n12305));
  NAND2xp33_ASAP7_75t_L     g12049(.A(new_n12305), .B(new_n12304), .Y(new_n12306));
  OAI21xp33_ASAP7_75t_L     g12050(.A1(new_n12210), .A2(new_n12213), .B(new_n12214), .Y(new_n12307));
  NAND2xp33_ASAP7_75t_L     g12051(.A(new_n1110), .B(new_n7341), .Y(new_n12308));
  OAI221xp5_ASAP7_75t_L     g12052(.A1(new_n1198), .A2(new_n7333), .B1(new_n7316), .B2(new_n1298), .C(new_n12308), .Y(new_n12309));
  AOI21xp33_ASAP7_75t_L     g12053(.A1(new_n1194), .A2(\b[46] ), .B(new_n12309), .Y(new_n12310));
  NAND2xp33_ASAP7_75t_L     g12054(.A(\a[17] ), .B(new_n12310), .Y(new_n12311));
  A2O1A1Ixp33_ASAP7_75t_L   g12055(.A1(\b[46] ), .A2(new_n1194), .B(new_n12309), .C(new_n1107), .Y(new_n12312));
  NAND2xp33_ASAP7_75t_L     g12056(.A(new_n12312), .B(new_n12311), .Y(new_n12313));
  INVx1_ASAP7_75t_L         g12057(.A(new_n12313), .Y(new_n12314));
  O2A1O1Ixp33_ASAP7_75t_L   g12058(.A1(new_n11856), .A2(new_n12204), .B(new_n12203), .C(new_n12192), .Y(new_n12315));
  NAND2xp33_ASAP7_75t_L     g12059(.A(new_n1404), .B(new_n6764), .Y(new_n12316));
  OAI221xp5_ASAP7_75t_L     g12060(.A1(new_n1412), .A2(new_n6756), .B1(new_n6220), .B2(new_n1398), .C(new_n12316), .Y(new_n12317));
  AOI21xp33_ASAP7_75t_L     g12061(.A1(new_n1548), .A2(\b[43] ), .B(new_n12317), .Y(new_n12318));
  NAND2xp33_ASAP7_75t_L     g12062(.A(\a[20] ), .B(new_n12318), .Y(new_n12319));
  A2O1A1Ixp33_ASAP7_75t_L   g12063(.A1(\b[43] ), .A2(new_n1548), .B(new_n12317), .C(new_n1401), .Y(new_n12320));
  NAND2xp33_ASAP7_75t_L     g12064(.A(new_n12320), .B(new_n12319), .Y(new_n12321));
  OAI22xp33_ASAP7_75t_L     g12065(.A1(new_n5687), .A2(new_n1771), .B1(new_n5680), .B2(new_n1772), .Y(new_n12322));
  AOI221xp5_ASAP7_75t_L     g12066(.A1(\b[40] ), .A2(new_n1910), .B1(\b[41] ), .B2(new_n1770), .C(new_n12322), .Y(new_n12323));
  XNOR2x2_ASAP7_75t_L       g12067(.A(new_n1761), .B(new_n12323), .Y(new_n12324));
  INVx1_ASAP7_75t_L         g12068(.A(new_n12324), .Y(new_n12325));
  INVx1_ASAP7_75t_L         g12069(.A(new_n12165), .Y(new_n12326));
  NOR3xp33_ASAP7_75t_L      g12070(.A(new_n12157), .B(new_n12326), .C(new_n12158), .Y(new_n12327));
  INVx1_ASAP7_75t_L         g12071(.A(new_n12327), .Y(new_n12328));
  NAND4xp25_ASAP7_75t_L     g12072(.A(new_n12154), .B(new_n12150), .C(new_n11977), .D(new_n11978), .Y(new_n12329));
  A2O1A1O1Ixp25_ASAP7_75t_L g12073(.A1(new_n11801), .A2(new_n11803), .B(new_n11972), .C(new_n12329), .D(new_n12155), .Y(new_n12330));
  AOI22xp33_ASAP7_75t_L     g12074(.A1(new_n2702), .A2(\b[36] ), .B1(new_n2700), .B2(new_n4473), .Y(new_n12331));
  OAI221xp5_ASAP7_75t_L     g12075(.A1(new_n2694), .A2(new_n4053), .B1(new_n3827), .B2(new_n2932), .C(new_n12331), .Y(new_n12332));
  XNOR2x2_ASAP7_75t_L       g12076(.A(\a[29] ), .B(new_n12332), .Y(new_n12333));
  A2O1A1Ixp33_ASAP7_75t_L   g12077(.A1(new_n11725), .A2(new_n11301), .B(new_n11617), .C(new_n11726), .Y(new_n12334));
  A2O1A1Ixp33_ASAP7_75t_L   g12078(.A1(new_n11727), .A2(new_n12334), .B(new_n12092), .C(new_n12084), .Y(new_n12335));
  AOI22xp33_ASAP7_75t_L     g12079(.A1(new_n6002), .A2(\b[21] ), .B1(new_n5999), .B2(new_n1715), .Y(new_n12336));
  OAI221xp5_ASAP7_75t_L     g12080(.A1(new_n6544), .A2(new_n1594), .B1(new_n1493), .B2(new_n6309), .C(new_n12336), .Y(new_n12337));
  XNOR2x2_ASAP7_75t_L       g12081(.A(\a[44] ), .B(new_n12337), .Y(new_n12338));
  INVx1_ASAP7_75t_L         g12082(.A(new_n12338), .Y(new_n12339));
  NAND3xp33_ASAP7_75t_L     g12083(.A(new_n12073), .B(new_n12074), .C(new_n12000), .Y(new_n12340));
  A2O1A1Ixp33_ASAP7_75t_L   g12084(.A1(new_n12071), .A2(new_n12075), .B(new_n12079), .C(new_n12340), .Y(new_n12341));
  NAND2xp33_ASAP7_75t_L     g12085(.A(new_n11683), .B(new_n12052), .Y(new_n12342));
  A2O1A1Ixp33_ASAP7_75t_L   g12086(.A1(new_n11701), .A2(new_n12342), .B(new_n12054), .C(new_n12050), .Y(new_n12343));
  AOI22xp33_ASAP7_75t_L     g12087(.A1(new_n8645), .A2(\b[12] ), .B1(new_n8642), .B2(new_n970), .Y(new_n12344));
  OAI221xp5_ASAP7_75t_L     g12088(.A1(new_n9322), .A2(new_n695), .B1(new_n631), .B2(new_n8965), .C(new_n12344), .Y(new_n12345));
  XNOR2x2_ASAP7_75t_L       g12089(.A(\a[53] ), .B(new_n12345), .Y(new_n12346));
  AOI22xp33_ASAP7_75t_L     g12090(.A1(new_n12014), .A2(new_n12015), .B1(new_n12036), .B2(new_n12040), .Y(new_n12347));
  A2O1A1O1Ixp25_ASAP7_75t_L g12091(.A1(new_n11675), .A2(new_n11672), .B(new_n11670), .C(new_n12041), .D(new_n12347), .Y(new_n12348));
  AOI22xp33_ASAP7_75t_L     g12092(.A1(new_n10594), .A2(\b[6] ), .B1(new_n10591), .B2(new_n389), .Y(new_n12349));
  OAI221xp5_ASAP7_75t_L     g12093(.A1(new_n11335), .A2(new_n353), .B1(new_n323), .B2(new_n11330), .C(new_n12349), .Y(new_n12350));
  OR2x4_ASAP7_75t_L         g12094(.A(new_n10588), .B(new_n12350), .Y(new_n12351));
  NAND2xp33_ASAP7_75t_L     g12095(.A(new_n10588), .B(new_n12350), .Y(new_n12352));
  NOR2xp33_ASAP7_75t_L      g12096(.A(\a[63] ), .B(new_n11651), .Y(new_n12353));
  INVx1_ASAP7_75t_L         g12097(.A(\a[63] ), .Y(new_n12354));
  NOR2xp33_ASAP7_75t_L      g12098(.A(\a[62] ), .B(new_n12354), .Y(new_n12355));
  NOR2xp33_ASAP7_75t_L      g12099(.A(new_n12353), .B(new_n12355), .Y(new_n12356));
  NOR2xp33_ASAP7_75t_L      g12100(.A(new_n11651), .B(new_n11658), .Y(new_n12357));
  A2O1A1Ixp33_ASAP7_75t_L   g12101(.A1(new_n11324), .A2(new_n11325), .B(new_n258), .C(new_n12357), .Y(new_n12358));
  INVx1_ASAP7_75t_L         g12102(.A(new_n12026), .Y(new_n12359));
  NOR2xp33_ASAP7_75t_L      g12103(.A(new_n12359), .B(new_n12358), .Y(new_n12360));
  OAI21xp33_ASAP7_75t_L     g12104(.A1(new_n258), .A2(new_n12356), .B(new_n12360), .Y(new_n12361));
  NOR2xp33_ASAP7_75t_L      g12105(.A(new_n258), .B(new_n12356), .Y(new_n12362));
  OAI21xp33_ASAP7_75t_L     g12106(.A1(new_n12359), .A2(new_n12358), .B(new_n12362), .Y(new_n12363));
  INVx1_ASAP7_75t_L         g12107(.A(new_n11647), .Y(new_n12364));
  NAND2xp33_ASAP7_75t_L     g12108(.A(\b[3] ), .B(new_n11656), .Y(new_n12365));
  OAI221xp5_ASAP7_75t_L     g12109(.A1(new_n12364), .A2(new_n278), .B1(new_n303), .B2(new_n12022), .C(new_n12365), .Y(new_n12366));
  AOI21xp33_ASAP7_75t_L     g12110(.A1(new_n12021), .A2(\b[1] ), .B(new_n12366), .Y(new_n12367));
  NAND2xp33_ASAP7_75t_L     g12111(.A(\a[62] ), .B(new_n12367), .Y(new_n12368));
  A2O1A1Ixp33_ASAP7_75t_L   g12112(.A1(\b[1] ), .A2(new_n12021), .B(new_n12366), .C(new_n11651), .Y(new_n12369));
  NAND2xp33_ASAP7_75t_L     g12113(.A(new_n12369), .B(new_n12368), .Y(new_n12370));
  INVx1_ASAP7_75t_L         g12114(.A(new_n12370), .Y(new_n12371));
  AOI21xp33_ASAP7_75t_L     g12115(.A1(new_n12361), .A2(new_n12363), .B(new_n12371), .Y(new_n12372));
  AND3x1_ASAP7_75t_L        g12116(.A(new_n12361), .B(new_n12371), .C(new_n12363), .Y(new_n12373));
  OAI211xp5_ASAP7_75t_L     g12117(.A1(new_n12372), .A2(new_n12373), .B(new_n12352), .C(new_n12351), .Y(new_n12374));
  NAND2xp33_ASAP7_75t_L     g12118(.A(new_n12352), .B(new_n12351), .Y(new_n12375));
  NOR2xp33_ASAP7_75t_L      g12119(.A(new_n12372), .B(new_n12373), .Y(new_n12376));
  NAND2xp33_ASAP7_75t_L     g12120(.A(new_n12375), .B(new_n12376), .Y(new_n12377));
  A2O1A1Ixp33_ASAP7_75t_L   g12121(.A1(new_n11663), .A2(new_n11662), .B(new_n12031), .C(new_n12038), .Y(new_n12378));
  NAND3xp33_ASAP7_75t_L     g12122(.A(new_n12377), .B(new_n12378), .C(new_n12374), .Y(new_n12379));
  AO21x2_ASAP7_75t_L        g12123(.A1(new_n12374), .A2(new_n12377), .B(new_n12378), .Y(new_n12380));
  AOI22xp33_ASAP7_75t_L     g12124(.A1(new_n9623), .A2(\b[9] ), .B1(new_n9620), .B2(new_n566), .Y(new_n12381));
  OAI221xp5_ASAP7_75t_L     g12125(.A1(new_n10280), .A2(new_n503), .B1(new_n421), .B2(new_n12010), .C(new_n12381), .Y(new_n12382));
  OR2x4_ASAP7_75t_L         g12126(.A(new_n9610), .B(new_n12382), .Y(new_n12383));
  NAND2xp33_ASAP7_75t_L     g12127(.A(new_n9610), .B(new_n12382), .Y(new_n12384));
  AND2x2_ASAP7_75t_L        g12128(.A(new_n12384), .B(new_n12383), .Y(new_n12385));
  NAND3xp33_ASAP7_75t_L     g12129(.A(new_n12385), .B(new_n12380), .C(new_n12379), .Y(new_n12386));
  AO22x1_ASAP7_75t_L        g12130(.A1(new_n12384), .A2(new_n12383), .B1(new_n12379), .B2(new_n12380), .Y(new_n12387));
  AOI21xp33_ASAP7_75t_L     g12131(.A1(new_n12387), .A2(new_n12386), .B(new_n12348), .Y(new_n12388));
  AND3x1_ASAP7_75t_L        g12132(.A(new_n12387), .B(new_n12386), .C(new_n12348), .Y(new_n12389));
  OAI21xp33_ASAP7_75t_L     g12133(.A1(new_n12388), .A2(new_n12389), .B(new_n12346), .Y(new_n12390));
  INVx1_ASAP7_75t_L         g12134(.A(new_n12346), .Y(new_n12391));
  AO21x2_ASAP7_75t_L        g12135(.A1(new_n12386), .A2(new_n12387), .B(new_n12348), .Y(new_n12392));
  NAND3xp33_ASAP7_75t_L     g12136(.A(new_n12387), .B(new_n12386), .C(new_n12348), .Y(new_n12393));
  NAND3xp33_ASAP7_75t_L     g12137(.A(new_n12392), .B(new_n12391), .C(new_n12393), .Y(new_n12394));
  NAND3xp33_ASAP7_75t_L     g12138(.A(new_n12343), .B(new_n12390), .C(new_n12394), .Y(new_n12395));
  A2O1A1O1Ixp25_ASAP7_75t_L g12139(.A1(new_n11683), .A2(new_n12052), .B(new_n11694), .C(new_n12049), .D(new_n12055), .Y(new_n12396));
  AOI21xp33_ASAP7_75t_L     g12140(.A1(new_n12392), .A2(new_n12393), .B(new_n12391), .Y(new_n12397));
  NOR3xp33_ASAP7_75t_L      g12141(.A(new_n12389), .B(new_n12388), .C(new_n12346), .Y(new_n12398));
  OAI21xp33_ASAP7_75t_L     g12142(.A1(new_n12397), .A2(new_n12398), .B(new_n12396), .Y(new_n12399));
  NAND2xp33_ASAP7_75t_L     g12143(.A(\b[13] ), .B(new_n7993), .Y(new_n12400));
  NAND2xp33_ASAP7_75t_L     g12144(.A(\b[14] ), .B(new_n7649), .Y(new_n12401));
  AOI22xp33_ASAP7_75t_L     g12145(.A1(new_n7659), .A2(\b[15] ), .B1(new_n7656), .B2(new_n959), .Y(new_n12402));
  NAND4xp25_ASAP7_75t_L     g12146(.A(new_n12402), .B(\a[50] ), .C(new_n12400), .D(new_n12401), .Y(new_n12403));
  NAND2xp33_ASAP7_75t_L     g12147(.A(new_n12401), .B(new_n12402), .Y(new_n12404));
  A2O1A1Ixp33_ASAP7_75t_L   g12148(.A1(\b[13] ), .A2(new_n7993), .B(new_n12404), .C(new_n7653), .Y(new_n12405));
  NAND4xp25_ASAP7_75t_L     g12149(.A(new_n12399), .B(new_n12395), .C(new_n12403), .D(new_n12405), .Y(new_n12406));
  NOR3xp33_ASAP7_75t_L      g12150(.A(new_n12396), .B(new_n12398), .C(new_n12397), .Y(new_n12407));
  AOI21xp33_ASAP7_75t_L     g12151(.A1(new_n12390), .A2(new_n12394), .B(new_n12343), .Y(new_n12408));
  NAND2xp33_ASAP7_75t_L     g12152(.A(new_n12403), .B(new_n12405), .Y(new_n12409));
  OAI21xp33_ASAP7_75t_L     g12153(.A1(new_n12408), .A2(new_n12407), .B(new_n12409), .Y(new_n12410));
  INVx1_ASAP7_75t_L         g12154(.A(new_n12062), .Y(new_n12411));
  NAND3xp33_ASAP7_75t_L     g12155(.A(new_n12056), .B(new_n12051), .C(new_n12411), .Y(new_n12412));
  AND4x1_ASAP7_75t_L        g12156(.A(new_n12073), .B(new_n12412), .C(new_n12410), .D(new_n12406), .Y(new_n12413));
  AOI22xp33_ASAP7_75t_L     g12157(.A1(new_n12406), .A2(new_n12410), .B1(new_n12412), .B2(new_n12073), .Y(new_n12414));
  AOI22xp33_ASAP7_75t_L     g12158(.A1(new_n6822), .A2(\b[18] ), .B1(new_n6819), .B2(new_n1363), .Y(new_n12415));
  OAI221xp5_ASAP7_75t_L     g12159(.A1(new_n7392), .A2(new_n1244), .B1(new_n1051), .B2(new_n7115), .C(new_n12415), .Y(new_n12416));
  XNOR2x2_ASAP7_75t_L       g12160(.A(\a[47] ), .B(new_n12416), .Y(new_n12417));
  OAI21xp33_ASAP7_75t_L     g12161(.A1(new_n12414), .A2(new_n12413), .B(new_n12417), .Y(new_n12418));
  NAND4xp25_ASAP7_75t_L     g12162(.A(new_n12073), .B(new_n12412), .C(new_n12410), .D(new_n12406), .Y(new_n12419));
  AO22x1_ASAP7_75t_L        g12163(.A1(new_n12406), .A2(new_n12410), .B1(new_n12412), .B2(new_n12073), .Y(new_n12420));
  XNOR2x2_ASAP7_75t_L       g12164(.A(new_n6816), .B(new_n12416), .Y(new_n12421));
  NAND3xp33_ASAP7_75t_L     g12165(.A(new_n12420), .B(new_n12419), .C(new_n12421), .Y(new_n12422));
  NAND3xp33_ASAP7_75t_L     g12166(.A(new_n12341), .B(new_n12418), .C(new_n12422), .Y(new_n12423));
  AOI21xp33_ASAP7_75t_L     g12167(.A1(new_n12422), .A2(new_n12418), .B(new_n12341), .Y(new_n12424));
  INVx1_ASAP7_75t_L         g12168(.A(new_n12424), .Y(new_n12425));
  NAND3xp33_ASAP7_75t_L     g12169(.A(new_n12425), .B(new_n12423), .C(new_n12339), .Y(new_n12426));
  INVx1_ASAP7_75t_L         g12170(.A(new_n12423), .Y(new_n12427));
  OAI21xp33_ASAP7_75t_L     g12171(.A1(new_n12424), .A2(new_n12427), .B(new_n12338), .Y(new_n12428));
  NAND3xp33_ASAP7_75t_L     g12172(.A(new_n12335), .B(new_n12426), .C(new_n12428), .Y(new_n12429));
  NOR3xp33_ASAP7_75t_L      g12173(.A(new_n12086), .B(new_n12088), .C(new_n12085), .Y(new_n12430));
  A2O1A1O1Ixp25_ASAP7_75t_L g12174(.A1(new_n11726), .A2(new_n11733), .B(new_n11722), .C(new_n12089), .D(new_n12430), .Y(new_n12431));
  NAND2xp33_ASAP7_75t_L     g12175(.A(new_n12426), .B(new_n12428), .Y(new_n12432));
  NAND2xp33_ASAP7_75t_L     g12176(.A(new_n12431), .B(new_n12432), .Y(new_n12433));
  AOI22xp33_ASAP7_75t_L     g12177(.A1(new_n5249), .A2(\b[24] ), .B1(new_n5247), .B2(new_n2027), .Y(new_n12434));
  OAI221xp5_ASAP7_75t_L     g12178(.A1(new_n5241), .A2(new_n1995), .B1(new_n1857), .B2(new_n5521), .C(new_n12434), .Y(new_n12435));
  XNOR2x2_ASAP7_75t_L       g12179(.A(\a[41] ), .B(new_n12435), .Y(new_n12436));
  NAND3xp33_ASAP7_75t_L     g12180(.A(new_n12433), .B(new_n12429), .C(new_n12436), .Y(new_n12437));
  NOR2xp33_ASAP7_75t_L      g12181(.A(new_n12431), .B(new_n12432), .Y(new_n12438));
  AOI21xp33_ASAP7_75t_L     g12182(.A1(new_n12428), .A2(new_n12426), .B(new_n12335), .Y(new_n12439));
  INVx1_ASAP7_75t_L         g12183(.A(new_n12436), .Y(new_n12440));
  OAI21xp33_ASAP7_75t_L     g12184(.A1(new_n12439), .A2(new_n12438), .B(new_n12440), .Y(new_n12441));
  A2O1A1O1Ixp25_ASAP7_75t_L g12185(.A1(new_n11981), .A2(new_n11738), .B(new_n11730), .C(new_n12099), .D(new_n12111), .Y(new_n12442));
  NAND3xp33_ASAP7_75t_L     g12186(.A(new_n12442), .B(new_n12441), .C(new_n12437), .Y(new_n12443));
  AOI21xp33_ASAP7_75t_L     g12187(.A1(new_n12441), .A2(new_n12437), .B(new_n12442), .Y(new_n12444));
  INVx1_ASAP7_75t_L         g12188(.A(new_n12444), .Y(new_n12445));
  NAND2xp33_ASAP7_75t_L     g12189(.A(new_n4542), .B(new_n2657), .Y(new_n12446));
  OAI221xp5_ASAP7_75t_L     g12190(.A1(new_n4550), .A2(new_n2650), .B1(new_n2477), .B2(new_n4536), .C(new_n12446), .Y(new_n12447));
  AOI21xp33_ASAP7_75t_L     g12191(.A1(new_n4780), .A2(\b[25] ), .B(new_n12447), .Y(new_n12448));
  NAND2xp33_ASAP7_75t_L     g12192(.A(\a[38] ), .B(new_n12448), .Y(new_n12449));
  A2O1A1Ixp33_ASAP7_75t_L   g12193(.A1(\b[25] ), .A2(new_n4780), .B(new_n12447), .C(new_n4539), .Y(new_n12450));
  NAND2xp33_ASAP7_75t_L     g12194(.A(new_n12450), .B(new_n12449), .Y(new_n12451));
  INVx1_ASAP7_75t_L         g12195(.A(new_n12451), .Y(new_n12452));
  NAND3xp33_ASAP7_75t_L     g12196(.A(new_n12445), .B(new_n12443), .C(new_n12452), .Y(new_n12453));
  INVx1_ASAP7_75t_L         g12197(.A(new_n12443), .Y(new_n12454));
  OAI21xp33_ASAP7_75t_L     g12198(.A1(new_n12444), .A2(new_n12454), .B(new_n12451), .Y(new_n12455));
  NAND2xp33_ASAP7_75t_L     g12199(.A(new_n12453), .B(new_n12455), .Y(new_n12456));
  NOR3xp33_ASAP7_75t_L      g12200(.A(new_n12103), .B(new_n12106), .C(new_n12100), .Y(new_n12457));
  INVx1_ASAP7_75t_L         g12201(.A(new_n12457), .Y(new_n12458));
  A2O1A1Ixp33_ASAP7_75t_L   g12202(.A1(new_n12122), .A2(new_n12121), .B(new_n12118), .C(new_n12458), .Y(new_n12459));
  NOR2xp33_ASAP7_75t_L      g12203(.A(new_n12459), .B(new_n12456), .Y(new_n12460));
  NOR3xp33_ASAP7_75t_L      g12204(.A(new_n12454), .B(new_n12444), .C(new_n12451), .Y(new_n12461));
  AOI21xp33_ASAP7_75t_L     g12205(.A1(new_n12445), .A2(new_n12443), .B(new_n12452), .Y(new_n12462));
  NOR2xp33_ASAP7_75t_L      g12206(.A(new_n12462), .B(new_n12461), .Y(new_n12463));
  O2A1O1Ixp33_ASAP7_75t_L   g12207(.A1(new_n11760), .A2(new_n12117), .B(new_n12123), .C(new_n12457), .Y(new_n12464));
  NOR2xp33_ASAP7_75t_L      g12208(.A(new_n12464), .B(new_n12463), .Y(new_n12465));
  AOI22xp33_ASAP7_75t_L     g12209(.A1(new_n3884), .A2(\b[30] ), .B1(new_n3881), .B2(new_n3219), .Y(new_n12466));
  OAI221xp5_ASAP7_75t_L     g12210(.A1(new_n4312), .A2(new_n2871), .B1(new_n2852), .B2(new_n4986), .C(new_n12466), .Y(new_n12467));
  XNOR2x2_ASAP7_75t_L       g12211(.A(\a[35] ), .B(new_n12467), .Y(new_n12468));
  OAI21xp33_ASAP7_75t_L     g12212(.A1(new_n12460), .A2(new_n12465), .B(new_n12468), .Y(new_n12469));
  NAND2xp33_ASAP7_75t_L     g12213(.A(new_n12464), .B(new_n12463), .Y(new_n12470));
  NAND2xp33_ASAP7_75t_L     g12214(.A(new_n12459), .B(new_n12456), .Y(new_n12471));
  INVx1_ASAP7_75t_L         g12215(.A(new_n12468), .Y(new_n12472));
  NAND3xp33_ASAP7_75t_L     g12216(.A(new_n12470), .B(new_n12471), .C(new_n12472), .Y(new_n12473));
  NAND3xp33_ASAP7_75t_L     g12217(.A(new_n12124), .B(new_n12119), .C(new_n12131), .Y(new_n12474));
  A2O1A1Ixp33_ASAP7_75t_L   g12218(.A1(new_n12135), .A2(new_n11782), .B(new_n12140), .C(new_n12474), .Y(new_n12475));
  NAND3xp33_ASAP7_75t_L     g12219(.A(new_n12475), .B(new_n12473), .C(new_n12469), .Y(new_n12476));
  INVx1_ASAP7_75t_L         g12220(.A(new_n12474), .Y(new_n12477));
  AOI221xp5_ASAP7_75t_L     g12221(.A1(new_n12136), .A2(new_n12133), .B1(new_n12473), .B2(new_n12469), .C(new_n12477), .Y(new_n12478));
  INVx1_ASAP7_75t_L         g12222(.A(new_n12478), .Y(new_n12479));
  AOI22xp33_ASAP7_75t_L     g12223(.A1(new_n3256), .A2(\b[33] ), .B1(new_n3254), .B2(new_n3813), .Y(new_n12480));
  OAI221xp5_ASAP7_75t_L     g12224(.A1(new_n3248), .A2(new_n3443), .B1(new_n3419), .B2(new_n3492), .C(new_n12480), .Y(new_n12481));
  XNOR2x2_ASAP7_75t_L       g12225(.A(\a[32] ), .B(new_n12481), .Y(new_n12482));
  NAND3xp33_ASAP7_75t_L     g12226(.A(new_n12476), .B(new_n12479), .C(new_n12482), .Y(new_n12483));
  NAND2xp33_ASAP7_75t_L     g12227(.A(new_n12473), .B(new_n12469), .Y(new_n12484));
  O2A1O1Ixp33_ASAP7_75t_L   g12228(.A1(new_n12138), .A2(new_n12139), .B(new_n12136), .C(new_n12477), .Y(new_n12485));
  NOR2xp33_ASAP7_75t_L      g12229(.A(new_n12485), .B(new_n12484), .Y(new_n12486));
  INVx1_ASAP7_75t_L         g12230(.A(new_n12482), .Y(new_n12487));
  OAI21xp33_ASAP7_75t_L     g12231(.A1(new_n12478), .A2(new_n12486), .B(new_n12487), .Y(new_n12488));
  AOI21xp33_ASAP7_75t_L     g12232(.A1(new_n12151), .A2(new_n12145), .B(new_n12153), .Y(new_n12489));
  AOI21xp33_ASAP7_75t_L     g12233(.A1(new_n12483), .A2(new_n12488), .B(new_n12489), .Y(new_n12490));
  NOR3xp33_ASAP7_75t_L      g12234(.A(new_n12486), .B(new_n12478), .C(new_n12487), .Y(new_n12491));
  AOI21xp33_ASAP7_75t_L     g12235(.A1(new_n12476), .A2(new_n12479), .B(new_n12482), .Y(new_n12492));
  A2O1A1Ixp33_ASAP7_75t_L   g12236(.A1(new_n11980), .A2(new_n11979), .B(new_n12152), .C(new_n12149), .Y(new_n12493));
  NOR3xp33_ASAP7_75t_L      g12237(.A(new_n12493), .B(new_n12492), .C(new_n12491), .Y(new_n12494));
  NOR3xp33_ASAP7_75t_L      g12238(.A(new_n12494), .B(new_n12490), .C(new_n12333), .Y(new_n12495));
  OA21x2_ASAP7_75t_L        g12239(.A1(new_n12490), .A2(new_n12494), .B(new_n12333), .Y(new_n12496));
  OAI21xp33_ASAP7_75t_L     g12240(.A1(new_n12495), .A2(new_n12496), .B(new_n12330), .Y(new_n12497));
  OR3x1_ASAP7_75t_L         g12241(.A(new_n12494), .B(new_n12333), .C(new_n12490), .Y(new_n12498));
  OAI21xp33_ASAP7_75t_L     g12242(.A1(new_n12490), .A2(new_n12494), .B(new_n12333), .Y(new_n12499));
  OAI211xp5_ASAP7_75t_L     g12243(.A1(new_n12155), .A2(new_n12158), .B(new_n12498), .C(new_n12499), .Y(new_n12500));
  NAND2xp33_ASAP7_75t_L     g12244(.A(new_n2226), .B(new_n5174), .Y(new_n12501));
  OAI221xp5_ASAP7_75t_L     g12245(.A1(new_n2234), .A2(new_n5166), .B1(new_n4915), .B2(new_n2220), .C(new_n12501), .Y(new_n12502));
  AOI21xp33_ASAP7_75t_L     g12246(.A1(new_n2386), .A2(\b[37] ), .B(new_n12502), .Y(new_n12503));
  NAND2xp33_ASAP7_75t_L     g12247(.A(\a[26] ), .B(new_n12503), .Y(new_n12504));
  A2O1A1Ixp33_ASAP7_75t_L   g12248(.A1(\b[37] ), .A2(new_n2386), .B(new_n12502), .C(new_n2223), .Y(new_n12505));
  NAND2xp33_ASAP7_75t_L     g12249(.A(new_n12505), .B(new_n12504), .Y(new_n12506));
  AO21x2_ASAP7_75t_L        g12250(.A1(new_n12497), .A2(new_n12500), .B(new_n12506), .Y(new_n12507));
  NAND3xp33_ASAP7_75t_L     g12251(.A(new_n12500), .B(new_n12497), .C(new_n12506), .Y(new_n12508));
  NAND2xp33_ASAP7_75t_L     g12252(.A(new_n12508), .B(new_n12507), .Y(new_n12509));
  O2A1O1Ixp33_ASAP7_75t_L   g12253(.A1(new_n12168), .A2(new_n12171), .B(new_n12328), .C(new_n12509), .Y(new_n12510));
  A2O1A1Ixp33_ASAP7_75t_L   g12254(.A1(new_n11832), .A2(new_n12169), .B(new_n12168), .C(new_n12328), .Y(new_n12511));
  AOI21xp33_ASAP7_75t_L     g12255(.A1(new_n12500), .A2(new_n12497), .B(new_n12506), .Y(new_n12512));
  AND3x1_ASAP7_75t_L        g12256(.A(new_n12500), .B(new_n12506), .C(new_n12497), .Y(new_n12513));
  NOR2xp33_ASAP7_75t_L      g12257(.A(new_n12512), .B(new_n12513), .Y(new_n12514));
  NOR2xp33_ASAP7_75t_L      g12258(.A(new_n12514), .B(new_n12511), .Y(new_n12515));
  OAI21xp33_ASAP7_75t_L     g12259(.A1(new_n12515), .A2(new_n12510), .B(new_n12325), .Y(new_n12516));
  A2O1A1Ixp33_ASAP7_75t_L   g12260(.A1(new_n12176), .A2(new_n12175), .B(new_n12327), .C(new_n12514), .Y(new_n12517));
  O2A1O1Ixp33_ASAP7_75t_L   g12261(.A1(new_n12166), .A2(new_n12167), .B(new_n12176), .C(new_n12327), .Y(new_n12518));
  NAND2xp33_ASAP7_75t_L     g12262(.A(new_n12518), .B(new_n12509), .Y(new_n12519));
  NAND3xp33_ASAP7_75t_L     g12263(.A(new_n12517), .B(new_n12324), .C(new_n12519), .Y(new_n12520));
  A2O1A1O1Ixp25_ASAP7_75t_L g12264(.A1(new_n11843), .A2(new_n11841), .B(new_n11970), .C(new_n12188), .D(new_n12185), .Y(new_n12521));
  AOI21xp33_ASAP7_75t_L     g12265(.A1(new_n12520), .A2(new_n12516), .B(new_n12521), .Y(new_n12522));
  AND3x1_ASAP7_75t_L        g12266(.A(new_n12521), .B(new_n12520), .C(new_n12516), .Y(new_n12523));
  OAI21xp33_ASAP7_75t_L     g12267(.A1(new_n12522), .A2(new_n12523), .B(new_n12321), .Y(new_n12524));
  NAND2xp33_ASAP7_75t_L     g12268(.A(new_n12520), .B(new_n12516), .Y(new_n12525));
  A2O1A1Ixp33_ASAP7_75t_L   g12269(.A1(new_n11844), .A2(new_n12193), .B(new_n12182), .C(new_n12189), .Y(new_n12526));
  NAND2xp33_ASAP7_75t_L     g12270(.A(new_n12525), .B(new_n12526), .Y(new_n12527));
  NAND3xp33_ASAP7_75t_L     g12271(.A(new_n12521), .B(new_n12520), .C(new_n12516), .Y(new_n12528));
  NAND4xp25_ASAP7_75t_L     g12272(.A(new_n12527), .B(new_n12319), .C(new_n12320), .D(new_n12528), .Y(new_n12529));
  AO21x2_ASAP7_75t_L        g12273(.A1(new_n12529), .A2(new_n12524), .B(new_n12315), .Y(new_n12530));
  NAND3xp33_ASAP7_75t_L     g12274(.A(new_n12315), .B(new_n12524), .C(new_n12529), .Y(new_n12531));
  AOI21xp33_ASAP7_75t_L     g12275(.A1(new_n12530), .A2(new_n12531), .B(new_n12314), .Y(new_n12532));
  AOI21xp33_ASAP7_75t_L     g12276(.A1(new_n12529), .A2(new_n12524), .B(new_n12315), .Y(new_n12533));
  INVx1_ASAP7_75t_L         g12277(.A(new_n11856), .Y(new_n12534));
  A2O1A1Ixp33_ASAP7_75t_L   g12278(.A1(new_n11838), .A2(new_n11844), .B(new_n11851), .C(new_n11606), .Y(new_n12535));
  A2O1A1Ixp33_ASAP7_75t_L   g12279(.A1(new_n12534), .A2(new_n12535), .B(new_n12197), .C(new_n12202), .Y(new_n12536));
  NAND2xp33_ASAP7_75t_L     g12280(.A(new_n12524), .B(new_n12529), .Y(new_n12537));
  NOR2xp33_ASAP7_75t_L      g12281(.A(new_n12536), .B(new_n12537), .Y(new_n12538));
  NOR3xp33_ASAP7_75t_L      g12282(.A(new_n12538), .B(new_n12533), .C(new_n12313), .Y(new_n12539));
  OAI21xp33_ASAP7_75t_L     g12283(.A1(new_n12532), .A2(new_n12539), .B(new_n12307), .Y(new_n12540));
  A2O1A1O1Ixp25_ASAP7_75t_L g12284(.A1(new_n11867), .A2(new_n11866), .B(new_n11863), .C(new_n12215), .D(new_n12206), .Y(new_n12541));
  OAI21xp33_ASAP7_75t_L     g12285(.A1(new_n12533), .A2(new_n12538), .B(new_n12313), .Y(new_n12542));
  NAND3xp33_ASAP7_75t_L     g12286(.A(new_n12530), .B(new_n12314), .C(new_n12531), .Y(new_n12543));
  NAND3xp33_ASAP7_75t_L     g12287(.A(new_n12542), .B(new_n12541), .C(new_n12543), .Y(new_n12544));
  NAND3xp33_ASAP7_75t_L     g12288(.A(new_n12540), .B(new_n12544), .C(new_n12306), .Y(new_n12545));
  AO21x2_ASAP7_75t_L        g12289(.A1(new_n12544), .A2(new_n12540), .B(new_n12306), .Y(new_n12546));
  NAND2xp33_ASAP7_75t_L     g12290(.A(new_n12545), .B(new_n12546), .Y(new_n12547));
  A2O1A1O1Ixp25_ASAP7_75t_L g12291(.A1(new_n12224), .A2(new_n12228), .B(new_n11955), .C(new_n12300), .D(new_n12547), .Y(new_n12548));
  A2O1A1Ixp33_ASAP7_75t_L   g12292(.A1(new_n12224), .A2(new_n12228), .B(new_n11955), .C(new_n12300), .Y(new_n12549));
  AOI21xp33_ASAP7_75t_L     g12293(.A1(new_n12546), .A2(new_n12545), .B(new_n12549), .Y(new_n12550));
  NAND2xp33_ASAP7_75t_L     g12294(.A(\b[54] ), .B(new_n600), .Y(new_n12551));
  OAI221xp5_ASAP7_75t_L     g12295(.A1(new_n8882), .A2(new_n721), .B1(new_n675), .B2(new_n9207), .C(new_n12551), .Y(new_n12552));
  AOI21xp33_ASAP7_75t_L     g12296(.A1(new_n674), .A2(\b[52] ), .B(new_n12552), .Y(new_n12553));
  NAND2xp33_ASAP7_75t_L     g12297(.A(\a[11] ), .B(new_n12553), .Y(new_n12554));
  A2O1A1Ixp33_ASAP7_75t_L   g12298(.A1(\b[52] ), .A2(new_n674), .B(new_n12552), .C(new_n594), .Y(new_n12555));
  NAND2xp33_ASAP7_75t_L     g12299(.A(new_n12555), .B(new_n12554), .Y(new_n12556));
  NOR3xp33_ASAP7_75t_L      g12300(.A(new_n12548), .B(new_n12550), .C(new_n12556), .Y(new_n12557));
  NAND3xp33_ASAP7_75t_L     g12301(.A(new_n12549), .B(new_n12545), .C(new_n12546), .Y(new_n12558));
  NAND3xp33_ASAP7_75t_L     g12302(.A(new_n12547), .B(new_n12233), .C(new_n12300), .Y(new_n12559));
  INVx1_ASAP7_75t_L         g12303(.A(new_n12556), .Y(new_n12560));
  AOI21xp33_ASAP7_75t_L     g12304(.A1(new_n12559), .A2(new_n12558), .B(new_n12560), .Y(new_n12561));
  OAI21xp33_ASAP7_75t_L     g12305(.A1(new_n12235), .A2(new_n11946), .B(new_n12238), .Y(new_n12562));
  NOR3xp33_ASAP7_75t_L      g12306(.A(new_n12562), .B(new_n12561), .C(new_n12557), .Y(new_n12563));
  NAND3xp33_ASAP7_75t_L     g12307(.A(new_n12559), .B(new_n12558), .C(new_n12560), .Y(new_n12564));
  OAI21xp33_ASAP7_75t_L     g12308(.A1(new_n12550), .A2(new_n12548), .B(new_n12556), .Y(new_n12565));
  A2O1A1O1Ixp25_ASAP7_75t_L g12309(.A1(new_n11885), .A2(new_n11895), .B(new_n11881), .C(new_n12239), .D(new_n12231), .Y(new_n12566));
  AOI21xp33_ASAP7_75t_L     g12310(.A1(new_n12565), .A2(new_n12564), .B(new_n12566), .Y(new_n12567));
  NAND2xp33_ASAP7_75t_L     g12311(.A(new_n448), .B(new_n10495), .Y(new_n12568));
  OAI221xp5_ASAP7_75t_L     g12312(.A1(new_n667), .A2(new_n10488), .B1(new_n10178), .B2(new_n529), .C(new_n12568), .Y(new_n12569));
  AOI21xp33_ASAP7_75t_L     g12313(.A1(new_n480), .A2(\b[55] ), .B(new_n12569), .Y(new_n12570));
  NAND2xp33_ASAP7_75t_L     g12314(.A(\a[8] ), .B(new_n12570), .Y(new_n12571));
  A2O1A1Ixp33_ASAP7_75t_L   g12315(.A1(\b[55] ), .A2(new_n480), .B(new_n12569), .C(new_n445), .Y(new_n12572));
  NAND2xp33_ASAP7_75t_L     g12316(.A(new_n12572), .B(new_n12571), .Y(new_n12573));
  NOR3xp33_ASAP7_75t_L      g12317(.A(new_n12563), .B(new_n12567), .C(new_n12573), .Y(new_n12574));
  NAND3xp33_ASAP7_75t_L     g12318(.A(new_n12566), .B(new_n12565), .C(new_n12564), .Y(new_n12575));
  OAI21xp33_ASAP7_75t_L     g12319(.A1(new_n12561), .A2(new_n12557), .B(new_n12562), .Y(new_n12576));
  INVx1_ASAP7_75t_L         g12320(.A(new_n12573), .Y(new_n12577));
  AOI21xp33_ASAP7_75t_L     g12321(.A1(new_n12575), .A2(new_n12576), .B(new_n12577), .Y(new_n12578));
  NOR2xp33_ASAP7_75t_L      g12322(.A(new_n10848), .B(new_n365), .Y(new_n12579));
  INVx1_ASAP7_75t_L         g12323(.A(new_n12579), .Y(new_n12580));
  NAND2xp33_ASAP7_75t_L     g12324(.A(\b[59] ), .B(new_n334), .Y(new_n12581));
  AOI22xp33_ASAP7_75t_L     g12325(.A1(new_n345), .A2(\b[60] ), .B1(new_n342), .B2(new_n11234), .Y(new_n12582));
  AND4x1_ASAP7_75t_L        g12326(.A(new_n12582), .B(new_n12581), .C(new_n12580), .D(\a[5] ), .Y(new_n12583));
  AOI31xp33_ASAP7_75t_L     g12327(.A1(new_n12582), .A2(new_n12581), .A3(new_n12580), .B(\a[5] ), .Y(new_n12584));
  NOR2xp33_ASAP7_75t_L      g12328(.A(new_n12584), .B(new_n12583), .Y(new_n12585));
  OAI21xp33_ASAP7_75t_L     g12329(.A1(new_n12578), .A2(new_n12574), .B(new_n12585), .Y(new_n12586));
  NAND3xp33_ASAP7_75t_L     g12330(.A(new_n12575), .B(new_n12576), .C(new_n12577), .Y(new_n12587));
  OAI21xp33_ASAP7_75t_L     g12331(.A1(new_n12567), .A2(new_n12563), .B(new_n12573), .Y(new_n12588));
  INVx1_ASAP7_75t_L         g12332(.A(new_n12585), .Y(new_n12589));
  NAND3xp33_ASAP7_75t_L     g12333(.A(new_n12588), .B(new_n12587), .C(new_n12589), .Y(new_n12590));
  A2O1A1Ixp33_ASAP7_75t_L   g12334(.A1(new_n12250), .A2(new_n12249), .B(new_n12251), .C(new_n12259), .Y(new_n12591));
  NAND3xp33_ASAP7_75t_L     g12335(.A(new_n12586), .B(new_n12591), .C(new_n12590), .Y(new_n12592));
  AOI21xp33_ASAP7_75t_L     g12336(.A1(new_n12588), .A2(new_n12587), .B(new_n12589), .Y(new_n12593));
  NOR3xp33_ASAP7_75t_L      g12337(.A(new_n12574), .B(new_n12578), .C(new_n12585), .Y(new_n12594));
  O2A1O1Ixp33_ASAP7_75t_L   g12338(.A1(new_n12236), .A2(new_n12240), .B(new_n12247), .C(new_n12267), .Y(new_n12595));
  OAI21xp33_ASAP7_75t_L     g12339(.A1(new_n12593), .A2(new_n12594), .B(new_n12595), .Y(new_n12596));
  A2O1A1O1Ixp25_ASAP7_75t_L g12340(.A1(new_n11913), .A2(new_n11916), .B(new_n11912), .C(new_n12275), .D(new_n12274), .Y(new_n12597));
  NOR2xp33_ASAP7_75t_L      g12341(.A(\b[63] ), .B(new_n12273), .Y(new_n12598));
  INVx1_ASAP7_75t_L         g12342(.A(\b[63] ), .Y(new_n12599));
  NOR2xp33_ASAP7_75t_L      g12343(.A(\b[62] ), .B(new_n12599), .Y(new_n12600));
  NOR2xp33_ASAP7_75t_L      g12344(.A(new_n12598), .B(new_n12600), .Y(new_n12601));
  INVx1_ASAP7_75t_L         g12345(.A(new_n12601), .Y(new_n12602));
  NAND2xp33_ASAP7_75t_L     g12346(.A(new_n12602), .B(new_n12597), .Y(new_n12603));
  O2A1O1Ixp33_ASAP7_75t_L   g12347(.A1(new_n11227), .A2(new_n11230), .B(new_n11913), .C(new_n11912), .Y(new_n12604));
  INVx1_ASAP7_75t_L         g12348(.A(new_n12274), .Y(new_n12605));
  O2A1O1Ixp33_ASAP7_75t_L   g12349(.A1(new_n12272), .A2(new_n12604), .B(new_n12605), .C(new_n12602), .Y(new_n12606));
  INVx1_ASAP7_75t_L         g12350(.A(new_n12606), .Y(new_n12607));
  AOI22xp33_ASAP7_75t_L     g12351(.A1(new_n380), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n272), .Y(new_n12608));
  A2O1A1Ixp33_ASAP7_75t_L   g12352(.A1(new_n12607), .A2(new_n12603), .B(new_n292), .C(new_n12608), .Y(new_n12609));
  AOI211xp5_ASAP7_75t_L     g12353(.A1(\b[61] ), .A2(new_n291), .B(new_n265), .C(new_n12609), .Y(new_n12610));
  INVx1_ASAP7_75t_L         g12354(.A(new_n12609), .Y(new_n12611));
  O2A1O1Ixp33_ASAP7_75t_L   g12355(.A1(new_n11911), .A2(new_n277), .B(new_n12611), .C(\a[2] ), .Y(new_n12612));
  NOR2xp33_ASAP7_75t_L      g12356(.A(new_n12610), .B(new_n12612), .Y(new_n12613));
  NAND3xp33_ASAP7_75t_L     g12357(.A(new_n12596), .B(new_n12592), .C(new_n12613), .Y(new_n12614));
  NOR3xp33_ASAP7_75t_L      g12358(.A(new_n12595), .B(new_n12594), .C(new_n12593), .Y(new_n12615));
  AOI21xp33_ASAP7_75t_L     g12359(.A1(new_n12586), .A2(new_n12590), .B(new_n12591), .Y(new_n12616));
  OAI22xp33_ASAP7_75t_L     g12360(.A1(new_n12615), .A2(new_n12616), .B1(new_n12612), .B2(new_n12610), .Y(new_n12617));
  O2A1O1Ixp33_ASAP7_75t_L   g12361(.A1(new_n12267), .A2(new_n12268), .B(new_n12270), .C(new_n12292), .Y(new_n12618));
  AO21x2_ASAP7_75t_L        g12362(.A1(new_n12614), .A2(new_n12617), .B(new_n12618), .Y(new_n12619));
  NAND3xp33_ASAP7_75t_L     g12363(.A(new_n12617), .B(new_n12618), .C(new_n12614), .Y(new_n12620));
  NAND2xp33_ASAP7_75t_L     g12364(.A(new_n12620), .B(new_n12619), .Y(new_n12621));
  INVx1_ASAP7_75t_L         g12365(.A(new_n12621), .Y(new_n12622));
  A2O1A1Ixp33_ASAP7_75t_L   g12366(.A1(new_n11945), .A2(new_n12298), .B(new_n12294), .C(new_n12622), .Y(new_n12623));
  A2O1A1O1Ixp25_ASAP7_75t_L g12367(.A1(new_n11938), .A2(new_n11941), .B(new_n11937), .C(new_n12298), .D(new_n12294), .Y(new_n12624));
  NAND2xp33_ASAP7_75t_L     g12368(.A(new_n12621), .B(new_n12624), .Y(new_n12625));
  AND2x2_ASAP7_75t_L        g12369(.A(new_n12625), .B(new_n12623), .Y(\f[63] ));
  INVx1_ASAP7_75t_L         g12370(.A(new_n12598), .Y(new_n12627));
  O2A1O1Ixp33_ASAP7_75t_L   g12371(.A1(new_n12272), .A2(new_n12604), .B(new_n12605), .C(new_n12627), .Y(new_n12628));
  A2O1A1Ixp33_ASAP7_75t_L   g12372(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n269), .Y(new_n12629));
  OAI221xp5_ASAP7_75t_L     g12373(.A1(new_n261), .A2(new_n12599), .B1(new_n12273), .B2(new_n277), .C(new_n12629), .Y(new_n12630));
  XNOR2x2_ASAP7_75t_L       g12374(.A(\a[2] ), .B(new_n12630), .Y(new_n12631));
  NOR3xp33_ASAP7_75t_L      g12375(.A(new_n12563), .B(new_n12567), .C(new_n12577), .Y(new_n12632));
  O2A1O1Ixp33_ASAP7_75t_L   g12376(.A1(new_n12578), .A2(new_n12574), .B(new_n12589), .C(new_n12632), .Y(new_n12633));
  NAND2xp33_ASAP7_75t_L     g12377(.A(new_n12558), .B(new_n12559), .Y(new_n12634));
  MAJIxp5_ASAP7_75t_L       g12378(.A(new_n12566), .B(new_n12560), .C(new_n12634), .Y(new_n12635));
  AOI22xp33_ASAP7_75t_L     g12379(.A1(new_n600), .A2(\b[55] ), .B1(new_n597), .B2(new_n9542), .Y(new_n12636));
  OAI221xp5_ASAP7_75t_L     g12380(.A1(new_n721), .A2(new_n9199), .B1(new_n8882), .B2(new_n1620), .C(new_n12636), .Y(new_n12637));
  XNOR2x2_ASAP7_75t_L       g12381(.A(\a[11] ), .B(new_n12637), .Y(new_n12638));
  INVx1_ASAP7_75t_L         g12382(.A(new_n12638), .Y(new_n12639));
  A2O1A1Ixp33_ASAP7_75t_L   g12383(.A1(new_n12233), .A2(new_n12300), .B(new_n12547), .C(new_n12545), .Y(new_n12640));
  NAND2xp33_ASAP7_75t_L     g12384(.A(\b[51] ), .B(new_n817), .Y(new_n12641));
  AOI22xp33_ASAP7_75t_L     g12385(.A1(new_n826), .A2(\b[52] ), .B1(new_n823), .B2(new_n8577), .Y(new_n12642));
  NAND2xp33_ASAP7_75t_L     g12386(.A(new_n12641), .B(new_n12642), .Y(new_n12643));
  AOI211xp5_ASAP7_75t_L     g12387(.A1(\b[50] ), .A2(new_n908), .B(new_n813), .C(new_n12643), .Y(new_n12644));
  INVx1_ASAP7_75t_L         g12388(.A(new_n12643), .Y(new_n12645));
  O2A1O1Ixp33_ASAP7_75t_L   g12389(.A1(new_n8228), .A2(new_n909), .B(new_n12645), .C(\a[14] ), .Y(new_n12646));
  NOR2xp33_ASAP7_75t_L      g12390(.A(new_n12644), .B(new_n12646), .Y(new_n12647));
  NOR2xp33_ASAP7_75t_L      g12391(.A(new_n12533), .B(new_n12538), .Y(new_n12648));
  NAND2xp33_ASAP7_75t_L     g12392(.A(new_n12313), .B(new_n12648), .Y(new_n12649));
  NAND2xp33_ASAP7_75t_L     g12393(.A(new_n1110), .B(new_n7914), .Y(new_n12650));
  OAI221xp5_ASAP7_75t_L     g12394(.A1(new_n1198), .A2(new_n7907), .B1(new_n7333), .B2(new_n1298), .C(new_n12650), .Y(new_n12651));
  AOI21xp33_ASAP7_75t_L     g12395(.A1(new_n1194), .A2(\b[47] ), .B(new_n12651), .Y(new_n12652));
  NAND2xp33_ASAP7_75t_L     g12396(.A(\a[17] ), .B(new_n12652), .Y(new_n12653));
  A2O1A1Ixp33_ASAP7_75t_L   g12397(.A1(\b[47] ), .A2(new_n1194), .B(new_n12651), .C(new_n1107), .Y(new_n12654));
  NAND2xp33_ASAP7_75t_L     g12398(.A(new_n12654), .B(new_n12653), .Y(new_n12655));
  NOR2xp33_ASAP7_75t_L      g12399(.A(new_n12522), .B(new_n12523), .Y(new_n12656));
  MAJIxp5_ASAP7_75t_L       g12400(.A(new_n12536), .B(new_n12321), .C(new_n12656), .Y(new_n12657));
  AOI22xp33_ASAP7_75t_L     g12401(.A1(new_n1406), .A2(\b[46] ), .B1(new_n1404), .B2(new_n7041), .Y(new_n12658));
  OAI221xp5_ASAP7_75t_L     g12402(.A1(new_n1398), .A2(new_n6756), .B1(new_n6220), .B2(new_n1549), .C(new_n12658), .Y(new_n12659));
  XNOR2x2_ASAP7_75t_L       g12403(.A(\a[20] ), .B(new_n12659), .Y(new_n12660));
  INVx1_ASAP7_75t_L         g12404(.A(new_n12660), .Y(new_n12661));
  NOR3xp33_ASAP7_75t_L      g12405(.A(new_n12510), .B(new_n12515), .C(new_n12324), .Y(new_n12662));
  INVx1_ASAP7_75t_L         g12406(.A(new_n12662), .Y(new_n12663));
  OAI21xp33_ASAP7_75t_L     g12407(.A1(new_n12491), .A2(new_n12492), .B(new_n12493), .Y(new_n12664));
  INVx1_ASAP7_75t_L         g12408(.A(new_n12473), .Y(new_n12665));
  AOI211xp5_ASAP7_75t_L     g12409(.A1(new_n12351), .A2(new_n12352), .B(new_n12372), .C(new_n12373), .Y(new_n12666));
  O2A1O1Ixp33_ASAP7_75t_L   g12410(.A1(new_n11665), .A2(new_n11660), .B(new_n11662), .C(new_n12031), .Y(new_n12667));
  O2A1O1Ixp33_ASAP7_75t_L   g12411(.A1(new_n12034), .A2(new_n12667), .B(new_n12374), .C(new_n12666), .Y(new_n12668));
  INVx1_ASAP7_75t_L         g12412(.A(new_n12356), .Y(new_n12669));
  NOR2xp33_ASAP7_75t_L      g12413(.A(new_n11651), .B(new_n12354), .Y(new_n12670));
  INVx1_ASAP7_75t_L         g12414(.A(new_n12670), .Y(new_n12671));
  NOR2xp33_ASAP7_75t_L      g12415(.A(new_n258), .B(new_n12671), .Y(new_n12672));
  NAND2xp33_ASAP7_75t_L     g12416(.A(new_n11654), .B(new_n328), .Y(new_n12673));
  OAI221xp5_ASAP7_75t_L     g12417(.A1(new_n12023), .A2(new_n323), .B1(new_n299), .B2(new_n12364), .C(new_n12673), .Y(new_n12674));
  AOI211xp5_ASAP7_75t_L     g12418(.A1(\b[2] ), .A2(new_n12021), .B(new_n11651), .C(new_n12674), .Y(new_n12675));
  AOI21xp33_ASAP7_75t_L     g12419(.A1(new_n12021), .A2(\b[2] ), .B(new_n12674), .Y(new_n12676));
  NOR2xp33_ASAP7_75t_L      g12420(.A(\a[62] ), .B(new_n12676), .Y(new_n12677));
  NOR2xp33_ASAP7_75t_L      g12421(.A(new_n12675), .B(new_n12677), .Y(new_n12678));
  A2O1A1Ixp33_ASAP7_75t_L   g12422(.A1(new_n12669), .A2(\b[1] ), .B(new_n12672), .C(new_n12678), .Y(new_n12679));
  O2A1O1Ixp33_ASAP7_75t_L   g12423(.A1(new_n12353), .A2(new_n12355), .B(\b[1] ), .C(new_n12672), .Y(new_n12680));
  OAI21xp33_ASAP7_75t_L     g12424(.A1(new_n12675), .A2(new_n12677), .B(new_n12680), .Y(new_n12681));
  MAJIxp5_ASAP7_75t_L       g12425(.A(new_n12360), .B(new_n12362), .C(new_n12370), .Y(new_n12682));
  NAND3xp33_ASAP7_75t_L     g12426(.A(new_n12679), .B(new_n12681), .C(new_n12682), .Y(new_n12683));
  AO21x2_ASAP7_75t_L        g12427(.A1(new_n12681), .A2(new_n12679), .B(new_n12682), .Y(new_n12684));
  AOI22xp33_ASAP7_75t_L     g12428(.A1(new_n10594), .A2(\b[7] ), .B1(new_n10591), .B2(new_n611), .Y(new_n12685));
  OAI221xp5_ASAP7_75t_L     g12429(.A1(new_n11335), .A2(new_n382), .B1(new_n353), .B2(new_n11330), .C(new_n12685), .Y(new_n12686));
  NOR2xp33_ASAP7_75t_L      g12430(.A(new_n10588), .B(new_n12686), .Y(new_n12687));
  NAND2xp33_ASAP7_75t_L     g12431(.A(new_n10588), .B(new_n12686), .Y(new_n12688));
  INVx1_ASAP7_75t_L         g12432(.A(new_n12688), .Y(new_n12689));
  AOI211xp5_ASAP7_75t_L     g12433(.A1(new_n12684), .A2(new_n12683), .B(new_n12687), .C(new_n12689), .Y(new_n12690));
  AND3x1_ASAP7_75t_L        g12434(.A(new_n12679), .B(new_n12682), .C(new_n12681), .Y(new_n12691));
  AOI21xp33_ASAP7_75t_L     g12435(.A1(new_n12679), .A2(new_n12681), .B(new_n12682), .Y(new_n12692));
  INVx1_ASAP7_75t_L         g12436(.A(new_n12687), .Y(new_n12693));
  AOI211xp5_ASAP7_75t_L     g12437(.A1(new_n12693), .A2(new_n12688), .B(new_n12692), .C(new_n12691), .Y(new_n12694));
  OR3x1_ASAP7_75t_L         g12438(.A(new_n12690), .B(new_n12668), .C(new_n12694), .Y(new_n12695));
  OAI21xp33_ASAP7_75t_L     g12439(.A1(new_n12694), .A2(new_n12690), .B(new_n12668), .Y(new_n12696));
  NAND2xp33_ASAP7_75t_L     g12440(.A(\b[10] ), .B(new_n9623), .Y(new_n12697));
  OAI221xp5_ASAP7_75t_L     g12441(.A1(new_n559), .A2(new_n10280), .B1(new_n9949), .B2(new_n641), .C(new_n12697), .Y(new_n12698));
  AOI21xp33_ASAP7_75t_L     g12442(.A1(new_n9948), .A2(\b[8] ), .B(new_n12698), .Y(new_n12699));
  NAND2xp33_ASAP7_75t_L     g12443(.A(\a[56] ), .B(new_n12699), .Y(new_n12700));
  A2O1A1Ixp33_ASAP7_75t_L   g12444(.A1(\b[8] ), .A2(new_n9948), .B(new_n12698), .C(new_n9610), .Y(new_n12701));
  NAND4xp25_ASAP7_75t_L     g12445(.A(new_n12695), .B(new_n12701), .C(new_n12700), .D(new_n12696), .Y(new_n12702));
  NOR3xp33_ASAP7_75t_L      g12446(.A(new_n12690), .B(new_n12668), .C(new_n12694), .Y(new_n12703));
  OA21x2_ASAP7_75t_L        g12447(.A1(new_n12694), .A2(new_n12690), .B(new_n12668), .Y(new_n12704));
  NAND2xp33_ASAP7_75t_L     g12448(.A(new_n12701), .B(new_n12700), .Y(new_n12705));
  OAI21xp33_ASAP7_75t_L     g12449(.A1(new_n12703), .A2(new_n12704), .B(new_n12705), .Y(new_n12706));
  NAND2xp33_ASAP7_75t_L     g12450(.A(new_n12706), .B(new_n12702), .Y(new_n12707));
  NAND2xp33_ASAP7_75t_L     g12451(.A(new_n12379), .B(new_n12380), .Y(new_n12708));
  MAJIxp5_ASAP7_75t_L       g12452(.A(new_n12348), .B(new_n12385), .C(new_n12708), .Y(new_n12709));
  NOR2xp33_ASAP7_75t_L      g12453(.A(new_n12709), .B(new_n12707), .Y(new_n12710));
  MAJx2_ASAP7_75t_L         g12454(.A(new_n12348), .B(new_n12708), .C(new_n12385), .Y(new_n12711));
  AOI21xp33_ASAP7_75t_L     g12455(.A1(new_n12706), .A2(new_n12702), .B(new_n12711), .Y(new_n12712));
  AOI22xp33_ASAP7_75t_L     g12456(.A1(new_n8645), .A2(\b[13] ), .B1(new_n8642), .B2(new_n800), .Y(new_n12713));
  OAI221xp5_ASAP7_75t_L     g12457(.A1(new_n9322), .A2(new_n763), .B1(new_n695), .B2(new_n8965), .C(new_n12713), .Y(new_n12714));
  XNOR2x2_ASAP7_75t_L       g12458(.A(\a[53] ), .B(new_n12714), .Y(new_n12715));
  OAI21xp33_ASAP7_75t_L     g12459(.A1(new_n12712), .A2(new_n12710), .B(new_n12715), .Y(new_n12716));
  NAND3xp33_ASAP7_75t_L     g12460(.A(new_n12711), .B(new_n12706), .C(new_n12702), .Y(new_n12717));
  NAND2xp33_ASAP7_75t_L     g12461(.A(new_n12709), .B(new_n12707), .Y(new_n12718));
  INVx1_ASAP7_75t_L         g12462(.A(new_n12715), .Y(new_n12719));
  NAND3xp33_ASAP7_75t_L     g12463(.A(new_n12717), .B(new_n12718), .C(new_n12719), .Y(new_n12720));
  A2O1A1Ixp33_ASAP7_75t_L   g12464(.A1(new_n12051), .A2(new_n12050), .B(new_n12397), .C(new_n12394), .Y(new_n12721));
  NAND3xp33_ASAP7_75t_L     g12465(.A(new_n12721), .B(new_n12716), .C(new_n12720), .Y(new_n12722));
  AOI21xp33_ASAP7_75t_L     g12466(.A1(new_n12717), .A2(new_n12718), .B(new_n12719), .Y(new_n12723));
  NOR3xp33_ASAP7_75t_L      g12467(.A(new_n12710), .B(new_n12712), .C(new_n12715), .Y(new_n12724));
  A2O1A1O1Ixp25_ASAP7_75t_L g12468(.A1(new_n12049), .A2(new_n12002), .B(new_n12055), .C(new_n12390), .D(new_n12398), .Y(new_n12725));
  OAI21xp33_ASAP7_75t_L     g12469(.A1(new_n12723), .A2(new_n12724), .B(new_n12725), .Y(new_n12726));
  AOI22xp33_ASAP7_75t_L     g12470(.A1(new_n7659), .A2(\b[16] ), .B1(new_n7656), .B2(new_n1058), .Y(new_n12727));
  OAI221xp5_ASAP7_75t_L     g12471(.A1(new_n8326), .A2(new_n952), .B1(new_n871), .B2(new_n7994), .C(new_n12727), .Y(new_n12728));
  XNOR2x2_ASAP7_75t_L       g12472(.A(\a[50] ), .B(new_n12728), .Y(new_n12729));
  NAND3xp33_ASAP7_75t_L     g12473(.A(new_n12726), .B(new_n12722), .C(new_n12729), .Y(new_n12730));
  NOR3xp33_ASAP7_75t_L      g12474(.A(new_n12725), .B(new_n12724), .C(new_n12723), .Y(new_n12731));
  AOI21xp33_ASAP7_75t_L     g12475(.A1(new_n12716), .A2(new_n12720), .B(new_n12721), .Y(new_n12732));
  INVx1_ASAP7_75t_L         g12476(.A(new_n12729), .Y(new_n12733));
  OAI21xp33_ASAP7_75t_L     g12477(.A1(new_n12732), .A2(new_n12731), .B(new_n12733), .Y(new_n12734));
  NAND2xp33_ASAP7_75t_L     g12478(.A(new_n12730), .B(new_n12734), .Y(new_n12735));
  A2O1A1Ixp33_ASAP7_75t_L   g12479(.A1(new_n11378), .A2(new_n11377), .B(new_n11708), .C(new_n11705), .Y(new_n12736));
  AND3x1_ASAP7_75t_L        g12480(.A(new_n12411), .B(new_n12056), .C(new_n12051), .Y(new_n12737));
  O2A1O1Ixp33_ASAP7_75t_L   g12481(.A1(new_n12067), .A2(new_n12068), .B(new_n12736), .C(new_n12737), .Y(new_n12738));
  NOR2xp33_ASAP7_75t_L      g12482(.A(new_n12408), .B(new_n12407), .Y(new_n12739));
  NAND2xp33_ASAP7_75t_L     g12483(.A(new_n12409), .B(new_n12739), .Y(new_n12740));
  A2O1A1Ixp33_ASAP7_75t_L   g12484(.A1(new_n12410), .A2(new_n12406), .B(new_n12738), .C(new_n12740), .Y(new_n12741));
  NOR2xp33_ASAP7_75t_L      g12485(.A(new_n12741), .B(new_n12735), .Y(new_n12742));
  AOI22xp33_ASAP7_75t_L     g12486(.A1(new_n12730), .A2(new_n12734), .B1(new_n12740), .B2(new_n12420), .Y(new_n12743));
  AOI22xp33_ASAP7_75t_L     g12487(.A1(new_n6822), .A2(\b[19] ), .B1(new_n6819), .B2(new_n1499), .Y(new_n12744));
  OAI221xp5_ASAP7_75t_L     g12488(.A1(new_n7392), .A2(new_n1356), .B1(new_n1244), .B2(new_n7115), .C(new_n12744), .Y(new_n12745));
  XNOR2x2_ASAP7_75t_L       g12489(.A(\a[47] ), .B(new_n12745), .Y(new_n12746));
  OAI21xp33_ASAP7_75t_L     g12490(.A1(new_n12743), .A2(new_n12742), .B(new_n12746), .Y(new_n12747));
  NAND4xp25_ASAP7_75t_L     g12491(.A(new_n12420), .B(new_n12740), .C(new_n12734), .D(new_n12730), .Y(new_n12748));
  NAND2xp33_ASAP7_75t_L     g12492(.A(new_n12741), .B(new_n12735), .Y(new_n12749));
  INVx1_ASAP7_75t_L         g12493(.A(new_n12746), .Y(new_n12750));
  NAND3xp33_ASAP7_75t_L     g12494(.A(new_n12749), .B(new_n12748), .C(new_n12750), .Y(new_n12751));
  INVx1_ASAP7_75t_L         g12495(.A(new_n12340), .Y(new_n12752));
  NOR3xp33_ASAP7_75t_L      g12496(.A(new_n12413), .B(new_n12414), .C(new_n12417), .Y(new_n12753));
  A2O1A1O1Ixp25_ASAP7_75t_L g12497(.A1(new_n12087), .A2(new_n12076), .B(new_n12752), .C(new_n12418), .D(new_n12753), .Y(new_n12754));
  INVx1_ASAP7_75t_L         g12498(.A(new_n12754), .Y(new_n12755));
  NAND3xp33_ASAP7_75t_L     g12499(.A(new_n12755), .B(new_n12751), .C(new_n12747), .Y(new_n12756));
  AOI21xp33_ASAP7_75t_L     g12500(.A1(new_n12749), .A2(new_n12748), .B(new_n12750), .Y(new_n12757));
  NOR3xp33_ASAP7_75t_L      g12501(.A(new_n12742), .B(new_n12743), .C(new_n12746), .Y(new_n12758));
  OAI21xp33_ASAP7_75t_L     g12502(.A1(new_n12757), .A2(new_n12758), .B(new_n12754), .Y(new_n12759));
  AOI22xp33_ASAP7_75t_L     g12503(.A1(new_n6002), .A2(\b[22] ), .B1(new_n5999), .B2(new_n1864), .Y(new_n12760));
  OAI221xp5_ASAP7_75t_L     g12504(.A1(new_n6544), .A2(new_n1709), .B1(new_n1594), .B2(new_n6309), .C(new_n12760), .Y(new_n12761));
  XNOR2x2_ASAP7_75t_L       g12505(.A(\a[44] ), .B(new_n12761), .Y(new_n12762));
  NAND3xp33_ASAP7_75t_L     g12506(.A(new_n12756), .B(new_n12759), .C(new_n12762), .Y(new_n12763));
  NOR3xp33_ASAP7_75t_L      g12507(.A(new_n12758), .B(new_n12757), .C(new_n12754), .Y(new_n12764));
  AOI21xp33_ASAP7_75t_L     g12508(.A1(new_n12751), .A2(new_n12747), .B(new_n12755), .Y(new_n12765));
  XNOR2x2_ASAP7_75t_L       g12509(.A(new_n5996), .B(new_n12761), .Y(new_n12766));
  OAI21xp33_ASAP7_75t_L     g12510(.A1(new_n12764), .A2(new_n12765), .B(new_n12766), .Y(new_n12767));
  NAND2xp33_ASAP7_75t_L     g12511(.A(new_n12763), .B(new_n12767), .Y(new_n12768));
  A2O1A1Ixp33_ASAP7_75t_L   g12512(.A1(new_n12084), .A2(new_n12091), .B(new_n12432), .C(new_n12426), .Y(new_n12769));
  NOR2xp33_ASAP7_75t_L      g12513(.A(new_n12768), .B(new_n12769), .Y(new_n12770));
  INVx1_ASAP7_75t_L         g12514(.A(new_n12426), .Y(new_n12771));
  A2O1A1O1Ixp25_ASAP7_75t_L g12515(.A1(new_n12089), .A2(new_n12090), .B(new_n12430), .C(new_n12428), .D(new_n12771), .Y(new_n12772));
  AOI21xp33_ASAP7_75t_L     g12516(.A1(new_n12767), .A2(new_n12763), .B(new_n12772), .Y(new_n12773));
  AOI22xp33_ASAP7_75t_L     g12517(.A1(new_n5249), .A2(\b[25] ), .B1(new_n5247), .B2(new_n2188), .Y(new_n12774));
  OAI221xp5_ASAP7_75t_L     g12518(.A1(new_n5241), .A2(new_n2019), .B1(new_n1995), .B2(new_n5521), .C(new_n12774), .Y(new_n12775));
  XNOR2x2_ASAP7_75t_L       g12519(.A(new_n5244), .B(new_n12775), .Y(new_n12776));
  NOR3xp33_ASAP7_75t_L      g12520(.A(new_n12770), .B(new_n12773), .C(new_n12776), .Y(new_n12777));
  NAND3xp33_ASAP7_75t_L     g12521(.A(new_n12772), .B(new_n12767), .C(new_n12763), .Y(new_n12778));
  A2O1A1Ixp33_ASAP7_75t_L   g12522(.A1(new_n12428), .A2(new_n12335), .B(new_n12771), .C(new_n12768), .Y(new_n12779));
  XNOR2x2_ASAP7_75t_L       g12523(.A(\a[41] ), .B(new_n12775), .Y(new_n12780));
  AOI21xp33_ASAP7_75t_L     g12524(.A1(new_n12779), .A2(new_n12778), .B(new_n12780), .Y(new_n12781));
  NOR2xp33_ASAP7_75t_L      g12525(.A(new_n12781), .B(new_n12777), .Y(new_n12782));
  NAND2xp33_ASAP7_75t_L     g12526(.A(new_n12437), .B(new_n12441), .Y(new_n12783));
  NOR3xp33_ASAP7_75t_L      g12527(.A(new_n12438), .B(new_n12439), .C(new_n12436), .Y(new_n12784));
  O2A1O1Ixp33_ASAP7_75t_L   g12528(.A1(new_n12111), .A2(new_n12103), .B(new_n12783), .C(new_n12784), .Y(new_n12785));
  NAND2xp33_ASAP7_75t_L     g12529(.A(new_n12782), .B(new_n12785), .Y(new_n12786));
  NOR2xp33_ASAP7_75t_L      g12530(.A(new_n12439), .B(new_n12438), .Y(new_n12787));
  NAND3xp33_ASAP7_75t_L     g12531(.A(new_n12779), .B(new_n12778), .C(new_n12780), .Y(new_n12788));
  OAI21xp33_ASAP7_75t_L     g12532(.A1(new_n12773), .A2(new_n12770), .B(new_n12776), .Y(new_n12789));
  NAND2xp33_ASAP7_75t_L     g12533(.A(new_n12788), .B(new_n12789), .Y(new_n12790));
  A2O1A1Ixp33_ASAP7_75t_L   g12534(.A1(new_n12440), .A2(new_n12787), .B(new_n12444), .C(new_n12790), .Y(new_n12791));
  AOI22xp33_ASAP7_75t_L     g12535(.A1(new_n4544), .A2(\b[28] ), .B1(new_n4542), .B2(new_n2858), .Y(new_n12792));
  OAI221xp5_ASAP7_75t_L     g12536(.A1(new_n4536), .A2(new_n2650), .B1(new_n2477), .B2(new_n4781), .C(new_n12792), .Y(new_n12793));
  XNOR2x2_ASAP7_75t_L       g12537(.A(\a[38] ), .B(new_n12793), .Y(new_n12794));
  NAND3xp33_ASAP7_75t_L     g12538(.A(new_n12786), .B(new_n12791), .C(new_n12794), .Y(new_n12795));
  NAND2xp33_ASAP7_75t_L     g12539(.A(new_n12440), .B(new_n12787), .Y(new_n12796));
  A2O1A1Ixp33_ASAP7_75t_L   g12540(.A1(new_n12441), .A2(new_n12437), .B(new_n12442), .C(new_n12796), .Y(new_n12797));
  NOR2xp33_ASAP7_75t_L      g12541(.A(new_n12797), .B(new_n12790), .Y(new_n12798));
  NOR2xp33_ASAP7_75t_L      g12542(.A(new_n12782), .B(new_n12785), .Y(new_n12799));
  INVx1_ASAP7_75t_L         g12543(.A(new_n12794), .Y(new_n12800));
  OAI21xp33_ASAP7_75t_L     g12544(.A1(new_n12798), .A2(new_n12799), .B(new_n12800), .Y(new_n12801));
  NAND2xp33_ASAP7_75t_L     g12545(.A(new_n12795), .B(new_n12801), .Y(new_n12802));
  NOR3xp33_ASAP7_75t_L      g12546(.A(new_n12454), .B(new_n12444), .C(new_n12452), .Y(new_n12803));
  INVx1_ASAP7_75t_L         g12547(.A(new_n12803), .Y(new_n12804));
  A2O1A1Ixp33_ASAP7_75t_L   g12548(.A1(new_n12455), .A2(new_n12453), .B(new_n12464), .C(new_n12804), .Y(new_n12805));
  NOR2xp33_ASAP7_75t_L      g12549(.A(new_n12802), .B(new_n12805), .Y(new_n12806));
  O2A1O1Ixp33_ASAP7_75t_L   g12550(.A1(new_n12461), .A2(new_n12462), .B(new_n12459), .C(new_n12803), .Y(new_n12807));
  AOI21xp33_ASAP7_75t_L     g12551(.A1(new_n12801), .A2(new_n12795), .B(new_n12807), .Y(new_n12808));
  AOI22xp33_ASAP7_75t_L     g12552(.A1(new_n3884), .A2(\b[31] ), .B1(new_n3881), .B2(new_n3426), .Y(new_n12809));
  OAI221xp5_ASAP7_75t_L     g12553(.A1(new_n4312), .A2(new_n3212), .B1(new_n2871), .B2(new_n4986), .C(new_n12809), .Y(new_n12810));
  XNOR2x2_ASAP7_75t_L       g12554(.A(\a[35] ), .B(new_n12810), .Y(new_n12811));
  OA21x2_ASAP7_75t_L        g12555(.A1(new_n12808), .A2(new_n12806), .B(new_n12811), .Y(new_n12812));
  NOR3xp33_ASAP7_75t_L      g12556(.A(new_n12806), .B(new_n12808), .C(new_n12811), .Y(new_n12813));
  NOR2xp33_ASAP7_75t_L      g12557(.A(new_n12813), .B(new_n12812), .Y(new_n12814));
  A2O1A1Ixp33_ASAP7_75t_L   g12558(.A1(new_n12475), .A2(new_n12469), .B(new_n12665), .C(new_n12814), .Y(new_n12815));
  A2O1A1O1Ixp25_ASAP7_75t_L g12559(.A1(new_n12136), .A2(new_n12133), .B(new_n12477), .C(new_n12469), .D(new_n12665), .Y(new_n12816));
  OAI21xp33_ASAP7_75t_L     g12560(.A1(new_n12813), .A2(new_n12812), .B(new_n12816), .Y(new_n12817));
  AOI22xp33_ASAP7_75t_L     g12561(.A1(new_n3256), .A2(\b[34] ), .B1(new_n3254), .B2(new_n3833), .Y(new_n12818));
  OAI221xp5_ASAP7_75t_L     g12562(.A1(new_n3248), .A2(new_n3807), .B1(new_n3443), .B2(new_n3492), .C(new_n12818), .Y(new_n12819));
  XNOR2x2_ASAP7_75t_L       g12563(.A(\a[32] ), .B(new_n12819), .Y(new_n12820));
  NAND3xp33_ASAP7_75t_L     g12564(.A(new_n12815), .B(new_n12817), .C(new_n12820), .Y(new_n12821));
  NOR3xp33_ASAP7_75t_L      g12565(.A(new_n12816), .B(new_n12812), .C(new_n12813), .Y(new_n12822));
  A2O1A1Ixp33_ASAP7_75t_L   g12566(.A1(new_n12147), .A2(new_n12474), .B(new_n12484), .C(new_n12473), .Y(new_n12823));
  NOR2xp33_ASAP7_75t_L      g12567(.A(new_n12823), .B(new_n12814), .Y(new_n12824));
  INVx1_ASAP7_75t_L         g12568(.A(new_n12820), .Y(new_n12825));
  OAI21xp33_ASAP7_75t_L     g12569(.A1(new_n12822), .A2(new_n12824), .B(new_n12825), .Y(new_n12826));
  NAND3xp33_ASAP7_75t_L     g12570(.A(new_n12476), .B(new_n12479), .C(new_n12487), .Y(new_n12827));
  NAND4xp25_ASAP7_75t_L     g12571(.A(new_n12821), .B(new_n12826), .C(new_n12664), .D(new_n12827), .Y(new_n12828));
  NOR3xp33_ASAP7_75t_L      g12572(.A(new_n12824), .B(new_n12825), .C(new_n12822), .Y(new_n12829));
  AOI21xp33_ASAP7_75t_L     g12573(.A1(new_n12815), .A2(new_n12817), .B(new_n12820), .Y(new_n12830));
  A2O1A1Ixp33_ASAP7_75t_L   g12574(.A1(new_n12483), .A2(new_n12488), .B(new_n12489), .C(new_n12827), .Y(new_n12831));
  OAI21xp33_ASAP7_75t_L     g12575(.A1(new_n12829), .A2(new_n12830), .B(new_n12831), .Y(new_n12832));
  AOI22xp33_ASAP7_75t_L     g12576(.A1(new_n2702), .A2(\b[37] ), .B1(new_n2700), .B2(new_n4709), .Y(new_n12833));
  OAI221xp5_ASAP7_75t_L     g12577(.A1(new_n2694), .A2(new_n4465), .B1(new_n4053), .B2(new_n2932), .C(new_n12833), .Y(new_n12834));
  XNOR2x2_ASAP7_75t_L       g12578(.A(\a[29] ), .B(new_n12834), .Y(new_n12835));
  AND3x1_ASAP7_75t_L        g12579(.A(new_n12832), .B(new_n12828), .C(new_n12835), .Y(new_n12836));
  AOI21xp33_ASAP7_75t_L     g12580(.A1(new_n12832), .A2(new_n12828), .B(new_n12835), .Y(new_n12837));
  OAI21xp33_ASAP7_75t_L     g12581(.A1(new_n12330), .A2(new_n12496), .B(new_n12498), .Y(new_n12838));
  OR3x1_ASAP7_75t_L         g12582(.A(new_n12836), .B(new_n12838), .C(new_n12837), .Y(new_n12839));
  OAI21xp33_ASAP7_75t_L     g12583(.A1(new_n12837), .A2(new_n12836), .B(new_n12838), .Y(new_n12840));
  AOI22xp33_ASAP7_75t_L     g12584(.A1(new_n2228), .A2(\b[40] ), .B1(new_n2226), .B2(new_n5194), .Y(new_n12841));
  OAI221xp5_ASAP7_75t_L     g12585(.A1(new_n2220), .A2(new_n5166), .B1(new_n4915), .B2(new_n2387), .C(new_n12841), .Y(new_n12842));
  XNOR2x2_ASAP7_75t_L       g12586(.A(\a[26] ), .B(new_n12842), .Y(new_n12843));
  NAND3xp33_ASAP7_75t_L     g12587(.A(new_n12839), .B(new_n12840), .C(new_n12843), .Y(new_n12844));
  NOR3xp33_ASAP7_75t_L      g12588(.A(new_n12836), .B(new_n12838), .C(new_n12837), .Y(new_n12845));
  OA21x2_ASAP7_75t_L        g12589(.A1(new_n12837), .A2(new_n12836), .B(new_n12838), .Y(new_n12846));
  INVx1_ASAP7_75t_L         g12590(.A(new_n12843), .Y(new_n12847));
  OAI21xp33_ASAP7_75t_L     g12591(.A1(new_n12845), .A2(new_n12846), .B(new_n12847), .Y(new_n12848));
  A2O1A1O1Ixp25_ASAP7_75t_L g12592(.A1(new_n12176), .A2(new_n12175), .B(new_n12327), .C(new_n12507), .D(new_n12513), .Y(new_n12849));
  INVx1_ASAP7_75t_L         g12593(.A(new_n12849), .Y(new_n12850));
  AOI21xp33_ASAP7_75t_L     g12594(.A1(new_n12848), .A2(new_n12844), .B(new_n12850), .Y(new_n12851));
  NAND2xp33_ASAP7_75t_L     g12595(.A(new_n12848), .B(new_n12844), .Y(new_n12852));
  O2A1O1Ixp33_ASAP7_75t_L   g12596(.A1(new_n12518), .A2(new_n12512), .B(new_n12508), .C(new_n12852), .Y(new_n12853));
  AOI22xp33_ASAP7_75t_L     g12597(.A1(new_n1766), .A2(\b[43] ), .B1(new_n1764), .B2(new_n6202), .Y(new_n12854));
  OAI221xp5_ASAP7_75t_L     g12598(.A1(new_n1758), .A2(new_n5680), .B1(new_n5666), .B2(new_n1911), .C(new_n12854), .Y(new_n12855));
  XNOR2x2_ASAP7_75t_L       g12599(.A(\a[23] ), .B(new_n12855), .Y(new_n12856));
  INVx1_ASAP7_75t_L         g12600(.A(new_n12856), .Y(new_n12857));
  OAI21xp33_ASAP7_75t_L     g12601(.A1(new_n12853), .A2(new_n12851), .B(new_n12857), .Y(new_n12858));
  NAND2xp33_ASAP7_75t_L     g12602(.A(new_n12849), .B(new_n12852), .Y(new_n12859));
  NAND3xp33_ASAP7_75t_L     g12603(.A(new_n12850), .B(new_n12848), .C(new_n12844), .Y(new_n12860));
  NAND3xp33_ASAP7_75t_L     g12604(.A(new_n12860), .B(new_n12859), .C(new_n12856), .Y(new_n12861));
  NAND2xp33_ASAP7_75t_L     g12605(.A(new_n12861), .B(new_n12858), .Y(new_n12862));
  A2O1A1O1Ixp25_ASAP7_75t_L g12606(.A1(new_n12520), .A2(new_n12516), .B(new_n12521), .C(new_n12663), .D(new_n12862), .Y(new_n12863));
  A2O1A1Ixp33_ASAP7_75t_L   g12607(.A1(new_n12520), .A2(new_n12516), .B(new_n12521), .C(new_n12663), .Y(new_n12864));
  AOI21xp33_ASAP7_75t_L     g12608(.A1(new_n12861), .A2(new_n12858), .B(new_n12864), .Y(new_n12865));
  OAI21xp33_ASAP7_75t_L     g12609(.A1(new_n12865), .A2(new_n12863), .B(new_n12661), .Y(new_n12866));
  NAND3xp33_ASAP7_75t_L     g12610(.A(new_n12864), .B(new_n12858), .C(new_n12861), .Y(new_n12867));
  A2O1A1O1Ixp25_ASAP7_75t_L g12611(.A1(new_n11840), .A2(new_n11839), .B(new_n11837), .C(new_n12193), .D(new_n12182), .Y(new_n12868));
  O2A1O1Ixp33_ASAP7_75t_L   g12612(.A1(new_n12185), .A2(new_n12868), .B(new_n12525), .C(new_n12662), .Y(new_n12869));
  NAND2xp33_ASAP7_75t_L     g12613(.A(new_n12869), .B(new_n12862), .Y(new_n12870));
  NAND3xp33_ASAP7_75t_L     g12614(.A(new_n12870), .B(new_n12867), .C(new_n12660), .Y(new_n12871));
  AOI21xp33_ASAP7_75t_L     g12615(.A1(new_n12866), .A2(new_n12871), .B(new_n12657), .Y(new_n12872));
  NAND2xp33_ASAP7_75t_L     g12616(.A(new_n12321), .B(new_n12656), .Y(new_n12873));
  A2O1A1Ixp33_ASAP7_75t_L   g12617(.A1(new_n12524), .A2(new_n12529), .B(new_n12315), .C(new_n12873), .Y(new_n12874));
  AOI21xp33_ASAP7_75t_L     g12618(.A1(new_n12870), .A2(new_n12867), .B(new_n12660), .Y(new_n12875));
  NOR3xp33_ASAP7_75t_L      g12619(.A(new_n12863), .B(new_n12865), .C(new_n12661), .Y(new_n12876));
  NOR3xp33_ASAP7_75t_L      g12620(.A(new_n12874), .B(new_n12876), .C(new_n12875), .Y(new_n12877));
  OAI21xp33_ASAP7_75t_L     g12621(.A1(new_n12872), .A2(new_n12877), .B(new_n12655), .Y(new_n12878));
  INVx1_ASAP7_75t_L         g12622(.A(new_n12655), .Y(new_n12879));
  OAI21xp33_ASAP7_75t_L     g12623(.A1(new_n12875), .A2(new_n12876), .B(new_n12874), .Y(new_n12880));
  NAND3xp33_ASAP7_75t_L     g12624(.A(new_n12866), .B(new_n12657), .C(new_n12871), .Y(new_n12881));
  NAND3xp33_ASAP7_75t_L     g12625(.A(new_n12880), .B(new_n12881), .C(new_n12879), .Y(new_n12882));
  AOI22xp33_ASAP7_75t_L     g12626(.A1(new_n12878), .A2(new_n12882), .B1(new_n12649), .B2(new_n12540), .Y(new_n12883));
  AND4x1_ASAP7_75t_L        g12627(.A(new_n12540), .B(new_n12882), .C(new_n12649), .D(new_n12878), .Y(new_n12884));
  NOR3xp33_ASAP7_75t_L      g12628(.A(new_n12884), .B(new_n12647), .C(new_n12883), .Y(new_n12885));
  INVx1_ASAP7_75t_L         g12629(.A(new_n12647), .Y(new_n12886));
  MAJx2_ASAP7_75t_L         g12630(.A(new_n12307), .B(new_n12313), .C(new_n12648), .Y(new_n12887));
  AOI21xp33_ASAP7_75t_L     g12631(.A1(new_n12880), .A2(new_n12881), .B(new_n12879), .Y(new_n12888));
  NOR3xp33_ASAP7_75t_L      g12632(.A(new_n12877), .B(new_n12872), .C(new_n12655), .Y(new_n12889));
  OAI21xp33_ASAP7_75t_L     g12633(.A1(new_n12888), .A2(new_n12889), .B(new_n12887), .Y(new_n12890));
  NAND4xp25_ASAP7_75t_L     g12634(.A(new_n12540), .B(new_n12882), .C(new_n12878), .D(new_n12649), .Y(new_n12891));
  AOI21xp33_ASAP7_75t_L     g12635(.A1(new_n12890), .A2(new_n12891), .B(new_n12886), .Y(new_n12892));
  NOR2xp33_ASAP7_75t_L      g12636(.A(new_n12892), .B(new_n12885), .Y(new_n12893));
  NAND2xp33_ASAP7_75t_L     g12637(.A(new_n12640), .B(new_n12893), .Y(new_n12894));
  INVx1_ASAP7_75t_L         g12638(.A(new_n12300), .Y(new_n12895));
  INVx1_ASAP7_75t_L         g12639(.A(new_n12545), .Y(new_n12896));
  O2A1O1Ixp33_ASAP7_75t_L   g12640(.A1(new_n12895), .A2(new_n12229), .B(new_n12546), .C(new_n12896), .Y(new_n12897));
  OAI21xp33_ASAP7_75t_L     g12641(.A1(new_n12885), .A2(new_n12892), .B(new_n12897), .Y(new_n12898));
  NAND3xp33_ASAP7_75t_L     g12642(.A(new_n12894), .B(new_n12898), .C(new_n12639), .Y(new_n12899));
  NOR3xp33_ASAP7_75t_L      g12643(.A(new_n12897), .B(new_n12885), .C(new_n12892), .Y(new_n12900));
  NAND3xp33_ASAP7_75t_L     g12644(.A(new_n12890), .B(new_n12886), .C(new_n12891), .Y(new_n12901));
  OAI21xp33_ASAP7_75t_L     g12645(.A1(new_n12883), .A2(new_n12884), .B(new_n12647), .Y(new_n12902));
  AOI221xp5_ASAP7_75t_L     g12646(.A1(new_n12549), .A2(new_n12546), .B1(new_n12901), .B2(new_n12902), .C(new_n12896), .Y(new_n12903));
  OAI21xp33_ASAP7_75t_L     g12647(.A1(new_n12903), .A2(new_n12900), .B(new_n12638), .Y(new_n12904));
  NAND3xp33_ASAP7_75t_L     g12648(.A(new_n12635), .B(new_n12899), .C(new_n12904), .Y(new_n12905));
  NOR2xp33_ASAP7_75t_L      g12649(.A(new_n12560), .B(new_n12634), .Y(new_n12906));
  O2A1O1Ixp33_ASAP7_75t_L   g12650(.A1(new_n12557), .A2(new_n12561), .B(new_n12562), .C(new_n12906), .Y(new_n12907));
  NAND2xp33_ASAP7_75t_L     g12651(.A(new_n12904), .B(new_n12899), .Y(new_n12908));
  NAND2xp33_ASAP7_75t_L     g12652(.A(new_n12907), .B(new_n12908), .Y(new_n12909));
  AOI22xp33_ASAP7_75t_L     g12653(.A1(new_n451), .A2(\b[58] ), .B1(new_n448), .B2(new_n10857), .Y(new_n12910));
  OAI221xp5_ASAP7_75t_L     g12654(.A1(new_n529), .A2(new_n10488), .B1(new_n10178), .B2(new_n481), .C(new_n12910), .Y(new_n12911));
  XNOR2x2_ASAP7_75t_L       g12655(.A(\a[8] ), .B(new_n12911), .Y(new_n12912));
  NAND3xp33_ASAP7_75t_L     g12656(.A(new_n12909), .B(new_n12905), .C(new_n12912), .Y(new_n12913));
  NOR2xp33_ASAP7_75t_L      g12657(.A(new_n12907), .B(new_n12908), .Y(new_n12914));
  AOI21xp33_ASAP7_75t_L     g12658(.A1(new_n12904), .A2(new_n12899), .B(new_n12635), .Y(new_n12915));
  INVx1_ASAP7_75t_L         g12659(.A(new_n12912), .Y(new_n12916));
  OAI21xp33_ASAP7_75t_L     g12660(.A1(new_n12915), .A2(new_n12914), .B(new_n12916), .Y(new_n12917));
  NAND2xp33_ASAP7_75t_L     g12661(.A(\b[59] ), .B(new_n366), .Y(new_n12918));
  NAND2xp33_ASAP7_75t_L     g12662(.A(\b[60] ), .B(new_n334), .Y(new_n12919));
  AOI22xp33_ASAP7_75t_L     g12663(.A1(new_n345), .A2(\b[61] ), .B1(new_n342), .B2(new_n11919), .Y(new_n12920));
  AND4x1_ASAP7_75t_L        g12664(.A(new_n12920), .B(new_n12919), .C(new_n12918), .D(\a[5] ), .Y(new_n12921));
  AOI31xp33_ASAP7_75t_L     g12665(.A1(new_n12920), .A2(new_n12919), .A3(new_n12918), .B(\a[5] ), .Y(new_n12922));
  NOR2xp33_ASAP7_75t_L      g12666(.A(new_n12922), .B(new_n12921), .Y(new_n12923));
  AOI21xp33_ASAP7_75t_L     g12667(.A1(new_n12917), .A2(new_n12913), .B(new_n12923), .Y(new_n12924));
  NOR3xp33_ASAP7_75t_L      g12668(.A(new_n12914), .B(new_n12915), .C(new_n12916), .Y(new_n12925));
  AOI21xp33_ASAP7_75t_L     g12669(.A1(new_n12909), .A2(new_n12905), .B(new_n12912), .Y(new_n12926));
  INVx1_ASAP7_75t_L         g12670(.A(new_n12923), .Y(new_n12927));
  NOR3xp33_ASAP7_75t_L      g12671(.A(new_n12925), .B(new_n12926), .C(new_n12927), .Y(new_n12928));
  NOR3xp33_ASAP7_75t_L      g12672(.A(new_n12928), .B(new_n12924), .C(new_n12633), .Y(new_n12929));
  INVx1_ASAP7_75t_L         g12673(.A(new_n12633), .Y(new_n12930));
  OAI21xp33_ASAP7_75t_L     g12674(.A1(new_n12926), .A2(new_n12925), .B(new_n12927), .Y(new_n12931));
  NAND3xp33_ASAP7_75t_L     g12675(.A(new_n12917), .B(new_n12913), .C(new_n12923), .Y(new_n12932));
  AOI21xp33_ASAP7_75t_L     g12676(.A1(new_n12931), .A2(new_n12932), .B(new_n12930), .Y(new_n12933));
  NOR3xp33_ASAP7_75t_L      g12677(.A(new_n12929), .B(new_n12933), .C(new_n12631), .Y(new_n12934));
  INVx1_ASAP7_75t_L         g12678(.A(new_n12631), .Y(new_n12935));
  NAND3xp33_ASAP7_75t_L     g12679(.A(new_n12931), .B(new_n12932), .C(new_n12930), .Y(new_n12936));
  OAI21xp33_ASAP7_75t_L     g12680(.A1(new_n12924), .A2(new_n12928), .B(new_n12633), .Y(new_n12937));
  AOI21xp33_ASAP7_75t_L     g12681(.A1(new_n12937), .A2(new_n12936), .B(new_n12935), .Y(new_n12938));
  AOI21xp33_ASAP7_75t_L     g12682(.A1(new_n12613), .A2(new_n12596), .B(new_n12615), .Y(new_n12939));
  INVx1_ASAP7_75t_L         g12683(.A(new_n12939), .Y(new_n12940));
  NOR3xp33_ASAP7_75t_L      g12684(.A(new_n12934), .B(new_n12938), .C(new_n12940), .Y(new_n12941));
  NAND3xp33_ASAP7_75t_L     g12685(.A(new_n12937), .B(new_n12936), .C(new_n12935), .Y(new_n12942));
  OAI21xp33_ASAP7_75t_L     g12686(.A1(new_n12933), .A2(new_n12929), .B(new_n12631), .Y(new_n12943));
  AOI21xp33_ASAP7_75t_L     g12687(.A1(new_n12943), .A2(new_n12942), .B(new_n12939), .Y(new_n12944));
  NOR2xp33_ASAP7_75t_L      g12688(.A(new_n12944), .B(new_n12941), .Y(new_n12945));
  INVx1_ASAP7_75t_L         g12689(.A(new_n12945), .Y(new_n12946));
  O2A1O1Ixp33_ASAP7_75t_L   g12690(.A1(new_n12624), .A2(new_n12621), .B(new_n12619), .C(new_n12946), .Y(new_n12947));
  INVx1_ASAP7_75t_L         g12691(.A(new_n12294), .Y(new_n12948));
  A2O1A1Ixp33_ASAP7_75t_L   g12692(.A1(new_n11941), .A2(new_n11938), .B(new_n11937), .C(new_n12298), .Y(new_n12949));
  A2O1A1Ixp33_ASAP7_75t_L   g12693(.A1(new_n12949), .A2(new_n12948), .B(new_n12621), .C(new_n12619), .Y(new_n12950));
  NOR2xp33_ASAP7_75t_L      g12694(.A(new_n12945), .B(new_n12950), .Y(new_n12951));
  NOR2xp33_ASAP7_75t_L      g12695(.A(new_n12951), .B(new_n12947), .Y(\f[64] ));
  NOR2xp33_ASAP7_75t_L      g12696(.A(new_n12888), .B(new_n12889), .Y(new_n12953));
  NOR3xp33_ASAP7_75t_L      g12697(.A(new_n12877), .B(new_n12872), .C(new_n12879), .Y(new_n12954));
  INVx1_ASAP7_75t_L         g12698(.A(new_n12954), .Y(new_n12955));
  A2O1A1Ixp33_ASAP7_75t_L   g12699(.A1(new_n12649), .A2(new_n12540), .B(new_n12953), .C(new_n12955), .Y(new_n12956));
  AOI22xp33_ASAP7_75t_L     g12700(.A1(new_n1113), .A2(\b[50] ), .B1(new_n1110), .B2(new_n8235), .Y(new_n12957));
  OAI221xp5_ASAP7_75t_L     g12701(.A1(new_n1298), .A2(new_n7907), .B1(new_n7333), .B2(new_n1195), .C(new_n12957), .Y(new_n12958));
  XNOR2x2_ASAP7_75t_L       g12702(.A(\a[17] ), .B(new_n12958), .Y(new_n12959));
  NAND3xp33_ASAP7_75t_L     g12703(.A(new_n12870), .B(new_n12867), .C(new_n12661), .Y(new_n12960));
  NAND2xp33_ASAP7_75t_L     g12704(.A(\b[45] ), .B(new_n1548), .Y(new_n12961));
  NAND2xp33_ASAP7_75t_L     g12705(.A(\b[46] ), .B(new_n1410), .Y(new_n12962));
  AOI22xp33_ASAP7_75t_L     g12706(.A1(new_n1406), .A2(\b[47] ), .B1(new_n1404), .B2(new_n7323), .Y(new_n12963));
  NAND4xp25_ASAP7_75t_L     g12707(.A(new_n12963), .B(\a[20] ), .C(new_n12961), .D(new_n12962), .Y(new_n12964));
  NAND2xp33_ASAP7_75t_L     g12708(.A(new_n12962), .B(new_n12963), .Y(new_n12965));
  A2O1A1Ixp33_ASAP7_75t_L   g12709(.A1(\b[45] ), .A2(new_n1548), .B(new_n12965), .C(new_n1401), .Y(new_n12966));
  NAND2xp33_ASAP7_75t_L     g12710(.A(new_n12964), .B(new_n12966), .Y(new_n12967));
  AOI22xp33_ASAP7_75t_L     g12711(.A1(new_n1766), .A2(\b[44] ), .B1(new_n1764), .B2(new_n7055), .Y(new_n12968));
  OAI221xp5_ASAP7_75t_L     g12712(.A1(new_n1758), .A2(new_n6195), .B1(new_n5680), .B2(new_n1911), .C(new_n12968), .Y(new_n12969));
  XNOR2x2_ASAP7_75t_L       g12713(.A(\a[23] ), .B(new_n12969), .Y(new_n12970));
  INVx1_ASAP7_75t_L         g12714(.A(new_n12970), .Y(new_n12971));
  NAND3xp33_ASAP7_75t_L     g12715(.A(new_n12839), .B(new_n12840), .C(new_n12847), .Y(new_n12972));
  A2O1A1Ixp33_ASAP7_75t_L   g12716(.A1(new_n12848), .A2(new_n12844), .B(new_n12849), .C(new_n12972), .Y(new_n12973));
  NOR3xp33_ASAP7_75t_L      g12717(.A(new_n12824), .B(new_n12820), .C(new_n12822), .Y(new_n12974));
  O2A1O1Ixp33_ASAP7_75t_L   g12718(.A1(new_n12829), .A2(new_n12830), .B(new_n12831), .C(new_n12974), .Y(new_n12975));
  AOI22xp33_ASAP7_75t_L     g12719(.A1(new_n3256), .A2(\b[35] ), .B1(new_n3254), .B2(new_n5649), .Y(new_n12976));
  OAI221xp5_ASAP7_75t_L     g12720(.A1(new_n3248), .A2(new_n3827), .B1(new_n3807), .B2(new_n3492), .C(new_n12976), .Y(new_n12977));
  XNOR2x2_ASAP7_75t_L       g12721(.A(\a[32] ), .B(new_n12977), .Y(new_n12978));
  INVx1_ASAP7_75t_L         g12722(.A(new_n12812), .Y(new_n12979));
  O2A1O1Ixp33_ASAP7_75t_L   g12723(.A1(new_n12665), .A2(new_n12486), .B(new_n12979), .C(new_n12813), .Y(new_n12980));
  NAND2xp33_ASAP7_75t_L     g12724(.A(new_n12759), .B(new_n12756), .Y(new_n12981));
  MAJIxp5_ASAP7_75t_L       g12725(.A(new_n12772), .B(new_n12762), .C(new_n12981), .Y(new_n12982));
  OAI22xp33_ASAP7_75t_L     g12726(.A1(new_n4860), .A2(new_n6311), .B1(new_n6312), .B2(new_n1995), .Y(new_n12983));
  AOI221xp5_ASAP7_75t_L     g12727(.A1(\b[21] ), .A2(new_n6308), .B1(\b[22] ), .B2(new_n5992), .C(new_n12983), .Y(new_n12984));
  XNOR2x2_ASAP7_75t_L       g12728(.A(new_n5996), .B(new_n12984), .Y(new_n12985));
  A2O1A1O1Ixp25_ASAP7_75t_L g12729(.A1(new_n12418), .A2(new_n12341), .B(new_n12753), .C(new_n12747), .D(new_n12758), .Y(new_n12986));
  NAND2xp33_ASAP7_75t_L     g12730(.A(new_n12722), .B(new_n12726), .Y(new_n12987));
  NOR2xp33_ASAP7_75t_L      g12731(.A(new_n12729), .B(new_n12987), .Y(new_n12988));
  A2O1A1O1Ixp25_ASAP7_75t_L g12732(.A1(new_n12409), .A2(new_n12739), .B(new_n12414), .C(new_n12735), .D(new_n12988), .Y(new_n12989));
  AOI22xp33_ASAP7_75t_L     g12733(.A1(new_n7659), .A2(\b[17] ), .B1(new_n7656), .B2(new_n1252), .Y(new_n12990));
  OAI221xp5_ASAP7_75t_L     g12734(.A1(new_n8326), .A2(new_n1051), .B1(new_n952), .B2(new_n7994), .C(new_n12990), .Y(new_n12991));
  XNOR2x2_ASAP7_75t_L       g12735(.A(new_n7653), .B(new_n12991), .Y(new_n12992));
  A2O1A1Ixp33_ASAP7_75t_L   g12736(.A1(new_n12395), .A2(new_n12394), .B(new_n12723), .C(new_n12720), .Y(new_n12993));
  NOR2xp33_ASAP7_75t_L      g12737(.A(new_n12703), .B(new_n12704), .Y(new_n12994));
  MAJIxp5_ASAP7_75t_L       g12738(.A(new_n12709), .B(new_n12994), .C(new_n12705), .Y(new_n12995));
  AOI22xp33_ASAP7_75t_L     g12739(.A1(new_n9623), .A2(\b[11] ), .B1(new_n9620), .B2(new_n702), .Y(new_n12996));
  OAI221xp5_ASAP7_75t_L     g12740(.A1(new_n10280), .A2(new_n631), .B1(new_n559), .B2(new_n12010), .C(new_n12996), .Y(new_n12997));
  XNOR2x2_ASAP7_75t_L       g12741(.A(\a[56] ), .B(new_n12997), .Y(new_n12998));
  INVx1_ASAP7_75t_L         g12742(.A(new_n12694), .Y(new_n12999));
  NOR2xp33_ASAP7_75t_L      g12743(.A(new_n276), .B(new_n12671), .Y(new_n13000));
  O2A1O1Ixp33_ASAP7_75t_L   g12744(.A1(new_n12353), .A2(new_n12355), .B(\b[2] ), .C(new_n13000), .Y(new_n13001));
  INVx1_ASAP7_75t_L         g12745(.A(new_n13001), .Y(new_n13002));
  INVx1_ASAP7_75t_L         g12746(.A(new_n12021), .Y(new_n13003));
  AOI22xp33_ASAP7_75t_L     g12747(.A1(new_n11656), .A2(\b[5] ), .B1(new_n11654), .B2(new_n360), .Y(new_n13004));
  OAI221xp5_ASAP7_75t_L     g12748(.A1(new_n12364), .A2(new_n323), .B1(new_n299), .B2(new_n13003), .C(new_n13004), .Y(new_n13005));
  XNOR2x2_ASAP7_75t_L       g12749(.A(new_n11651), .B(new_n13005), .Y(new_n13006));
  XNOR2x2_ASAP7_75t_L       g12750(.A(new_n13002), .B(new_n13006), .Y(new_n13007));
  MAJIxp5_ASAP7_75t_L       g12751(.A(new_n12682), .B(new_n12680), .C(new_n12678), .Y(new_n13008));
  INVx1_ASAP7_75t_L         g12752(.A(new_n13008), .Y(new_n13009));
  NAND2xp33_ASAP7_75t_L     g12753(.A(new_n13007), .B(new_n13009), .Y(new_n13010));
  INVx1_ASAP7_75t_L         g12754(.A(new_n13000), .Y(new_n13011));
  O2A1O1Ixp33_ASAP7_75t_L   g12755(.A1(new_n278), .A2(new_n12356), .B(new_n13011), .C(new_n13006), .Y(new_n13012));
  AND2x2_ASAP7_75t_L        g12756(.A(new_n13001), .B(new_n13006), .Y(new_n13013));
  OAI21xp33_ASAP7_75t_L     g12757(.A1(new_n13012), .A2(new_n13013), .B(new_n13008), .Y(new_n13014));
  NAND2xp33_ASAP7_75t_L     g12758(.A(new_n13014), .B(new_n13010), .Y(new_n13015));
  AOI22xp33_ASAP7_75t_L     g12759(.A1(new_n10594), .A2(\b[8] ), .B1(new_n10591), .B2(new_n510), .Y(new_n13016));
  OAI221xp5_ASAP7_75t_L     g12760(.A1(new_n11335), .A2(new_n421), .B1(new_n382), .B2(new_n11330), .C(new_n13016), .Y(new_n13017));
  XNOR2x2_ASAP7_75t_L       g12761(.A(\a[59] ), .B(new_n13017), .Y(new_n13018));
  NAND2xp33_ASAP7_75t_L     g12762(.A(new_n13018), .B(new_n13015), .Y(new_n13019));
  INVx1_ASAP7_75t_L         g12763(.A(new_n13018), .Y(new_n13020));
  NAND3xp33_ASAP7_75t_L     g12764(.A(new_n13020), .B(new_n13014), .C(new_n13010), .Y(new_n13021));
  NAND4xp25_ASAP7_75t_L     g12765(.A(new_n12695), .B(new_n13019), .C(new_n13021), .D(new_n12999), .Y(new_n13022));
  A2O1A1Ixp33_ASAP7_75t_L   g12766(.A1(new_n12379), .A2(new_n12377), .B(new_n12690), .C(new_n12999), .Y(new_n13023));
  AOI21xp33_ASAP7_75t_L     g12767(.A1(new_n13014), .A2(new_n13010), .B(new_n13020), .Y(new_n13024));
  NOR2xp33_ASAP7_75t_L      g12768(.A(new_n13018), .B(new_n13015), .Y(new_n13025));
  OAI21xp33_ASAP7_75t_L     g12769(.A1(new_n13024), .A2(new_n13025), .B(new_n13023), .Y(new_n13026));
  NAND3xp33_ASAP7_75t_L     g12770(.A(new_n13022), .B(new_n13026), .C(new_n12998), .Y(new_n13027));
  AO21x2_ASAP7_75t_L        g12771(.A1(new_n13026), .A2(new_n13022), .B(new_n12998), .Y(new_n13028));
  NAND2xp33_ASAP7_75t_L     g12772(.A(new_n13027), .B(new_n13028), .Y(new_n13029));
  NOR2xp33_ASAP7_75t_L      g12773(.A(new_n12995), .B(new_n13029), .Y(new_n13030));
  AOI221xp5_ASAP7_75t_L     g12774(.A1(new_n13028), .A2(new_n13027), .B1(new_n12994), .B2(new_n12705), .C(new_n12712), .Y(new_n13031));
  AOI22xp33_ASAP7_75t_L     g12775(.A1(new_n8645), .A2(\b[14] ), .B1(new_n8642), .B2(new_n879), .Y(new_n13032));
  OAI221xp5_ASAP7_75t_L     g12776(.A1(new_n9322), .A2(new_n793), .B1(new_n763), .B2(new_n8965), .C(new_n13032), .Y(new_n13033));
  XNOR2x2_ASAP7_75t_L       g12777(.A(\a[53] ), .B(new_n13033), .Y(new_n13034));
  INVx1_ASAP7_75t_L         g12778(.A(new_n13034), .Y(new_n13035));
  NOR3xp33_ASAP7_75t_L      g12779(.A(new_n13030), .B(new_n13031), .C(new_n13035), .Y(new_n13036));
  INVx1_ASAP7_75t_L         g12780(.A(new_n13027), .Y(new_n13037));
  AOI21xp33_ASAP7_75t_L     g12781(.A1(new_n13022), .A2(new_n13026), .B(new_n12998), .Y(new_n13038));
  OR3x1_ASAP7_75t_L         g12782(.A(new_n13037), .B(new_n12995), .C(new_n13038), .Y(new_n13039));
  NAND2xp33_ASAP7_75t_L     g12783(.A(new_n12995), .B(new_n13029), .Y(new_n13040));
  AOI21xp33_ASAP7_75t_L     g12784(.A1(new_n13039), .A2(new_n13040), .B(new_n13034), .Y(new_n13041));
  OAI21xp33_ASAP7_75t_L     g12785(.A1(new_n13036), .A2(new_n13041), .B(new_n12993), .Y(new_n13042));
  A2O1A1O1Ixp25_ASAP7_75t_L g12786(.A1(new_n12390), .A2(new_n12343), .B(new_n12398), .C(new_n12716), .D(new_n12724), .Y(new_n13043));
  NAND3xp33_ASAP7_75t_L     g12787(.A(new_n13039), .B(new_n13040), .C(new_n13034), .Y(new_n13044));
  OAI21xp33_ASAP7_75t_L     g12788(.A1(new_n13031), .A2(new_n13030), .B(new_n13035), .Y(new_n13045));
  NAND3xp33_ASAP7_75t_L     g12789(.A(new_n13044), .B(new_n13043), .C(new_n13045), .Y(new_n13046));
  NAND3xp33_ASAP7_75t_L     g12790(.A(new_n13042), .B(new_n13046), .C(new_n12992), .Y(new_n13047));
  AO21x2_ASAP7_75t_L        g12791(.A1(new_n13046), .A2(new_n13042), .B(new_n12992), .Y(new_n13048));
  NAND2xp33_ASAP7_75t_L     g12792(.A(new_n13047), .B(new_n13048), .Y(new_n13049));
  NAND2xp33_ASAP7_75t_L     g12793(.A(new_n12989), .B(new_n13049), .Y(new_n13050));
  OAI211xp5_ASAP7_75t_L     g12794(.A1(new_n12988), .A2(new_n12743), .B(new_n13047), .C(new_n13048), .Y(new_n13051));
  AOI22xp33_ASAP7_75t_L     g12795(.A1(new_n6822), .A2(\b[20] ), .B1(new_n6819), .B2(new_n1600), .Y(new_n13052));
  OAI221xp5_ASAP7_75t_L     g12796(.A1(new_n7392), .A2(new_n1493), .B1(new_n1356), .B2(new_n7115), .C(new_n13052), .Y(new_n13053));
  XNOR2x2_ASAP7_75t_L       g12797(.A(\a[47] ), .B(new_n13053), .Y(new_n13054));
  NAND3xp33_ASAP7_75t_L     g12798(.A(new_n13050), .B(new_n13051), .C(new_n13054), .Y(new_n13055));
  AOI211xp5_ASAP7_75t_L     g12799(.A1(new_n13047), .A2(new_n13048), .B(new_n12988), .C(new_n12743), .Y(new_n13056));
  O2A1O1Ixp33_ASAP7_75t_L   g12800(.A1(new_n12987), .A2(new_n12729), .B(new_n12749), .C(new_n13049), .Y(new_n13057));
  INVx1_ASAP7_75t_L         g12801(.A(new_n13054), .Y(new_n13058));
  OAI21xp33_ASAP7_75t_L     g12802(.A1(new_n13056), .A2(new_n13057), .B(new_n13058), .Y(new_n13059));
  AOI21xp33_ASAP7_75t_L     g12803(.A1(new_n13059), .A2(new_n13055), .B(new_n12986), .Y(new_n13060));
  A2O1A1Ixp33_ASAP7_75t_L   g12804(.A1(new_n12423), .A2(new_n12422), .B(new_n12757), .C(new_n12751), .Y(new_n13061));
  NOR3xp33_ASAP7_75t_L      g12805(.A(new_n13057), .B(new_n13058), .C(new_n13056), .Y(new_n13062));
  AOI21xp33_ASAP7_75t_L     g12806(.A1(new_n13050), .A2(new_n13051), .B(new_n13054), .Y(new_n13063));
  NOR3xp33_ASAP7_75t_L      g12807(.A(new_n13062), .B(new_n13063), .C(new_n13061), .Y(new_n13064));
  NOR3xp33_ASAP7_75t_L      g12808(.A(new_n13064), .B(new_n13060), .C(new_n12985), .Y(new_n13065));
  INVx1_ASAP7_75t_L         g12809(.A(new_n12985), .Y(new_n13066));
  OAI21xp33_ASAP7_75t_L     g12810(.A1(new_n13063), .A2(new_n13062), .B(new_n13061), .Y(new_n13067));
  NAND3xp33_ASAP7_75t_L     g12811(.A(new_n13059), .B(new_n13055), .C(new_n12986), .Y(new_n13068));
  AOI21xp33_ASAP7_75t_L     g12812(.A1(new_n13067), .A2(new_n13068), .B(new_n13066), .Y(new_n13069));
  NOR2xp33_ASAP7_75t_L      g12813(.A(new_n13069), .B(new_n13065), .Y(new_n13070));
  NOR2xp33_ASAP7_75t_L      g12814(.A(new_n12982), .B(new_n13070), .Y(new_n13071));
  NAND3xp33_ASAP7_75t_L     g12815(.A(new_n13067), .B(new_n13068), .C(new_n13066), .Y(new_n13072));
  OAI21xp33_ASAP7_75t_L     g12816(.A1(new_n13060), .A2(new_n13064), .B(new_n12985), .Y(new_n13073));
  NAND2xp33_ASAP7_75t_L     g12817(.A(new_n13072), .B(new_n13073), .Y(new_n13074));
  O2A1O1Ixp33_ASAP7_75t_L   g12818(.A1(new_n12981), .A2(new_n12762), .B(new_n12779), .C(new_n13074), .Y(new_n13075));
  AOI22xp33_ASAP7_75t_L     g12819(.A1(new_n5249), .A2(\b[26] ), .B1(new_n5247), .B2(new_n2888), .Y(new_n13076));
  OAI221xp5_ASAP7_75t_L     g12820(.A1(new_n5241), .A2(new_n2180), .B1(new_n2019), .B2(new_n5521), .C(new_n13076), .Y(new_n13077));
  XNOR2x2_ASAP7_75t_L       g12821(.A(\a[41] ), .B(new_n13077), .Y(new_n13078));
  INVx1_ASAP7_75t_L         g12822(.A(new_n13078), .Y(new_n13079));
  NOR3xp33_ASAP7_75t_L      g12823(.A(new_n13075), .B(new_n13071), .C(new_n13079), .Y(new_n13080));
  INVx1_ASAP7_75t_L         g12824(.A(new_n12981), .Y(new_n13081));
  NAND2xp33_ASAP7_75t_L     g12825(.A(new_n12766), .B(new_n13081), .Y(new_n13082));
  NAND3xp33_ASAP7_75t_L     g12826(.A(new_n13074), .B(new_n12779), .C(new_n13082), .Y(new_n13083));
  A2O1A1Ixp33_ASAP7_75t_L   g12827(.A1(new_n12766), .A2(new_n13081), .B(new_n12773), .C(new_n13070), .Y(new_n13084));
  AOI21xp33_ASAP7_75t_L     g12828(.A1(new_n13084), .A2(new_n13083), .B(new_n13078), .Y(new_n13085));
  NOR2xp33_ASAP7_75t_L      g12829(.A(new_n13080), .B(new_n13085), .Y(new_n13086));
  NOR3xp33_ASAP7_75t_L      g12830(.A(new_n12770), .B(new_n12773), .C(new_n12780), .Y(new_n13087));
  O2A1O1Ixp33_ASAP7_75t_L   g12831(.A1(new_n12777), .A2(new_n12781), .B(new_n12797), .C(new_n13087), .Y(new_n13088));
  NAND2xp33_ASAP7_75t_L     g12832(.A(new_n13088), .B(new_n13086), .Y(new_n13089));
  NAND3xp33_ASAP7_75t_L     g12833(.A(new_n13084), .B(new_n13083), .C(new_n13078), .Y(new_n13090));
  OAI21xp33_ASAP7_75t_L     g12834(.A1(new_n13071), .A2(new_n13075), .B(new_n13079), .Y(new_n13091));
  NAND2xp33_ASAP7_75t_L     g12835(.A(new_n13091), .B(new_n13090), .Y(new_n13092));
  A2O1A1Ixp33_ASAP7_75t_L   g12836(.A1(new_n12790), .A2(new_n12797), .B(new_n13087), .C(new_n13092), .Y(new_n13093));
  AOI22xp33_ASAP7_75t_L     g12837(.A1(new_n4544), .A2(\b[29] ), .B1(new_n4542), .B2(new_n5472), .Y(new_n13094));
  OAI221xp5_ASAP7_75t_L     g12838(.A1(new_n4536), .A2(new_n2852), .B1(new_n2650), .B2(new_n4781), .C(new_n13094), .Y(new_n13095));
  XNOR2x2_ASAP7_75t_L       g12839(.A(\a[38] ), .B(new_n13095), .Y(new_n13096));
  NAND3xp33_ASAP7_75t_L     g12840(.A(new_n13093), .B(new_n13089), .C(new_n13096), .Y(new_n13097));
  NOR3xp33_ASAP7_75t_L      g12841(.A(new_n13092), .B(new_n12799), .C(new_n13087), .Y(new_n13098));
  NOR2xp33_ASAP7_75t_L      g12842(.A(new_n13088), .B(new_n13086), .Y(new_n13099));
  INVx1_ASAP7_75t_L         g12843(.A(new_n13096), .Y(new_n13100));
  OAI21xp33_ASAP7_75t_L     g12844(.A1(new_n13099), .A2(new_n13098), .B(new_n13100), .Y(new_n13101));
  NAND2xp33_ASAP7_75t_L     g12845(.A(new_n13097), .B(new_n13101), .Y(new_n13102));
  NOR2xp33_ASAP7_75t_L      g12846(.A(new_n12798), .B(new_n12799), .Y(new_n13103));
  NAND2xp33_ASAP7_75t_L     g12847(.A(new_n12800), .B(new_n13103), .Y(new_n13104));
  A2O1A1Ixp33_ASAP7_75t_L   g12848(.A1(new_n12801), .A2(new_n12795), .B(new_n12807), .C(new_n13104), .Y(new_n13105));
  NOR2xp33_ASAP7_75t_L      g12849(.A(new_n13105), .B(new_n13102), .Y(new_n13106));
  NAND2xp33_ASAP7_75t_L     g12850(.A(new_n12791), .B(new_n12786), .Y(new_n13107));
  A2O1A1Ixp33_ASAP7_75t_L   g12851(.A1(new_n12456), .A2(new_n12459), .B(new_n12803), .C(new_n12802), .Y(new_n13108));
  NOR3xp33_ASAP7_75t_L      g12852(.A(new_n13098), .B(new_n13099), .C(new_n13100), .Y(new_n13109));
  AOI21xp33_ASAP7_75t_L     g12853(.A1(new_n13093), .A2(new_n13089), .B(new_n13096), .Y(new_n13110));
  NOR2xp33_ASAP7_75t_L      g12854(.A(new_n13110), .B(new_n13109), .Y(new_n13111));
  O2A1O1Ixp33_ASAP7_75t_L   g12855(.A1(new_n13107), .A2(new_n12794), .B(new_n13108), .C(new_n13111), .Y(new_n13112));
  AOI22xp33_ASAP7_75t_L     g12856(.A1(new_n3884), .A2(\b[32] ), .B1(new_n3881), .B2(new_n3450), .Y(new_n13113));
  OAI221xp5_ASAP7_75t_L     g12857(.A1(new_n4312), .A2(new_n3419), .B1(new_n3212), .B2(new_n4986), .C(new_n13113), .Y(new_n13114));
  XNOR2x2_ASAP7_75t_L       g12858(.A(\a[35] ), .B(new_n13114), .Y(new_n13115));
  OAI21xp33_ASAP7_75t_L     g12859(.A1(new_n13106), .A2(new_n13112), .B(new_n13115), .Y(new_n13116));
  NAND3xp33_ASAP7_75t_L     g12860(.A(new_n13111), .B(new_n13108), .C(new_n13104), .Y(new_n13117));
  A2O1A1Ixp33_ASAP7_75t_L   g12861(.A1(new_n12800), .A2(new_n13103), .B(new_n12808), .C(new_n13102), .Y(new_n13118));
  INVx1_ASAP7_75t_L         g12862(.A(new_n13115), .Y(new_n13119));
  NAND3xp33_ASAP7_75t_L     g12863(.A(new_n13117), .B(new_n13118), .C(new_n13119), .Y(new_n13120));
  NAND3xp33_ASAP7_75t_L     g12864(.A(new_n12980), .B(new_n13116), .C(new_n13120), .Y(new_n13121));
  OR3x1_ASAP7_75t_L         g12865(.A(new_n12806), .B(new_n12808), .C(new_n12811), .Y(new_n13122));
  A2O1A1Ixp33_ASAP7_75t_L   g12866(.A1(new_n12476), .A2(new_n12473), .B(new_n12812), .C(new_n13122), .Y(new_n13123));
  NAND2xp33_ASAP7_75t_L     g12867(.A(new_n13120), .B(new_n13116), .Y(new_n13124));
  NAND2xp33_ASAP7_75t_L     g12868(.A(new_n13123), .B(new_n13124), .Y(new_n13125));
  AOI21xp33_ASAP7_75t_L     g12869(.A1(new_n13125), .A2(new_n13121), .B(new_n12978), .Y(new_n13126));
  INVx1_ASAP7_75t_L         g12870(.A(new_n12978), .Y(new_n13127));
  NOR2xp33_ASAP7_75t_L      g12871(.A(new_n13123), .B(new_n13124), .Y(new_n13128));
  AOI21xp33_ASAP7_75t_L     g12872(.A1(new_n13120), .A2(new_n13116), .B(new_n12980), .Y(new_n13129));
  NOR3xp33_ASAP7_75t_L      g12873(.A(new_n13128), .B(new_n13129), .C(new_n13127), .Y(new_n13130));
  OAI21xp33_ASAP7_75t_L     g12874(.A1(new_n13126), .A2(new_n13130), .B(new_n12975), .Y(new_n13131));
  AOI22xp33_ASAP7_75t_L     g12875(.A1(new_n12827), .A2(new_n12664), .B1(new_n12826), .B2(new_n12821), .Y(new_n13132));
  OAI21xp33_ASAP7_75t_L     g12876(.A1(new_n13129), .A2(new_n13128), .B(new_n13127), .Y(new_n13133));
  NAND3xp33_ASAP7_75t_L     g12877(.A(new_n13125), .B(new_n13121), .C(new_n12978), .Y(new_n13134));
  OAI211xp5_ASAP7_75t_L     g12878(.A1(new_n12974), .A2(new_n13132), .B(new_n13133), .C(new_n13134), .Y(new_n13135));
  AOI22xp33_ASAP7_75t_L     g12879(.A1(new_n2702), .A2(\b[38] ), .B1(new_n2700), .B2(new_n4923), .Y(new_n13136));
  OAI221xp5_ASAP7_75t_L     g12880(.A1(new_n2694), .A2(new_n4701), .B1(new_n4465), .B2(new_n2932), .C(new_n13136), .Y(new_n13137));
  XNOR2x2_ASAP7_75t_L       g12881(.A(\a[29] ), .B(new_n13137), .Y(new_n13138));
  NAND3xp33_ASAP7_75t_L     g12882(.A(new_n13135), .B(new_n13131), .C(new_n13138), .Y(new_n13139));
  AO21x2_ASAP7_75t_L        g12883(.A1(new_n13131), .A2(new_n13135), .B(new_n13138), .Y(new_n13140));
  NOR3xp33_ASAP7_75t_L      g12884(.A(new_n12830), .B(new_n12831), .C(new_n12829), .Y(new_n13141));
  NOR3xp33_ASAP7_75t_L      g12885(.A(new_n13141), .B(new_n13132), .C(new_n12835), .Y(new_n13142));
  O2A1O1Ixp33_ASAP7_75t_L   g12886(.A1(new_n12837), .A2(new_n12836), .B(new_n12838), .C(new_n13142), .Y(new_n13143));
  AND3x1_ASAP7_75t_L        g12887(.A(new_n13143), .B(new_n13140), .C(new_n13139), .Y(new_n13144));
  AOI21xp33_ASAP7_75t_L     g12888(.A1(new_n13140), .A2(new_n13139), .B(new_n13143), .Y(new_n13145));
  AOI22xp33_ASAP7_75t_L     g12889(.A1(new_n2228), .A2(\b[41] ), .B1(new_n2226), .B2(new_n5669), .Y(new_n13146));
  OAI221xp5_ASAP7_75t_L     g12890(.A1(new_n2220), .A2(new_n5186), .B1(new_n5166), .B2(new_n2387), .C(new_n13146), .Y(new_n13147));
  XNOR2x2_ASAP7_75t_L       g12891(.A(\a[26] ), .B(new_n13147), .Y(new_n13148));
  OAI21xp33_ASAP7_75t_L     g12892(.A1(new_n13145), .A2(new_n13144), .B(new_n13148), .Y(new_n13149));
  NAND3xp33_ASAP7_75t_L     g12893(.A(new_n13143), .B(new_n13140), .C(new_n13139), .Y(new_n13150));
  AO21x2_ASAP7_75t_L        g12894(.A1(new_n13139), .A2(new_n13140), .B(new_n13143), .Y(new_n13151));
  INVx1_ASAP7_75t_L         g12895(.A(new_n13148), .Y(new_n13152));
  NAND3xp33_ASAP7_75t_L     g12896(.A(new_n13151), .B(new_n13150), .C(new_n13152), .Y(new_n13153));
  NAND2xp33_ASAP7_75t_L     g12897(.A(new_n13153), .B(new_n13149), .Y(new_n13154));
  NOR2xp33_ASAP7_75t_L      g12898(.A(new_n12973), .B(new_n13154), .Y(new_n13155));
  NAND2xp33_ASAP7_75t_L     g12899(.A(new_n12840), .B(new_n12839), .Y(new_n13156));
  A2O1A1Ixp33_ASAP7_75t_L   g12900(.A1(new_n12507), .A2(new_n12511), .B(new_n12513), .C(new_n12852), .Y(new_n13157));
  AOI21xp33_ASAP7_75t_L     g12901(.A1(new_n13151), .A2(new_n13150), .B(new_n13152), .Y(new_n13158));
  NOR3xp33_ASAP7_75t_L      g12902(.A(new_n13144), .B(new_n13145), .C(new_n13148), .Y(new_n13159));
  NOR2xp33_ASAP7_75t_L      g12903(.A(new_n13158), .B(new_n13159), .Y(new_n13160));
  O2A1O1Ixp33_ASAP7_75t_L   g12904(.A1(new_n13156), .A2(new_n12843), .B(new_n13157), .C(new_n13160), .Y(new_n13161));
  OAI21xp33_ASAP7_75t_L     g12905(.A1(new_n13155), .A2(new_n13161), .B(new_n12971), .Y(new_n13162));
  NAND3xp33_ASAP7_75t_L     g12906(.A(new_n13160), .B(new_n13157), .C(new_n12972), .Y(new_n13163));
  NOR2xp33_ASAP7_75t_L      g12907(.A(new_n12843), .B(new_n13156), .Y(new_n13164));
  A2O1A1Ixp33_ASAP7_75t_L   g12908(.A1(new_n12850), .A2(new_n12852), .B(new_n13164), .C(new_n13154), .Y(new_n13165));
  NAND3xp33_ASAP7_75t_L     g12909(.A(new_n13163), .B(new_n13165), .C(new_n12970), .Y(new_n13166));
  NAND2xp33_ASAP7_75t_L     g12910(.A(new_n13166), .B(new_n13162), .Y(new_n13167));
  O2A1O1Ixp33_ASAP7_75t_L   g12911(.A1(new_n12869), .A2(new_n12862), .B(new_n12858), .C(new_n13167), .Y(new_n13168));
  A2O1A1Ixp33_ASAP7_75t_L   g12912(.A1(new_n12527), .A2(new_n12663), .B(new_n12862), .C(new_n12858), .Y(new_n13169));
  AOI21xp33_ASAP7_75t_L     g12913(.A1(new_n13163), .A2(new_n13165), .B(new_n12970), .Y(new_n13170));
  NOR3xp33_ASAP7_75t_L      g12914(.A(new_n13161), .B(new_n13155), .C(new_n12971), .Y(new_n13171));
  NOR2xp33_ASAP7_75t_L      g12915(.A(new_n13170), .B(new_n13171), .Y(new_n13172));
  NOR2xp33_ASAP7_75t_L      g12916(.A(new_n13169), .B(new_n13172), .Y(new_n13173));
  OAI21xp33_ASAP7_75t_L     g12917(.A1(new_n13173), .A2(new_n13168), .B(new_n12967), .Y(new_n13174));
  INVx1_ASAP7_75t_L         g12918(.A(new_n12967), .Y(new_n13175));
  INVx1_ASAP7_75t_L         g12919(.A(new_n12858), .Y(new_n13176));
  A2O1A1Ixp33_ASAP7_75t_L   g12920(.A1(new_n12861), .A2(new_n12864), .B(new_n13176), .C(new_n13172), .Y(new_n13177));
  O2A1O1Ixp33_ASAP7_75t_L   g12921(.A1(new_n12662), .A2(new_n12522), .B(new_n12861), .C(new_n13176), .Y(new_n13178));
  NAND2xp33_ASAP7_75t_L     g12922(.A(new_n13178), .B(new_n13167), .Y(new_n13179));
  NAND3xp33_ASAP7_75t_L     g12923(.A(new_n13177), .B(new_n13175), .C(new_n13179), .Y(new_n13180));
  AOI22xp33_ASAP7_75t_L     g12924(.A1(new_n13174), .A2(new_n13180), .B1(new_n12960), .B2(new_n12880), .Y(new_n13181));
  A2O1A1Ixp33_ASAP7_75t_L   g12925(.A1(new_n12866), .A2(new_n12871), .B(new_n12657), .C(new_n12960), .Y(new_n13182));
  NAND2xp33_ASAP7_75t_L     g12926(.A(new_n13180), .B(new_n13174), .Y(new_n13183));
  NOR2xp33_ASAP7_75t_L      g12927(.A(new_n13182), .B(new_n13183), .Y(new_n13184));
  OAI21xp33_ASAP7_75t_L     g12928(.A1(new_n13181), .A2(new_n13184), .B(new_n12959), .Y(new_n13185));
  INVx1_ASAP7_75t_L         g12929(.A(new_n12959), .Y(new_n13186));
  NAND2xp33_ASAP7_75t_L     g12930(.A(new_n13182), .B(new_n13183), .Y(new_n13187));
  NAND4xp25_ASAP7_75t_L     g12931(.A(new_n12880), .B(new_n13180), .C(new_n13174), .D(new_n12960), .Y(new_n13188));
  NAND3xp33_ASAP7_75t_L     g12932(.A(new_n13187), .B(new_n13186), .C(new_n13188), .Y(new_n13189));
  NAND3xp33_ASAP7_75t_L     g12933(.A(new_n12956), .B(new_n13185), .C(new_n13189), .Y(new_n13190));
  O2A1O1Ixp33_ASAP7_75t_L   g12934(.A1(new_n12888), .A2(new_n12889), .B(new_n12887), .C(new_n12954), .Y(new_n13191));
  NAND2xp33_ASAP7_75t_L     g12935(.A(new_n13189), .B(new_n13185), .Y(new_n13192));
  NAND2xp33_ASAP7_75t_L     g12936(.A(new_n13191), .B(new_n13192), .Y(new_n13193));
  AOI22xp33_ASAP7_75t_L     g12937(.A1(new_n826), .A2(\b[53] ), .B1(new_n823), .B2(new_n8889), .Y(new_n13194));
  OAI221xp5_ASAP7_75t_L     g12938(.A1(new_n994), .A2(new_n8569), .B1(new_n8249), .B2(new_n909), .C(new_n13194), .Y(new_n13195));
  XNOR2x2_ASAP7_75t_L       g12939(.A(\a[14] ), .B(new_n13195), .Y(new_n13196));
  NAND3xp33_ASAP7_75t_L     g12940(.A(new_n13193), .B(new_n13190), .C(new_n13196), .Y(new_n13197));
  NOR2xp33_ASAP7_75t_L      g12941(.A(new_n13191), .B(new_n13192), .Y(new_n13198));
  AOI21xp33_ASAP7_75t_L     g12942(.A1(new_n13189), .A2(new_n13185), .B(new_n12956), .Y(new_n13199));
  INVx1_ASAP7_75t_L         g12943(.A(new_n13196), .Y(new_n13200));
  OAI21xp33_ASAP7_75t_L     g12944(.A1(new_n13199), .A2(new_n13198), .B(new_n13200), .Y(new_n13201));
  A2O1A1O1Ixp25_ASAP7_75t_L g12945(.A1(new_n12546), .A2(new_n12549), .B(new_n12896), .C(new_n12902), .D(new_n12885), .Y(new_n13202));
  AND3x1_ASAP7_75t_L        g12946(.A(new_n13201), .B(new_n13202), .C(new_n13197), .Y(new_n13203));
  AOI21xp33_ASAP7_75t_L     g12947(.A1(new_n13201), .A2(new_n13197), .B(new_n13202), .Y(new_n13204));
  AOI22xp33_ASAP7_75t_L     g12948(.A1(new_n600), .A2(\b[56] ), .B1(new_n597), .B2(new_n10185), .Y(new_n13205));
  OAI221xp5_ASAP7_75t_L     g12949(.A1(new_n721), .A2(new_n9534), .B1(new_n9199), .B2(new_n1620), .C(new_n13205), .Y(new_n13206));
  XNOR2x2_ASAP7_75t_L       g12950(.A(\a[11] ), .B(new_n13206), .Y(new_n13207));
  OAI21xp33_ASAP7_75t_L     g12951(.A1(new_n13204), .A2(new_n13203), .B(new_n13207), .Y(new_n13208));
  NAND3xp33_ASAP7_75t_L     g12952(.A(new_n13201), .B(new_n13197), .C(new_n13202), .Y(new_n13209));
  AO21x2_ASAP7_75t_L        g12953(.A1(new_n13197), .A2(new_n13201), .B(new_n13202), .Y(new_n13210));
  INVx1_ASAP7_75t_L         g12954(.A(new_n13207), .Y(new_n13211));
  NAND3xp33_ASAP7_75t_L     g12955(.A(new_n13210), .B(new_n13209), .C(new_n13211), .Y(new_n13212));
  NAND2xp33_ASAP7_75t_L     g12956(.A(\b[59] ), .B(new_n451), .Y(new_n13213));
  OAI221xp5_ASAP7_75t_L     g12957(.A1(new_n10848), .A2(new_n529), .B1(new_n482), .B2(new_n10888), .C(new_n13213), .Y(new_n13214));
  AOI21xp33_ASAP7_75t_L     g12958(.A1(new_n480), .A2(\b[57] ), .B(new_n13214), .Y(new_n13215));
  NAND2xp33_ASAP7_75t_L     g12959(.A(\a[8] ), .B(new_n13215), .Y(new_n13216));
  A2O1A1Ixp33_ASAP7_75t_L   g12960(.A1(\b[57] ), .A2(new_n480), .B(new_n13214), .C(new_n445), .Y(new_n13217));
  NAND2xp33_ASAP7_75t_L     g12961(.A(new_n13217), .B(new_n13216), .Y(new_n13218));
  INVx1_ASAP7_75t_L         g12962(.A(new_n13218), .Y(new_n13219));
  NAND3xp33_ASAP7_75t_L     g12963(.A(new_n13208), .B(new_n13212), .C(new_n13219), .Y(new_n13220));
  AOI21xp33_ASAP7_75t_L     g12964(.A1(new_n13210), .A2(new_n13209), .B(new_n13211), .Y(new_n13221));
  NOR3xp33_ASAP7_75t_L      g12965(.A(new_n13203), .B(new_n13204), .C(new_n13207), .Y(new_n13222));
  OAI21xp33_ASAP7_75t_L     g12966(.A1(new_n13221), .A2(new_n13222), .B(new_n13218), .Y(new_n13223));
  NOR3xp33_ASAP7_75t_L      g12967(.A(new_n12900), .B(new_n12903), .C(new_n12638), .Y(new_n13224));
  O2A1O1Ixp33_ASAP7_75t_L   g12968(.A1(new_n12906), .A2(new_n12567), .B(new_n12904), .C(new_n13224), .Y(new_n13225));
  NAND3xp33_ASAP7_75t_L     g12969(.A(new_n13223), .B(new_n13220), .C(new_n13225), .Y(new_n13226));
  NOR3xp33_ASAP7_75t_L      g12970(.A(new_n13222), .B(new_n13221), .C(new_n13218), .Y(new_n13227));
  AOI21xp33_ASAP7_75t_L     g12971(.A1(new_n13208), .A2(new_n13212), .B(new_n13219), .Y(new_n13228));
  INVx1_ASAP7_75t_L         g12972(.A(new_n13225), .Y(new_n13229));
  OAI21xp33_ASAP7_75t_L     g12973(.A1(new_n13228), .A2(new_n13227), .B(new_n13229), .Y(new_n13230));
  NAND2xp33_ASAP7_75t_L     g12974(.A(\b[60] ), .B(new_n366), .Y(new_n13231));
  NAND2xp33_ASAP7_75t_L     g12975(.A(\b[61] ), .B(new_n334), .Y(new_n13232));
  AOI22xp33_ASAP7_75t_L     g12976(.A1(new_n345), .A2(\b[62] ), .B1(new_n342), .B2(new_n12280), .Y(new_n13233));
  AND4x1_ASAP7_75t_L        g12977(.A(new_n13233), .B(new_n13232), .C(new_n13231), .D(\a[5] ), .Y(new_n13234));
  AOI31xp33_ASAP7_75t_L     g12978(.A1(new_n13233), .A2(new_n13232), .A3(new_n13231), .B(\a[5] ), .Y(new_n13235));
  NOR2xp33_ASAP7_75t_L      g12979(.A(new_n13235), .B(new_n13234), .Y(new_n13236));
  NAND3xp33_ASAP7_75t_L     g12980(.A(new_n13230), .B(new_n13236), .C(new_n13226), .Y(new_n13237));
  NOR3xp33_ASAP7_75t_L      g12981(.A(new_n13227), .B(new_n13228), .C(new_n13229), .Y(new_n13238));
  AOI21xp33_ASAP7_75t_L     g12982(.A1(new_n13223), .A2(new_n13220), .B(new_n13225), .Y(new_n13239));
  INVx1_ASAP7_75t_L         g12983(.A(new_n13236), .Y(new_n13240));
  OAI21xp33_ASAP7_75t_L     g12984(.A1(new_n13239), .A2(new_n13238), .B(new_n13240), .Y(new_n13241));
  NOR2xp33_ASAP7_75t_L      g12985(.A(new_n12915), .B(new_n12914), .Y(new_n13242));
  O2A1O1Ixp33_ASAP7_75t_L   g12986(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n12599), .Y(new_n13243));
  NOR2xp33_ASAP7_75t_L      g12987(.A(new_n12599), .B(new_n277), .Y(new_n13244));
  A2O1A1Ixp33_ASAP7_75t_L   g12988(.A1(new_n13243), .A2(new_n269), .B(new_n13244), .C(\a[2] ), .Y(new_n13245));
  A2O1A1Ixp33_ASAP7_75t_L   g12989(.A1(new_n269), .A2(new_n13243), .B(\a[2] ), .C(new_n13245), .Y(new_n13246));
  INVx1_ASAP7_75t_L         g12990(.A(new_n13246), .Y(new_n13247));
  A2O1A1Ixp33_ASAP7_75t_L   g12991(.A1(new_n12916), .A2(new_n13242), .B(new_n12924), .C(new_n13247), .Y(new_n13248));
  INVx1_ASAP7_75t_L         g12992(.A(new_n13242), .Y(new_n13249));
  OAI211xp5_ASAP7_75t_L     g12993(.A1(new_n12912), .A2(new_n13249), .B(new_n12931), .C(new_n13246), .Y(new_n13250));
  AOI22xp33_ASAP7_75t_L     g12994(.A1(new_n13237), .A2(new_n13241), .B1(new_n13248), .B2(new_n13250), .Y(new_n13251));
  AND4x1_ASAP7_75t_L        g12995(.A(new_n13250), .B(new_n13248), .C(new_n13241), .D(new_n13237), .Y(new_n13252));
  OAI21xp33_ASAP7_75t_L     g12996(.A1(new_n12631), .A2(new_n12933), .B(new_n12936), .Y(new_n13253));
  NOR3xp33_ASAP7_75t_L      g12997(.A(new_n13252), .B(new_n13253), .C(new_n13251), .Y(new_n13254));
  NAND2xp33_ASAP7_75t_L     g12998(.A(new_n13237), .B(new_n13241), .Y(new_n13255));
  O2A1O1Ixp33_ASAP7_75t_L   g12999(.A1(new_n13249), .A2(new_n12912), .B(new_n12931), .C(new_n13246), .Y(new_n13256));
  AOI211xp5_ASAP7_75t_L     g13000(.A1(new_n12916), .A2(new_n13242), .B(new_n13247), .C(new_n12924), .Y(new_n13257));
  OAI21xp33_ASAP7_75t_L     g13001(.A1(new_n13256), .A2(new_n13257), .B(new_n13255), .Y(new_n13258));
  NAND4xp25_ASAP7_75t_L     g13002(.A(new_n13250), .B(new_n13248), .C(new_n13237), .D(new_n13241), .Y(new_n13259));
  AOI21xp33_ASAP7_75t_L     g13003(.A1(new_n12937), .A2(new_n12935), .B(new_n12929), .Y(new_n13260));
  AOI21xp33_ASAP7_75t_L     g13004(.A1(new_n13258), .A2(new_n13259), .B(new_n13260), .Y(new_n13261));
  NOR2xp33_ASAP7_75t_L      g13005(.A(new_n13261), .B(new_n13254), .Y(new_n13262));
  A2O1A1Ixp33_ASAP7_75t_L   g13006(.A1(new_n12950), .A2(new_n12945), .B(new_n12941), .C(new_n13262), .Y(new_n13263));
  INVx1_ASAP7_75t_L         g13007(.A(new_n13263), .Y(new_n13264));
  NOR3xp33_ASAP7_75t_L      g13008(.A(new_n12947), .B(new_n13262), .C(new_n12941), .Y(new_n13265));
  NOR2xp33_ASAP7_75t_L      g13009(.A(new_n13264), .B(new_n13265), .Y(\f[65] ));
  NAND2xp33_ASAP7_75t_L     g13010(.A(new_n13250), .B(new_n13259), .Y(new_n13267));
  AOI22xp33_ASAP7_75t_L     g13011(.A1(new_n600), .A2(\b[57] ), .B1(new_n597), .B2(new_n10495), .Y(new_n13268));
  OAI221xp5_ASAP7_75t_L     g13012(.A1(new_n721), .A2(new_n10178), .B1(new_n9534), .B2(new_n1620), .C(new_n13268), .Y(new_n13269));
  XNOR2x2_ASAP7_75t_L       g13013(.A(\a[11] ), .B(new_n13269), .Y(new_n13270));
  NAND2xp33_ASAP7_75t_L     g13014(.A(new_n13197), .B(new_n13201), .Y(new_n13271));
  NOR3xp33_ASAP7_75t_L      g13015(.A(new_n13198), .B(new_n13199), .C(new_n13196), .Y(new_n13272));
  O2A1O1Ixp33_ASAP7_75t_L   g13016(.A1(new_n12885), .A2(new_n12900), .B(new_n13271), .C(new_n13272), .Y(new_n13273));
  NAND2xp33_ASAP7_75t_L     g13017(.A(new_n13270), .B(new_n13273), .Y(new_n13274));
  INVx1_ASAP7_75t_L         g13018(.A(new_n13272), .Y(new_n13275));
  A2O1A1O1Ixp25_ASAP7_75t_L g13019(.A1(new_n13201), .A2(new_n13197), .B(new_n13202), .C(new_n13275), .D(new_n13270), .Y(new_n13276));
  INVx1_ASAP7_75t_L         g13020(.A(new_n13276), .Y(new_n13277));
  AOI22xp33_ASAP7_75t_L     g13021(.A1(new_n817), .A2(\b[53] ), .B1(\b[54] ), .B2(new_n826), .Y(new_n13278));
  OAI221xp5_ASAP7_75t_L     g13022(.A1(new_n909), .A2(new_n8569), .B1(new_n911), .B2(new_n9207), .C(new_n13278), .Y(new_n13279));
  XNOR2x2_ASAP7_75t_L       g13023(.A(\a[14] ), .B(new_n13279), .Y(new_n13280));
  INVx1_ASAP7_75t_L         g13024(.A(new_n13280), .Y(new_n13281));
  O2A1O1Ixp33_ASAP7_75t_L   g13025(.A1(new_n13191), .A2(new_n13192), .B(new_n13189), .C(new_n13281), .Y(new_n13282));
  INVx1_ASAP7_75t_L         g13026(.A(new_n13282), .Y(new_n13283));
  INVx1_ASAP7_75t_L         g13027(.A(new_n13189), .Y(new_n13284));
  O2A1O1Ixp33_ASAP7_75t_L   g13028(.A1(new_n12883), .A2(new_n12954), .B(new_n13185), .C(new_n13284), .Y(new_n13285));
  NAND2xp33_ASAP7_75t_L     g13029(.A(new_n13281), .B(new_n13285), .Y(new_n13286));
  AOI22xp33_ASAP7_75t_L     g13030(.A1(new_n1113), .A2(\b[51] ), .B1(new_n1110), .B2(new_n8257), .Y(new_n13287));
  OAI221xp5_ASAP7_75t_L     g13031(.A1(new_n1298), .A2(new_n8228), .B1(new_n7907), .B2(new_n1195), .C(new_n13287), .Y(new_n13288));
  XNOR2x2_ASAP7_75t_L       g13032(.A(\a[17] ), .B(new_n13288), .Y(new_n13289));
  INVx1_ASAP7_75t_L         g13033(.A(new_n13289), .Y(new_n13290));
  NAND2xp33_ASAP7_75t_L     g13034(.A(new_n13179), .B(new_n13177), .Y(new_n13291));
  A2O1A1Ixp33_ASAP7_75t_L   g13035(.A1(new_n12966), .A2(new_n12964), .B(new_n13291), .C(new_n13187), .Y(new_n13292));
  NOR2xp33_ASAP7_75t_L      g13036(.A(new_n13290), .B(new_n13292), .Y(new_n13293));
  O2A1O1Ixp33_ASAP7_75t_L   g13037(.A1(new_n13175), .A2(new_n13291), .B(new_n13187), .C(new_n13289), .Y(new_n13294));
  AOI22xp33_ASAP7_75t_L     g13038(.A1(new_n1406), .A2(\b[48] ), .B1(new_n1404), .B2(new_n7341), .Y(new_n13295));
  OAI221xp5_ASAP7_75t_L     g13039(.A1(new_n1398), .A2(new_n7316), .B1(new_n7033), .B2(new_n1549), .C(new_n13295), .Y(new_n13296));
  XNOR2x2_ASAP7_75t_L       g13040(.A(\a[20] ), .B(new_n13296), .Y(new_n13297));
  A2O1A1O1Ixp25_ASAP7_75t_L g13041(.A1(new_n12864), .A2(new_n12861), .B(new_n13176), .C(new_n13166), .D(new_n13170), .Y(new_n13298));
  NAND2xp33_ASAP7_75t_L     g13042(.A(new_n13297), .B(new_n13298), .Y(new_n13299));
  O2A1O1Ixp33_ASAP7_75t_L   g13043(.A1(new_n13171), .A2(new_n13178), .B(new_n13162), .C(new_n13297), .Y(new_n13300));
  INVx1_ASAP7_75t_L         g13044(.A(new_n13300), .Y(new_n13301));
  NAND2xp33_ASAP7_75t_L     g13045(.A(new_n13299), .B(new_n13301), .Y(new_n13302));
  AOI22xp33_ASAP7_75t_L     g13046(.A1(new_n1766), .A2(\b[45] ), .B1(new_n1764), .B2(new_n6764), .Y(new_n13303));
  OAI221xp5_ASAP7_75t_L     g13047(.A1(new_n1758), .A2(new_n6220), .B1(new_n6195), .B2(new_n1911), .C(new_n13303), .Y(new_n13304));
  XNOR2x2_ASAP7_75t_L       g13048(.A(\a[23] ), .B(new_n13304), .Y(new_n13305));
  INVx1_ASAP7_75t_L         g13049(.A(new_n13305), .Y(new_n13306));
  A2O1A1O1Ixp25_ASAP7_75t_L g13050(.A1(new_n13157), .A2(new_n12972), .B(new_n13158), .C(new_n13153), .D(new_n13306), .Y(new_n13307));
  A2O1A1O1Ixp25_ASAP7_75t_L g13051(.A1(new_n12848), .A2(new_n12844), .B(new_n12849), .C(new_n12972), .D(new_n13158), .Y(new_n13308));
  NOR3xp33_ASAP7_75t_L      g13052(.A(new_n13308), .B(new_n13305), .C(new_n13159), .Y(new_n13309));
  NOR2xp33_ASAP7_75t_L      g13053(.A(new_n13309), .B(new_n13307), .Y(new_n13310));
  NAND2xp33_ASAP7_75t_L     g13054(.A(new_n13131), .B(new_n13135), .Y(new_n13311));
  AOI22xp33_ASAP7_75t_L     g13055(.A1(new_n2228), .A2(\b[42] ), .B1(new_n2226), .B2(new_n5688), .Y(new_n13312));
  OAI221xp5_ASAP7_75t_L     g13056(.A1(new_n2220), .A2(new_n5666), .B1(new_n5186), .B2(new_n2387), .C(new_n13312), .Y(new_n13313));
  XNOR2x2_ASAP7_75t_L       g13057(.A(\a[26] ), .B(new_n13313), .Y(new_n13314));
  OA211x2_ASAP7_75t_L       g13058(.A1(new_n13311), .A2(new_n13138), .B(new_n13151), .C(new_n13314), .Y(new_n13315));
  O2A1O1Ixp33_ASAP7_75t_L   g13059(.A1(new_n13311), .A2(new_n13138), .B(new_n13151), .C(new_n13314), .Y(new_n13316));
  NOR2xp33_ASAP7_75t_L      g13060(.A(new_n13316), .B(new_n13315), .Y(new_n13317));
  NAND2xp33_ASAP7_75t_L     g13061(.A(new_n2700), .B(new_n5174), .Y(new_n13318));
  AOI22xp33_ASAP7_75t_L     g13062(.A1(new_n2706), .A2(\b[38] ), .B1(\b[39] ), .B2(new_n2702), .Y(new_n13319));
  OAI211xp5_ASAP7_75t_L     g13063(.A1(new_n2932), .A2(new_n4701), .B(new_n13318), .C(new_n13319), .Y(new_n13320));
  XNOR2x2_ASAP7_75t_L       g13064(.A(\a[29] ), .B(new_n13320), .Y(new_n13321));
  O2A1O1Ixp33_ASAP7_75t_L   g13065(.A1(new_n13130), .A2(new_n12975), .B(new_n13133), .C(new_n13321), .Y(new_n13322));
  O2A1O1Ixp33_ASAP7_75t_L   g13066(.A1(new_n12974), .A2(new_n13132), .B(new_n13134), .C(new_n13126), .Y(new_n13323));
  AND2x2_ASAP7_75t_L        g13067(.A(new_n13321), .B(new_n13323), .Y(new_n13324));
  AOI22xp33_ASAP7_75t_L     g13068(.A1(new_n9623), .A2(\b[12] ), .B1(new_n9620), .B2(new_n970), .Y(new_n13325));
  OAI221xp5_ASAP7_75t_L     g13069(.A1(new_n10280), .A2(new_n695), .B1(new_n631), .B2(new_n12010), .C(new_n13325), .Y(new_n13326));
  XNOR2x2_ASAP7_75t_L       g13070(.A(\a[56] ), .B(new_n13326), .Y(new_n13327));
  INVx1_ASAP7_75t_L         g13071(.A(new_n13327), .Y(new_n13328));
  INVx1_ASAP7_75t_L         g13072(.A(new_n13014), .Y(new_n13329));
  NOR2xp33_ASAP7_75t_L      g13073(.A(new_n278), .B(new_n12671), .Y(new_n13330));
  A2O1A1Ixp33_ASAP7_75t_L   g13074(.A1(new_n12669), .A2(\b[3] ), .B(new_n13330), .C(\a[2] ), .Y(new_n13331));
  O2A1O1Ixp33_ASAP7_75t_L   g13075(.A1(new_n12353), .A2(new_n12355), .B(\b[3] ), .C(new_n13330), .Y(new_n13332));
  NAND2xp33_ASAP7_75t_L     g13076(.A(new_n265), .B(new_n13332), .Y(new_n13333));
  NAND2xp33_ASAP7_75t_L     g13077(.A(new_n13331), .B(new_n13333), .Y(new_n13334));
  AOI22xp33_ASAP7_75t_L     g13078(.A1(new_n11647), .A2(\b[5] ), .B1(\b[6] ), .B2(new_n11656), .Y(new_n13335));
  OAI221xp5_ASAP7_75t_L     g13079(.A1(new_n13003), .A2(new_n323), .B1(new_n12022), .B2(new_n540), .C(new_n13335), .Y(new_n13336));
  XNOR2x2_ASAP7_75t_L       g13080(.A(\a[62] ), .B(new_n13336), .Y(new_n13337));
  NOR2xp33_ASAP7_75t_L      g13081(.A(new_n13334), .B(new_n13337), .Y(new_n13338));
  INVx1_ASAP7_75t_L         g13082(.A(new_n13338), .Y(new_n13339));
  NAND2xp33_ASAP7_75t_L     g13083(.A(new_n13334), .B(new_n13337), .Y(new_n13340));
  NAND2xp33_ASAP7_75t_L     g13084(.A(new_n13340), .B(new_n13339), .Y(new_n13341));
  INVx1_ASAP7_75t_L         g13085(.A(new_n13341), .Y(new_n13342));
  A2O1A1Ixp33_ASAP7_75t_L   g13086(.A1(new_n13006), .A2(new_n13002), .B(new_n13329), .C(new_n13342), .Y(new_n13343));
  A2O1A1Ixp33_ASAP7_75t_L   g13087(.A1(new_n12669), .A2(\b[2] ), .B(new_n13000), .C(new_n13006), .Y(new_n13344));
  AND3x1_ASAP7_75t_L        g13088(.A(new_n13341), .B(new_n13344), .C(new_n13014), .Y(new_n13345));
  INVx1_ASAP7_75t_L         g13089(.A(new_n13345), .Y(new_n13346));
  AOI22xp33_ASAP7_75t_L     g13090(.A1(new_n10594), .A2(\b[9] ), .B1(new_n10591), .B2(new_n566), .Y(new_n13347));
  OAI221xp5_ASAP7_75t_L     g13091(.A1(new_n11335), .A2(new_n503), .B1(new_n421), .B2(new_n11330), .C(new_n13347), .Y(new_n13348));
  XNOR2x2_ASAP7_75t_L       g13092(.A(\a[59] ), .B(new_n13348), .Y(new_n13349));
  AND3x1_ASAP7_75t_L        g13093(.A(new_n13346), .B(new_n13349), .C(new_n13343), .Y(new_n13350));
  AOI21xp33_ASAP7_75t_L     g13094(.A1(new_n13346), .A2(new_n13343), .B(new_n13349), .Y(new_n13351));
  NOR2xp33_ASAP7_75t_L      g13095(.A(new_n13351), .B(new_n13350), .Y(new_n13352));
  A2O1A1Ixp33_ASAP7_75t_L   g13096(.A1(new_n13010), .A2(new_n13014), .B(new_n13020), .C(new_n13023), .Y(new_n13353));
  O2A1O1Ixp33_ASAP7_75t_L   g13097(.A1(new_n13018), .A2(new_n13015), .B(new_n13353), .C(new_n13352), .Y(new_n13354));
  A2O1A1Ixp33_ASAP7_75t_L   g13098(.A1(new_n12695), .A2(new_n12999), .B(new_n13024), .C(new_n13021), .Y(new_n13355));
  NOR3xp33_ASAP7_75t_L      g13099(.A(new_n13355), .B(new_n13351), .C(new_n13350), .Y(new_n13356));
  NOR2xp33_ASAP7_75t_L      g13100(.A(new_n13356), .B(new_n13354), .Y(new_n13357));
  XNOR2x2_ASAP7_75t_L       g13101(.A(new_n13328), .B(new_n13357), .Y(new_n13358));
  O2A1O1Ixp33_ASAP7_75t_L   g13102(.A1(new_n12995), .A2(new_n13037), .B(new_n13028), .C(new_n13358), .Y(new_n13359));
  A2O1A1O1Ixp25_ASAP7_75t_L g13103(.A1(new_n12705), .A2(new_n12994), .B(new_n12712), .C(new_n13027), .D(new_n13038), .Y(new_n13360));
  AND2x2_ASAP7_75t_L        g13104(.A(new_n13360), .B(new_n13358), .Y(new_n13361));
  AOI22xp33_ASAP7_75t_L     g13105(.A1(new_n8645), .A2(\b[15] ), .B1(new_n8642), .B2(new_n959), .Y(new_n13362));
  OAI221xp5_ASAP7_75t_L     g13106(.A1(new_n9322), .A2(new_n871), .B1(new_n793), .B2(new_n8965), .C(new_n13362), .Y(new_n13363));
  XNOR2x2_ASAP7_75t_L       g13107(.A(new_n8639), .B(new_n13363), .Y(new_n13364));
  NOR3xp33_ASAP7_75t_L      g13108(.A(new_n13361), .B(new_n13364), .C(new_n13359), .Y(new_n13365));
  OA21x2_ASAP7_75t_L        g13109(.A1(new_n13359), .A2(new_n13361), .B(new_n13364), .Y(new_n13366));
  NAND3xp33_ASAP7_75t_L     g13110(.A(new_n13039), .B(new_n13040), .C(new_n13035), .Y(new_n13367));
  A2O1A1Ixp33_ASAP7_75t_L   g13111(.A1(new_n13044), .A2(new_n13045), .B(new_n13043), .C(new_n13367), .Y(new_n13368));
  OR3x1_ASAP7_75t_L         g13112(.A(new_n13366), .B(new_n13365), .C(new_n13368), .Y(new_n13369));
  OAI21xp33_ASAP7_75t_L     g13113(.A1(new_n13365), .A2(new_n13366), .B(new_n13368), .Y(new_n13370));
  AOI22xp33_ASAP7_75t_L     g13114(.A1(new_n7659), .A2(\b[18] ), .B1(new_n7656), .B2(new_n1363), .Y(new_n13371));
  OAI221xp5_ASAP7_75t_L     g13115(.A1(new_n8326), .A2(new_n1244), .B1(new_n1051), .B2(new_n7994), .C(new_n13371), .Y(new_n13372));
  XNOR2x2_ASAP7_75t_L       g13116(.A(\a[50] ), .B(new_n13372), .Y(new_n13373));
  NAND3xp33_ASAP7_75t_L     g13117(.A(new_n13369), .B(new_n13370), .C(new_n13373), .Y(new_n13374));
  AO21x2_ASAP7_75t_L        g13118(.A1(new_n13370), .A2(new_n13369), .B(new_n13373), .Y(new_n13375));
  INVx1_ASAP7_75t_L         g13119(.A(new_n13047), .Y(new_n13376));
  O2A1O1Ixp33_ASAP7_75t_L   g13120(.A1(new_n12988), .A2(new_n12743), .B(new_n13048), .C(new_n13376), .Y(new_n13377));
  AND3x1_ASAP7_75t_L        g13121(.A(new_n13375), .B(new_n13377), .C(new_n13374), .Y(new_n13378));
  AND2x2_ASAP7_75t_L        g13122(.A(new_n13374), .B(new_n13375), .Y(new_n13379));
  O2A1O1Ixp33_ASAP7_75t_L   g13123(.A1(new_n12989), .A2(new_n13049), .B(new_n13047), .C(new_n13379), .Y(new_n13380));
  AOI22xp33_ASAP7_75t_L     g13124(.A1(new_n6822), .A2(\b[21] ), .B1(new_n6819), .B2(new_n1715), .Y(new_n13381));
  OAI221xp5_ASAP7_75t_L     g13125(.A1(new_n7392), .A2(new_n1594), .B1(new_n1493), .B2(new_n7115), .C(new_n13381), .Y(new_n13382));
  XNOR2x2_ASAP7_75t_L       g13126(.A(\a[47] ), .B(new_n13382), .Y(new_n13383));
  OAI21xp33_ASAP7_75t_L     g13127(.A1(new_n13378), .A2(new_n13380), .B(new_n13383), .Y(new_n13384));
  NOR2xp33_ASAP7_75t_L      g13128(.A(new_n13378), .B(new_n13380), .Y(new_n13385));
  INVx1_ASAP7_75t_L         g13129(.A(new_n13383), .Y(new_n13386));
  NAND2xp33_ASAP7_75t_L     g13130(.A(new_n13386), .B(new_n13385), .Y(new_n13387));
  NAND2xp33_ASAP7_75t_L     g13131(.A(new_n13384), .B(new_n13387), .Y(new_n13388));
  NOR2xp33_ASAP7_75t_L      g13132(.A(new_n13056), .B(new_n13057), .Y(new_n13389));
  NAND2xp33_ASAP7_75t_L     g13133(.A(new_n13058), .B(new_n13389), .Y(new_n13390));
  A2O1A1O1Ixp25_ASAP7_75t_L g13134(.A1(new_n13055), .A2(new_n13059), .B(new_n12986), .C(new_n13390), .D(new_n13388), .Y(new_n13391));
  A2O1A1Ixp33_ASAP7_75t_L   g13135(.A1(new_n13055), .A2(new_n13059), .B(new_n12986), .C(new_n13390), .Y(new_n13392));
  AOI21xp33_ASAP7_75t_L     g13136(.A1(new_n13387), .A2(new_n13384), .B(new_n13392), .Y(new_n13393));
  AOI22xp33_ASAP7_75t_L     g13137(.A1(new_n6002), .A2(\b[24] ), .B1(new_n5999), .B2(new_n2027), .Y(new_n13394));
  OAI221xp5_ASAP7_75t_L     g13138(.A1(new_n6544), .A2(new_n1995), .B1(new_n1857), .B2(new_n6309), .C(new_n13394), .Y(new_n13395));
  XNOR2x2_ASAP7_75t_L       g13139(.A(\a[44] ), .B(new_n13395), .Y(new_n13396));
  INVx1_ASAP7_75t_L         g13140(.A(new_n13396), .Y(new_n13397));
  OR3x1_ASAP7_75t_L         g13141(.A(new_n13391), .B(new_n13393), .C(new_n13397), .Y(new_n13398));
  OAI21xp33_ASAP7_75t_L     g13142(.A1(new_n13393), .A2(new_n13391), .B(new_n13397), .Y(new_n13399));
  NAND2xp33_ASAP7_75t_L     g13143(.A(new_n13399), .B(new_n13398), .Y(new_n13400));
  NOR3xp33_ASAP7_75t_L      g13144(.A(new_n13400), .B(new_n13075), .C(new_n13065), .Y(new_n13401));
  INVx1_ASAP7_75t_L         g13145(.A(new_n13401), .Y(new_n13402));
  A2O1A1Ixp33_ASAP7_75t_L   g13146(.A1(new_n13073), .A2(new_n12982), .B(new_n13065), .C(new_n13400), .Y(new_n13403));
  AOI22xp33_ASAP7_75t_L     g13147(.A1(new_n5249), .A2(\b[27] ), .B1(new_n5247), .B2(new_n2657), .Y(new_n13404));
  OAI221xp5_ASAP7_75t_L     g13148(.A1(new_n5241), .A2(new_n2477), .B1(new_n2180), .B2(new_n5521), .C(new_n13404), .Y(new_n13405));
  XNOR2x2_ASAP7_75t_L       g13149(.A(\a[41] ), .B(new_n13405), .Y(new_n13406));
  NAND3xp33_ASAP7_75t_L     g13150(.A(new_n13402), .B(new_n13403), .C(new_n13406), .Y(new_n13407));
  AO21x2_ASAP7_75t_L        g13151(.A1(new_n13403), .A2(new_n13402), .B(new_n13406), .Y(new_n13408));
  NOR2xp33_ASAP7_75t_L      g13152(.A(new_n13071), .B(new_n13075), .Y(new_n13409));
  NAND2xp33_ASAP7_75t_L     g13153(.A(new_n13079), .B(new_n13409), .Y(new_n13410));
  A2O1A1Ixp33_ASAP7_75t_L   g13154(.A1(new_n13091), .A2(new_n13090), .B(new_n13088), .C(new_n13410), .Y(new_n13411));
  INVx1_ASAP7_75t_L         g13155(.A(new_n13411), .Y(new_n13412));
  NAND3xp33_ASAP7_75t_L     g13156(.A(new_n13408), .B(new_n13407), .C(new_n13412), .Y(new_n13413));
  NAND2xp33_ASAP7_75t_L     g13157(.A(new_n13407), .B(new_n13408), .Y(new_n13414));
  A2O1A1Ixp33_ASAP7_75t_L   g13158(.A1(new_n13079), .A2(new_n13409), .B(new_n13099), .C(new_n13414), .Y(new_n13415));
  AOI22xp33_ASAP7_75t_L     g13159(.A1(new_n4544), .A2(\b[30] ), .B1(new_n4542), .B2(new_n3219), .Y(new_n13416));
  OAI221xp5_ASAP7_75t_L     g13160(.A1(new_n4536), .A2(new_n2871), .B1(new_n2852), .B2(new_n4781), .C(new_n13416), .Y(new_n13417));
  XNOR2x2_ASAP7_75t_L       g13161(.A(new_n4539), .B(new_n13417), .Y(new_n13418));
  AO21x2_ASAP7_75t_L        g13162(.A1(new_n13413), .A2(new_n13415), .B(new_n13418), .Y(new_n13419));
  NAND3xp33_ASAP7_75t_L     g13163(.A(new_n13415), .B(new_n13413), .C(new_n13418), .Y(new_n13420));
  NAND3xp33_ASAP7_75t_L     g13164(.A(new_n13093), .B(new_n13089), .C(new_n13100), .Y(new_n13421));
  A2O1A1Ixp33_ASAP7_75t_L   g13165(.A1(new_n13104), .A2(new_n13108), .B(new_n13111), .C(new_n13421), .Y(new_n13422));
  NAND3xp33_ASAP7_75t_L     g13166(.A(new_n13419), .B(new_n13420), .C(new_n13422), .Y(new_n13423));
  INVx1_ASAP7_75t_L         g13167(.A(new_n13423), .Y(new_n13424));
  AOI21xp33_ASAP7_75t_L     g13168(.A1(new_n13419), .A2(new_n13420), .B(new_n13422), .Y(new_n13425));
  AOI22xp33_ASAP7_75t_L     g13169(.A1(new_n3884), .A2(\b[33] ), .B1(new_n3881), .B2(new_n3813), .Y(new_n13426));
  OAI221xp5_ASAP7_75t_L     g13170(.A1(new_n4312), .A2(new_n3443), .B1(new_n3419), .B2(new_n4986), .C(new_n13426), .Y(new_n13427));
  XNOR2x2_ASAP7_75t_L       g13171(.A(\a[35] ), .B(new_n13427), .Y(new_n13428));
  INVx1_ASAP7_75t_L         g13172(.A(new_n13428), .Y(new_n13429));
  NOR3xp33_ASAP7_75t_L      g13173(.A(new_n13424), .B(new_n13425), .C(new_n13429), .Y(new_n13430));
  INVx1_ASAP7_75t_L         g13174(.A(new_n13425), .Y(new_n13431));
  AOI21xp33_ASAP7_75t_L     g13175(.A1(new_n13431), .A2(new_n13423), .B(new_n13428), .Y(new_n13432));
  NOR2xp33_ASAP7_75t_L      g13176(.A(new_n13430), .B(new_n13432), .Y(new_n13433));
  NAND2xp33_ASAP7_75t_L     g13177(.A(new_n3254), .B(new_n4473), .Y(new_n13434));
  AOI22xp33_ASAP7_75t_L     g13178(.A1(new_n3260), .A2(\b[35] ), .B1(\b[36] ), .B2(new_n3256), .Y(new_n13435));
  OAI211xp5_ASAP7_75t_L     g13179(.A1(new_n3492), .A2(new_n3827), .B(new_n13434), .C(new_n13435), .Y(new_n13436));
  XNOR2x2_ASAP7_75t_L       g13180(.A(\a[32] ), .B(new_n13436), .Y(new_n13437));
  INVx1_ASAP7_75t_L         g13181(.A(new_n13437), .Y(new_n13438));
  A2O1A1Ixp33_ASAP7_75t_L   g13182(.A1(new_n12823), .A2(new_n12979), .B(new_n12813), .C(new_n13116), .Y(new_n13439));
  NAND2xp33_ASAP7_75t_L     g13183(.A(new_n13120), .B(new_n13439), .Y(new_n13440));
  XNOR2x2_ASAP7_75t_L       g13184(.A(new_n13438), .B(new_n13440), .Y(new_n13441));
  XNOR2x2_ASAP7_75t_L       g13185(.A(new_n13441), .B(new_n13433), .Y(new_n13442));
  OR3x1_ASAP7_75t_L         g13186(.A(new_n13442), .B(new_n13322), .C(new_n13324), .Y(new_n13443));
  NOR2xp33_ASAP7_75t_L      g13187(.A(new_n13322), .B(new_n13324), .Y(new_n13444));
  INVx1_ASAP7_75t_L         g13188(.A(new_n13444), .Y(new_n13445));
  NAND2xp33_ASAP7_75t_L     g13189(.A(new_n13445), .B(new_n13442), .Y(new_n13446));
  AND2x2_ASAP7_75t_L        g13190(.A(new_n13446), .B(new_n13443), .Y(new_n13447));
  XNOR2x2_ASAP7_75t_L       g13191(.A(new_n13317), .B(new_n13447), .Y(new_n13448));
  XNOR2x2_ASAP7_75t_L       g13192(.A(new_n13310), .B(new_n13448), .Y(new_n13449));
  NOR2xp33_ASAP7_75t_L      g13193(.A(new_n13302), .B(new_n13449), .Y(new_n13450));
  INVx1_ASAP7_75t_L         g13194(.A(new_n13450), .Y(new_n13451));
  NAND2xp33_ASAP7_75t_L     g13195(.A(new_n13302), .B(new_n13449), .Y(new_n13452));
  NAND2xp33_ASAP7_75t_L     g13196(.A(new_n13452), .B(new_n13451), .Y(new_n13453));
  OR3x1_ASAP7_75t_L         g13197(.A(new_n13293), .B(new_n13294), .C(new_n13453), .Y(new_n13454));
  OAI21xp33_ASAP7_75t_L     g13198(.A1(new_n13294), .A2(new_n13293), .B(new_n13453), .Y(new_n13455));
  AND4x1_ASAP7_75t_L        g13199(.A(new_n13455), .B(new_n13454), .C(new_n13286), .D(new_n13283), .Y(new_n13456));
  AOI22xp33_ASAP7_75t_L     g13200(.A1(new_n13286), .A2(new_n13283), .B1(new_n13455), .B2(new_n13454), .Y(new_n13457));
  NOR2xp33_ASAP7_75t_L      g13201(.A(new_n13457), .B(new_n13456), .Y(new_n13458));
  NAND3xp33_ASAP7_75t_L     g13202(.A(new_n13274), .B(new_n13277), .C(new_n13458), .Y(new_n13459));
  INVx1_ASAP7_75t_L         g13203(.A(new_n13270), .Y(new_n13460));
  A2O1A1Ixp33_ASAP7_75t_L   g13204(.A1(new_n13201), .A2(new_n13197), .B(new_n13202), .C(new_n13275), .Y(new_n13461));
  NOR2xp33_ASAP7_75t_L      g13205(.A(new_n13460), .B(new_n13461), .Y(new_n13462));
  INVx1_ASAP7_75t_L         g13206(.A(new_n13458), .Y(new_n13463));
  OAI21xp33_ASAP7_75t_L     g13207(.A1(new_n13276), .A2(new_n13462), .B(new_n13463), .Y(new_n13464));
  NAND2xp33_ASAP7_75t_L     g13208(.A(new_n13459), .B(new_n13464), .Y(new_n13465));
  OAI32xp33_ASAP7_75t_L     g13209(.A1(new_n11233), .A2(new_n11230), .A3(new_n482), .B1(new_n667), .B2(new_n11226), .Y(new_n13466));
  AOI221xp5_ASAP7_75t_L     g13210(.A1(\b[58] ), .A2(new_n480), .B1(\b[59] ), .B2(new_n441), .C(new_n13466), .Y(new_n13467));
  XNOR2x2_ASAP7_75t_L       g13211(.A(new_n445), .B(new_n13467), .Y(new_n13468));
  INVx1_ASAP7_75t_L         g13212(.A(new_n13468), .Y(new_n13469));
  O2A1O1Ixp33_ASAP7_75t_L   g13213(.A1(new_n13203), .A2(new_n13204), .B(new_n13207), .C(new_n13227), .Y(new_n13470));
  NAND2xp33_ASAP7_75t_L     g13214(.A(new_n13469), .B(new_n13470), .Y(new_n13471));
  O2A1O1Ixp33_ASAP7_75t_L   g13215(.A1(new_n13218), .A2(new_n13222), .B(new_n13208), .C(new_n13469), .Y(new_n13472));
  INVx1_ASAP7_75t_L         g13216(.A(new_n13472), .Y(new_n13473));
  NAND3xp33_ASAP7_75t_L     g13217(.A(new_n13471), .B(new_n13465), .C(new_n13473), .Y(new_n13474));
  INVx1_ASAP7_75t_L         g13218(.A(new_n13459), .Y(new_n13475));
  AOI21xp33_ASAP7_75t_L     g13219(.A1(new_n13274), .A2(new_n13277), .B(new_n13458), .Y(new_n13476));
  NOR2xp33_ASAP7_75t_L      g13220(.A(new_n13476), .B(new_n13475), .Y(new_n13477));
  A2O1A1Ixp33_ASAP7_75t_L   g13221(.A1(new_n13210), .A2(new_n13209), .B(new_n13211), .C(new_n13220), .Y(new_n13478));
  NOR2xp33_ASAP7_75t_L      g13222(.A(new_n13468), .B(new_n13478), .Y(new_n13479));
  OAI21xp33_ASAP7_75t_L     g13223(.A1(new_n13472), .A2(new_n13479), .B(new_n13477), .Y(new_n13480));
  NAND2xp33_ASAP7_75t_L     g13224(.A(new_n13480), .B(new_n13474), .Y(new_n13481));
  NAND2xp33_ASAP7_75t_L     g13225(.A(\b[63] ), .B(new_n345), .Y(new_n13482));
  A2O1A1Ixp33_ASAP7_75t_L   g13226(.A1(new_n12607), .A2(new_n12603), .B(new_n367), .C(new_n13482), .Y(new_n13483));
  AOI221xp5_ASAP7_75t_L     g13227(.A1(\b[61] ), .A2(new_n366), .B1(\b[62] ), .B2(new_n334), .C(new_n13483), .Y(new_n13484));
  XNOR2x2_ASAP7_75t_L       g13228(.A(new_n339), .B(new_n13484), .Y(new_n13485));
  INVx1_ASAP7_75t_L         g13229(.A(new_n13485), .Y(new_n13486));
  AOI21xp33_ASAP7_75t_L     g13230(.A1(new_n13230), .A2(new_n13236), .B(new_n13238), .Y(new_n13487));
  NAND2xp33_ASAP7_75t_L     g13231(.A(new_n13486), .B(new_n13487), .Y(new_n13488));
  A2O1A1Ixp33_ASAP7_75t_L   g13232(.A1(new_n13230), .A2(new_n13236), .B(new_n13238), .C(new_n13485), .Y(new_n13489));
  NAND2xp33_ASAP7_75t_L     g13233(.A(new_n13489), .B(new_n13488), .Y(new_n13490));
  NOR2xp33_ASAP7_75t_L      g13234(.A(new_n13481), .B(new_n13490), .Y(new_n13491));
  AND2x2_ASAP7_75t_L        g13235(.A(new_n13480), .B(new_n13474), .Y(new_n13492));
  AOI21xp33_ASAP7_75t_L     g13236(.A1(new_n13489), .A2(new_n13488), .B(new_n13492), .Y(new_n13493));
  OAI21xp33_ASAP7_75t_L     g13237(.A1(new_n13491), .A2(new_n13493), .B(new_n13267), .Y(new_n13494));
  NOR2xp33_ASAP7_75t_L      g13238(.A(new_n13257), .B(new_n13252), .Y(new_n13495));
  NAND3xp33_ASAP7_75t_L     g13239(.A(new_n13492), .B(new_n13488), .C(new_n13489), .Y(new_n13496));
  NAND2xp33_ASAP7_75t_L     g13240(.A(new_n13481), .B(new_n13490), .Y(new_n13497));
  NAND3xp33_ASAP7_75t_L     g13241(.A(new_n13496), .B(new_n13495), .C(new_n13497), .Y(new_n13498));
  NAND2xp33_ASAP7_75t_L     g13242(.A(new_n13498), .B(new_n13494), .Y(new_n13499));
  A2O1A1O1Ixp25_ASAP7_75t_L g13243(.A1(new_n13259), .A2(new_n13258), .B(new_n13260), .C(new_n13263), .D(new_n13499), .Y(new_n13500));
  INVx1_ASAP7_75t_L         g13244(.A(new_n13261), .Y(new_n13501));
  AND3x1_ASAP7_75t_L        g13245(.A(new_n13499), .B(new_n13263), .C(new_n13501), .Y(new_n13502));
  NOR2xp33_ASAP7_75t_L      g13246(.A(new_n13500), .B(new_n13502), .Y(\f[66] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g13247(.A1(new_n12945), .A2(new_n12950), .B(new_n12941), .C(new_n13262), .D(new_n13261), .Y(new_n13504));
  AOI21xp33_ASAP7_75t_L     g13248(.A1(new_n13487), .A2(new_n13486), .B(new_n13491), .Y(new_n13505));
  INVx1_ASAP7_75t_L         g13249(.A(new_n12628), .Y(new_n13506));
  NAND2xp33_ASAP7_75t_L     g13250(.A(new_n12600), .B(new_n12597), .Y(new_n13507));
  AOI22xp33_ASAP7_75t_L     g13251(.A1(new_n334), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n366), .Y(new_n13508));
  A2O1A1Ixp33_ASAP7_75t_L   g13252(.A1(new_n13506), .A2(new_n13507), .B(new_n367), .C(new_n13508), .Y(new_n13509));
  NOR2xp33_ASAP7_75t_L      g13253(.A(new_n339), .B(new_n13509), .Y(new_n13510));
  A2O1A1O1Ixp25_ASAP7_75t_L g13254(.A1(new_n13507), .A2(new_n13506), .B(new_n367), .C(new_n13508), .D(\a[5] ), .Y(new_n13511));
  NOR2xp33_ASAP7_75t_L      g13255(.A(new_n13511), .B(new_n13510), .Y(new_n13512));
  A2O1A1Ixp33_ASAP7_75t_L   g13256(.A1(new_n13465), .A2(new_n13473), .B(new_n13479), .C(new_n13512), .Y(new_n13513));
  O2A1O1Ixp33_ASAP7_75t_L   g13257(.A1(new_n13476), .A2(new_n13475), .B(new_n13473), .C(new_n13479), .Y(new_n13514));
  INVx1_ASAP7_75t_L         g13258(.A(new_n13512), .Y(new_n13515));
  NAND2xp33_ASAP7_75t_L     g13259(.A(new_n13515), .B(new_n13514), .Y(new_n13516));
  NAND2xp33_ASAP7_75t_L     g13260(.A(new_n13455), .B(new_n13454), .Y(new_n13517));
  A2O1A1Ixp33_ASAP7_75t_L   g13261(.A1(new_n12956), .A2(new_n13185), .B(new_n13284), .C(new_n13281), .Y(new_n13518));
  A2O1A1Ixp33_ASAP7_75t_L   g13262(.A1(new_n13286), .A2(new_n13283), .B(new_n13517), .C(new_n13518), .Y(new_n13519));
  AOI22xp33_ASAP7_75t_L     g13263(.A1(new_n590), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n600), .Y(new_n13520));
  OAI221xp5_ASAP7_75t_L     g13264(.A1(new_n1620), .A2(new_n10178), .B1(new_n675), .B2(new_n10856), .C(new_n13520), .Y(new_n13521));
  XNOR2x2_ASAP7_75t_L       g13265(.A(\a[11] ), .B(new_n13521), .Y(new_n13522));
  XNOR2x2_ASAP7_75t_L       g13266(.A(new_n13522), .B(new_n13519), .Y(new_n13523));
  AOI22xp33_ASAP7_75t_L     g13267(.A1(new_n826), .A2(\b[55] ), .B1(new_n823), .B2(new_n9542), .Y(new_n13524));
  OAI221xp5_ASAP7_75t_L     g13268(.A1(new_n994), .A2(new_n9199), .B1(new_n8882), .B2(new_n909), .C(new_n13524), .Y(new_n13525));
  XNOR2x2_ASAP7_75t_L       g13269(.A(\a[14] ), .B(new_n13525), .Y(new_n13526));
  INVx1_ASAP7_75t_L         g13270(.A(new_n13294), .Y(new_n13527));
  OA21x2_ASAP7_75t_L        g13271(.A1(new_n13453), .A2(new_n13293), .B(new_n13527), .Y(new_n13528));
  AND2x2_ASAP7_75t_L        g13272(.A(new_n13526), .B(new_n13528), .Y(new_n13529));
  O2A1O1Ixp33_ASAP7_75t_L   g13273(.A1(new_n13293), .A2(new_n13453), .B(new_n13527), .C(new_n13526), .Y(new_n13530));
  AOI22xp33_ASAP7_75t_L     g13274(.A1(new_n1406), .A2(\b[49] ), .B1(new_n1404), .B2(new_n7914), .Y(new_n13531));
  OAI221xp5_ASAP7_75t_L     g13275(.A1(new_n1398), .A2(new_n7333), .B1(new_n7316), .B2(new_n1549), .C(new_n13531), .Y(new_n13532));
  XNOR2x2_ASAP7_75t_L       g13276(.A(\a[20] ), .B(new_n13532), .Y(new_n13533));
  INVx1_ASAP7_75t_L         g13277(.A(new_n13533), .Y(new_n13534));
  A2O1A1Ixp33_ASAP7_75t_L   g13278(.A1(new_n13149), .A2(new_n12973), .B(new_n13159), .C(new_n13305), .Y(new_n13535));
  A2O1A1O1Ixp25_ASAP7_75t_L g13279(.A1(new_n12852), .A2(new_n12850), .B(new_n13164), .C(new_n13149), .D(new_n13159), .Y(new_n13536));
  NAND2xp33_ASAP7_75t_L     g13280(.A(new_n13536), .B(new_n13306), .Y(new_n13537));
  A2O1A1Ixp33_ASAP7_75t_L   g13281(.A1(new_n13149), .A2(new_n12973), .B(new_n13159), .C(new_n13306), .Y(new_n13538));
  A2O1A1Ixp33_ASAP7_75t_L   g13282(.A1(new_n13537), .A2(new_n13535), .B(new_n13448), .C(new_n13538), .Y(new_n13539));
  NOR2xp33_ASAP7_75t_L      g13283(.A(new_n13534), .B(new_n13539), .Y(new_n13540));
  O2A1O1Ixp33_ASAP7_75t_L   g13284(.A1(new_n13310), .A2(new_n13448), .B(new_n13538), .C(new_n13533), .Y(new_n13541));
  NOR2xp33_ASAP7_75t_L      g13285(.A(new_n13541), .B(new_n13540), .Y(new_n13542));
  AOI22xp33_ASAP7_75t_L     g13286(.A1(new_n1766), .A2(\b[46] ), .B1(new_n1764), .B2(new_n7041), .Y(new_n13543));
  OAI221xp5_ASAP7_75t_L     g13287(.A1(new_n1758), .A2(new_n6756), .B1(new_n6220), .B2(new_n1911), .C(new_n13543), .Y(new_n13544));
  XNOR2x2_ASAP7_75t_L       g13288(.A(\a[23] ), .B(new_n13544), .Y(new_n13545));
  INVx1_ASAP7_75t_L         g13289(.A(new_n13545), .Y(new_n13546));
  AOI21xp33_ASAP7_75t_L     g13290(.A1(new_n13447), .A2(new_n13317), .B(new_n13316), .Y(new_n13547));
  NAND2xp33_ASAP7_75t_L     g13291(.A(new_n13546), .B(new_n13547), .Y(new_n13548));
  A2O1A1Ixp33_ASAP7_75t_L   g13292(.A1(new_n13447), .A2(new_n13317), .B(new_n13316), .C(new_n13545), .Y(new_n13549));
  AOI22xp33_ASAP7_75t_L     g13293(.A1(new_n2228), .A2(\b[43] ), .B1(new_n2226), .B2(new_n6202), .Y(new_n13550));
  OAI221xp5_ASAP7_75t_L     g13294(.A1(new_n2220), .A2(new_n5680), .B1(new_n5666), .B2(new_n2387), .C(new_n13550), .Y(new_n13551));
  XNOR2x2_ASAP7_75t_L       g13295(.A(\a[26] ), .B(new_n13551), .Y(new_n13552));
  INVx1_ASAP7_75t_L         g13296(.A(new_n13552), .Y(new_n13553));
  INVx1_ASAP7_75t_L         g13297(.A(new_n13322), .Y(new_n13554));
  OAI21xp33_ASAP7_75t_L     g13298(.A1(new_n13324), .A2(new_n13442), .B(new_n13554), .Y(new_n13555));
  NOR2xp33_ASAP7_75t_L      g13299(.A(new_n13553), .B(new_n13555), .Y(new_n13556));
  O2A1O1Ixp33_ASAP7_75t_L   g13300(.A1(new_n13445), .A2(new_n13442), .B(new_n13554), .C(new_n13552), .Y(new_n13557));
  NOR2xp33_ASAP7_75t_L      g13301(.A(new_n13557), .B(new_n13556), .Y(new_n13558));
  INVx1_ASAP7_75t_L         g13302(.A(new_n4709), .Y(new_n13559));
  AOI22xp33_ASAP7_75t_L     g13303(.A1(new_n3260), .A2(\b[36] ), .B1(\b[37] ), .B2(new_n3256), .Y(new_n13560));
  OAI221xp5_ASAP7_75t_L     g13304(.A1(new_n3492), .A2(new_n4053), .B1(new_n3261), .B2(new_n13559), .C(new_n13560), .Y(new_n13561));
  XNOR2x2_ASAP7_75t_L       g13305(.A(new_n3251), .B(new_n13561), .Y(new_n13562));
  AOI21xp33_ASAP7_75t_L     g13306(.A1(new_n13423), .A2(new_n13428), .B(new_n13425), .Y(new_n13563));
  XNOR2x2_ASAP7_75t_L       g13307(.A(new_n13562), .B(new_n13563), .Y(new_n13564));
  AOI22xp33_ASAP7_75t_L     g13308(.A1(new_n3884), .A2(\b[34] ), .B1(new_n3881), .B2(new_n3833), .Y(new_n13565));
  OAI221xp5_ASAP7_75t_L     g13309(.A1(new_n4312), .A2(new_n3807), .B1(new_n3443), .B2(new_n4986), .C(new_n13565), .Y(new_n13566));
  XNOR2x2_ASAP7_75t_L       g13310(.A(\a[35] ), .B(new_n13566), .Y(new_n13567));
  A2O1A1Ixp33_ASAP7_75t_L   g13311(.A1(new_n13408), .A2(new_n13407), .B(new_n13412), .C(new_n13420), .Y(new_n13568));
  AOI22xp33_ASAP7_75t_L     g13312(.A1(new_n6002), .A2(\b[25] ), .B1(new_n5999), .B2(new_n2188), .Y(new_n13569));
  OAI221xp5_ASAP7_75t_L     g13313(.A1(new_n6544), .A2(new_n2019), .B1(new_n1995), .B2(new_n6309), .C(new_n13569), .Y(new_n13570));
  XNOR2x2_ASAP7_75t_L       g13314(.A(\a[44] ), .B(new_n13570), .Y(new_n13571));
  AOI22xp33_ASAP7_75t_L     g13315(.A1(new_n11656), .A2(\b[7] ), .B1(new_n11654), .B2(new_n611), .Y(new_n13572));
  OAI221xp5_ASAP7_75t_L     g13316(.A1(new_n12364), .A2(new_n382), .B1(new_n353), .B2(new_n13003), .C(new_n13572), .Y(new_n13573));
  XNOR2x2_ASAP7_75t_L       g13317(.A(\a[62] ), .B(new_n13573), .Y(new_n13574));
  NOR2xp33_ASAP7_75t_L      g13318(.A(new_n299), .B(new_n12671), .Y(new_n13575));
  O2A1O1Ixp33_ASAP7_75t_L   g13319(.A1(new_n12353), .A2(new_n12355), .B(\b[4] ), .C(new_n13575), .Y(new_n13576));
  NAND2xp33_ASAP7_75t_L     g13320(.A(\a[2] ), .B(new_n13576), .Y(new_n13577));
  A2O1A1Ixp33_ASAP7_75t_L   g13321(.A1(new_n12669), .A2(\b[4] ), .B(new_n13575), .C(new_n265), .Y(new_n13578));
  AND2x2_ASAP7_75t_L        g13322(.A(new_n13578), .B(new_n13577), .Y(new_n13579));
  XNOR2x2_ASAP7_75t_L       g13323(.A(new_n13579), .B(new_n13574), .Y(new_n13580));
  A2O1A1O1Ixp25_ASAP7_75t_L g13324(.A1(new_n12669), .A2(\b[3] ), .B(new_n13330), .C(\a[2] ), .D(new_n13338), .Y(new_n13581));
  NAND2xp33_ASAP7_75t_L     g13325(.A(new_n13581), .B(new_n13580), .Y(new_n13582));
  O2A1O1Ixp33_ASAP7_75t_L   g13326(.A1(new_n13334), .A2(new_n13337), .B(new_n13331), .C(new_n13580), .Y(new_n13583));
  INVx1_ASAP7_75t_L         g13327(.A(new_n13583), .Y(new_n13584));
  AOI22xp33_ASAP7_75t_L     g13328(.A1(new_n10594), .A2(\b[10] ), .B1(new_n10591), .B2(new_n852), .Y(new_n13585));
  OAI221xp5_ASAP7_75t_L     g13329(.A1(new_n11335), .A2(new_n559), .B1(new_n503), .B2(new_n11330), .C(new_n13585), .Y(new_n13586));
  XNOR2x2_ASAP7_75t_L       g13330(.A(\a[59] ), .B(new_n13586), .Y(new_n13587));
  NAND3xp33_ASAP7_75t_L     g13331(.A(new_n13584), .B(new_n13582), .C(new_n13587), .Y(new_n13588));
  AO21x2_ASAP7_75t_L        g13332(.A1(new_n13582), .A2(new_n13584), .B(new_n13587), .Y(new_n13589));
  NAND2xp33_ASAP7_75t_L     g13333(.A(new_n13588), .B(new_n13589), .Y(new_n13590));
  INVx1_ASAP7_75t_L         g13334(.A(new_n13590), .Y(new_n13591));
  A2O1A1Ixp33_ASAP7_75t_L   g13335(.A1(new_n13349), .A2(new_n13343), .B(new_n13345), .C(new_n13591), .Y(new_n13592));
  NOR2xp33_ASAP7_75t_L      g13336(.A(new_n13345), .B(new_n13350), .Y(new_n13593));
  NAND2xp33_ASAP7_75t_L     g13337(.A(new_n13593), .B(new_n13590), .Y(new_n13594));
  NAND2xp33_ASAP7_75t_L     g13338(.A(new_n13594), .B(new_n13592), .Y(new_n13595));
  AOI22xp33_ASAP7_75t_L     g13339(.A1(new_n9623), .A2(\b[13] ), .B1(new_n9620), .B2(new_n800), .Y(new_n13596));
  OAI221xp5_ASAP7_75t_L     g13340(.A1(new_n10280), .A2(new_n763), .B1(new_n695), .B2(new_n12010), .C(new_n13596), .Y(new_n13597));
  XNOR2x2_ASAP7_75t_L       g13341(.A(\a[56] ), .B(new_n13597), .Y(new_n13598));
  XOR2x2_ASAP7_75t_L        g13342(.A(new_n13598), .B(new_n13595), .Y(new_n13599));
  A2O1A1Ixp33_ASAP7_75t_L   g13343(.A1(new_n13357), .A2(new_n13328), .B(new_n13354), .C(new_n13599), .Y(new_n13600));
  NOR3xp33_ASAP7_75t_L      g13344(.A(new_n13354), .B(new_n13356), .C(new_n13327), .Y(new_n13601));
  OR3x1_ASAP7_75t_L         g13345(.A(new_n13599), .B(new_n13354), .C(new_n13601), .Y(new_n13602));
  AOI22xp33_ASAP7_75t_L     g13346(.A1(new_n8645), .A2(\b[16] ), .B1(new_n8642), .B2(new_n1058), .Y(new_n13603));
  OAI221xp5_ASAP7_75t_L     g13347(.A1(new_n9322), .A2(new_n952), .B1(new_n871), .B2(new_n8965), .C(new_n13603), .Y(new_n13604));
  XNOR2x2_ASAP7_75t_L       g13348(.A(\a[53] ), .B(new_n13604), .Y(new_n13605));
  NAND3xp33_ASAP7_75t_L     g13349(.A(new_n13600), .B(new_n13602), .C(new_n13605), .Y(new_n13606));
  AO21x2_ASAP7_75t_L        g13350(.A1(new_n13600), .A2(new_n13602), .B(new_n13605), .Y(new_n13607));
  OAI211xp5_ASAP7_75t_L     g13351(.A1(new_n13361), .A2(new_n13365), .B(new_n13607), .C(new_n13606), .Y(new_n13608));
  AO221x2_ASAP7_75t_L       g13352(.A1(new_n13360), .A2(new_n13358), .B1(new_n13607), .B2(new_n13606), .C(new_n13365), .Y(new_n13609));
  NAND2xp33_ASAP7_75t_L     g13353(.A(\b[19] ), .B(new_n7659), .Y(new_n13610));
  OAI221xp5_ASAP7_75t_L     g13354(.A1(new_n1356), .A2(new_n8326), .B1(new_n7996), .B2(new_n2793), .C(new_n13610), .Y(new_n13611));
  AOI21xp33_ASAP7_75t_L     g13355(.A1(new_n7993), .A2(\b[17] ), .B(new_n13611), .Y(new_n13612));
  NAND2xp33_ASAP7_75t_L     g13356(.A(\a[50] ), .B(new_n13612), .Y(new_n13613));
  A2O1A1Ixp33_ASAP7_75t_L   g13357(.A1(\b[17] ), .A2(new_n7993), .B(new_n13611), .C(new_n7653), .Y(new_n13614));
  AND2x2_ASAP7_75t_L        g13358(.A(new_n13614), .B(new_n13613), .Y(new_n13615));
  NAND3xp33_ASAP7_75t_L     g13359(.A(new_n13609), .B(new_n13608), .C(new_n13615), .Y(new_n13616));
  NAND2xp33_ASAP7_75t_L     g13360(.A(new_n13608), .B(new_n13609), .Y(new_n13617));
  INVx1_ASAP7_75t_L         g13361(.A(new_n13615), .Y(new_n13618));
  NAND2xp33_ASAP7_75t_L     g13362(.A(new_n13618), .B(new_n13617), .Y(new_n13619));
  NAND2xp33_ASAP7_75t_L     g13363(.A(new_n13369), .B(new_n13374), .Y(new_n13620));
  NAND3xp33_ASAP7_75t_L     g13364(.A(new_n13619), .B(new_n13616), .C(new_n13620), .Y(new_n13621));
  NAND2xp33_ASAP7_75t_L     g13365(.A(new_n13616), .B(new_n13619), .Y(new_n13622));
  NAND3xp33_ASAP7_75t_L     g13366(.A(new_n13622), .B(new_n13374), .C(new_n13369), .Y(new_n13623));
  AOI22xp33_ASAP7_75t_L     g13367(.A1(new_n6822), .A2(\b[22] ), .B1(new_n6819), .B2(new_n1864), .Y(new_n13624));
  OAI221xp5_ASAP7_75t_L     g13368(.A1(new_n7392), .A2(new_n1709), .B1(new_n1594), .B2(new_n7115), .C(new_n13624), .Y(new_n13625));
  XNOR2x2_ASAP7_75t_L       g13369(.A(\a[47] ), .B(new_n13625), .Y(new_n13626));
  NAND3xp33_ASAP7_75t_L     g13370(.A(new_n13623), .B(new_n13621), .C(new_n13626), .Y(new_n13627));
  AO21x2_ASAP7_75t_L        g13371(.A1(new_n13621), .A2(new_n13623), .B(new_n13626), .Y(new_n13628));
  NAND2xp33_ASAP7_75t_L     g13372(.A(new_n13627), .B(new_n13628), .Y(new_n13629));
  AOI21xp33_ASAP7_75t_L     g13373(.A1(new_n13385), .A2(new_n13386), .B(new_n13380), .Y(new_n13630));
  XOR2x2_ASAP7_75t_L        g13374(.A(new_n13630), .B(new_n13629), .Y(new_n13631));
  NOR2xp33_ASAP7_75t_L      g13375(.A(new_n13571), .B(new_n13631), .Y(new_n13632));
  NAND2xp33_ASAP7_75t_L     g13376(.A(new_n13571), .B(new_n13631), .Y(new_n13633));
  INVx1_ASAP7_75t_L         g13377(.A(new_n13633), .Y(new_n13634));
  A2O1A1Ixp33_ASAP7_75t_L   g13378(.A1(new_n13387), .A2(new_n13384), .B(new_n13392), .C(new_n13398), .Y(new_n13635));
  OA21x2_ASAP7_75t_L        g13379(.A1(new_n13632), .A2(new_n13634), .B(new_n13635), .Y(new_n13636));
  NOR3xp33_ASAP7_75t_L      g13380(.A(new_n13634), .B(new_n13635), .C(new_n13632), .Y(new_n13637));
  AOI22xp33_ASAP7_75t_L     g13381(.A1(new_n5249), .A2(\b[28] ), .B1(new_n5247), .B2(new_n2858), .Y(new_n13638));
  OAI221xp5_ASAP7_75t_L     g13382(.A1(new_n5241), .A2(new_n2650), .B1(new_n2477), .B2(new_n5521), .C(new_n13638), .Y(new_n13639));
  XNOR2x2_ASAP7_75t_L       g13383(.A(\a[41] ), .B(new_n13639), .Y(new_n13640));
  INVx1_ASAP7_75t_L         g13384(.A(new_n13640), .Y(new_n13641));
  NOR3xp33_ASAP7_75t_L      g13385(.A(new_n13636), .B(new_n13637), .C(new_n13641), .Y(new_n13642));
  OA21x2_ASAP7_75t_L        g13386(.A1(new_n13637), .A2(new_n13636), .B(new_n13641), .Y(new_n13643));
  AOI21xp33_ASAP7_75t_L     g13387(.A1(new_n13403), .A2(new_n13406), .B(new_n13401), .Y(new_n13644));
  NOR3xp33_ASAP7_75t_L      g13388(.A(new_n13643), .B(new_n13644), .C(new_n13642), .Y(new_n13645));
  OAI21xp33_ASAP7_75t_L     g13389(.A1(new_n13642), .A2(new_n13643), .B(new_n13644), .Y(new_n13646));
  INVx1_ASAP7_75t_L         g13390(.A(new_n13646), .Y(new_n13647));
  AOI22xp33_ASAP7_75t_L     g13391(.A1(new_n4544), .A2(\b[31] ), .B1(new_n4542), .B2(new_n3426), .Y(new_n13648));
  OAI221xp5_ASAP7_75t_L     g13392(.A1(new_n4536), .A2(new_n3212), .B1(new_n2871), .B2(new_n4781), .C(new_n13648), .Y(new_n13649));
  XNOR2x2_ASAP7_75t_L       g13393(.A(\a[38] ), .B(new_n13649), .Y(new_n13650));
  OAI21xp33_ASAP7_75t_L     g13394(.A1(new_n13645), .A2(new_n13647), .B(new_n13650), .Y(new_n13651));
  INVx1_ASAP7_75t_L         g13395(.A(new_n13645), .Y(new_n13652));
  INVx1_ASAP7_75t_L         g13396(.A(new_n13650), .Y(new_n13653));
  NAND3xp33_ASAP7_75t_L     g13397(.A(new_n13652), .B(new_n13646), .C(new_n13653), .Y(new_n13654));
  NAND3xp33_ASAP7_75t_L     g13398(.A(new_n13568), .B(new_n13651), .C(new_n13654), .Y(new_n13655));
  AOI21xp33_ASAP7_75t_L     g13399(.A1(new_n13654), .A2(new_n13651), .B(new_n13568), .Y(new_n13656));
  INVx1_ASAP7_75t_L         g13400(.A(new_n13656), .Y(new_n13657));
  AO21x2_ASAP7_75t_L        g13401(.A1(new_n13655), .A2(new_n13657), .B(new_n13567), .Y(new_n13658));
  NAND3xp33_ASAP7_75t_L     g13402(.A(new_n13657), .B(new_n13655), .C(new_n13567), .Y(new_n13659));
  NAND3xp33_ASAP7_75t_L     g13403(.A(new_n13564), .B(new_n13658), .C(new_n13659), .Y(new_n13660));
  AO21x2_ASAP7_75t_L        g13404(.A1(new_n13659), .A2(new_n13658), .B(new_n13564), .Y(new_n13661));
  NAND2xp33_ASAP7_75t_L     g13405(.A(new_n13660), .B(new_n13661), .Y(new_n13662));
  NOR2xp33_ASAP7_75t_L      g13406(.A(new_n13441), .B(new_n13433), .Y(new_n13663));
  AOI22xp33_ASAP7_75t_L     g13407(.A1(new_n2706), .A2(\b[39] ), .B1(\b[40] ), .B2(new_n2702), .Y(new_n13664));
  OAI221xp5_ASAP7_75t_L     g13408(.A1(new_n2932), .A2(new_n4915), .B1(new_n2707), .B2(new_n11823), .C(new_n13664), .Y(new_n13665));
  XNOR2x2_ASAP7_75t_L       g13409(.A(\a[29] ), .B(new_n13665), .Y(new_n13666));
  A2O1A1Ixp33_ASAP7_75t_L   g13410(.A1(new_n13440), .A2(new_n13438), .B(new_n13663), .C(new_n13666), .Y(new_n13667));
  AOI21xp33_ASAP7_75t_L     g13411(.A1(new_n13117), .A2(new_n13118), .B(new_n13119), .Y(new_n13668));
  O2A1O1Ixp33_ASAP7_75t_L   g13412(.A1(new_n13668), .A2(new_n12980), .B(new_n13120), .C(new_n13437), .Y(new_n13669));
  NOR3xp33_ASAP7_75t_L      g13413(.A(new_n13663), .B(new_n13669), .C(new_n13666), .Y(new_n13670));
  INVx1_ASAP7_75t_L         g13414(.A(new_n13670), .Y(new_n13671));
  AO21x2_ASAP7_75t_L        g13415(.A1(new_n13667), .A2(new_n13671), .B(new_n13662), .Y(new_n13672));
  NAND3xp33_ASAP7_75t_L     g13416(.A(new_n13671), .B(new_n13667), .C(new_n13662), .Y(new_n13673));
  NAND2xp33_ASAP7_75t_L     g13417(.A(new_n13673), .B(new_n13672), .Y(new_n13674));
  XNOR2x2_ASAP7_75t_L       g13418(.A(new_n13558), .B(new_n13674), .Y(new_n13675));
  NAND3xp33_ASAP7_75t_L     g13419(.A(new_n13675), .B(new_n13548), .C(new_n13549), .Y(new_n13676));
  NAND2xp33_ASAP7_75t_L     g13420(.A(new_n13549), .B(new_n13548), .Y(new_n13677));
  INVx1_ASAP7_75t_L         g13421(.A(new_n13675), .Y(new_n13678));
  NAND2xp33_ASAP7_75t_L     g13422(.A(new_n13678), .B(new_n13677), .Y(new_n13679));
  NAND3xp33_ASAP7_75t_L     g13423(.A(new_n13542), .B(new_n13676), .C(new_n13679), .Y(new_n13680));
  AO21x2_ASAP7_75t_L        g13424(.A1(new_n13679), .A2(new_n13676), .B(new_n13542), .Y(new_n13681));
  NAND2xp33_ASAP7_75t_L     g13425(.A(new_n13680), .B(new_n13681), .Y(new_n13682));
  AOI22xp33_ASAP7_75t_L     g13426(.A1(new_n1113), .A2(\b[52] ), .B1(new_n1110), .B2(new_n8577), .Y(new_n13683));
  OAI221xp5_ASAP7_75t_L     g13427(.A1(new_n1298), .A2(new_n8249), .B1(new_n8228), .B2(new_n1195), .C(new_n13683), .Y(new_n13684));
  XNOR2x2_ASAP7_75t_L       g13428(.A(new_n1107), .B(new_n13684), .Y(new_n13685));
  NOR2xp33_ASAP7_75t_L      g13429(.A(new_n13300), .B(new_n13450), .Y(new_n13686));
  NAND2xp33_ASAP7_75t_L     g13430(.A(new_n13685), .B(new_n13686), .Y(new_n13687));
  INVx1_ASAP7_75t_L         g13431(.A(new_n13687), .Y(new_n13688));
  O2A1O1Ixp33_ASAP7_75t_L   g13432(.A1(new_n13302), .A2(new_n13449), .B(new_n13301), .C(new_n13685), .Y(new_n13689));
  OAI21xp33_ASAP7_75t_L     g13433(.A1(new_n13689), .A2(new_n13688), .B(new_n13682), .Y(new_n13690));
  AND2x2_ASAP7_75t_L        g13434(.A(new_n13680), .B(new_n13681), .Y(new_n13691));
  INVx1_ASAP7_75t_L         g13435(.A(new_n13689), .Y(new_n13692));
  NAND3xp33_ASAP7_75t_L     g13436(.A(new_n13691), .B(new_n13687), .C(new_n13692), .Y(new_n13693));
  NAND2xp33_ASAP7_75t_L     g13437(.A(new_n13690), .B(new_n13693), .Y(new_n13694));
  NOR3xp33_ASAP7_75t_L      g13438(.A(new_n13694), .B(new_n13530), .C(new_n13529), .Y(new_n13695));
  OA21x2_ASAP7_75t_L        g13439(.A1(new_n13530), .A2(new_n13529), .B(new_n13694), .Y(new_n13696));
  NOR2xp33_ASAP7_75t_L      g13440(.A(new_n13695), .B(new_n13696), .Y(new_n13697));
  XNOR2x2_ASAP7_75t_L       g13441(.A(new_n13697), .B(new_n13523), .Y(new_n13698));
  AOI22xp33_ASAP7_75t_L     g13442(.A1(new_n441), .A2(\b[60] ), .B1(\b[61] ), .B2(new_n451), .Y(new_n13699));
  OAI221xp5_ASAP7_75t_L     g13443(.A1(new_n481), .A2(new_n10881), .B1(new_n482), .B2(new_n11920), .C(new_n13699), .Y(new_n13700));
  XNOR2x2_ASAP7_75t_L       g13444(.A(\a[8] ), .B(new_n13700), .Y(new_n13701));
  NOR3xp33_ASAP7_75t_L      g13445(.A(new_n13475), .B(new_n13701), .C(new_n13462), .Y(new_n13702));
  A2O1A1Ixp33_ASAP7_75t_L   g13446(.A1(new_n13277), .A2(new_n13458), .B(new_n13462), .C(new_n13701), .Y(new_n13703));
  INVx1_ASAP7_75t_L         g13447(.A(new_n13703), .Y(new_n13704));
  NOR3xp33_ASAP7_75t_L      g13448(.A(new_n13702), .B(new_n13704), .C(new_n13698), .Y(new_n13705));
  INVx1_ASAP7_75t_L         g13449(.A(new_n13705), .Y(new_n13706));
  OAI21xp33_ASAP7_75t_L     g13450(.A1(new_n13704), .A2(new_n13702), .B(new_n13698), .Y(new_n13707));
  NAND2xp33_ASAP7_75t_L     g13451(.A(new_n13707), .B(new_n13706), .Y(new_n13708));
  AOI21xp33_ASAP7_75t_L     g13452(.A1(new_n13516), .A2(new_n13513), .B(new_n13708), .Y(new_n13709));
  NAND2xp33_ASAP7_75t_L     g13453(.A(new_n13513), .B(new_n13516), .Y(new_n13710));
  INVx1_ASAP7_75t_L         g13454(.A(new_n13707), .Y(new_n13711));
  NOR2xp33_ASAP7_75t_L      g13455(.A(new_n13705), .B(new_n13711), .Y(new_n13712));
  NOR2xp33_ASAP7_75t_L      g13456(.A(new_n13710), .B(new_n13712), .Y(new_n13713));
  NOR3xp33_ASAP7_75t_L      g13457(.A(new_n13505), .B(new_n13709), .C(new_n13713), .Y(new_n13714));
  OA21x2_ASAP7_75t_L        g13458(.A1(new_n13713), .A2(new_n13709), .B(new_n13505), .Y(new_n13715));
  NOR2xp33_ASAP7_75t_L      g13459(.A(new_n13714), .B(new_n13715), .Y(new_n13716));
  INVx1_ASAP7_75t_L         g13460(.A(new_n13716), .Y(new_n13717));
  O2A1O1Ixp33_ASAP7_75t_L   g13461(.A1(new_n13499), .A2(new_n13504), .B(new_n13498), .C(new_n13717), .Y(new_n13718));
  A2O1A1Ixp33_ASAP7_75t_L   g13462(.A1(new_n13263), .A2(new_n13501), .B(new_n13499), .C(new_n13498), .Y(new_n13719));
  NOR2xp33_ASAP7_75t_L      g13463(.A(new_n13716), .B(new_n13719), .Y(new_n13720));
  NOR2xp33_ASAP7_75t_L      g13464(.A(new_n13720), .B(new_n13718), .Y(\f[67] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g13465(.A1(new_n13464), .A2(new_n13459), .B(new_n13472), .C(new_n13471), .D(new_n13512), .Y(new_n13722));
  INVx1_ASAP7_75t_L         g13466(.A(new_n13722), .Y(new_n13723));
  A2O1A1Ixp33_ASAP7_75t_L   g13467(.A1(new_n13516), .A2(new_n13513), .B(new_n13708), .C(new_n13723), .Y(new_n13724));
  A2O1A1O1Ixp25_ASAP7_75t_L g13468(.A1(new_n13286), .A2(new_n13283), .B(new_n13517), .C(new_n13518), .D(new_n13522), .Y(new_n13725));
  AOI22xp33_ASAP7_75t_L     g13469(.A1(new_n441), .A2(\b[61] ), .B1(\b[62] ), .B2(new_n451), .Y(new_n13726));
  OAI221xp5_ASAP7_75t_L     g13470(.A1(new_n481), .A2(new_n11226), .B1(new_n482), .B2(new_n12281), .C(new_n13726), .Y(new_n13727));
  XNOR2x2_ASAP7_75t_L       g13471(.A(\a[8] ), .B(new_n13727), .Y(new_n13728));
  A2O1A1Ixp33_ASAP7_75t_L   g13472(.A1(new_n13523), .A2(new_n13697), .B(new_n13725), .C(new_n13728), .Y(new_n13729));
  AOI211xp5_ASAP7_75t_L     g13473(.A1(new_n13523), .A2(new_n13697), .B(new_n13725), .C(new_n13728), .Y(new_n13730));
  INVx1_ASAP7_75t_L         g13474(.A(new_n13730), .Y(new_n13731));
  AOI22xp33_ASAP7_75t_L     g13475(.A1(new_n600), .A2(\b[59] ), .B1(new_n597), .B2(new_n10887), .Y(new_n13732));
  OAI221xp5_ASAP7_75t_L     g13476(.A1(new_n721), .A2(new_n10848), .B1(new_n10488), .B2(new_n1620), .C(new_n13732), .Y(new_n13733));
  XNOR2x2_ASAP7_75t_L       g13477(.A(\a[11] ), .B(new_n13733), .Y(new_n13734));
  MAJIxp5_ASAP7_75t_L       g13478(.A(new_n13694), .B(new_n13526), .C(new_n13528), .Y(new_n13735));
  INVx1_ASAP7_75t_L         g13479(.A(new_n13735), .Y(new_n13736));
  NAND2xp33_ASAP7_75t_L     g13480(.A(new_n13734), .B(new_n13736), .Y(new_n13737));
  INVx1_ASAP7_75t_L         g13481(.A(new_n13734), .Y(new_n13738));
  NAND2xp33_ASAP7_75t_L     g13482(.A(new_n13738), .B(new_n13735), .Y(new_n13739));
  AOI22xp33_ASAP7_75t_L     g13483(.A1(new_n826), .A2(\b[56] ), .B1(new_n823), .B2(new_n10185), .Y(new_n13740));
  OAI221xp5_ASAP7_75t_L     g13484(.A1(new_n994), .A2(new_n9534), .B1(new_n9199), .B2(new_n909), .C(new_n13740), .Y(new_n13741));
  INVx1_ASAP7_75t_L         g13485(.A(new_n13741), .Y(new_n13742));
  NAND2xp33_ASAP7_75t_L     g13486(.A(\a[14] ), .B(new_n13742), .Y(new_n13743));
  NAND2xp33_ASAP7_75t_L     g13487(.A(new_n813), .B(new_n13741), .Y(new_n13744));
  NAND2xp33_ASAP7_75t_L     g13488(.A(new_n13744), .B(new_n13743), .Y(new_n13745));
  INVx1_ASAP7_75t_L         g13489(.A(new_n13685), .Y(new_n13746));
  O2A1O1Ixp33_ASAP7_75t_L   g13490(.A1(new_n13302), .A2(new_n13449), .B(new_n13301), .C(new_n13746), .Y(new_n13747));
  O2A1O1Ixp33_ASAP7_75t_L   g13491(.A1(new_n13689), .A2(new_n13688), .B(new_n13682), .C(new_n13747), .Y(new_n13748));
  NAND2xp33_ASAP7_75t_L     g13492(.A(new_n13745), .B(new_n13748), .Y(new_n13749));
  INVx1_ASAP7_75t_L         g13493(.A(new_n13747), .Y(new_n13750));
  A2O1A1O1Ixp25_ASAP7_75t_L g13494(.A1(new_n13687), .A2(new_n13692), .B(new_n13691), .C(new_n13750), .D(new_n13745), .Y(new_n13751));
  INVx1_ASAP7_75t_L         g13495(.A(new_n13751), .Y(new_n13752));
  AOI22xp33_ASAP7_75t_L     g13496(.A1(new_n1103), .A2(\b[52] ), .B1(\b[53] ), .B2(new_n1113), .Y(new_n13753));
  OAI221xp5_ASAP7_75t_L     g13497(.A1(new_n1195), .A2(new_n8249), .B1(new_n1197), .B2(new_n8888), .C(new_n13753), .Y(new_n13754));
  XNOR2x2_ASAP7_75t_L       g13498(.A(\a[17] ), .B(new_n13754), .Y(new_n13755));
  INVx1_ASAP7_75t_L         g13499(.A(new_n13755), .Y(new_n13756));
  AOI31xp33_ASAP7_75t_L     g13500(.A1(new_n13542), .A2(new_n13676), .A3(new_n13679), .B(new_n13540), .Y(new_n13757));
  NAND2xp33_ASAP7_75t_L     g13501(.A(new_n13756), .B(new_n13757), .Y(new_n13758));
  O2A1O1Ixp33_ASAP7_75t_L   g13502(.A1(new_n13534), .A2(new_n13539), .B(new_n13680), .C(new_n13756), .Y(new_n13759));
  INVx1_ASAP7_75t_L         g13503(.A(new_n13759), .Y(new_n13760));
  OAI22xp33_ASAP7_75t_L     g13504(.A1(new_n8234), .A2(new_n1411), .B1(new_n8228), .B2(new_n1412), .Y(new_n13761));
  AOI221xp5_ASAP7_75t_L     g13505(.A1(\b[48] ), .A2(new_n1548), .B1(\b[49] ), .B2(new_n1410), .C(new_n13761), .Y(new_n13762));
  AND2x2_ASAP7_75t_L        g13506(.A(\a[20] ), .B(new_n13762), .Y(new_n13763));
  NOR2xp33_ASAP7_75t_L      g13507(.A(\a[20] ), .B(new_n13762), .Y(new_n13764));
  NOR2xp33_ASAP7_75t_L      g13508(.A(new_n13764), .B(new_n13763), .Y(new_n13765));
  A2O1A1Ixp33_ASAP7_75t_L   g13509(.A1(new_n13447), .A2(new_n13317), .B(new_n13316), .C(new_n13546), .Y(new_n13766));
  A2O1A1Ixp33_ASAP7_75t_L   g13510(.A1(new_n13549), .A2(new_n13548), .B(new_n13678), .C(new_n13766), .Y(new_n13767));
  NOR2xp33_ASAP7_75t_L      g13511(.A(new_n13765), .B(new_n13767), .Y(new_n13768));
  INVx1_ASAP7_75t_L         g13512(.A(new_n13766), .Y(new_n13769));
  A2O1A1Ixp33_ASAP7_75t_L   g13513(.A1(new_n13677), .A2(new_n13675), .B(new_n13769), .C(new_n13765), .Y(new_n13770));
  INVx1_ASAP7_75t_L         g13514(.A(new_n13770), .Y(new_n13771));
  INVx1_ASAP7_75t_L         g13515(.A(new_n13557), .Y(new_n13772));
  AOI22xp33_ASAP7_75t_L     g13516(.A1(new_n1766), .A2(\b[47] ), .B1(new_n1764), .B2(new_n7323), .Y(new_n13773));
  OAI221xp5_ASAP7_75t_L     g13517(.A1(new_n1758), .A2(new_n7033), .B1(new_n6756), .B2(new_n1911), .C(new_n13773), .Y(new_n13774));
  XNOR2x2_ASAP7_75t_L       g13518(.A(\a[23] ), .B(new_n13774), .Y(new_n13775));
  OAI211xp5_ASAP7_75t_L     g13519(.A1(new_n13556), .A2(new_n13674), .B(new_n13775), .C(new_n13772), .Y(new_n13776));
  O2A1O1Ixp33_ASAP7_75t_L   g13520(.A1(new_n13556), .A2(new_n13674), .B(new_n13772), .C(new_n13775), .Y(new_n13777));
  INVx1_ASAP7_75t_L         g13521(.A(new_n13777), .Y(new_n13778));
  AOI22xp33_ASAP7_75t_L     g13522(.A1(new_n2702), .A2(\b[41] ), .B1(new_n2700), .B2(new_n5669), .Y(new_n13779));
  OAI221xp5_ASAP7_75t_L     g13523(.A1(new_n2694), .A2(new_n5186), .B1(new_n5166), .B2(new_n2932), .C(new_n13779), .Y(new_n13780));
  XNOR2x2_ASAP7_75t_L       g13524(.A(\a[29] ), .B(new_n13780), .Y(new_n13781));
  INVx1_ASAP7_75t_L         g13525(.A(new_n13781), .Y(new_n13782));
  NAND2xp33_ASAP7_75t_L     g13526(.A(new_n13562), .B(new_n13563), .Y(new_n13783));
  O2A1O1Ixp33_ASAP7_75t_L   g13527(.A1(new_n13429), .A2(new_n13424), .B(new_n13431), .C(new_n13562), .Y(new_n13784));
  A2O1A1Ixp33_ASAP7_75t_L   g13528(.A1(new_n13658), .A2(new_n13659), .B(new_n13784), .C(new_n13783), .Y(new_n13785));
  NOR2xp33_ASAP7_75t_L      g13529(.A(new_n13782), .B(new_n13785), .Y(new_n13786));
  A2O1A1O1Ixp25_ASAP7_75t_L g13530(.A1(new_n13659), .A2(new_n13658), .B(new_n13784), .C(new_n13783), .D(new_n13781), .Y(new_n13787));
  NOR2xp33_ASAP7_75t_L      g13531(.A(new_n13787), .B(new_n13786), .Y(new_n13788));
  AOI22xp33_ASAP7_75t_L     g13532(.A1(new_n8645), .A2(\b[17] ), .B1(new_n8642), .B2(new_n1252), .Y(new_n13789));
  OAI221xp5_ASAP7_75t_L     g13533(.A1(new_n9322), .A2(new_n1051), .B1(new_n952), .B2(new_n8965), .C(new_n13789), .Y(new_n13790));
  XNOR2x2_ASAP7_75t_L       g13534(.A(\a[53] ), .B(new_n13790), .Y(new_n13791));
  INVx1_ASAP7_75t_L         g13535(.A(new_n13791), .Y(new_n13792));
  NOR2xp33_ASAP7_75t_L      g13536(.A(new_n382), .B(new_n13003), .Y(new_n13793));
  NAND2xp33_ASAP7_75t_L     g13537(.A(\b[8] ), .B(new_n11656), .Y(new_n13794));
  OAI221xp5_ASAP7_75t_L     g13538(.A1(new_n421), .A2(new_n12364), .B1(new_n12022), .B2(new_n509), .C(new_n13794), .Y(new_n13795));
  OR3x1_ASAP7_75t_L         g13539(.A(new_n13795), .B(new_n11651), .C(new_n13793), .Y(new_n13796));
  A2O1A1Ixp33_ASAP7_75t_L   g13540(.A1(\b[6] ), .A2(new_n12021), .B(new_n13795), .C(new_n11651), .Y(new_n13797));
  NAND2xp33_ASAP7_75t_L     g13541(.A(new_n13797), .B(new_n13796), .Y(new_n13798));
  NOR2xp33_ASAP7_75t_L      g13542(.A(new_n323), .B(new_n12671), .Y(new_n13799));
  O2A1O1Ixp33_ASAP7_75t_L   g13543(.A1(new_n12353), .A2(new_n12355), .B(\b[5] ), .C(new_n13799), .Y(new_n13800));
  NAND2xp33_ASAP7_75t_L     g13544(.A(\a[2] ), .B(new_n13800), .Y(new_n13801));
  INVx1_ASAP7_75t_L         g13545(.A(new_n13801), .Y(new_n13802));
  INVx1_ASAP7_75t_L         g13546(.A(new_n13799), .Y(new_n13803));
  O2A1O1Ixp33_ASAP7_75t_L   g13547(.A1(new_n353), .A2(new_n12356), .B(new_n13803), .C(\a[2] ), .Y(new_n13804));
  NOR2xp33_ASAP7_75t_L      g13548(.A(new_n13804), .B(new_n13802), .Y(new_n13805));
  XNOR2x2_ASAP7_75t_L       g13549(.A(new_n13805), .B(new_n13798), .Y(new_n13806));
  A2O1A1Ixp33_ASAP7_75t_L   g13550(.A1(new_n12669), .A2(\b[4] ), .B(new_n13575), .C(\a[2] ), .Y(new_n13807));
  A2O1A1Ixp33_ASAP7_75t_L   g13551(.A1(new_n13577), .A2(new_n13578), .B(new_n13574), .C(new_n13807), .Y(new_n13808));
  XNOR2x2_ASAP7_75t_L       g13552(.A(new_n13808), .B(new_n13806), .Y(new_n13809));
  AOI22xp33_ASAP7_75t_L     g13553(.A1(new_n10594), .A2(\b[11] ), .B1(new_n10591), .B2(new_n702), .Y(new_n13810));
  OAI221xp5_ASAP7_75t_L     g13554(.A1(new_n11335), .A2(new_n631), .B1(new_n559), .B2(new_n11330), .C(new_n13810), .Y(new_n13811));
  XNOR2x2_ASAP7_75t_L       g13555(.A(new_n10588), .B(new_n13811), .Y(new_n13812));
  INVx1_ASAP7_75t_L         g13556(.A(new_n13812), .Y(new_n13813));
  NAND2xp33_ASAP7_75t_L     g13557(.A(new_n13809), .B(new_n13813), .Y(new_n13814));
  NOR2xp33_ASAP7_75t_L      g13558(.A(new_n13809), .B(new_n13813), .Y(new_n13815));
  INVx1_ASAP7_75t_L         g13559(.A(new_n13815), .Y(new_n13816));
  AND2x2_ASAP7_75t_L        g13560(.A(new_n13814), .B(new_n13816), .Y(new_n13817));
  NAND3xp33_ASAP7_75t_L     g13561(.A(new_n13817), .B(new_n13588), .C(new_n13582), .Y(new_n13818));
  INVx1_ASAP7_75t_L         g13562(.A(new_n13582), .Y(new_n13819));
  INVx1_ASAP7_75t_L         g13563(.A(new_n13817), .Y(new_n13820));
  A2O1A1Ixp33_ASAP7_75t_L   g13564(.A1(new_n13584), .A2(new_n13587), .B(new_n13819), .C(new_n13820), .Y(new_n13821));
  AOI22xp33_ASAP7_75t_L     g13565(.A1(new_n9623), .A2(\b[14] ), .B1(new_n9620), .B2(new_n879), .Y(new_n13822));
  OAI221xp5_ASAP7_75t_L     g13566(.A1(new_n10280), .A2(new_n793), .B1(new_n763), .B2(new_n12010), .C(new_n13822), .Y(new_n13823));
  XNOR2x2_ASAP7_75t_L       g13567(.A(\a[56] ), .B(new_n13823), .Y(new_n13824));
  NAND3xp33_ASAP7_75t_L     g13568(.A(new_n13821), .B(new_n13818), .C(new_n13824), .Y(new_n13825));
  AO21x2_ASAP7_75t_L        g13569(.A1(new_n13818), .A2(new_n13821), .B(new_n13824), .Y(new_n13826));
  NAND2xp33_ASAP7_75t_L     g13570(.A(new_n13825), .B(new_n13826), .Y(new_n13827));
  OA21x2_ASAP7_75t_L        g13571(.A1(new_n13598), .A2(new_n13595), .B(new_n13594), .Y(new_n13828));
  XNOR2x2_ASAP7_75t_L       g13572(.A(new_n13828), .B(new_n13827), .Y(new_n13829));
  XNOR2x2_ASAP7_75t_L       g13573(.A(new_n13792), .B(new_n13829), .Y(new_n13830));
  NAND2xp33_ASAP7_75t_L     g13574(.A(new_n13602), .B(new_n13606), .Y(new_n13831));
  XNOR2x2_ASAP7_75t_L       g13575(.A(new_n13831), .B(new_n13830), .Y(new_n13832));
  AOI22xp33_ASAP7_75t_L     g13576(.A1(new_n7659), .A2(\b[20] ), .B1(new_n7656), .B2(new_n1600), .Y(new_n13833));
  OAI221xp5_ASAP7_75t_L     g13577(.A1(new_n8326), .A2(new_n1493), .B1(new_n1356), .B2(new_n7994), .C(new_n13833), .Y(new_n13834));
  XNOR2x2_ASAP7_75t_L       g13578(.A(\a[50] ), .B(new_n13834), .Y(new_n13835));
  XOR2x2_ASAP7_75t_L        g13579(.A(new_n13835), .B(new_n13832), .Y(new_n13836));
  NAND2xp33_ASAP7_75t_L     g13580(.A(new_n13608), .B(new_n13616), .Y(new_n13837));
  XNOR2x2_ASAP7_75t_L       g13581(.A(new_n13837), .B(new_n13836), .Y(new_n13838));
  AOI22xp33_ASAP7_75t_L     g13582(.A1(new_n6822), .A2(\b[23] ), .B1(new_n6819), .B2(new_n2002), .Y(new_n13839));
  OAI221xp5_ASAP7_75t_L     g13583(.A1(new_n7392), .A2(new_n1857), .B1(new_n1709), .B2(new_n7115), .C(new_n13839), .Y(new_n13840));
  XNOR2x2_ASAP7_75t_L       g13584(.A(\a[47] ), .B(new_n13840), .Y(new_n13841));
  XNOR2x2_ASAP7_75t_L       g13585(.A(new_n13841), .B(new_n13838), .Y(new_n13842));
  A2O1A1Ixp33_ASAP7_75t_L   g13586(.A1(new_n13374), .A2(new_n13369), .B(new_n13622), .C(new_n13627), .Y(new_n13843));
  XNOR2x2_ASAP7_75t_L       g13587(.A(new_n13843), .B(new_n13842), .Y(new_n13844));
  AOI22xp33_ASAP7_75t_L     g13588(.A1(new_n6002), .A2(\b[26] ), .B1(new_n5999), .B2(new_n2888), .Y(new_n13845));
  OAI221xp5_ASAP7_75t_L     g13589(.A1(new_n6544), .A2(new_n2180), .B1(new_n2019), .B2(new_n6309), .C(new_n13845), .Y(new_n13846));
  XNOR2x2_ASAP7_75t_L       g13590(.A(\a[44] ), .B(new_n13846), .Y(new_n13847));
  XOR2x2_ASAP7_75t_L        g13591(.A(new_n13847), .B(new_n13844), .Y(new_n13848));
  A2O1A1O1Ixp25_ASAP7_75t_L g13592(.A1(new_n13385), .A2(new_n13386), .B(new_n13380), .C(new_n13629), .D(new_n13632), .Y(new_n13849));
  NAND2xp33_ASAP7_75t_L     g13593(.A(new_n13849), .B(new_n13848), .Y(new_n13850));
  INVx1_ASAP7_75t_L         g13594(.A(new_n13630), .Y(new_n13851));
  XNOR2x2_ASAP7_75t_L       g13595(.A(new_n13847), .B(new_n13844), .Y(new_n13852));
  A2O1A1Ixp33_ASAP7_75t_L   g13596(.A1(new_n13851), .A2(new_n13629), .B(new_n13632), .C(new_n13852), .Y(new_n13853));
  NAND2xp33_ASAP7_75t_L     g13597(.A(new_n13850), .B(new_n13853), .Y(new_n13854));
  AOI22xp33_ASAP7_75t_L     g13598(.A1(new_n5249), .A2(\b[29] ), .B1(new_n5247), .B2(new_n5472), .Y(new_n13855));
  OAI221xp5_ASAP7_75t_L     g13599(.A1(new_n5241), .A2(new_n2852), .B1(new_n2650), .B2(new_n5521), .C(new_n13855), .Y(new_n13856));
  XNOR2x2_ASAP7_75t_L       g13600(.A(\a[41] ), .B(new_n13856), .Y(new_n13857));
  INVx1_ASAP7_75t_L         g13601(.A(new_n13857), .Y(new_n13858));
  NOR2xp33_ASAP7_75t_L      g13602(.A(new_n13858), .B(new_n13854), .Y(new_n13859));
  XNOR2x2_ASAP7_75t_L       g13603(.A(new_n13849), .B(new_n13852), .Y(new_n13860));
  NOR2xp33_ASAP7_75t_L      g13604(.A(new_n13857), .B(new_n13860), .Y(new_n13861));
  O2A1O1Ixp33_ASAP7_75t_L   g13605(.A1(new_n13632), .A2(new_n13634), .B(new_n13635), .C(new_n13642), .Y(new_n13862));
  NOR3xp33_ASAP7_75t_L      g13606(.A(new_n13859), .B(new_n13861), .C(new_n13862), .Y(new_n13863));
  NAND2xp33_ASAP7_75t_L     g13607(.A(new_n13857), .B(new_n13860), .Y(new_n13864));
  NAND2xp33_ASAP7_75t_L     g13608(.A(new_n13858), .B(new_n13854), .Y(new_n13865));
  INVx1_ASAP7_75t_L         g13609(.A(new_n13862), .Y(new_n13866));
  AOI21xp33_ASAP7_75t_L     g13610(.A1(new_n13865), .A2(new_n13864), .B(new_n13866), .Y(new_n13867));
  AOI22xp33_ASAP7_75t_L     g13611(.A1(new_n4544), .A2(\b[32] ), .B1(new_n4542), .B2(new_n3450), .Y(new_n13868));
  OAI221xp5_ASAP7_75t_L     g13612(.A1(new_n4536), .A2(new_n3419), .B1(new_n3212), .B2(new_n4781), .C(new_n13868), .Y(new_n13869));
  XNOR2x2_ASAP7_75t_L       g13613(.A(\a[38] ), .B(new_n13869), .Y(new_n13870));
  OAI21xp33_ASAP7_75t_L     g13614(.A1(new_n13867), .A2(new_n13863), .B(new_n13870), .Y(new_n13871));
  NAND3xp33_ASAP7_75t_L     g13615(.A(new_n13865), .B(new_n13864), .C(new_n13866), .Y(new_n13872));
  OAI21xp33_ASAP7_75t_L     g13616(.A1(new_n13861), .A2(new_n13859), .B(new_n13862), .Y(new_n13873));
  INVx1_ASAP7_75t_L         g13617(.A(new_n13870), .Y(new_n13874));
  NAND3xp33_ASAP7_75t_L     g13618(.A(new_n13873), .B(new_n13872), .C(new_n13874), .Y(new_n13875));
  NAND2xp33_ASAP7_75t_L     g13619(.A(new_n13646), .B(new_n13654), .Y(new_n13876));
  NAND3xp33_ASAP7_75t_L     g13620(.A(new_n13871), .B(new_n13875), .C(new_n13876), .Y(new_n13877));
  AOI21xp33_ASAP7_75t_L     g13621(.A1(new_n13873), .A2(new_n13872), .B(new_n13874), .Y(new_n13878));
  NOR3xp33_ASAP7_75t_L      g13622(.A(new_n13863), .B(new_n13867), .C(new_n13870), .Y(new_n13879));
  INVx1_ASAP7_75t_L         g13623(.A(new_n13876), .Y(new_n13880));
  OAI21xp33_ASAP7_75t_L     g13624(.A1(new_n13878), .A2(new_n13879), .B(new_n13880), .Y(new_n13881));
  AOI22xp33_ASAP7_75t_L     g13625(.A1(new_n3884), .A2(\b[35] ), .B1(new_n3881), .B2(new_n5649), .Y(new_n13882));
  OAI221xp5_ASAP7_75t_L     g13626(.A1(new_n4312), .A2(new_n3827), .B1(new_n3807), .B2(new_n4986), .C(new_n13882), .Y(new_n13883));
  XNOR2x2_ASAP7_75t_L       g13627(.A(\a[35] ), .B(new_n13883), .Y(new_n13884));
  AND3x1_ASAP7_75t_L        g13628(.A(new_n13881), .B(new_n13884), .C(new_n13877), .Y(new_n13885));
  AOI21xp33_ASAP7_75t_L     g13629(.A1(new_n13881), .A2(new_n13877), .B(new_n13884), .Y(new_n13886));
  NOR2xp33_ASAP7_75t_L      g13630(.A(new_n13886), .B(new_n13885), .Y(new_n13887));
  AOI22xp33_ASAP7_75t_L     g13631(.A1(new_n3260), .A2(\b[37] ), .B1(\b[38] ), .B2(new_n3256), .Y(new_n13888));
  OAI221xp5_ASAP7_75t_L     g13632(.A1(new_n3492), .A2(new_n4465), .B1(new_n3261), .B2(new_n8160), .C(new_n13888), .Y(new_n13889));
  XNOR2x2_ASAP7_75t_L       g13633(.A(\a[32] ), .B(new_n13889), .Y(new_n13890));
  AOI21xp33_ASAP7_75t_L     g13634(.A1(new_n13655), .A2(new_n13567), .B(new_n13656), .Y(new_n13891));
  XNOR2x2_ASAP7_75t_L       g13635(.A(new_n13890), .B(new_n13891), .Y(new_n13892));
  XNOR2x2_ASAP7_75t_L       g13636(.A(new_n13892), .B(new_n13887), .Y(new_n13893));
  XNOR2x2_ASAP7_75t_L       g13637(.A(new_n13893), .B(new_n13788), .Y(new_n13894));
  NOR2xp33_ASAP7_75t_L      g13638(.A(new_n13669), .B(new_n13663), .Y(new_n13895));
  MAJIxp5_ASAP7_75t_L       g13639(.A(new_n13662), .B(new_n13666), .C(new_n13895), .Y(new_n13896));
  AOI22xp33_ASAP7_75t_L     g13640(.A1(new_n2232), .A2(\b[43] ), .B1(\b[44] ), .B2(new_n2228), .Y(new_n13897));
  OAI221xp5_ASAP7_75t_L     g13641(.A1(new_n2387), .A2(new_n5680), .B1(new_n2233), .B2(new_n6229), .C(new_n13897), .Y(new_n13898));
  XNOR2x2_ASAP7_75t_L       g13642(.A(new_n2223), .B(new_n13898), .Y(new_n13899));
  XNOR2x2_ASAP7_75t_L       g13643(.A(new_n13899), .B(new_n13896), .Y(new_n13900));
  NOR2xp33_ASAP7_75t_L      g13644(.A(new_n13900), .B(new_n13894), .Y(new_n13901));
  AND2x2_ASAP7_75t_L        g13645(.A(new_n13900), .B(new_n13894), .Y(new_n13902));
  NOR2xp33_ASAP7_75t_L      g13646(.A(new_n13901), .B(new_n13902), .Y(new_n13903));
  NAND3xp33_ASAP7_75t_L     g13647(.A(new_n13903), .B(new_n13778), .C(new_n13776), .Y(new_n13904));
  AO21x2_ASAP7_75t_L        g13648(.A1(new_n13776), .A2(new_n13778), .B(new_n13903), .Y(new_n13905));
  NAND2xp33_ASAP7_75t_L     g13649(.A(new_n13904), .B(new_n13905), .Y(new_n13906));
  OAI21xp33_ASAP7_75t_L     g13650(.A1(new_n13768), .A2(new_n13771), .B(new_n13906), .Y(new_n13907));
  AOI21xp33_ASAP7_75t_L     g13651(.A1(new_n13677), .A2(new_n13675), .B(new_n13769), .Y(new_n13908));
  OAI21xp33_ASAP7_75t_L     g13652(.A1(new_n13763), .A2(new_n13764), .B(new_n13908), .Y(new_n13909));
  NAND2xp33_ASAP7_75t_L     g13653(.A(new_n13776), .B(new_n13778), .Y(new_n13910));
  XNOR2x2_ASAP7_75t_L       g13654(.A(new_n13903), .B(new_n13910), .Y(new_n13911));
  NAND3xp33_ASAP7_75t_L     g13655(.A(new_n13911), .B(new_n13770), .C(new_n13909), .Y(new_n13912));
  NAND2xp33_ASAP7_75t_L     g13656(.A(new_n13912), .B(new_n13907), .Y(new_n13913));
  INVx1_ASAP7_75t_L         g13657(.A(new_n13913), .Y(new_n13914));
  NAND3xp33_ASAP7_75t_L     g13658(.A(new_n13914), .B(new_n13760), .C(new_n13758), .Y(new_n13915));
  INVx1_ASAP7_75t_L         g13659(.A(new_n13758), .Y(new_n13916));
  OAI21xp33_ASAP7_75t_L     g13660(.A1(new_n13759), .A2(new_n13916), .B(new_n13913), .Y(new_n13917));
  AND2x2_ASAP7_75t_L        g13661(.A(new_n13917), .B(new_n13915), .Y(new_n13918));
  AOI21xp33_ASAP7_75t_L     g13662(.A1(new_n13752), .A2(new_n13749), .B(new_n13918), .Y(new_n13919));
  INVx1_ASAP7_75t_L         g13663(.A(new_n13745), .Y(new_n13920));
  A2O1A1Ixp33_ASAP7_75t_L   g13664(.A1(new_n13692), .A2(new_n13687), .B(new_n13691), .C(new_n13750), .Y(new_n13921));
  NOR2xp33_ASAP7_75t_L      g13665(.A(new_n13920), .B(new_n13921), .Y(new_n13922));
  NAND2xp33_ASAP7_75t_L     g13666(.A(new_n13917), .B(new_n13915), .Y(new_n13923));
  NOR3xp33_ASAP7_75t_L      g13667(.A(new_n13923), .B(new_n13751), .C(new_n13922), .Y(new_n13924));
  NOR2xp33_ASAP7_75t_L      g13668(.A(new_n13924), .B(new_n13919), .Y(new_n13925));
  NAND3xp33_ASAP7_75t_L     g13669(.A(new_n13737), .B(new_n13925), .C(new_n13739), .Y(new_n13926));
  AO21x2_ASAP7_75t_L        g13670(.A1(new_n13739), .A2(new_n13737), .B(new_n13925), .Y(new_n13927));
  NAND2xp33_ASAP7_75t_L     g13671(.A(new_n13926), .B(new_n13927), .Y(new_n13928));
  AO21x2_ASAP7_75t_L        g13672(.A1(new_n13729), .A2(new_n13731), .B(new_n13928), .Y(new_n13929));
  NAND3xp33_ASAP7_75t_L     g13673(.A(new_n13928), .B(new_n13731), .C(new_n13729), .Y(new_n13930));
  INVx1_ASAP7_75t_L         g13674(.A(new_n13698), .Y(new_n13931));
  A2O1A1Ixp33_ASAP7_75t_L   g13675(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n342), .Y(new_n13932));
  A2O1A1Ixp33_ASAP7_75t_L   g13676(.A1(new_n13932), .A2(new_n365), .B(new_n12599), .C(\a[5] ), .Y(new_n13933));
  O2A1O1Ixp33_ASAP7_75t_L   g13677(.A1(\b[60] ), .A2(new_n11916), .B(\b[61] ), .C(\b[62] ), .Y(new_n13934));
  O2A1O1Ixp33_ASAP7_75t_L   g13678(.A1(new_n367), .A2(new_n13934), .B(new_n365), .C(new_n12599), .Y(new_n13935));
  NAND2xp33_ASAP7_75t_L     g13679(.A(new_n339), .B(new_n13935), .Y(new_n13936));
  AND2x2_ASAP7_75t_L        g13680(.A(new_n13936), .B(new_n13933), .Y(new_n13937));
  INVx1_ASAP7_75t_L         g13681(.A(new_n13937), .Y(new_n13938));
  A2O1A1Ixp33_ASAP7_75t_L   g13682(.A1(new_n13931), .A2(new_n13703), .B(new_n13702), .C(new_n13938), .Y(new_n13939));
  INVx1_ASAP7_75t_L         g13683(.A(new_n13702), .Y(new_n13940));
  OAI211xp5_ASAP7_75t_L     g13684(.A1(new_n13698), .A2(new_n13704), .B(new_n13940), .C(new_n13937), .Y(new_n13941));
  NAND4xp25_ASAP7_75t_L     g13685(.A(new_n13941), .B(new_n13939), .C(new_n13929), .D(new_n13930), .Y(new_n13942));
  AO22x1_ASAP7_75t_L        g13686(.A1(new_n13929), .A2(new_n13930), .B1(new_n13939), .B2(new_n13941), .Y(new_n13943));
  NAND2xp33_ASAP7_75t_L     g13687(.A(new_n13942), .B(new_n13943), .Y(new_n13944));
  XNOR2x2_ASAP7_75t_L       g13688(.A(new_n13724), .B(new_n13944), .Y(new_n13945));
  A2O1A1Ixp33_ASAP7_75t_L   g13689(.A1(new_n13719), .A2(new_n13716), .B(new_n13714), .C(new_n13945), .Y(new_n13946));
  INVx1_ASAP7_75t_L         g13690(.A(new_n13946), .Y(new_n13947));
  NOR3xp33_ASAP7_75t_L      g13691(.A(new_n13718), .B(new_n13945), .C(new_n13714), .Y(new_n13948));
  NOR2xp33_ASAP7_75t_L      g13692(.A(new_n13947), .B(new_n13948), .Y(\f[68] ));
  INVx1_ASAP7_75t_L         g13693(.A(new_n13944), .Y(new_n13950));
  A2O1A1Ixp33_ASAP7_75t_L   g13694(.A1(new_n13706), .A2(new_n13940), .B(new_n13937), .C(new_n13942), .Y(new_n13951));
  INVx1_ASAP7_75t_L         g13695(.A(new_n13728), .Y(new_n13952));
  A2O1A1Ixp33_ASAP7_75t_L   g13696(.A1(new_n13523), .A2(new_n13697), .B(new_n13725), .C(new_n13952), .Y(new_n13953));
  NAND2xp33_ASAP7_75t_L     g13697(.A(\b[63] ), .B(new_n451), .Y(new_n13954));
  A2O1A1Ixp33_ASAP7_75t_L   g13698(.A1(new_n12607), .A2(new_n12603), .B(new_n482), .C(new_n13954), .Y(new_n13955));
  AOI221xp5_ASAP7_75t_L     g13699(.A1(\b[61] ), .A2(new_n480), .B1(\b[62] ), .B2(new_n441), .C(new_n13955), .Y(new_n13956));
  XNOR2x2_ASAP7_75t_L       g13700(.A(new_n445), .B(new_n13956), .Y(new_n13957));
  INVx1_ASAP7_75t_L         g13701(.A(new_n13957), .Y(new_n13958));
  A2O1A1O1Ixp25_ASAP7_75t_L g13702(.A1(new_n13731), .A2(new_n13729), .B(new_n13928), .C(new_n13953), .D(new_n13958), .Y(new_n13959));
  A2O1A1Ixp33_ASAP7_75t_L   g13703(.A1(new_n13731), .A2(new_n13729), .B(new_n13928), .C(new_n13953), .Y(new_n13960));
  NOR2xp33_ASAP7_75t_L      g13704(.A(new_n13957), .B(new_n13960), .Y(new_n13961));
  NOR2xp33_ASAP7_75t_L      g13705(.A(new_n13959), .B(new_n13961), .Y(new_n13962));
  INVx1_ASAP7_75t_L         g13706(.A(new_n13962), .Y(new_n13963));
  AOI22xp33_ASAP7_75t_L     g13707(.A1(new_n600), .A2(\b[60] ), .B1(new_n597), .B2(new_n11234), .Y(new_n13964));
  OAI221xp5_ASAP7_75t_L     g13708(.A1(new_n721), .A2(new_n10881), .B1(new_n10848), .B2(new_n1620), .C(new_n13964), .Y(new_n13965));
  XNOR2x2_ASAP7_75t_L       g13709(.A(\a[11] ), .B(new_n13965), .Y(new_n13966));
  AND3x1_ASAP7_75t_L        g13710(.A(new_n13737), .B(new_n13925), .C(new_n13739), .Y(new_n13967));
  O2A1O1Ixp33_ASAP7_75t_L   g13711(.A1(new_n13530), .A2(new_n13695), .B(new_n13738), .C(new_n13967), .Y(new_n13968));
  NAND2xp33_ASAP7_75t_L     g13712(.A(new_n13966), .B(new_n13968), .Y(new_n13969));
  O2A1O1Ixp33_ASAP7_75t_L   g13713(.A1(new_n13734), .A2(new_n13736), .B(new_n13926), .C(new_n13966), .Y(new_n13970));
  INVx1_ASAP7_75t_L         g13714(.A(new_n13970), .Y(new_n13971));
  NAND2xp33_ASAP7_75t_L     g13715(.A(new_n13971), .B(new_n13969), .Y(new_n13972));
  AOI22xp33_ASAP7_75t_L     g13716(.A1(new_n826), .A2(\b[57] ), .B1(new_n823), .B2(new_n10495), .Y(new_n13973));
  OAI221xp5_ASAP7_75t_L     g13717(.A1(new_n994), .A2(new_n10178), .B1(new_n9534), .B2(new_n909), .C(new_n13973), .Y(new_n13974));
  XNOR2x2_ASAP7_75t_L       g13718(.A(\a[14] ), .B(new_n13974), .Y(new_n13975));
  A2O1A1O1Ixp25_ASAP7_75t_L g13719(.A1(new_n13687), .A2(new_n13692), .B(new_n13691), .C(new_n13750), .D(new_n13920), .Y(new_n13976));
  INVx1_ASAP7_75t_L         g13720(.A(new_n13976), .Y(new_n13977));
  A2O1A1O1Ixp25_ASAP7_75t_L g13721(.A1(new_n13752), .A2(new_n13749), .B(new_n13918), .C(new_n13977), .D(new_n13975), .Y(new_n13978));
  INVx1_ASAP7_75t_L         g13722(.A(new_n13978), .Y(new_n13979));
  O2A1O1Ixp33_ASAP7_75t_L   g13723(.A1(new_n13751), .A2(new_n13922), .B(new_n13923), .C(new_n13976), .Y(new_n13980));
  NAND2xp33_ASAP7_75t_L     g13724(.A(new_n13975), .B(new_n13980), .Y(new_n13981));
  NAND2xp33_ASAP7_75t_L     g13725(.A(new_n1764), .B(new_n7341), .Y(new_n13982));
  OAI221xp5_ASAP7_75t_L     g13726(.A1(new_n1772), .A2(new_n7333), .B1(new_n7316), .B2(new_n1758), .C(new_n13982), .Y(new_n13983));
  AOI21xp33_ASAP7_75t_L     g13727(.A1(new_n1910), .A2(\b[46] ), .B(new_n13983), .Y(new_n13984));
  NAND2xp33_ASAP7_75t_L     g13728(.A(\a[23] ), .B(new_n13984), .Y(new_n13985));
  A2O1A1Ixp33_ASAP7_75t_L   g13729(.A1(\b[46] ), .A2(new_n1910), .B(new_n13983), .C(new_n1761), .Y(new_n13986));
  NAND2xp33_ASAP7_75t_L     g13730(.A(new_n13986), .B(new_n13985), .Y(new_n13987));
  AOI211xp5_ASAP7_75t_L     g13731(.A1(new_n13903), .A2(new_n13776), .B(new_n13987), .C(new_n13777), .Y(new_n13988));
  A2O1A1Ixp33_ASAP7_75t_L   g13732(.A1(new_n13903), .A2(new_n13776), .B(new_n13777), .C(new_n13987), .Y(new_n13989));
  INVx1_ASAP7_75t_L         g13733(.A(new_n13989), .Y(new_n13990));
  NOR2xp33_ASAP7_75t_L      g13734(.A(new_n13988), .B(new_n13990), .Y(new_n13991));
  AOI22xp33_ASAP7_75t_L     g13735(.A1(new_n2228), .A2(\b[45] ), .B1(new_n2226), .B2(new_n6764), .Y(new_n13992));
  OAI221xp5_ASAP7_75t_L     g13736(.A1(new_n2220), .A2(new_n6220), .B1(new_n6195), .B2(new_n2387), .C(new_n13992), .Y(new_n13993));
  XNOR2x2_ASAP7_75t_L       g13737(.A(\a[26] ), .B(new_n13993), .Y(new_n13994));
  A2O1A1Ixp33_ASAP7_75t_L   g13738(.A1(new_n13899), .A2(new_n13896), .B(new_n13901), .C(new_n13994), .Y(new_n13995));
  AOI21xp33_ASAP7_75t_L     g13739(.A1(new_n13899), .A2(new_n13896), .B(new_n13901), .Y(new_n13996));
  INVx1_ASAP7_75t_L         g13740(.A(new_n13994), .Y(new_n13997));
  NAND2xp33_ASAP7_75t_L     g13741(.A(new_n13997), .B(new_n13996), .Y(new_n13998));
  NAND2xp33_ASAP7_75t_L     g13742(.A(new_n13995), .B(new_n13998), .Y(new_n13999));
  AOI22xp33_ASAP7_75t_L     g13743(.A1(new_n2702), .A2(\b[42] ), .B1(new_n2700), .B2(new_n5688), .Y(new_n14000));
  OAI221xp5_ASAP7_75t_L     g13744(.A1(new_n2694), .A2(new_n5666), .B1(new_n5186), .B2(new_n2932), .C(new_n14000), .Y(new_n14001));
  XNOR2x2_ASAP7_75t_L       g13745(.A(\a[29] ), .B(new_n14001), .Y(new_n14002));
  MAJIxp5_ASAP7_75t_L       g13746(.A(new_n13893), .B(new_n13782), .C(new_n13785), .Y(new_n14003));
  NAND2xp33_ASAP7_75t_L     g13747(.A(new_n14002), .B(new_n14003), .Y(new_n14004));
  NOR2xp33_ASAP7_75t_L      g13748(.A(new_n14002), .B(new_n14003), .Y(new_n14005));
  INVx1_ASAP7_75t_L         g13749(.A(new_n14005), .Y(new_n14006));
  NAND2xp33_ASAP7_75t_L     g13750(.A(new_n14004), .B(new_n14006), .Y(new_n14007));
  AOI22xp33_ASAP7_75t_L     g13751(.A1(new_n3884), .A2(\b[36] ), .B1(new_n3881), .B2(new_n4473), .Y(new_n14008));
  OAI221xp5_ASAP7_75t_L     g13752(.A1(new_n4312), .A2(new_n4053), .B1(new_n3827), .B2(new_n4986), .C(new_n14008), .Y(new_n14009));
  XNOR2x2_ASAP7_75t_L       g13753(.A(\a[35] ), .B(new_n14009), .Y(new_n14010));
  O2A1O1Ixp33_ASAP7_75t_L   g13754(.A1(new_n13859), .A2(new_n13861), .B(new_n13862), .C(new_n13879), .Y(new_n14011));
  AOI22xp33_ASAP7_75t_L     g13755(.A1(new_n4544), .A2(\b[33] ), .B1(new_n4542), .B2(new_n3813), .Y(new_n14012));
  OAI221xp5_ASAP7_75t_L     g13756(.A1(new_n4536), .A2(new_n3443), .B1(new_n3419), .B2(new_n4781), .C(new_n14012), .Y(new_n14013));
  XNOR2x2_ASAP7_75t_L       g13757(.A(\a[38] ), .B(new_n14013), .Y(new_n14014));
  A2O1A1O1Ixp25_ASAP7_75t_L g13758(.A1(new_n13374), .A2(new_n13369), .B(new_n13622), .C(new_n13627), .D(new_n13842), .Y(new_n14015));
  AOI22xp33_ASAP7_75t_L     g13759(.A1(new_n6822), .A2(\b[24] ), .B1(new_n6819), .B2(new_n2027), .Y(new_n14016));
  OAI221xp5_ASAP7_75t_L     g13760(.A1(new_n7392), .A2(new_n1995), .B1(new_n1857), .B2(new_n7115), .C(new_n14016), .Y(new_n14017));
  XNOR2x2_ASAP7_75t_L       g13761(.A(new_n6816), .B(new_n14017), .Y(new_n14018));
  MAJx2_ASAP7_75t_L         g13762(.A(new_n13830), .B(new_n13831), .C(new_n13835), .Y(new_n14019));
  INVx1_ASAP7_75t_L         g13763(.A(new_n13827), .Y(new_n14020));
  NAND2xp33_ASAP7_75t_L     g13764(.A(new_n13828), .B(new_n14020), .Y(new_n14021));
  INVx1_ASAP7_75t_L         g13765(.A(new_n14021), .Y(new_n14022));
  INVx1_ASAP7_75t_L         g13766(.A(new_n13821), .Y(new_n14023));
  AOI22xp33_ASAP7_75t_L     g13767(.A1(new_n9623), .A2(\b[15] ), .B1(new_n9620), .B2(new_n959), .Y(new_n14024));
  OAI221xp5_ASAP7_75t_L     g13768(.A1(new_n10280), .A2(new_n871), .B1(new_n793), .B2(new_n12010), .C(new_n14024), .Y(new_n14025));
  XNOR2x2_ASAP7_75t_L       g13769(.A(\a[56] ), .B(new_n14025), .Y(new_n14026));
  INVx1_ASAP7_75t_L         g13770(.A(new_n14026), .Y(new_n14027));
  INVx1_ASAP7_75t_L         g13771(.A(new_n13576), .Y(new_n14028));
  NOR2xp33_ASAP7_75t_L      g13772(.A(new_n13579), .B(new_n13574), .Y(new_n14029));
  A2O1A1Ixp33_ASAP7_75t_L   g13773(.A1(\a[2] ), .A2(new_n14028), .B(new_n14029), .C(new_n13806), .Y(new_n14030));
  AOI22xp33_ASAP7_75t_L     g13774(.A1(new_n10594), .A2(\b[12] ), .B1(new_n10591), .B2(new_n970), .Y(new_n14031));
  OAI221xp5_ASAP7_75t_L     g13775(.A1(new_n11335), .A2(new_n695), .B1(new_n631), .B2(new_n11330), .C(new_n14031), .Y(new_n14032));
  XNOR2x2_ASAP7_75t_L       g13776(.A(\a[59] ), .B(new_n14032), .Y(new_n14033));
  O2A1O1Ixp33_ASAP7_75t_L   g13777(.A1(new_n353), .A2(new_n12356), .B(new_n13803), .C(new_n265), .Y(new_n14034));
  O2A1O1Ixp33_ASAP7_75t_L   g13778(.A1(new_n13802), .A2(new_n13804), .B(new_n13798), .C(new_n14034), .Y(new_n14035));
  NOR2xp33_ASAP7_75t_L      g13779(.A(new_n353), .B(new_n12671), .Y(new_n14036));
  INVx1_ASAP7_75t_L         g13780(.A(new_n14036), .Y(new_n14037));
  XNOR2x2_ASAP7_75t_L       g13781(.A(\a[5] ), .B(\a[2] ), .Y(new_n14038));
  O2A1O1Ixp33_ASAP7_75t_L   g13782(.A1(new_n382), .A2(new_n12356), .B(new_n14037), .C(new_n14038), .Y(new_n14039));
  INVx1_ASAP7_75t_L         g13783(.A(new_n14039), .Y(new_n14040));
  O2A1O1Ixp33_ASAP7_75t_L   g13784(.A1(new_n12353), .A2(new_n12355), .B(\b[6] ), .C(new_n14036), .Y(new_n14041));
  NAND2xp33_ASAP7_75t_L     g13785(.A(new_n14038), .B(new_n14041), .Y(new_n14042));
  AND2x2_ASAP7_75t_L        g13786(.A(new_n14042), .B(new_n14040), .Y(new_n14043));
  INVx1_ASAP7_75t_L         g13787(.A(new_n14043), .Y(new_n14044));
  NAND2xp33_ASAP7_75t_L     g13788(.A(new_n14044), .B(new_n14035), .Y(new_n14045));
  INVx1_ASAP7_75t_L         g13789(.A(new_n13805), .Y(new_n14046));
  A2O1A1Ixp33_ASAP7_75t_L   g13790(.A1(new_n13798), .A2(new_n14046), .B(new_n14034), .C(new_n14043), .Y(new_n14047));
  NAND2xp33_ASAP7_75t_L     g13791(.A(new_n14047), .B(new_n14045), .Y(new_n14048));
  AOI22xp33_ASAP7_75t_L     g13792(.A1(new_n11656), .A2(\b[9] ), .B1(new_n11654), .B2(new_n566), .Y(new_n14049));
  OAI221xp5_ASAP7_75t_L     g13793(.A1(new_n12364), .A2(new_n503), .B1(new_n421), .B2(new_n13003), .C(new_n14049), .Y(new_n14050));
  XNOR2x2_ASAP7_75t_L       g13794(.A(\a[62] ), .B(new_n14050), .Y(new_n14051));
  AND2x2_ASAP7_75t_L        g13795(.A(new_n14051), .B(new_n14048), .Y(new_n14052));
  NOR2xp33_ASAP7_75t_L      g13796(.A(new_n14051), .B(new_n14048), .Y(new_n14053));
  NOR2xp33_ASAP7_75t_L      g13797(.A(new_n14053), .B(new_n14052), .Y(new_n14054));
  XNOR2x2_ASAP7_75t_L       g13798(.A(new_n14033), .B(new_n14054), .Y(new_n14055));
  INVx1_ASAP7_75t_L         g13799(.A(new_n14055), .Y(new_n14056));
  O2A1O1Ixp33_ASAP7_75t_L   g13800(.A1(new_n13809), .A2(new_n13813), .B(new_n14030), .C(new_n14056), .Y(new_n14057));
  AOI211xp5_ASAP7_75t_L     g13801(.A1(new_n13806), .A2(new_n13808), .B(new_n13815), .C(new_n14055), .Y(new_n14058));
  NOR2xp33_ASAP7_75t_L      g13802(.A(new_n14057), .B(new_n14058), .Y(new_n14059));
  XNOR2x2_ASAP7_75t_L       g13803(.A(new_n14027), .B(new_n14059), .Y(new_n14060));
  A2O1A1Ixp33_ASAP7_75t_L   g13804(.A1(new_n13824), .A2(new_n13818), .B(new_n14023), .C(new_n14060), .Y(new_n14061));
  A2O1A1Ixp33_ASAP7_75t_L   g13805(.A1(new_n13588), .A2(new_n13582), .B(new_n13817), .C(new_n13825), .Y(new_n14062));
  NOR2xp33_ASAP7_75t_L      g13806(.A(new_n14062), .B(new_n14060), .Y(new_n14063));
  INVx1_ASAP7_75t_L         g13807(.A(new_n14063), .Y(new_n14064));
  NAND2xp33_ASAP7_75t_L     g13808(.A(new_n14064), .B(new_n14061), .Y(new_n14065));
  AOI22xp33_ASAP7_75t_L     g13809(.A1(new_n8645), .A2(\b[18] ), .B1(new_n8642), .B2(new_n1363), .Y(new_n14066));
  OAI221xp5_ASAP7_75t_L     g13810(.A1(new_n9322), .A2(new_n1244), .B1(new_n1051), .B2(new_n8965), .C(new_n14066), .Y(new_n14067));
  XNOR2x2_ASAP7_75t_L       g13811(.A(\a[53] ), .B(new_n14067), .Y(new_n14068));
  XNOR2x2_ASAP7_75t_L       g13812(.A(new_n14068), .B(new_n14065), .Y(new_n14069));
  A2O1A1Ixp33_ASAP7_75t_L   g13813(.A1(new_n13829), .A2(new_n13791), .B(new_n14022), .C(new_n14069), .Y(new_n14070));
  O2A1O1Ixp33_ASAP7_75t_L   g13814(.A1(new_n13595), .A2(new_n13598), .B(new_n13594), .C(new_n14020), .Y(new_n14071));
  XOR2x2_ASAP7_75t_L        g13815(.A(new_n14068), .B(new_n14065), .Y(new_n14072));
  OAI211xp5_ASAP7_75t_L     g13816(.A1(new_n13792), .A2(new_n14071), .B(new_n14072), .C(new_n14021), .Y(new_n14073));
  AND2x2_ASAP7_75t_L        g13817(.A(new_n14070), .B(new_n14073), .Y(new_n14074));
  AOI22xp33_ASAP7_75t_L     g13818(.A1(new_n7659), .A2(\b[21] ), .B1(new_n7656), .B2(new_n1715), .Y(new_n14075));
  OAI221xp5_ASAP7_75t_L     g13819(.A1(new_n8326), .A2(new_n1594), .B1(new_n1493), .B2(new_n7994), .C(new_n14075), .Y(new_n14076));
  XNOR2x2_ASAP7_75t_L       g13820(.A(\a[50] ), .B(new_n14076), .Y(new_n14077));
  NAND2xp33_ASAP7_75t_L     g13821(.A(new_n14077), .B(new_n14074), .Y(new_n14078));
  NAND2xp33_ASAP7_75t_L     g13822(.A(new_n14070), .B(new_n14073), .Y(new_n14079));
  INVx1_ASAP7_75t_L         g13823(.A(new_n14077), .Y(new_n14080));
  NAND2xp33_ASAP7_75t_L     g13824(.A(new_n14080), .B(new_n14079), .Y(new_n14081));
  AOI21xp33_ASAP7_75t_L     g13825(.A1(new_n14078), .A2(new_n14081), .B(new_n14019), .Y(new_n14082));
  AND3x1_ASAP7_75t_L        g13826(.A(new_n14078), .B(new_n14081), .C(new_n14019), .Y(new_n14083));
  NOR2xp33_ASAP7_75t_L      g13827(.A(new_n14082), .B(new_n14083), .Y(new_n14084));
  XOR2x2_ASAP7_75t_L        g13828(.A(new_n14018), .B(new_n14084), .Y(new_n14085));
  O2A1O1Ixp33_ASAP7_75t_L   g13829(.A1(new_n13617), .A2(new_n13618), .B(new_n13608), .C(new_n13836), .Y(new_n14086));
  AOI21xp33_ASAP7_75t_L     g13830(.A1(new_n13838), .A2(new_n13841), .B(new_n14086), .Y(new_n14087));
  XNOR2x2_ASAP7_75t_L       g13831(.A(new_n14087), .B(new_n14085), .Y(new_n14088));
  AOI22xp33_ASAP7_75t_L     g13832(.A1(new_n6002), .A2(\b[27] ), .B1(new_n5999), .B2(new_n2657), .Y(new_n14089));
  OAI221xp5_ASAP7_75t_L     g13833(.A1(new_n6544), .A2(new_n2477), .B1(new_n2180), .B2(new_n6309), .C(new_n14089), .Y(new_n14090));
  XNOR2x2_ASAP7_75t_L       g13834(.A(\a[44] ), .B(new_n14090), .Y(new_n14091));
  XNOR2x2_ASAP7_75t_L       g13835(.A(new_n14091), .B(new_n14088), .Y(new_n14092));
  A2O1A1Ixp33_ASAP7_75t_L   g13836(.A1(new_n13844), .A2(new_n13847), .B(new_n14015), .C(new_n14092), .Y(new_n14093));
  NAND2xp33_ASAP7_75t_L     g13837(.A(new_n13847), .B(new_n13844), .Y(new_n14094));
  A2O1A1Ixp33_ASAP7_75t_L   g13838(.A1(new_n13627), .A2(new_n13621), .B(new_n13842), .C(new_n14094), .Y(new_n14095));
  OR2x4_ASAP7_75t_L         g13839(.A(new_n14095), .B(new_n14092), .Y(new_n14096));
  NAND2xp33_ASAP7_75t_L     g13840(.A(new_n14093), .B(new_n14096), .Y(new_n14097));
  AOI22xp33_ASAP7_75t_L     g13841(.A1(new_n5249), .A2(\b[30] ), .B1(new_n5247), .B2(new_n3219), .Y(new_n14098));
  OAI221xp5_ASAP7_75t_L     g13842(.A1(new_n5241), .A2(new_n2871), .B1(new_n2852), .B2(new_n5521), .C(new_n14098), .Y(new_n14099));
  XNOR2x2_ASAP7_75t_L       g13843(.A(\a[41] ), .B(new_n14099), .Y(new_n14100));
  INVx1_ASAP7_75t_L         g13844(.A(new_n14100), .Y(new_n14101));
  XNOR2x2_ASAP7_75t_L       g13845(.A(new_n14101), .B(new_n14097), .Y(new_n14102));
  NAND3xp33_ASAP7_75t_L     g13846(.A(new_n14102), .B(new_n13864), .C(new_n13850), .Y(new_n14103));
  AND2x2_ASAP7_75t_L        g13847(.A(new_n14093), .B(new_n14096), .Y(new_n14104));
  NAND2xp33_ASAP7_75t_L     g13848(.A(new_n14101), .B(new_n14104), .Y(new_n14105));
  NAND2xp33_ASAP7_75t_L     g13849(.A(new_n14100), .B(new_n14097), .Y(new_n14106));
  NAND2xp33_ASAP7_75t_L     g13850(.A(new_n14106), .B(new_n14105), .Y(new_n14107));
  A2O1A1Ixp33_ASAP7_75t_L   g13851(.A1(new_n13849), .A2(new_n13848), .B(new_n13859), .C(new_n14107), .Y(new_n14108));
  NAND3xp33_ASAP7_75t_L     g13852(.A(new_n14108), .B(new_n14103), .C(new_n14014), .Y(new_n14109));
  INVx1_ASAP7_75t_L         g13853(.A(new_n14014), .Y(new_n14110));
  NAND2xp33_ASAP7_75t_L     g13854(.A(new_n13850), .B(new_n13864), .Y(new_n14111));
  NOR2xp33_ASAP7_75t_L      g13855(.A(new_n14111), .B(new_n14107), .Y(new_n14112));
  O2A1O1Ixp33_ASAP7_75t_L   g13856(.A1(new_n13854), .A2(new_n13858), .B(new_n13850), .C(new_n14102), .Y(new_n14113));
  OAI21xp33_ASAP7_75t_L     g13857(.A1(new_n14113), .A2(new_n14112), .B(new_n14110), .Y(new_n14114));
  AOI21xp33_ASAP7_75t_L     g13858(.A1(new_n14109), .A2(new_n14114), .B(new_n14011), .Y(new_n14115));
  INVx1_ASAP7_75t_L         g13859(.A(new_n14011), .Y(new_n14116));
  NOR3xp33_ASAP7_75t_L      g13860(.A(new_n14112), .B(new_n14113), .C(new_n14110), .Y(new_n14117));
  AOI21xp33_ASAP7_75t_L     g13861(.A1(new_n14108), .A2(new_n14103), .B(new_n14014), .Y(new_n14118));
  NOR3xp33_ASAP7_75t_L      g13862(.A(new_n14118), .B(new_n14117), .C(new_n14116), .Y(new_n14119));
  NOR3xp33_ASAP7_75t_L      g13863(.A(new_n14119), .B(new_n14115), .C(new_n14010), .Y(new_n14120));
  INVx1_ASAP7_75t_L         g13864(.A(new_n14010), .Y(new_n14121));
  OAI21xp33_ASAP7_75t_L     g13865(.A1(new_n14117), .A2(new_n14118), .B(new_n14116), .Y(new_n14122));
  NAND3xp33_ASAP7_75t_L     g13866(.A(new_n14109), .B(new_n14114), .C(new_n14011), .Y(new_n14123));
  AOI21xp33_ASAP7_75t_L     g13867(.A1(new_n14122), .A2(new_n14123), .B(new_n14121), .Y(new_n14124));
  NOR3xp33_ASAP7_75t_L      g13868(.A(new_n13879), .B(new_n13880), .C(new_n13878), .Y(new_n14125));
  INVx1_ASAP7_75t_L         g13869(.A(new_n13884), .Y(new_n14126));
  OAI21xp33_ASAP7_75t_L     g13870(.A1(new_n14126), .A2(new_n14125), .B(new_n13881), .Y(new_n14127));
  OAI21xp33_ASAP7_75t_L     g13871(.A1(new_n14124), .A2(new_n14120), .B(new_n14127), .Y(new_n14128));
  NAND3xp33_ASAP7_75t_L     g13872(.A(new_n14122), .B(new_n14123), .C(new_n14121), .Y(new_n14129));
  OAI21xp33_ASAP7_75t_L     g13873(.A1(new_n14115), .A2(new_n14119), .B(new_n14010), .Y(new_n14130));
  INVx1_ASAP7_75t_L         g13874(.A(new_n14127), .Y(new_n14131));
  NAND3xp33_ASAP7_75t_L     g13875(.A(new_n14130), .B(new_n14129), .C(new_n14131), .Y(new_n14132));
  NAND2xp33_ASAP7_75t_L     g13876(.A(new_n14132), .B(new_n14128), .Y(new_n14133));
  AOI22xp33_ASAP7_75t_L     g13877(.A1(new_n3256), .A2(\b[39] ), .B1(new_n3254), .B2(new_n5174), .Y(new_n14134));
  OAI221xp5_ASAP7_75t_L     g13878(.A1(new_n3248), .A2(new_n4915), .B1(new_n4701), .B2(new_n3492), .C(new_n14134), .Y(new_n14135));
  XNOR2x2_ASAP7_75t_L       g13879(.A(\a[32] ), .B(new_n14135), .Y(new_n14136));
  INVx1_ASAP7_75t_L         g13880(.A(new_n13890), .Y(new_n14137));
  NAND2xp33_ASAP7_75t_L     g13881(.A(new_n13892), .B(new_n13887), .Y(new_n14138));
  A2O1A1Ixp33_ASAP7_75t_L   g13882(.A1(new_n13659), .A2(new_n13657), .B(new_n14137), .C(new_n14138), .Y(new_n14139));
  XNOR2x2_ASAP7_75t_L       g13883(.A(new_n14136), .B(new_n14139), .Y(new_n14140));
  XNOR2x2_ASAP7_75t_L       g13884(.A(new_n14133), .B(new_n14140), .Y(new_n14141));
  XNOR2x2_ASAP7_75t_L       g13885(.A(new_n14007), .B(new_n14141), .Y(new_n14142));
  XOR2x2_ASAP7_75t_L        g13886(.A(new_n13999), .B(new_n14142), .Y(new_n14143));
  XNOR2x2_ASAP7_75t_L       g13887(.A(new_n13991), .B(new_n14143), .Y(new_n14144));
  NAND2xp33_ASAP7_75t_L     g13888(.A(new_n13770), .B(new_n13909), .Y(new_n14145));
  AOI22xp33_ASAP7_75t_L     g13889(.A1(new_n1406), .A2(\b[51] ), .B1(new_n1404), .B2(new_n8257), .Y(new_n14146));
  OAI221xp5_ASAP7_75t_L     g13890(.A1(new_n1398), .A2(new_n8228), .B1(new_n7907), .B2(new_n1549), .C(new_n14146), .Y(new_n14147));
  XNOR2x2_ASAP7_75t_L       g13891(.A(\a[20] ), .B(new_n14147), .Y(new_n14148));
  INVx1_ASAP7_75t_L         g13892(.A(new_n14148), .Y(new_n14149));
  A2O1A1O1Ixp25_ASAP7_75t_L g13893(.A1(new_n13549), .A2(new_n13548), .B(new_n13678), .C(new_n13766), .D(new_n13765), .Y(new_n14150));
  A2O1A1Ixp33_ASAP7_75t_L   g13894(.A1(new_n14145), .A2(new_n13911), .B(new_n14150), .C(new_n14149), .Y(new_n14151));
  INVx1_ASAP7_75t_L         g13895(.A(new_n14150), .Y(new_n14152));
  A2O1A1Ixp33_ASAP7_75t_L   g13896(.A1(new_n13770), .A2(new_n13909), .B(new_n13906), .C(new_n14152), .Y(new_n14153));
  NOR2xp33_ASAP7_75t_L      g13897(.A(new_n14149), .B(new_n14153), .Y(new_n14154));
  INVx1_ASAP7_75t_L         g13898(.A(new_n14154), .Y(new_n14155));
  NAND2xp33_ASAP7_75t_L     g13899(.A(new_n14151), .B(new_n14155), .Y(new_n14156));
  XOR2x2_ASAP7_75t_L        g13900(.A(new_n14144), .B(new_n14156), .Y(new_n14157));
  AOI22xp33_ASAP7_75t_L     g13901(.A1(new_n1113), .A2(\b[54] ), .B1(new_n1110), .B2(new_n9208), .Y(new_n14158));
  OAI221xp5_ASAP7_75t_L     g13902(.A1(new_n1298), .A2(new_n8882), .B1(new_n8569), .B2(new_n1195), .C(new_n14158), .Y(new_n14159));
  XNOR2x2_ASAP7_75t_L       g13903(.A(\a[17] ), .B(new_n14159), .Y(new_n14160));
  NAND2xp33_ASAP7_75t_L     g13904(.A(new_n13760), .B(new_n13915), .Y(new_n14161));
  NOR2xp33_ASAP7_75t_L      g13905(.A(new_n14160), .B(new_n14161), .Y(new_n14162));
  A2O1A1Ixp33_ASAP7_75t_L   g13906(.A1(new_n13914), .A2(new_n13758), .B(new_n13759), .C(new_n14160), .Y(new_n14163));
  INVx1_ASAP7_75t_L         g13907(.A(new_n14163), .Y(new_n14164));
  NOR3xp33_ASAP7_75t_L      g13908(.A(new_n14157), .B(new_n14162), .C(new_n14164), .Y(new_n14165));
  XNOR2x2_ASAP7_75t_L       g13909(.A(new_n14144), .B(new_n14156), .Y(new_n14166));
  OR2x4_ASAP7_75t_L         g13910(.A(new_n14160), .B(new_n14161), .Y(new_n14167));
  AOI21xp33_ASAP7_75t_L     g13911(.A1(new_n14167), .A2(new_n14163), .B(new_n14166), .Y(new_n14168));
  NOR2xp33_ASAP7_75t_L      g13912(.A(new_n14165), .B(new_n14168), .Y(new_n14169));
  NAND3xp33_ASAP7_75t_L     g13913(.A(new_n14169), .B(new_n13981), .C(new_n13979), .Y(new_n14170));
  NAND2xp33_ASAP7_75t_L     g13914(.A(new_n13981), .B(new_n13979), .Y(new_n14171));
  INVx1_ASAP7_75t_L         g13915(.A(new_n14169), .Y(new_n14172));
  NAND2xp33_ASAP7_75t_L     g13916(.A(new_n14171), .B(new_n14172), .Y(new_n14173));
  AND2x2_ASAP7_75t_L        g13917(.A(new_n14170), .B(new_n14173), .Y(new_n14174));
  XNOR2x2_ASAP7_75t_L       g13918(.A(new_n14174), .B(new_n13972), .Y(new_n14175));
  NAND2xp33_ASAP7_75t_L     g13919(.A(new_n13963), .B(new_n14175), .Y(new_n14176));
  NOR2xp33_ASAP7_75t_L      g13920(.A(new_n14174), .B(new_n13972), .Y(new_n14177));
  AND2x2_ASAP7_75t_L        g13921(.A(new_n14174), .B(new_n13972), .Y(new_n14178));
  OR4x2_ASAP7_75t_L         g13922(.A(new_n14178), .B(new_n14177), .C(new_n13961), .D(new_n13959), .Y(new_n14179));
  NAND3xp33_ASAP7_75t_L     g13923(.A(new_n14179), .B(new_n14176), .C(new_n13951), .Y(new_n14180));
  AO21x2_ASAP7_75t_L        g13924(.A1(new_n14176), .A2(new_n14179), .B(new_n13951), .Y(new_n14181));
  NAND2xp33_ASAP7_75t_L     g13925(.A(new_n14180), .B(new_n14181), .Y(new_n14182));
  INVx1_ASAP7_75t_L         g13926(.A(new_n14182), .Y(new_n14183));
  A2O1A1Ixp33_ASAP7_75t_L   g13927(.A1(new_n13950), .A2(new_n13724), .B(new_n13947), .C(new_n14183), .Y(new_n14184));
  A2O1A1Ixp33_ASAP7_75t_L   g13928(.A1(new_n13712), .A2(new_n13710), .B(new_n13722), .C(new_n13950), .Y(new_n14185));
  INVx1_ASAP7_75t_L         g13929(.A(new_n14185), .Y(new_n14186));
  A2O1A1O1Ixp25_ASAP7_75t_L g13930(.A1(new_n13719), .A2(new_n13716), .B(new_n13714), .C(new_n13945), .D(new_n14186), .Y(new_n14187));
  NAND2xp33_ASAP7_75t_L     g13931(.A(new_n14182), .B(new_n14187), .Y(new_n14188));
  AND2x2_ASAP7_75t_L        g13932(.A(new_n14188), .B(new_n14184), .Y(\f[69] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13933(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n448), .Y(new_n14190));
  AOI22xp33_ASAP7_75t_L     g13934(.A1(new_n441), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n480), .Y(new_n14191));
  NAND3xp33_ASAP7_75t_L     g13935(.A(new_n14190), .B(\a[8] ), .C(new_n14191), .Y(new_n14192));
  A2O1A1O1Ixp25_ASAP7_75t_L g13936(.A1(new_n13507), .A2(new_n13506), .B(new_n482), .C(new_n14191), .D(\a[8] ), .Y(new_n14193));
  INVx1_ASAP7_75t_L         g13937(.A(new_n14193), .Y(new_n14194));
  AND2x2_ASAP7_75t_L        g13938(.A(new_n14192), .B(new_n14194), .Y(new_n14195));
  INVx1_ASAP7_75t_L         g13939(.A(new_n14195), .Y(new_n14196));
  OAI211xp5_ASAP7_75t_L     g13940(.A1(new_n13970), .A2(new_n14174), .B(new_n13969), .C(new_n14196), .Y(new_n14197));
  A2O1A1O1Ixp25_ASAP7_75t_L g13941(.A1(new_n14173), .A2(new_n14170), .B(new_n13970), .C(new_n13969), .D(new_n14196), .Y(new_n14198));
  INVx1_ASAP7_75t_L         g13942(.A(new_n14198), .Y(new_n14199));
  AOI22xp33_ASAP7_75t_L     g13943(.A1(new_n600), .A2(\b[61] ), .B1(new_n597), .B2(new_n11919), .Y(new_n14200));
  OAI221xp5_ASAP7_75t_L     g13944(.A1(new_n721), .A2(new_n11226), .B1(new_n10881), .B2(new_n1620), .C(new_n14200), .Y(new_n14201));
  XNOR2x2_ASAP7_75t_L       g13945(.A(\a[11] ), .B(new_n14201), .Y(new_n14202));
  AOI21xp33_ASAP7_75t_L     g13946(.A1(new_n14169), .A2(new_n13981), .B(new_n13978), .Y(new_n14203));
  NAND2xp33_ASAP7_75t_L     g13947(.A(new_n14202), .B(new_n14203), .Y(new_n14204));
  O2A1O1Ixp33_ASAP7_75t_L   g13948(.A1(new_n14171), .A2(new_n14172), .B(new_n13979), .C(new_n14202), .Y(new_n14205));
  INVx1_ASAP7_75t_L         g13949(.A(new_n14205), .Y(new_n14206));
  AOI22xp33_ASAP7_75t_L     g13950(.A1(new_n817), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n826), .Y(new_n14207));
  OAI221xp5_ASAP7_75t_L     g13951(.A1(new_n909), .A2(new_n10178), .B1(new_n911), .B2(new_n10856), .C(new_n14207), .Y(new_n14208));
  XNOR2x2_ASAP7_75t_L       g13952(.A(\a[14] ), .B(new_n14208), .Y(new_n14209));
  INVx1_ASAP7_75t_L         g13953(.A(new_n14209), .Y(new_n14210));
  A2O1A1Ixp33_ASAP7_75t_L   g13954(.A1(new_n14166), .A2(new_n14163), .B(new_n14162), .C(new_n14210), .Y(new_n14211));
  OAI211xp5_ASAP7_75t_L     g13955(.A1(new_n14164), .A2(new_n14157), .B(new_n14167), .C(new_n14209), .Y(new_n14212));
  NAND2xp33_ASAP7_75t_L     g13956(.A(new_n14211), .B(new_n14212), .Y(new_n14213));
  A2O1A1O1Ixp25_ASAP7_75t_L g13957(.A1(new_n13770), .A2(new_n13909), .B(new_n13906), .C(new_n14152), .D(new_n14148), .Y(new_n14214));
  AOI22xp33_ASAP7_75t_L     g13958(.A1(new_n1113), .A2(\b[55] ), .B1(new_n1110), .B2(new_n9542), .Y(new_n14215));
  OAI221xp5_ASAP7_75t_L     g13959(.A1(new_n1298), .A2(new_n9199), .B1(new_n8882), .B2(new_n1195), .C(new_n14215), .Y(new_n14216));
  XNOR2x2_ASAP7_75t_L       g13960(.A(\a[17] ), .B(new_n14216), .Y(new_n14217));
  INVx1_ASAP7_75t_L         g13961(.A(new_n14217), .Y(new_n14218));
  O2A1O1Ixp33_ASAP7_75t_L   g13962(.A1(new_n14214), .A2(new_n14144), .B(new_n14155), .C(new_n14218), .Y(new_n14219));
  OA211x2_ASAP7_75t_L       g13963(.A1(new_n14214), .A2(new_n14144), .B(new_n14218), .C(new_n14155), .Y(new_n14220));
  NOR2xp33_ASAP7_75t_L      g13964(.A(new_n14219), .B(new_n14220), .Y(new_n14221));
  AOI22xp33_ASAP7_75t_L     g13965(.A1(new_n1406), .A2(\b[52] ), .B1(new_n1404), .B2(new_n8577), .Y(new_n14222));
  OAI221xp5_ASAP7_75t_L     g13966(.A1(new_n1398), .A2(new_n8249), .B1(new_n8228), .B2(new_n1549), .C(new_n14222), .Y(new_n14223));
  XNOR2x2_ASAP7_75t_L       g13967(.A(new_n1401), .B(new_n14223), .Y(new_n14224));
  AOI21xp33_ASAP7_75t_L     g13968(.A1(new_n14143), .A2(new_n13989), .B(new_n13988), .Y(new_n14225));
  XOR2x2_ASAP7_75t_L        g13969(.A(new_n14224), .B(new_n14225), .Y(new_n14226));
  AOI22xp33_ASAP7_75t_L     g13970(.A1(new_n1766), .A2(\b[49] ), .B1(new_n1764), .B2(new_n7914), .Y(new_n14227));
  OAI221xp5_ASAP7_75t_L     g13971(.A1(new_n1758), .A2(new_n7333), .B1(new_n7316), .B2(new_n1911), .C(new_n14227), .Y(new_n14228));
  XNOR2x2_ASAP7_75t_L       g13972(.A(\a[23] ), .B(new_n14228), .Y(new_n14229));
  A2O1A1Ixp33_ASAP7_75t_L   g13973(.A1(new_n13899), .A2(new_n13896), .B(new_n13901), .C(new_n13997), .Y(new_n14230));
  A2O1A1Ixp33_ASAP7_75t_L   g13974(.A1(new_n13998), .A2(new_n13995), .B(new_n14142), .C(new_n14230), .Y(new_n14231));
  NOR2xp33_ASAP7_75t_L      g13975(.A(new_n14229), .B(new_n14231), .Y(new_n14232));
  INVx1_ASAP7_75t_L         g13976(.A(new_n14229), .Y(new_n14233));
  A2O1A1O1Ixp25_ASAP7_75t_L g13977(.A1(new_n13995), .A2(new_n13998), .B(new_n14142), .C(new_n14230), .D(new_n14233), .Y(new_n14234));
  NOR2xp33_ASAP7_75t_L      g13978(.A(new_n14234), .B(new_n14232), .Y(new_n14235));
  AOI22xp33_ASAP7_75t_L     g13979(.A1(new_n2232), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n2228), .Y(new_n14236));
  OAI221xp5_ASAP7_75t_L     g13980(.A1(new_n2387), .A2(new_n6220), .B1(new_n2233), .B2(new_n7887), .C(new_n14236), .Y(new_n14237));
  XNOR2x2_ASAP7_75t_L       g13981(.A(\a[26] ), .B(new_n14237), .Y(new_n14238));
  O2A1O1Ixp33_ASAP7_75t_L   g13982(.A1(new_n14007), .A2(new_n14141), .B(new_n14006), .C(new_n14238), .Y(new_n14239));
  INVx1_ASAP7_75t_L         g13983(.A(new_n14239), .Y(new_n14240));
  OAI211xp5_ASAP7_75t_L     g13984(.A1(new_n14007), .A2(new_n14141), .B(new_n14006), .C(new_n14238), .Y(new_n14241));
  AND2x2_ASAP7_75t_L        g13985(.A(new_n14241), .B(new_n14240), .Y(new_n14242));
  AOI22xp33_ASAP7_75t_L     g13986(.A1(new_n2702), .A2(\b[43] ), .B1(new_n2700), .B2(new_n6202), .Y(new_n14243));
  OAI221xp5_ASAP7_75t_L     g13987(.A1(new_n2694), .A2(new_n5680), .B1(new_n5666), .B2(new_n2932), .C(new_n14243), .Y(new_n14244));
  XNOR2x2_ASAP7_75t_L       g13988(.A(\a[29] ), .B(new_n14244), .Y(new_n14245));
  MAJx2_ASAP7_75t_L         g13989(.A(new_n14133), .B(new_n14136), .C(new_n14139), .Y(new_n14246));
  INVx1_ASAP7_75t_L         g13990(.A(new_n14246), .Y(new_n14247));
  NOR2xp33_ASAP7_75t_L      g13991(.A(new_n14245), .B(new_n14247), .Y(new_n14248));
  INVx1_ASAP7_75t_L         g13992(.A(new_n14245), .Y(new_n14249));
  NOR2xp33_ASAP7_75t_L      g13993(.A(new_n14249), .B(new_n14246), .Y(new_n14250));
  AOI22xp33_ASAP7_75t_L     g13994(.A1(new_n3256), .A2(\b[40] ), .B1(new_n3254), .B2(new_n5194), .Y(new_n14251));
  OAI221xp5_ASAP7_75t_L     g13995(.A1(new_n3248), .A2(new_n5166), .B1(new_n4915), .B2(new_n3492), .C(new_n14251), .Y(new_n14252));
  XNOR2x2_ASAP7_75t_L       g13996(.A(\a[32] ), .B(new_n14252), .Y(new_n14253));
  AOI21xp33_ASAP7_75t_L     g13997(.A1(new_n14130), .A2(new_n14131), .B(new_n14120), .Y(new_n14254));
  NAND2xp33_ASAP7_75t_L     g13998(.A(new_n14253), .B(new_n14254), .Y(new_n14255));
  INVx1_ASAP7_75t_L         g13999(.A(new_n14255), .Y(new_n14256));
  O2A1O1Ixp33_ASAP7_75t_L   g14000(.A1(new_n14127), .A2(new_n14124), .B(new_n14129), .C(new_n14253), .Y(new_n14257));
  NAND2xp33_ASAP7_75t_L     g14001(.A(\b[37] ), .B(new_n3884), .Y(new_n14258));
  OAI221xp5_ASAP7_75t_L     g14002(.A1(new_n4465), .A2(new_n4312), .B1(new_n4114), .B2(new_n13559), .C(new_n14258), .Y(new_n14259));
  AOI21xp33_ASAP7_75t_L     g14003(.A1(new_n4111), .A2(\b[35] ), .B(new_n14259), .Y(new_n14260));
  NAND2xp33_ASAP7_75t_L     g14004(.A(\a[35] ), .B(new_n14260), .Y(new_n14261));
  A2O1A1Ixp33_ASAP7_75t_L   g14005(.A1(\b[35] ), .A2(new_n4111), .B(new_n14259), .C(new_n3878), .Y(new_n14262));
  NAND2xp33_ASAP7_75t_L     g14006(.A(new_n14262), .B(new_n14261), .Y(new_n14263));
  INVx1_ASAP7_75t_L         g14007(.A(new_n14263), .Y(new_n14264));
  NOR2xp33_ASAP7_75t_L      g14008(.A(new_n14113), .B(new_n14112), .Y(new_n14265));
  NAND2xp33_ASAP7_75t_L     g14009(.A(new_n14110), .B(new_n14265), .Y(new_n14266));
  A2O1A1Ixp33_ASAP7_75t_L   g14010(.A1(new_n14109), .A2(new_n14114), .B(new_n14011), .C(new_n14266), .Y(new_n14267));
  AOI22xp33_ASAP7_75t_L     g14011(.A1(new_n4544), .A2(\b[34] ), .B1(new_n4542), .B2(new_n3833), .Y(new_n14268));
  OAI221xp5_ASAP7_75t_L     g14012(.A1(new_n4536), .A2(new_n3807), .B1(new_n3443), .B2(new_n4781), .C(new_n14268), .Y(new_n14269));
  XNOR2x2_ASAP7_75t_L       g14013(.A(\a[38] ), .B(new_n14269), .Y(new_n14270));
  INVx1_ASAP7_75t_L         g14014(.A(new_n14270), .Y(new_n14271));
  INVx1_ASAP7_75t_L         g14015(.A(new_n14057), .Y(new_n14272));
  NOR2xp33_ASAP7_75t_L      g14016(.A(new_n382), .B(new_n12671), .Y(new_n14273));
  O2A1O1Ixp33_ASAP7_75t_L   g14017(.A1(new_n12353), .A2(new_n12355), .B(\b[7] ), .C(new_n14273), .Y(new_n14274));
  INVx1_ASAP7_75t_L         g14018(.A(new_n14274), .Y(new_n14275));
  O2A1O1Ixp33_ASAP7_75t_L   g14019(.A1(\a[2] ), .A2(\a[5] ), .B(new_n14040), .C(new_n14275), .Y(new_n14276));
  INVx1_ASAP7_75t_L         g14020(.A(new_n14276), .Y(new_n14277));
  AOI21xp33_ASAP7_75t_L     g14021(.A1(new_n339), .A2(new_n265), .B(new_n14039), .Y(new_n14278));
  A2O1A1Ixp33_ASAP7_75t_L   g14022(.A1(\b[7] ), .A2(new_n12669), .B(new_n14273), .C(new_n14278), .Y(new_n14279));
  AOI22xp33_ASAP7_75t_L     g14023(.A1(new_n11647), .A2(\b[9] ), .B1(\b[10] ), .B2(new_n11656), .Y(new_n14280));
  OAI221xp5_ASAP7_75t_L     g14024(.A1(new_n13003), .A2(new_n503), .B1(new_n12022), .B2(new_n641), .C(new_n14280), .Y(new_n14281));
  XNOR2x2_ASAP7_75t_L       g14025(.A(new_n11651), .B(new_n14281), .Y(new_n14282));
  NAND3xp33_ASAP7_75t_L     g14026(.A(new_n14282), .B(new_n14279), .C(new_n14277), .Y(new_n14283));
  AO21x2_ASAP7_75t_L        g14027(.A1(new_n14277), .A2(new_n14279), .B(new_n14282), .Y(new_n14284));
  AND2x2_ASAP7_75t_L        g14028(.A(new_n14283), .B(new_n14284), .Y(new_n14285));
  INVx1_ASAP7_75t_L         g14029(.A(new_n14285), .Y(new_n14286));
  O2A1O1Ixp33_ASAP7_75t_L   g14030(.A1(new_n14048), .A2(new_n14051), .B(new_n14047), .C(new_n14286), .Y(new_n14287));
  INVx1_ASAP7_75t_L         g14031(.A(new_n14287), .Y(new_n14288));
  A2O1A1O1Ixp25_ASAP7_75t_L g14032(.A1(new_n14046), .A2(new_n13798), .B(new_n14034), .C(new_n14043), .D(new_n14053), .Y(new_n14289));
  NAND2xp33_ASAP7_75t_L     g14033(.A(new_n14286), .B(new_n14289), .Y(new_n14290));
  AOI22xp33_ASAP7_75t_L     g14034(.A1(new_n10594), .A2(\b[13] ), .B1(new_n10591), .B2(new_n800), .Y(new_n14291));
  OAI221xp5_ASAP7_75t_L     g14035(.A1(new_n11335), .A2(new_n763), .B1(new_n695), .B2(new_n11330), .C(new_n14291), .Y(new_n14292));
  XNOR2x2_ASAP7_75t_L       g14036(.A(\a[59] ), .B(new_n14292), .Y(new_n14293));
  NAND3xp33_ASAP7_75t_L     g14037(.A(new_n14288), .B(new_n14290), .C(new_n14293), .Y(new_n14294));
  AO21x2_ASAP7_75t_L        g14038(.A1(new_n14290), .A2(new_n14288), .B(new_n14293), .Y(new_n14295));
  NAND2xp33_ASAP7_75t_L     g14039(.A(new_n14294), .B(new_n14295), .Y(new_n14296));
  INVx1_ASAP7_75t_L         g14040(.A(new_n14296), .Y(new_n14297));
  INVx1_ASAP7_75t_L         g14041(.A(new_n14033), .Y(new_n14298));
  NAND2xp33_ASAP7_75t_L     g14042(.A(new_n14298), .B(new_n14054), .Y(new_n14299));
  NAND3xp33_ASAP7_75t_L     g14043(.A(new_n14297), .B(new_n14272), .C(new_n14299), .Y(new_n14300));
  A2O1A1Ixp33_ASAP7_75t_L   g14044(.A1(new_n14054), .A2(new_n14298), .B(new_n14057), .C(new_n14296), .Y(new_n14301));
  AOI22xp33_ASAP7_75t_L     g14045(.A1(new_n9623), .A2(\b[16] ), .B1(new_n9620), .B2(new_n1058), .Y(new_n14302));
  OAI221xp5_ASAP7_75t_L     g14046(.A1(new_n10280), .A2(new_n952), .B1(new_n871), .B2(new_n12010), .C(new_n14302), .Y(new_n14303));
  XNOR2x2_ASAP7_75t_L       g14047(.A(\a[56] ), .B(new_n14303), .Y(new_n14304));
  NAND3xp33_ASAP7_75t_L     g14048(.A(new_n14300), .B(new_n14301), .C(new_n14304), .Y(new_n14305));
  AO21x2_ASAP7_75t_L        g14049(.A1(new_n14301), .A2(new_n14300), .B(new_n14304), .Y(new_n14306));
  AOI21xp33_ASAP7_75t_L     g14050(.A1(new_n14059), .A2(new_n14027), .B(new_n14063), .Y(new_n14307));
  NAND3xp33_ASAP7_75t_L     g14051(.A(new_n14307), .B(new_n14306), .C(new_n14305), .Y(new_n14308));
  NAND2xp33_ASAP7_75t_L     g14052(.A(new_n14305), .B(new_n14306), .Y(new_n14309));
  A2O1A1Ixp33_ASAP7_75t_L   g14053(.A1(new_n14059), .A2(new_n14027), .B(new_n14063), .C(new_n14309), .Y(new_n14310));
  AOI22xp33_ASAP7_75t_L     g14054(.A1(new_n8645), .A2(\b[19] ), .B1(new_n8642), .B2(new_n1499), .Y(new_n14311));
  OAI221xp5_ASAP7_75t_L     g14055(.A1(new_n9322), .A2(new_n1356), .B1(new_n1244), .B2(new_n8965), .C(new_n14311), .Y(new_n14312));
  XNOR2x2_ASAP7_75t_L       g14056(.A(\a[53] ), .B(new_n14312), .Y(new_n14313));
  NAND3xp33_ASAP7_75t_L     g14057(.A(new_n14308), .B(new_n14310), .C(new_n14313), .Y(new_n14314));
  AO21x2_ASAP7_75t_L        g14058(.A1(new_n14310), .A2(new_n14308), .B(new_n14313), .Y(new_n14315));
  NAND2xp33_ASAP7_75t_L     g14059(.A(new_n14314), .B(new_n14315), .Y(new_n14316));
  OAI21xp33_ASAP7_75t_L     g14060(.A1(new_n14065), .A2(new_n14068), .B(new_n14073), .Y(new_n14317));
  NOR2xp33_ASAP7_75t_L      g14061(.A(new_n14316), .B(new_n14317), .Y(new_n14318));
  INVx1_ASAP7_75t_L         g14062(.A(new_n14316), .Y(new_n14319));
  O2A1O1Ixp33_ASAP7_75t_L   g14063(.A1(new_n14065), .A2(new_n14068), .B(new_n14073), .C(new_n14319), .Y(new_n14320));
  NOR2xp33_ASAP7_75t_L      g14064(.A(new_n14320), .B(new_n14318), .Y(new_n14321));
  AOI22xp33_ASAP7_75t_L     g14065(.A1(new_n7659), .A2(\b[22] ), .B1(new_n7656), .B2(new_n1864), .Y(new_n14322));
  OAI221xp5_ASAP7_75t_L     g14066(.A1(new_n8326), .A2(new_n1709), .B1(new_n1594), .B2(new_n7994), .C(new_n14322), .Y(new_n14323));
  XNOR2x2_ASAP7_75t_L       g14067(.A(\a[50] ), .B(new_n14323), .Y(new_n14324));
  XOR2x2_ASAP7_75t_L        g14068(.A(new_n14324), .B(new_n14321), .Y(new_n14325));
  AOI21xp33_ASAP7_75t_L     g14069(.A1(new_n14080), .A2(new_n14074), .B(new_n14082), .Y(new_n14326));
  XOR2x2_ASAP7_75t_L        g14070(.A(new_n14326), .B(new_n14325), .Y(new_n14327));
  AOI22xp33_ASAP7_75t_L     g14071(.A1(new_n6822), .A2(\b[25] ), .B1(new_n6819), .B2(new_n2188), .Y(new_n14328));
  OAI221xp5_ASAP7_75t_L     g14072(.A1(new_n7392), .A2(new_n2019), .B1(new_n1995), .B2(new_n7115), .C(new_n14328), .Y(new_n14329));
  XNOR2x2_ASAP7_75t_L       g14073(.A(\a[47] ), .B(new_n14329), .Y(new_n14330));
  XNOR2x2_ASAP7_75t_L       g14074(.A(new_n14330), .B(new_n14327), .Y(new_n14331));
  MAJx2_ASAP7_75t_L         g14075(.A(new_n14087), .B(new_n14018), .C(new_n14084), .Y(new_n14332));
  OR2x4_ASAP7_75t_L         g14076(.A(new_n14332), .B(new_n14331), .Y(new_n14333));
  NAND2xp33_ASAP7_75t_L     g14077(.A(new_n14332), .B(new_n14331), .Y(new_n14334));
  NAND2xp33_ASAP7_75t_L     g14078(.A(\b[28] ), .B(new_n6002), .Y(new_n14335));
  OAI221xp5_ASAP7_75t_L     g14079(.A1(new_n2650), .A2(new_n6544), .B1(new_n6311), .B2(new_n5212), .C(new_n14335), .Y(new_n14336));
  AOI21xp33_ASAP7_75t_L     g14080(.A1(new_n6308), .A2(\b[26] ), .B(new_n14336), .Y(new_n14337));
  NAND2xp33_ASAP7_75t_L     g14081(.A(\a[44] ), .B(new_n14337), .Y(new_n14338));
  A2O1A1Ixp33_ASAP7_75t_L   g14082(.A1(\b[26] ), .A2(new_n6308), .B(new_n14336), .C(new_n5996), .Y(new_n14339));
  AND2x2_ASAP7_75t_L        g14083(.A(new_n14339), .B(new_n14338), .Y(new_n14340));
  NAND3xp33_ASAP7_75t_L     g14084(.A(new_n14333), .B(new_n14334), .C(new_n14340), .Y(new_n14341));
  AO21x2_ASAP7_75t_L        g14085(.A1(new_n14334), .A2(new_n14333), .B(new_n14340), .Y(new_n14342));
  NAND2xp33_ASAP7_75t_L     g14086(.A(new_n14341), .B(new_n14342), .Y(new_n14343));
  OAI21xp33_ASAP7_75t_L     g14087(.A1(new_n14088), .A2(new_n14091), .B(new_n14096), .Y(new_n14344));
  XNOR2x2_ASAP7_75t_L       g14088(.A(new_n14343), .B(new_n14344), .Y(new_n14345));
  AOI22xp33_ASAP7_75t_L     g14089(.A1(new_n5249), .A2(\b[31] ), .B1(new_n5247), .B2(new_n3426), .Y(new_n14346));
  OAI221xp5_ASAP7_75t_L     g14090(.A1(new_n5241), .A2(new_n3212), .B1(new_n2871), .B2(new_n5521), .C(new_n14346), .Y(new_n14347));
  XNOR2x2_ASAP7_75t_L       g14091(.A(\a[41] ), .B(new_n14347), .Y(new_n14348));
  NAND2xp33_ASAP7_75t_L     g14092(.A(new_n14348), .B(new_n14345), .Y(new_n14349));
  INVx1_ASAP7_75t_L         g14093(.A(new_n14349), .Y(new_n14350));
  NOR2xp33_ASAP7_75t_L      g14094(.A(new_n14348), .B(new_n14345), .Y(new_n14351));
  NOR2xp33_ASAP7_75t_L      g14095(.A(new_n14351), .B(new_n14350), .Y(new_n14352));
  A2O1A1Ixp33_ASAP7_75t_L   g14096(.A1(new_n14101), .A2(new_n14104), .B(new_n14112), .C(new_n14352), .Y(new_n14353));
  INVx1_ASAP7_75t_L         g14097(.A(new_n14351), .Y(new_n14354));
  NAND2xp33_ASAP7_75t_L     g14098(.A(new_n14349), .B(new_n14354), .Y(new_n14355));
  NAND3xp33_ASAP7_75t_L     g14099(.A(new_n14355), .B(new_n14103), .C(new_n14105), .Y(new_n14356));
  NAND3xp33_ASAP7_75t_L     g14100(.A(new_n14353), .B(new_n14356), .C(new_n14271), .Y(new_n14357));
  O2A1O1Ixp33_ASAP7_75t_L   g14101(.A1(new_n14097), .A2(new_n14100), .B(new_n14103), .C(new_n14355), .Y(new_n14358));
  NAND2xp33_ASAP7_75t_L     g14102(.A(new_n14105), .B(new_n14103), .Y(new_n14359));
  NOR2xp33_ASAP7_75t_L      g14103(.A(new_n14359), .B(new_n14352), .Y(new_n14360));
  OAI21xp33_ASAP7_75t_L     g14104(.A1(new_n14360), .A2(new_n14358), .B(new_n14270), .Y(new_n14361));
  NAND3xp33_ASAP7_75t_L     g14105(.A(new_n14361), .B(new_n14357), .C(new_n14267), .Y(new_n14362));
  INVx1_ASAP7_75t_L         g14106(.A(new_n14267), .Y(new_n14363));
  NOR3xp33_ASAP7_75t_L      g14107(.A(new_n14358), .B(new_n14360), .C(new_n14270), .Y(new_n14364));
  AOI21xp33_ASAP7_75t_L     g14108(.A1(new_n14353), .A2(new_n14356), .B(new_n14271), .Y(new_n14365));
  OAI21xp33_ASAP7_75t_L     g14109(.A1(new_n14365), .A2(new_n14364), .B(new_n14363), .Y(new_n14366));
  AOI21xp33_ASAP7_75t_L     g14110(.A1(new_n14366), .A2(new_n14362), .B(new_n14264), .Y(new_n14367));
  AND3x1_ASAP7_75t_L        g14111(.A(new_n14366), .B(new_n14362), .C(new_n14264), .Y(new_n14368));
  NOR2xp33_ASAP7_75t_L      g14112(.A(new_n14367), .B(new_n14368), .Y(new_n14369));
  NOR3xp33_ASAP7_75t_L      g14113(.A(new_n14369), .B(new_n14257), .C(new_n14256), .Y(new_n14370));
  INVx1_ASAP7_75t_L         g14114(.A(new_n14257), .Y(new_n14371));
  AOI211xp5_ASAP7_75t_L     g14115(.A1(new_n14255), .A2(new_n14371), .B(new_n14367), .C(new_n14368), .Y(new_n14372));
  NOR2xp33_ASAP7_75t_L      g14116(.A(new_n14372), .B(new_n14370), .Y(new_n14373));
  OA21x2_ASAP7_75t_L        g14117(.A1(new_n14248), .A2(new_n14250), .B(new_n14373), .Y(new_n14374));
  NOR3xp33_ASAP7_75t_L      g14118(.A(new_n14373), .B(new_n14250), .C(new_n14248), .Y(new_n14375));
  NOR2xp33_ASAP7_75t_L      g14119(.A(new_n14375), .B(new_n14374), .Y(new_n14376));
  NAND2xp33_ASAP7_75t_L     g14120(.A(new_n14242), .B(new_n14376), .Y(new_n14377));
  NAND2xp33_ASAP7_75t_L     g14121(.A(new_n14241), .B(new_n14240), .Y(new_n14378));
  OAI21xp33_ASAP7_75t_L     g14122(.A1(new_n14374), .A2(new_n14375), .B(new_n14378), .Y(new_n14379));
  NAND2xp33_ASAP7_75t_L     g14123(.A(new_n14379), .B(new_n14377), .Y(new_n14380));
  XOR2x2_ASAP7_75t_L        g14124(.A(new_n14235), .B(new_n14380), .Y(new_n14381));
  XNOR2x2_ASAP7_75t_L       g14125(.A(new_n14226), .B(new_n14381), .Y(new_n14382));
  XOR2x2_ASAP7_75t_L        g14126(.A(new_n14221), .B(new_n14382), .Y(new_n14383));
  NOR2xp33_ASAP7_75t_L      g14127(.A(new_n14213), .B(new_n14383), .Y(new_n14384));
  AND2x2_ASAP7_75t_L        g14128(.A(new_n14213), .B(new_n14383), .Y(new_n14385));
  NOR2xp33_ASAP7_75t_L      g14129(.A(new_n14384), .B(new_n14385), .Y(new_n14386));
  NAND3xp33_ASAP7_75t_L     g14130(.A(new_n14206), .B(new_n14386), .C(new_n14204), .Y(new_n14387));
  AO21x2_ASAP7_75t_L        g14131(.A1(new_n14204), .A2(new_n14206), .B(new_n14386), .Y(new_n14388));
  NAND2xp33_ASAP7_75t_L     g14132(.A(new_n14387), .B(new_n14388), .Y(new_n14389));
  NAND3xp33_ASAP7_75t_L     g14133(.A(new_n14389), .B(new_n14199), .C(new_n14197), .Y(new_n14390));
  AO21x2_ASAP7_75t_L        g14134(.A1(new_n14197), .A2(new_n14199), .B(new_n14389), .Y(new_n14391));
  NAND2xp33_ASAP7_75t_L     g14135(.A(new_n14390), .B(new_n14391), .Y(new_n14392));
  A2O1A1O1Ixp25_ASAP7_75t_L g14136(.A1(new_n13731), .A2(new_n13729), .B(new_n13928), .C(new_n13953), .D(new_n13957), .Y(new_n14393));
  O2A1O1Ixp33_ASAP7_75t_L   g14137(.A1(new_n14177), .A2(new_n14178), .B(new_n13963), .C(new_n14393), .Y(new_n14394));
  XNOR2x2_ASAP7_75t_L       g14138(.A(new_n14394), .B(new_n14392), .Y(new_n14395));
  INVx1_ASAP7_75t_L         g14139(.A(new_n14395), .Y(new_n14396));
  O2A1O1Ixp33_ASAP7_75t_L   g14140(.A1(new_n14187), .A2(new_n14182), .B(new_n14180), .C(new_n14396), .Y(new_n14397));
  A2O1A1Ixp33_ASAP7_75t_L   g14141(.A1(new_n13946), .A2(new_n14185), .B(new_n14182), .C(new_n14180), .Y(new_n14398));
  NOR2xp33_ASAP7_75t_L      g14142(.A(new_n14395), .B(new_n14398), .Y(new_n14399));
  NOR2xp33_ASAP7_75t_L      g14143(.A(new_n14399), .B(new_n14397), .Y(\f[70] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14144(.A1(new_n13963), .A2(new_n14175), .B(new_n14393), .C(new_n14392), .Y(new_n14401));
  INVx1_ASAP7_75t_L         g14145(.A(new_n14401), .Y(new_n14402));
  AOI22xp33_ASAP7_75t_L     g14146(.A1(new_n590), .A2(\b[61] ), .B1(\b[62] ), .B2(new_n600), .Y(new_n14403));
  OAI221xp5_ASAP7_75t_L     g14147(.A1(new_n1620), .A2(new_n11226), .B1(new_n675), .B2(new_n12281), .C(new_n14403), .Y(new_n14404));
  NOR2xp33_ASAP7_75t_L      g14148(.A(new_n594), .B(new_n14404), .Y(new_n14405));
  AND2x2_ASAP7_75t_L        g14149(.A(new_n594), .B(new_n14404), .Y(new_n14406));
  NOR2xp33_ASAP7_75t_L      g14150(.A(new_n14405), .B(new_n14406), .Y(new_n14407));
  INVx1_ASAP7_75t_L         g14151(.A(new_n14407), .Y(new_n14408));
  O2A1O1Ixp33_ASAP7_75t_L   g14152(.A1(new_n14213), .A2(new_n14383), .B(new_n14211), .C(new_n14408), .Y(new_n14409));
  INVx1_ASAP7_75t_L         g14153(.A(new_n14409), .Y(new_n14410));
  O2A1O1Ixp33_ASAP7_75t_L   g14154(.A1(new_n14162), .A2(new_n14165), .B(new_n14210), .C(new_n14384), .Y(new_n14411));
  NAND2xp33_ASAP7_75t_L     g14155(.A(new_n14408), .B(new_n14411), .Y(new_n14412));
  NAND2xp33_ASAP7_75t_L     g14156(.A(new_n14410), .B(new_n14412), .Y(new_n14413));
  AOI22xp33_ASAP7_75t_L     g14157(.A1(new_n1113), .A2(\b[56] ), .B1(new_n1110), .B2(new_n10185), .Y(new_n14414));
  OAI221xp5_ASAP7_75t_L     g14158(.A1(new_n1298), .A2(new_n9534), .B1(new_n9199), .B2(new_n1195), .C(new_n14414), .Y(new_n14415));
  XNOR2x2_ASAP7_75t_L       g14159(.A(\a[17] ), .B(new_n14415), .Y(new_n14416));
  INVx1_ASAP7_75t_L         g14160(.A(new_n14416), .Y(new_n14417));
  MAJIxp5_ASAP7_75t_L       g14161(.A(new_n14381), .B(new_n14224), .C(new_n14225), .Y(new_n14418));
  XNOR2x2_ASAP7_75t_L       g14162(.A(new_n14417), .B(new_n14418), .Y(new_n14419));
  AOI22xp33_ASAP7_75t_L     g14163(.A1(new_n1766), .A2(\b[50] ), .B1(new_n1764), .B2(new_n8235), .Y(new_n14420));
  OAI221xp5_ASAP7_75t_L     g14164(.A1(new_n1758), .A2(new_n7907), .B1(new_n7333), .B2(new_n1911), .C(new_n14420), .Y(new_n14421));
  XNOR2x2_ASAP7_75t_L       g14165(.A(\a[23] ), .B(new_n14421), .Y(new_n14422));
  AOI21xp33_ASAP7_75t_L     g14166(.A1(new_n14376), .A2(new_n14241), .B(new_n14239), .Y(new_n14423));
  NAND2xp33_ASAP7_75t_L     g14167(.A(new_n14422), .B(new_n14423), .Y(new_n14424));
  NOR2xp33_ASAP7_75t_L      g14168(.A(new_n14422), .B(new_n14423), .Y(new_n14425));
  INVx1_ASAP7_75t_L         g14169(.A(new_n14425), .Y(new_n14426));
  AOI22xp33_ASAP7_75t_L     g14170(.A1(new_n2228), .A2(\b[47] ), .B1(new_n2226), .B2(new_n7323), .Y(new_n14427));
  OAI221xp5_ASAP7_75t_L     g14171(.A1(new_n2220), .A2(new_n7033), .B1(new_n6756), .B2(new_n2387), .C(new_n14427), .Y(new_n14428));
  XNOR2x2_ASAP7_75t_L       g14172(.A(\a[26] ), .B(new_n14428), .Y(new_n14429));
  MAJx2_ASAP7_75t_L         g14173(.A(new_n14373), .B(new_n14247), .C(new_n14249), .Y(new_n14430));
  XNOR2x2_ASAP7_75t_L       g14174(.A(new_n14429), .B(new_n14430), .Y(new_n14431));
  AOI22xp33_ASAP7_75t_L     g14175(.A1(new_n2706), .A2(\b[43] ), .B1(\b[44] ), .B2(new_n2702), .Y(new_n14432));
  OAI221xp5_ASAP7_75t_L     g14176(.A1(new_n2932), .A2(new_n5680), .B1(new_n2707), .B2(new_n6229), .C(new_n14432), .Y(new_n14433));
  NOR2xp33_ASAP7_75t_L      g14177(.A(new_n2697), .B(new_n14433), .Y(new_n14434));
  AND2x2_ASAP7_75t_L        g14178(.A(new_n2697), .B(new_n14433), .Y(new_n14435));
  NOR2xp33_ASAP7_75t_L      g14179(.A(new_n14434), .B(new_n14435), .Y(new_n14436));
  AOI21xp33_ASAP7_75t_L     g14180(.A1(new_n14369), .A2(new_n14371), .B(new_n14256), .Y(new_n14437));
  NAND2xp33_ASAP7_75t_L     g14181(.A(new_n14436), .B(new_n14437), .Y(new_n14438));
  INVx1_ASAP7_75t_L         g14182(.A(new_n14436), .Y(new_n14439));
  A2O1A1Ixp33_ASAP7_75t_L   g14183(.A1(new_n14369), .A2(new_n14371), .B(new_n14256), .C(new_n14439), .Y(new_n14440));
  NAND2xp33_ASAP7_75t_L     g14184(.A(new_n14440), .B(new_n14438), .Y(new_n14441));
  NOR2xp33_ASAP7_75t_L      g14185(.A(new_n14365), .B(new_n14364), .Y(new_n14442));
  NAND3xp33_ASAP7_75t_L     g14186(.A(new_n14366), .B(new_n14362), .C(new_n14264), .Y(new_n14443));
  AOI22xp33_ASAP7_75t_L     g14187(.A1(new_n3256), .A2(\b[41] ), .B1(new_n3254), .B2(new_n5669), .Y(new_n14444));
  OAI221xp5_ASAP7_75t_L     g14188(.A1(new_n3248), .A2(new_n5186), .B1(new_n5166), .B2(new_n3492), .C(new_n14444), .Y(new_n14445));
  XNOR2x2_ASAP7_75t_L       g14189(.A(\a[32] ), .B(new_n14445), .Y(new_n14446));
  INVx1_ASAP7_75t_L         g14190(.A(new_n14446), .Y(new_n14447));
  O2A1O1Ixp33_ASAP7_75t_L   g14191(.A1(new_n14267), .A2(new_n14442), .B(new_n14443), .C(new_n14447), .Y(new_n14448));
  MAJIxp5_ASAP7_75t_L       g14192(.A(new_n14442), .B(new_n14263), .C(new_n14267), .Y(new_n14449));
  NOR2xp33_ASAP7_75t_L      g14193(.A(new_n14446), .B(new_n14449), .Y(new_n14450));
  AOI22xp33_ASAP7_75t_L     g14194(.A1(new_n7659), .A2(\b[23] ), .B1(new_n7656), .B2(new_n2002), .Y(new_n14451));
  OAI221xp5_ASAP7_75t_L     g14195(.A1(new_n8326), .A2(new_n1857), .B1(new_n1709), .B2(new_n7994), .C(new_n14451), .Y(new_n14452));
  XNOR2x2_ASAP7_75t_L       g14196(.A(\a[50] ), .B(new_n14452), .Y(new_n14453));
  INVx1_ASAP7_75t_L         g14197(.A(new_n14453), .Y(new_n14454));
  INVx1_ASAP7_75t_L         g14198(.A(new_n14300), .Y(new_n14455));
  INVx1_ASAP7_75t_L         g14199(.A(new_n14289), .Y(new_n14456));
  AOI22xp33_ASAP7_75t_L     g14200(.A1(new_n10594), .A2(\b[14] ), .B1(new_n10591), .B2(new_n879), .Y(new_n14457));
  OAI221xp5_ASAP7_75t_L     g14201(.A1(new_n11335), .A2(new_n793), .B1(new_n763), .B2(new_n11330), .C(new_n14457), .Y(new_n14458));
  XNOR2x2_ASAP7_75t_L       g14202(.A(\a[59] ), .B(new_n14458), .Y(new_n14459));
  INVx1_ASAP7_75t_L         g14203(.A(new_n14459), .Y(new_n14460));
  AOI22xp33_ASAP7_75t_L     g14204(.A1(new_n11656), .A2(\b[11] ), .B1(new_n11654), .B2(new_n702), .Y(new_n14461));
  OAI221xp5_ASAP7_75t_L     g14205(.A1(new_n12364), .A2(new_n631), .B1(new_n559), .B2(new_n13003), .C(new_n14461), .Y(new_n14462));
  XNOR2x2_ASAP7_75t_L       g14206(.A(\a[62] ), .B(new_n14462), .Y(new_n14463));
  INVx1_ASAP7_75t_L         g14207(.A(new_n14463), .Y(new_n14464));
  AOI21xp33_ASAP7_75t_L     g14208(.A1(new_n14282), .A2(new_n14279), .B(new_n14276), .Y(new_n14465));
  NOR2xp33_ASAP7_75t_L      g14209(.A(new_n421), .B(new_n12671), .Y(new_n14466));
  INVx1_ASAP7_75t_L         g14210(.A(new_n14466), .Y(new_n14467));
  O2A1O1Ixp33_ASAP7_75t_L   g14211(.A1(new_n12356), .A2(new_n503), .B(new_n14467), .C(new_n14275), .Y(new_n14468));
  O2A1O1Ixp33_ASAP7_75t_L   g14212(.A1(new_n12353), .A2(new_n12355), .B(\b[8] ), .C(new_n14466), .Y(new_n14469));
  A2O1A1Ixp33_ASAP7_75t_L   g14213(.A1(new_n12669), .A2(\b[7] ), .B(new_n14273), .C(new_n14469), .Y(new_n14470));
  INVx1_ASAP7_75t_L         g14214(.A(new_n14470), .Y(new_n14471));
  OAI21xp33_ASAP7_75t_L     g14215(.A1(new_n14468), .A2(new_n14471), .B(new_n14465), .Y(new_n14472));
  NOR2xp33_ASAP7_75t_L      g14216(.A(new_n14471), .B(new_n14468), .Y(new_n14473));
  A2O1A1Ixp33_ASAP7_75t_L   g14217(.A1(new_n14282), .A2(new_n14279), .B(new_n14276), .C(new_n14473), .Y(new_n14474));
  NAND3xp33_ASAP7_75t_L     g14218(.A(new_n14464), .B(new_n14472), .C(new_n14474), .Y(new_n14475));
  AO21x2_ASAP7_75t_L        g14219(.A1(new_n14474), .A2(new_n14472), .B(new_n14464), .Y(new_n14476));
  NAND3xp33_ASAP7_75t_L     g14220(.A(new_n14460), .B(new_n14475), .C(new_n14476), .Y(new_n14477));
  NAND2xp33_ASAP7_75t_L     g14221(.A(new_n14475), .B(new_n14476), .Y(new_n14478));
  NAND2xp33_ASAP7_75t_L     g14222(.A(new_n14459), .B(new_n14478), .Y(new_n14479));
  AND2x2_ASAP7_75t_L        g14223(.A(new_n14479), .B(new_n14477), .Y(new_n14480));
  O2A1O1Ixp33_ASAP7_75t_L   g14224(.A1(new_n14456), .A2(new_n14285), .B(new_n14294), .C(new_n14480), .Y(new_n14481));
  INVx1_ASAP7_75t_L         g14225(.A(new_n14481), .Y(new_n14482));
  NAND3xp33_ASAP7_75t_L     g14226(.A(new_n14480), .B(new_n14294), .C(new_n14290), .Y(new_n14483));
  AOI22xp33_ASAP7_75t_L     g14227(.A1(new_n9623), .A2(\b[17] ), .B1(new_n9620), .B2(new_n1252), .Y(new_n14484));
  OAI221xp5_ASAP7_75t_L     g14228(.A1(new_n10280), .A2(new_n1051), .B1(new_n952), .B2(new_n12010), .C(new_n14484), .Y(new_n14485));
  XNOR2x2_ASAP7_75t_L       g14229(.A(\a[56] ), .B(new_n14485), .Y(new_n14486));
  AND3x1_ASAP7_75t_L        g14230(.A(new_n14482), .B(new_n14486), .C(new_n14483), .Y(new_n14487));
  AOI21xp33_ASAP7_75t_L     g14231(.A1(new_n14482), .A2(new_n14483), .B(new_n14486), .Y(new_n14488));
  NOR2xp33_ASAP7_75t_L      g14232(.A(new_n14488), .B(new_n14487), .Y(new_n14489));
  A2O1A1Ixp33_ASAP7_75t_L   g14233(.A1(new_n14301), .A2(new_n14304), .B(new_n14455), .C(new_n14489), .Y(new_n14490));
  INVx1_ASAP7_75t_L         g14234(.A(new_n14489), .Y(new_n14491));
  NAND3xp33_ASAP7_75t_L     g14235(.A(new_n14491), .B(new_n14305), .C(new_n14300), .Y(new_n14492));
  NAND2xp33_ASAP7_75t_L     g14236(.A(new_n14490), .B(new_n14492), .Y(new_n14493));
  AOI22xp33_ASAP7_75t_L     g14237(.A1(new_n8645), .A2(\b[20] ), .B1(new_n8642), .B2(new_n1600), .Y(new_n14494));
  OAI221xp5_ASAP7_75t_L     g14238(.A1(new_n9322), .A2(new_n1493), .B1(new_n1356), .B2(new_n8965), .C(new_n14494), .Y(new_n14495));
  XNOR2x2_ASAP7_75t_L       g14239(.A(\a[53] ), .B(new_n14495), .Y(new_n14496));
  INVx1_ASAP7_75t_L         g14240(.A(new_n14496), .Y(new_n14497));
  XNOR2x2_ASAP7_75t_L       g14241(.A(new_n14497), .B(new_n14493), .Y(new_n14498));
  NAND2xp33_ASAP7_75t_L     g14242(.A(new_n14308), .B(new_n14314), .Y(new_n14499));
  XNOR2x2_ASAP7_75t_L       g14243(.A(new_n14499), .B(new_n14498), .Y(new_n14500));
  NAND2xp33_ASAP7_75t_L     g14244(.A(new_n14454), .B(new_n14500), .Y(new_n14501));
  INVx1_ASAP7_75t_L         g14245(.A(new_n14500), .Y(new_n14502));
  NAND2xp33_ASAP7_75t_L     g14246(.A(new_n14453), .B(new_n14502), .Y(new_n14503));
  NAND2xp33_ASAP7_75t_L     g14247(.A(new_n14501), .B(new_n14503), .Y(new_n14504));
  AO21x2_ASAP7_75t_L        g14248(.A1(new_n14324), .A2(new_n14321), .B(new_n14318), .Y(new_n14505));
  XNOR2x2_ASAP7_75t_L       g14249(.A(new_n14505), .B(new_n14504), .Y(new_n14506));
  AOI22xp33_ASAP7_75t_L     g14250(.A1(new_n6822), .A2(\b[26] ), .B1(new_n6819), .B2(new_n2888), .Y(new_n14507));
  OAI221xp5_ASAP7_75t_L     g14251(.A1(new_n7392), .A2(new_n2180), .B1(new_n2019), .B2(new_n7115), .C(new_n14507), .Y(new_n14508));
  XNOR2x2_ASAP7_75t_L       g14252(.A(\a[47] ), .B(new_n14508), .Y(new_n14509));
  XNOR2x2_ASAP7_75t_L       g14253(.A(new_n14509), .B(new_n14506), .Y(new_n14510));
  NAND2xp33_ASAP7_75t_L     g14254(.A(new_n14326), .B(new_n14325), .Y(new_n14511));
  INVx1_ASAP7_75t_L         g14255(.A(new_n14511), .Y(new_n14512));
  AO21x2_ASAP7_75t_L        g14256(.A1(new_n14330), .A2(new_n14327), .B(new_n14512), .Y(new_n14513));
  AND2x2_ASAP7_75t_L        g14257(.A(new_n14513), .B(new_n14510), .Y(new_n14514));
  NOR2xp33_ASAP7_75t_L      g14258(.A(new_n14513), .B(new_n14510), .Y(new_n14515));
  NOR2xp33_ASAP7_75t_L      g14259(.A(new_n14515), .B(new_n14514), .Y(new_n14516));
  AOI22xp33_ASAP7_75t_L     g14260(.A1(new_n6002), .A2(\b[29] ), .B1(new_n5999), .B2(new_n5472), .Y(new_n14517));
  OAI221xp5_ASAP7_75t_L     g14261(.A1(new_n6544), .A2(new_n2852), .B1(new_n2650), .B2(new_n6309), .C(new_n14517), .Y(new_n14518));
  XNOR2x2_ASAP7_75t_L       g14262(.A(\a[44] ), .B(new_n14518), .Y(new_n14519));
  NAND2xp33_ASAP7_75t_L     g14263(.A(new_n14519), .B(new_n14516), .Y(new_n14520));
  INVx1_ASAP7_75t_L         g14264(.A(new_n14519), .Y(new_n14521));
  OAI21xp33_ASAP7_75t_L     g14265(.A1(new_n14515), .A2(new_n14514), .B(new_n14521), .Y(new_n14522));
  NAND2xp33_ASAP7_75t_L     g14266(.A(new_n14522), .B(new_n14520), .Y(new_n14523));
  NAND2xp33_ASAP7_75t_L     g14267(.A(new_n14333), .B(new_n14341), .Y(new_n14524));
  XOR2x2_ASAP7_75t_L        g14268(.A(new_n14524), .B(new_n14523), .Y(new_n14525));
  AOI22xp33_ASAP7_75t_L     g14269(.A1(new_n5249), .A2(\b[32] ), .B1(new_n5247), .B2(new_n3450), .Y(new_n14526));
  OAI221xp5_ASAP7_75t_L     g14270(.A1(new_n5241), .A2(new_n3419), .B1(new_n3212), .B2(new_n5521), .C(new_n14526), .Y(new_n14527));
  XNOR2x2_ASAP7_75t_L       g14271(.A(\a[41] ), .B(new_n14527), .Y(new_n14528));
  AND2x2_ASAP7_75t_L        g14272(.A(new_n14528), .B(new_n14525), .Y(new_n14529));
  NOR2xp33_ASAP7_75t_L      g14273(.A(new_n14528), .B(new_n14525), .Y(new_n14530));
  NOR2xp33_ASAP7_75t_L      g14274(.A(new_n14530), .B(new_n14529), .Y(new_n14531));
  NAND2xp33_ASAP7_75t_L     g14275(.A(new_n14343), .B(new_n14344), .Y(new_n14532));
  NAND2xp33_ASAP7_75t_L     g14276(.A(new_n14532), .B(new_n14354), .Y(new_n14533));
  XNOR2x2_ASAP7_75t_L       g14277(.A(new_n14531), .B(new_n14533), .Y(new_n14534));
  AOI22xp33_ASAP7_75t_L     g14278(.A1(new_n4544), .A2(\b[35] ), .B1(new_n4542), .B2(new_n5649), .Y(new_n14535));
  OAI221xp5_ASAP7_75t_L     g14279(.A1(new_n4536), .A2(new_n3827), .B1(new_n3807), .B2(new_n4781), .C(new_n14535), .Y(new_n14536));
  XNOR2x2_ASAP7_75t_L       g14280(.A(\a[38] ), .B(new_n14536), .Y(new_n14537));
  INVx1_ASAP7_75t_L         g14281(.A(new_n14537), .Y(new_n14538));
  NOR2xp33_ASAP7_75t_L      g14282(.A(new_n14538), .B(new_n14534), .Y(new_n14539));
  XNOR2x2_ASAP7_75t_L       g14283(.A(new_n14528), .B(new_n14525), .Y(new_n14540));
  O2A1O1Ixp33_ASAP7_75t_L   g14284(.A1(new_n14345), .A2(new_n14348), .B(new_n14532), .C(new_n14540), .Y(new_n14541));
  NOR2xp33_ASAP7_75t_L      g14285(.A(new_n14531), .B(new_n14533), .Y(new_n14542));
  NOR2xp33_ASAP7_75t_L      g14286(.A(new_n14541), .B(new_n14542), .Y(new_n14543));
  NOR2xp33_ASAP7_75t_L      g14287(.A(new_n14537), .B(new_n14543), .Y(new_n14544));
  NOR2xp33_ASAP7_75t_L      g14288(.A(new_n14539), .B(new_n14544), .Y(new_n14545));
  A2O1A1O1Ixp25_ASAP7_75t_L g14289(.A1(new_n14101), .A2(new_n14104), .B(new_n14112), .C(new_n14352), .D(new_n14364), .Y(new_n14546));
  NAND2xp33_ASAP7_75t_L     g14290(.A(new_n14546), .B(new_n14545), .Y(new_n14547));
  NAND2xp33_ASAP7_75t_L     g14291(.A(new_n14537), .B(new_n14543), .Y(new_n14548));
  NAND2xp33_ASAP7_75t_L     g14292(.A(new_n14538), .B(new_n14534), .Y(new_n14549));
  NAND2xp33_ASAP7_75t_L     g14293(.A(new_n14549), .B(new_n14548), .Y(new_n14550));
  A2O1A1Ixp33_ASAP7_75t_L   g14294(.A1(new_n14359), .A2(new_n14352), .B(new_n14364), .C(new_n14550), .Y(new_n14551));
  AOI22xp33_ASAP7_75t_L     g14295(.A1(new_n3884), .A2(\b[38] ), .B1(new_n3881), .B2(new_n4923), .Y(new_n14552));
  OAI221xp5_ASAP7_75t_L     g14296(.A1(new_n4312), .A2(new_n4701), .B1(new_n4465), .B2(new_n4986), .C(new_n14552), .Y(new_n14553));
  XNOR2x2_ASAP7_75t_L       g14297(.A(\a[35] ), .B(new_n14553), .Y(new_n14554));
  INVx1_ASAP7_75t_L         g14298(.A(new_n14554), .Y(new_n14555));
  NAND3xp33_ASAP7_75t_L     g14299(.A(new_n14551), .B(new_n14547), .C(new_n14555), .Y(new_n14556));
  A2O1A1Ixp33_ASAP7_75t_L   g14300(.A1(new_n14103), .A2(new_n14105), .B(new_n14355), .C(new_n14357), .Y(new_n14557));
  NOR2xp33_ASAP7_75t_L      g14301(.A(new_n14557), .B(new_n14550), .Y(new_n14558));
  AOI21xp33_ASAP7_75t_L     g14302(.A1(new_n14549), .A2(new_n14548), .B(new_n14546), .Y(new_n14559));
  OAI21xp33_ASAP7_75t_L     g14303(.A1(new_n14559), .A2(new_n14558), .B(new_n14554), .Y(new_n14560));
  NAND2xp33_ASAP7_75t_L     g14304(.A(new_n14560), .B(new_n14556), .Y(new_n14561));
  NOR3xp33_ASAP7_75t_L      g14305(.A(new_n14561), .B(new_n14450), .C(new_n14448), .Y(new_n14562));
  NOR2xp33_ASAP7_75t_L      g14306(.A(new_n14450), .B(new_n14448), .Y(new_n14563));
  AOI21xp33_ASAP7_75t_L     g14307(.A1(new_n14560), .A2(new_n14556), .B(new_n14563), .Y(new_n14564));
  NOR2xp33_ASAP7_75t_L      g14308(.A(new_n14564), .B(new_n14562), .Y(new_n14565));
  XNOR2x2_ASAP7_75t_L       g14309(.A(new_n14441), .B(new_n14565), .Y(new_n14566));
  XNOR2x2_ASAP7_75t_L       g14310(.A(new_n14566), .B(new_n14431), .Y(new_n14567));
  AOI21xp33_ASAP7_75t_L     g14311(.A1(new_n14426), .A2(new_n14424), .B(new_n14567), .Y(new_n14568));
  INVx1_ASAP7_75t_L         g14312(.A(new_n14424), .Y(new_n14569));
  XOR2x2_ASAP7_75t_L        g14313(.A(new_n14441), .B(new_n14565), .Y(new_n14570));
  XNOR2x2_ASAP7_75t_L       g14314(.A(new_n14570), .B(new_n14431), .Y(new_n14571));
  NOR3xp33_ASAP7_75t_L      g14315(.A(new_n14571), .B(new_n14425), .C(new_n14569), .Y(new_n14572));
  NOR2xp33_ASAP7_75t_L      g14316(.A(new_n14568), .B(new_n14572), .Y(new_n14573));
  NAND2xp33_ASAP7_75t_L     g14317(.A(new_n14233), .B(new_n14231), .Y(new_n14574));
  AOI22xp33_ASAP7_75t_L     g14318(.A1(new_n1410), .A2(\b[52] ), .B1(\b[53] ), .B2(new_n1406), .Y(new_n14575));
  OAI221xp5_ASAP7_75t_L     g14319(.A1(new_n1549), .A2(new_n8249), .B1(new_n1411), .B2(new_n8888), .C(new_n14575), .Y(new_n14576));
  NOR2xp33_ASAP7_75t_L      g14320(.A(new_n1401), .B(new_n14576), .Y(new_n14577));
  AND2x2_ASAP7_75t_L        g14321(.A(new_n1401), .B(new_n14576), .Y(new_n14578));
  NOR2xp33_ASAP7_75t_L      g14322(.A(new_n14577), .B(new_n14578), .Y(new_n14579));
  INVx1_ASAP7_75t_L         g14323(.A(new_n14579), .Y(new_n14580));
  O2A1O1Ixp33_ASAP7_75t_L   g14324(.A1(new_n14235), .A2(new_n14380), .B(new_n14574), .C(new_n14580), .Y(new_n14581));
  OAI21xp33_ASAP7_75t_L     g14325(.A1(new_n14235), .A2(new_n14380), .B(new_n14574), .Y(new_n14582));
  NOR2xp33_ASAP7_75t_L      g14326(.A(new_n14579), .B(new_n14582), .Y(new_n14583));
  NOR2xp33_ASAP7_75t_L      g14327(.A(new_n14581), .B(new_n14583), .Y(new_n14584));
  XNOR2x2_ASAP7_75t_L       g14328(.A(new_n14584), .B(new_n14573), .Y(new_n14585));
  XNOR2x2_ASAP7_75t_L       g14329(.A(new_n14419), .B(new_n14585), .Y(new_n14586));
  AOI22xp33_ASAP7_75t_L     g14330(.A1(new_n826), .A2(\b[59] ), .B1(new_n823), .B2(new_n10887), .Y(new_n14587));
  OAI221xp5_ASAP7_75t_L     g14331(.A1(new_n994), .A2(new_n10848), .B1(new_n10488), .B2(new_n909), .C(new_n14587), .Y(new_n14588));
  XNOR2x2_ASAP7_75t_L       g14332(.A(\a[14] ), .B(new_n14588), .Y(new_n14589));
  NOR3xp33_ASAP7_75t_L      g14333(.A(new_n14382), .B(new_n14220), .C(new_n14219), .Y(new_n14590));
  NOR2xp33_ASAP7_75t_L      g14334(.A(new_n14220), .B(new_n14590), .Y(new_n14591));
  XNOR2x2_ASAP7_75t_L       g14335(.A(new_n14589), .B(new_n14591), .Y(new_n14592));
  XOR2x2_ASAP7_75t_L        g14336(.A(new_n14586), .B(new_n14592), .Y(new_n14593));
  NAND2xp33_ASAP7_75t_L     g14337(.A(new_n14413), .B(new_n14593), .Y(new_n14594));
  NOR2xp33_ASAP7_75t_L      g14338(.A(new_n14413), .B(new_n14593), .Y(new_n14595));
  INVx1_ASAP7_75t_L         g14339(.A(new_n14595), .Y(new_n14596));
  A2O1A1Ixp33_ASAP7_75t_L   g14340(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n448), .Y(new_n14597));
  A2O1A1Ixp33_ASAP7_75t_L   g14341(.A1(new_n14597), .A2(new_n481), .B(new_n12599), .C(\a[8] ), .Y(new_n14598));
  O2A1O1Ixp33_ASAP7_75t_L   g14342(.A1(new_n482), .A2(new_n13934), .B(new_n481), .C(new_n12599), .Y(new_n14599));
  NAND2xp33_ASAP7_75t_L     g14343(.A(new_n445), .B(new_n14599), .Y(new_n14600));
  AND2x2_ASAP7_75t_L        g14344(.A(new_n14600), .B(new_n14598), .Y(new_n14601));
  O2A1O1Ixp33_ASAP7_75t_L   g14345(.A1(new_n14202), .A2(new_n14203), .B(new_n14387), .C(new_n14601), .Y(new_n14602));
  INVx1_ASAP7_75t_L         g14346(.A(new_n14602), .Y(new_n14603));
  AOI21xp33_ASAP7_75t_L     g14347(.A1(new_n14386), .A2(new_n14204), .B(new_n14205), .Y(new_n14604));
  NAND2xp33_ASAP7_75t_L     g14348(.A(new_n14601), .B(new_n14604), .Y(new_n14605));
  NAND4xp25_ASAP7_75t_L     g14349(.A(new_n14596), .B(new_n14594), .C(new_n14603), .D(new_n14605), .Y(new_n14606));
  INVx1_ASAP7_75t_L         g14350(.A(new_n14594), .Y(new_n14607));
  INVx1_ASAP7_75t_L         g14351(.A(new_n14605), .Y(new_n14608));
  OAI22xp33_ASAP7_75t_L     g14352(.A1(new_n14607), .A2(new_n14595), .B1(new_n14608), .B2(new_n14602), .Y(new_n14609));
  AOI21xp33_ASAP7_75t_L     g14353(.A1(new_n14389), .A2(new_n14197), .B(new_n14198), .Y(new_n14610));
  AND3x1_ASAP7_75t_L        g14354(.A(new_n14609), .B(new_n14606), .C(new_n14610), .Y(new_n14611));
  AOI21xp33_ASAP7_75t_L     g14355(.A1(new_n14609), .A2(new_n14606), .B(new_n14610), .Y(new_n14612));
  NOR2xp33_ASAP7_75t_L      g14356(.A(new_n14612), .B(new_n14611), .Y(new_n14613));
  A2O1A1Ixp33_ASAP7_75t_L   g14357(.A1(new_n14398), .A2(new_n14395), .B(new_n14402), .C(new_n14613), .Y(new_n14614));
  INVx1_ASAP7_75t_L         g14358(.A(new_n14614), .Y(new_n14615));
  A2O1A1Ixp33_ASAP7_75t_L   g14359(.A1(new_n14184), .A2(new_n14180), .B(new_n14396), .C(new_n14401), .Y(new_n14616));
  NOR2xp33_ASAP7_75t_L      g14360(.A(new_n14613), .B(new_n14616), .Y(new_n14617));
  NOR2xp33_ASAP7_75t_L      g14361(.A(new_n14615), .B(new_n14617), .Y(\f[71] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14362(.A1(new_n14598), .A2(new_n14600), .B(new_n14604), .C(new_n14606), .Y(new_n14619));
  NAND2xp33_ASAP7_75t_L     g14363(.A(\b[63] ), .B(new_n600), .Y(new_n14620));
  A2O1A1Ixp33_ASAP7_75t_L   g14364(.A1(new_n12607), .A2(new_n12603), .B(new_n675), .C(new_n14620), .Y(new_n14621));
  AOI221xp5_ASAP7_75t_L     g14365(.A1(\b[61] ), .A2(new_n674), .B1(\b[62] ), .B2(new_n590), .C(new_n14621), .Y(new_n14622));
  XNOR2x2_ASAP7_75t_L       g14366(.A(new_n594), .B(new_n14622), .Y(new_n14623));
  INVx1_ASAP7_75t_L         g14367(.A(new_n14623), .Y(new_n14624));
  O2A1O1Ixp33_ASAP7_75t_L   g14368(.A1(new_n14411), .A2(new_n14407), .B(new_n14594), .C(new_n14624), .Y(new_n14625));
  O2A1O1Ixp33_ASAP7_75t_L   g14369(.A1(new_n14213), .A2(new_n14383), .B(new_n14211), .C(new_n14407), .Y(new_n14626));
  INVx1_ASAP7_75t_L         g14370(.A(new_n14626), .Y(new_n14627));
  NAND3xp33_ASAP7_75t_L     g14371(.A(new_n14594), .B(new_n14627), .C(new_n14624), .Y(new_n14628));
  INVx1_ASAP7_75t_L         g14372(.A(new_n14628), .Y(new_n14629));
  MAJIxp5_ASAP7_75t_L       g14373(.A(new_n14586), .B(new_n14589), .C(new_n14591), .Y(new_n14630));
  INVx1_ASAP7_75t_L         g14374(.A(new_n14630), .Y(new_n14631));
  AOI22xp33_ASAP7_75t_L     g14375(.A1(new_n826), .A2(\b[60] ), .B1(new_n823), .B2(new_n11234), .Y(new_n14632));
  OAI221xp5_ASAP7_75t_L     g14376(.A1(new_n994), .A2(new_n10881), .B1(new_n10848), .B2(new_n909), .C(new_n14632), .Y(new_n14633));
  XNOR2x2_ASAP7_75t_L       g14377(.A(\a[14] ), .B(new_n14633), .Y(new_n14634));
  INVx1_ASAP7_75t_L         g14378(.A(new_n14634), .Y(new_n14635));
  NOR2xp33_ASAP7_75t_L      g14379(.A(new_n14635), .B(new_n14631), .Y(new_n14636));
  INVx1_ASAP7_75t_L         g14380(.A(new_n14636), .Y(new_n14637));
  NOR2xp33_ASAP7_75t_L      g14381(.A(new_n14634), .B(new_n14630), .Y(new_n14638));
  INVx1_ASAP7_75t_L         g14382(.A(new_n14638), .Y(new_n14639));
  AOI22xp33_ASAP7_75t_L     g14383(.A1(new_n1113), .A2(\b[57] ), .B1(new_n1110), .B2(new_n10495), .Y(new_n14640));
  OAI221xp5_ASAP7_75t_L     g14384(.A1(new_n1298), .A2(new_n10178), .B1(new_n9534), .B2(new_n1195), .C(new_n14640), .Y(new_n14641));
  XNOR2x2_ASAP7_75t_L       g14385(.A(\a[17] ), .B(new_n14641), .Y(new_n14642));
  INVx1_ASAP7_75t_L         g14386(.A(new_n14418), .Y(new_n14643));
  MAJIxp5_ASAP7_75t_L       g14387(.A(new_n14585), .B(new_n14417), .C(new_n14643), .Y(new_n14644));
  NAND2xp33_ASAP7_75t_L     g14388(.A(new_n14642), .B(new_n14644), .Y(new_n14645));
  INVx1_ASAP7_75t_L         g14389(.A(new_n14645), .Y(new_n14646));
  NOR2xp33_ASAP7_75t_L      g14390(.A(new_n14642), .B(new_n14644), .Y(new_n14647));
  NOR3xp33_ASAP7_75t_L      g14391(.A(new_n14584), .B(new_n14572), .C(new_n14568), .Y(new_n14648));
  AOI22xp33_ASAP7_75t_L     g14392(.A1(new_n1406), .A2(\b[54] ), .B1(new_n1404), .B2(new_n9208), .Y(new_n14649));
  OAI221xp5_ASAP7_75t_L     g14393(.A1(new_n1398), .A2(new_n8882), .B1(new_n8569), .B2(new_n1549), .C(new_n14649), .Y(new_n14650));
  XNOR2x2_ASAP7_75t_L       g14394(.A(\a[20] ), .B(new_n14650), .Y(new_n14651));
  A2O1A1Ixp33_ASAP7_75t_L   g14395(.A1(new_n14580), .A2(new_n14582), .B(new_n14648), .C(new_n14651), .Y(new_n14652));
  O2A1O1Ixp33_ASAP7_75t_L   g14396(.A1(new_n14235), .A2(new_n14380), .B(new_n14574), .C(new_n14579), .Y(new_n14653));
  O2A1O1Ixp33_ASAP7_75t_L   g14397(.A1(new_n14581), .A2(new_n14583), .B(new_n14573), .C(new_n14653), .Y(new_n14654));
  INVx1_ASAP7_75t_L         g14398(.A(new_n14651), .Y(new_n14655));
  NAND2xp33_ASAP7_75t_L     g14399(.A(new_n14655), .B(new_n14654), .Y(new_n14656));
  AOI22xp33_ASAP7_75t_L     g14400(.A1(new_n1766), .A2(\b[51] ), .B1(new_n1764), .B2(new_n8257), .Y(new_n14657));
  OAI221xp5_ASAP7_75t_L     g14401(.A1(new_n1758), .A2(new_n8228), .B1(new_n7907), .B2(new_n1911), .C(new_n14657), .Y(new_n14658));
  XNOR2x2_ASAP7_75t_L       g14402(.A(new_n1761), .B(new_n14658), .Y(new_n14659));
  A2O1A1Ixp33_ASAP7_75t_L   g14403(.A1(new_n14567), .A2(new_n14424), .B(new_n14425), .C(new_n14659), .Y(new_n14660));
  INVx1_ASAP7_75t_L         g14404(.A(new_n14660), .Y(new_n14661));
  NOR3xp33_ASAP7_75t_L      g14405(.A(new_n14572), .B(new_n14659), .C(new_n14425), .Y(new_n14662));
  AOI22xp33_ASAP7_75t_L     g14406(.A1(new_n2228), .A2(\b[48] ), .B1(new_n2226), .B2(new_n7341), .Y(new_n14663));
  OAI221xp5_ASAP7_75t_L     g14407(.A1(new_n2220), .A2(new_n7316), .B1(new_n7033), .B2(new_n2387), .C(new_n14663), .Y(new_n14664));
  XNOR2x2_ASAP7_75t_L       g14408(.A(\a[26] ), .B(new_n14664), .Y(new_n14665));
  INVx1_ASAP7_75t_L         g14409(.A(new_n14429), .Y(new_n14666));
  MAJIxp5_ASAP7_75t_L       g14410(.A(new_n14570), .B(new_n14666), .C(new_n14430), .Y(new_n14667));
  XOR2x2_ASAP7_75t_L        g14411(.A(new_n14665), .B(new_n14667), .Y(new_n14668));
  AOI211xp5_ASAP7_75t_L     g14412(.A1(new_n14440), .A2(new_n14438), .B(new_n14564), .C(new_n14562), .Y(new_n14669));
  O2A1O1Ixp33_ASAP7_75t_L   g14413(.A1(new_n14434), .A2(new_n14435), .B(new_n14437), .C(new_n14669), .Y(new_n14670));
  AOI22xp33_ASAP7_75t_L     g14414(.A1(new_n2702), .A2(\b[45] ), .B1(new_n2700), .B2(new_n6764), .Y(new_n14671));
  OAI221xp5_ASAP7_75t_L     g14415(.A1(new_n2694), .A2(new_n6220), .B1(new_n6195), .B2(new_n2932), .C(new_n14671), .Y(new_n14672));
  XNOR2x2_ASAP7_75t_L       g14416(.A(\a[29] ), .B(new_n14672), .Y(new_n14673));
  INVx1_ASAP7_75t_L         g14417(.A(new_n14673), .Y(new_n14674));
  NOR2xp33_ASAP7_75t_L      g14418(.A(new_n14674), .B(new_n14670), .Y(new_n14675));
  AO21x2_ASAP7_75t_L        g14419(.A1(new_n14439), .A2(new_n14437), .B(new_n14669), .Y(new_n14676));
  NOR2xp33_ASAP7_75t_L      g14420(.A(new_n14673), .B(new_n14676), .Y(new_n14677));
  INVx1_ASAP7_75t_L         g14421(.A(new_n14450), .Y(new_n14678));
  AOI22xp33_ASAP7_75t_L     g14422(.A1(new_n3256), .A2(\b[42] ), .B1(new_n3254), .B2(new_n5688), .Y(new_n14679));
  OAI221xp5_ASAP7_75t_L     g14423(.A1(new_n3248), .A2(new_n5666), .B1(new_n5186), .B2(new_n3492), .C(new_n14679), .Y(new_n14680));
  XNOR2x2_ASAP7_75t_L       g14424(.A(\a[32] ), .B(new_n14680), .Y(new_n14681));
  INVx1_ASAP7_75t_L         g14425(.A(new_n14681), .Y(new_n14682));
  O2A1O1Ixp33_ASAP7_75t_L   g14426(.A1(new_n14448), .A2(new_n14561), .B(new_n14678), .C(new_n14682), .Y(new_n14683));
  OAI211xp5_ASAP7_75t_L     g14427(.A1(new_n14448), .A2(new_n14561), .B(new_n14682), .C(new_n14678), .Y(new_n14684));
  INVx1_ASAP7_75t_L         g14428(.A(new_n14684), .Y(new_n14685));
  AOI22xp33_ASAP7_75t_L     g14429(.A1(new_n4544), .A2(\b[36] ), .B1(new_n4542), .B2(new_n4473), .Y(new_n14686));
  OAI221xp5_ASAP7_75t_L     g14430(.A1(new_n4536), .A2(new_n4053), .B1(new_n3827), .B2(new_n4781), .C(new_n14686), .Y(new_n14687));
  XNOR2x2_ASAP7_75t_L       g14431(.A(\a[38] ), .B(new_n14687), .Y(new_n14688));
  AOI31xp33_ASAP7_75t_L     g14432(.A1(new_n14341), .A2(new_n14333), .A3(new_n14523), .B(new_n14530), .Y(new_n14689));
  AOI22xp33_ASAP7_75t_L     g14433(.A1(new_n5249), .A2(\b[33] ), .B1(new_n5247), .B2(new_n3813), .Y(new_n14690));
  OAI221xp5_ASAP7_75t_L     g14434(.A1(new_n5241), .A2(new_n3443), .B1(new_n3419), .B2(new_n5521), .C(new_n14690), .Y(new_n14691));
  XNOR2x2_ASAP7_75t_L       g14435(.A(\a[41] ), .B(new_n14691), .Y(new_n14692));
  INVx1_ASAP7_75t_L         g14436(.A(new_n14692), .Y(new_n14693));
  INVx1_ASAP7_75t_L         g14437(.A(new_n14514), .Y(new_n14694));
  INVx1_ASAP7_75t_L         g14438(.A(new_n14498), .Y(new_n14695));
  OAI21xp33_ASAP7_75t_L     g14439(.A1(new_n14695), .A2(new_n14499), .B(new_n14501), .Y(new_n14696));
  AOI22xp33_ASAP7_75t_L     g14440(.A1(new_n7659), .A2(\b[24] ), .B1(new_n7656), .B2(new_n2027), .Y(new_n14697));
  OAI221xp5_ASAP7_75t_L     g14441(.A1(new_n8326), .A2(new_n1995), .B1(new_n1857), .B2(new_n7994), .C(new_n14697), .Y(new_n14698));
  XNOR2x2_ASAP7_75t_L       g14442(.A(\a[50] ), .B(new_n14698), .Y(new_n14699));
  INVx1_ASAP7_75t_L         g14443(.A(new_n14487), .Y(new_n14700));
  NAND2xp33_ASAP7_75t_L     g14444(.A(new_n14475), .B(new_n14477), .Y(new_n14701));
  AOI22xp33_ASAP7_75t_L     g14445(.A1(new_n11656), .A2(\b[12] ), .B1(new_n11654), .B2(new_n970), .Y(new_n14702));
  OAI221xp5_ASAP7_75t_L     g14446(.A1(new_n12364), .A2(new_n695), .B1(new_n631), .B2(new_n13003), .C(new_n14702), .Y(new_n14703));
  XNOR2x2_ASAP7_75t_L       g14447(.A(\a[62] ), .B(new_n14703), .Y(new_n14704));
  NOR2xp33_ASAP7_75t_L      g14448(.A(new_n503), .B(new_n12671), .Y(new_n14705));
  O2A1O1Ixp33_ASAP7_75t_L   g14449(.A1(new_n503), .A2(new_n12356), .B(new_n14467), .C(new_n445), .Y(new_n14706));
  AOI211xp5_ASAP7_75t_L     g14450(.A1(new_n12669), .A2(\b[8] ), .B(new_n14466), .C(\a[8] ), .Y(new_n14707));
  NOR2xp33_ASAP7_75t_L      g14451(.A(new_n14707), .B(new_n14706), .Y(new_n14708));
  INVx1_ASAP7_75t_L         g14452(.A(new_n14708), .Y(new_n14709));
  A2O1A1Ixp33_ASAP7_75t_L   g14453(.A1(new_n12669), .A2(\b[9] ), .B(new_n14705), .C(new_n14709), .Y(new_n14710));
  O2A1O1Ixp33_ASAP7_75t_L   g14454(.A1(new_n12353), .A2(new_n12355), .B(\b[9] ), .C(new_n14705), .Y(new_n14711));
  NAND2xp33_ASAP7_75t_L     g14455(.A(new_n14711), .B(new_n14708), .Y(new_n14712));
  AND2x2_ASAP7_75t_L        g14456(.A(new_n14712), .B(new_n14710), .Y(new_n14713));
  NAND2xp33_ASAP7_75t_L     g14457(.A(new_n14470), .B(new_n14465), .Y(new_n14714));
  OAI211xp5_ASAP7_75t_L     g14458(.A1(new_n14275), .A2(new_n14469), .B(new_n14714), .C(new_n14713), .Y(new_n14715));
  INVx1_ASAP7_75t_L         g14459(.A(new_n14713), .Y(new_n14716));
  A2O1A1Ixp33_ASAP7_75t_L   g14460(.A1(new_n14465), .A2(new_n14470), .B(new_n14468), .C(new_n14716), .Y(new_n14717));
  NAND3xp33_ASAP7_75t_L     g14461(.A(new_n14715), .B(new_n14704), .C(new_n14717), .Y(new_n14718));
  INVx1_ASAP7_75t_L         g14462(.A(new_n14704), .Y(new_n14719));
  NAND2xp33_ASAP7_75t_L     g14463(.A(new_n14717), .B(new_n14715), .Y(new_n14720));
  NAND2xp33_ASAP7_75t_L     g14464(.A(new_n14719), .B(new_n14720), .Y(new_n14721));
  NAND2xp33_ASAP7_75t_L     g14465(.A(new_n14718), .B(new_n14721), .Y(new_n14722));
  AOI22xp33_ASAP7_75t_L     g14466(.A1(new_n10594), .A2(\b[15] ), .B1(new_n10591), .B2(new_n959), .Y(new_n14723));
  OAI221xp5_ASAP7_75t_L     g14467(.A1(new_n11335), .A2(new_n871), .B1(new_n793), .B2(new_n11330), .C(new_n14723), .Y(new_n14724));
  XNOR2x2_ASAP7_75t_L       g14468(.A(\a[59] ), .B(new_n14724), .Y(new_n14725));
  INVx1_ASAP7_75t_L         g14469(.A(new_n14725), .Y(new_n14726));
  NAND2xp33_ASAP7_75t_L     g14470(.A(new_n14726), .B(new_n14722), .Y(new_n14727));
  NAND3xp33_ASAP7_75t_L     g14471(.A(new_n14725), .B(new_n14721), .C(new_n14718), .Y(new_n14728));
  NAND3xp33_ASAP7_75t_L     g14472(.A(new_n14701), .B(new_n14727), .C(new_n14728), .Y(new_n14729));
  INVx1_ASAP7_75t_L         g14473(.A(new_n14729), .Y(new_n14730));
  AOI21xp33_ASAP7_75t_L     g14474(.A1(new_n14728), .A2(new_n14727), .B(new_n14701), .Y(new_n14731));
  NOR2xp33_ASAP7_75t_L      g14475(.A(new_n14731), .B(new_n14730), .Y(new_n14732));
  AOI22xp33_ASAP7_75t_L     g14476(.A1(new_n9623), .A2(\b[18] ), .B1(new_n9620), .B2(new_n1363), .Y(new_n14733));
  OAI221xp5_ASAP7_75t_L     g14477(.A1(new_n10280), .A2(new_n1244), .B1(new_n1051), .B2(new_n12010), .C(new_n14733), .Y(new_n14734));
  XNOR2x2_ASAP7_75t_L       g14478(.A(\a[56] ), .B(new_n14734), .Y(new_n14735));
  XNOR2x2_ASAP7_75t_L       g14479(.A(new_n14735), .B(new_n14732), .Y(new_n14736));
  A2O1A1O1Ixp25_ASAP7_75t_L g14480(.A1(new_n14294), .A2(new_n14290), .B(new_n14480), .C(new_n14700), .D(new_n14736), .Y(new_n14737));
  INVx1_ASAP7_75t_L         g14481(.A(new_n14737), .Y(new_n14738));
  NAND3xp33_ASAP7_75t_L     g14482(.A(new_n14736), .B(new_n14700), .C(new_n14482), .Y(new_n14739));
  NAND2xp33_ASAP7_75t_L     g14483(.A(new_n14739), .B(new_n14738), .Y(new_n14740));
  AOI22xp33_ASAP7_75t_L     g14484(.A1(new_n8645), .A2(\b[21] ), .B1(new_n8642), .B2(new_n1715), .Y(new_n14741));
  OAI221xp5_ASAP7_75t_L     g14485(.A1(new_n9322), .A2(new_n1594), .B1(new_n1493), .B2(new_n8965), .C(new_n14741), .Y(new_n14742));
  XNOR2x2_ASAP7_75t_L       g14486(.A(\a[53] ), .B(new_n14742), .Y(new_n14743));
  XNOR2x2_ASAP7_75t_L       g14487(.A(new_n14743), .B(new_n14740), .Y(new_n14744));
  INVx1_ASAP7_75t_L         g14488(.A(new_n14488), .Y(new_n14745));
  NAND2xp33_ASAP7_75t_L     g14489(.A(new_n14300), .B(new_n14305), .Y(new_n14746));
  INVx1_ASAP7_75t_L         g14490(.A(new_n14493), .Y(new_n14747));
  NAND2xp33_ASAP7_75t_L     g14491(.A(new_n14497), .B(new_n14747), .Y(new_n14748));
  A2O1A1Ixp33_ASAP7_75t_L   g14492(.A1(new_n14745), .A2(new_n14700), .B(new_n14746), .C(new_n14748), .Y(new_n14749));
  XNOR2x2_ASAP7_75t_L       g14493(.A(new_n14744), .B(new_n14749), .Y(new_n14750));
  XNOR2x2_ASAP7_75t_L       g14494(.A(new_n14699), .B(new_n14750), .Y(new_n14751));
  XNOR2x2_ASAP7_75t_L       g14495(.A(new_n14696), .B(new_n14751), .Y(new_n14752));
  AOI22xp33_ASAP7_75t_L     g14496(.A1(new_n6822), .A2(\b[27] ), .B1(new_n6819), .B2(new_n2657), .Y(new_n14753));
  OAI221xp5_ASAP7_75t_L     g14497(.A1(new_n7392), .A2(new_n2477), .B1(new_n2180), .B2(new_n7115), .C(new_n14753), .Y(new_n14754));
  XNOR2x2_ASAP7_75t_L       g14498(.A(\a[47] ), .B(new_n14754), .Y(new_n14755));
  XNOR2x2_ASAP7_75t_L       g14499(.A(new_n14755), .B(new_n14752), .Y(new_n14756));
  MAJx2_ASAP7_75t_L         g14500(.A(new_n14504), .B(new_n14509), .C(new_n14505), .Y(new_n14757));
  XOR2x2_ASAP7_75t_L        g14501(.A(new_n14757), .B(new_n14756), .Y(new_n14758));
  AOI22xp33_ASAP7_75t_L     g14502(.A1(new_n6002), .A2(\b[30] ), .B1(new_n5999), .B2(new_n3219), .Y(new_n14759));
  OAI221xp5_ASAP7_75t_L     g14503(.A1(new_n6544), .A2(new_n2871), .B1(new_n2852), .B2(new_n6309), .C(new_n14759), .Y(new_n14760));
  XNOR2x2_ASAP7_75t_L       g14504(.A(new_n5996), .B(new_n14760), .Y(new_n14761));
  NAND2xp33_ASAP7_75t_L     g14505(.A(new_n14761), .B(new_n14758), .Y(new_n14762));
  OR2x4_ASAP7_75t_L         g14506(.A(new_n14761), .B(new_n14758), .Y(new_n14763));
  NAND4xp25_ASAP7_75t_L     g14507(.A(new_n14763), .B(new_n14694), .C(new_n14520), .D(new_n14762), .Y(new_n14764));
  AO22x1_ASAP7_75t_L        g14508(.A1(new_n14694), .A2(new_n14520), .B1(new_n14762), .B2(new_n14763), .Y(new_n14765));
  AND2x2_ASAP7_75t_L        g14509(.A(new_n14764), .B(new_n14765), .Y(new_n14766));
  XNOR2x2_ASAP7_75t_L       g14510(.A(new_n14693), .B(new_n14766), .Y(new_n14767));
  NOR2xp33_ASAP7_75t_L      g14511(.A(new_n14689), .B(new_n14767), .Y(new_n14768));
  AND2x2_ASAP7_75t_L        g14512(.A(new_n14689), .B(new_n14767), .Y(new_n14769));
  NOR2xp33_ASAP7_75t_L      g14513(.A(new_n14768), .B(new_n14769), .Y(new_n14770));
  XNOR2x2_ASAP7_75t_L       g14514(.A(new_n14688), .B(new_n14770), .Y(new_n14771));
  O2A1O1Ixp33_ASAP7_75t_L   g14515(.A1(new_n14531), .A2(new_n14533), .B(new_n14548), .C(new_n14771), .Y(new_n14772));
  INVx1_ASAP7_75t_L         g14516(.A(new_n14688), .Y(new_n14773));
  NAND2xp33_ASAP7_75t_L     g14517(.A(new_n14773), .B(new_n14770), .Y(new_n14774));
  OAI21xp33_ASAP7_75t_L     g14518(.A1(new_n14768), .A2(new_n14769), .B(new_n14688), .Y(new_n14775));
  NAND2xp33_ASAP7_75t_L     g14519(.A(new_n14775), .B(new_n14774), .Y(new_n14776));
  NOR3xp33_ASAP7_75t_L      g14520(.A(new_n14776), .B(new_n14539), .C(new_n14542), .Y(new_n14777));
  NOR2xp33_ASAP7_75t_L      g14521(.A(new_n14777), .B(new_n14772), .Y(new_n14778));
  AOI22xp33_ASAP7_75t_L     g14522(.A1(new_n3884), .A2(\b[39] ), .B1(new_n3881), .B2(new_n5174), .Y(new_n14779));
  OAI221xp5_ASAP7_75t_L     g14523(.A1(new_n4312), .A2(new_n4915), .B1(new_n4701), .B2(new_n4986), .C(new_n14779), .Y(new_n14780));
  XNOR2x2_ASAP7_75t_L       g14524(.A(\a[35] ), .B(new_n14780), .Y(new_n14781));
  NAND2xp33_ASAP7_75t_L     g14525(.A(new_n14781), .B(new_n14778), .Y(new_n14782));
  INVx1_ASAP7_75t_L         g14526(.A(new_n14533), .Y(new_n14783));
  A2O1A1Ixp33_ASAP7_75t_L   g14527(.A1(new_n14783), .A2(new_n14540), .B(new_n14539), .C(new_n14776), .Y(new_n14784));
  O2A1O1Ixp33_ASAP7_75t_L   g14528(.A1(new_n14529), .A2(new_n14530), .B(new_n14783), .C(new_n14539), .Y(new_n14785));
  NAND2xp33_ASAP7_75t_L     g14529(.A(new_n14785), .B(new_n14771), .Y(new_n14786));
  NAND2xp33_ASAP7_75t_L     g14530(.A(new_n14786), .B(new_n14784), .Y(new_n14787));
  INVx1_ASAP7_75t_L         g14531(.A(new_n14781), .Y(new_n14788));
  NAND2xp33_ASAP7_75t_L     g14532(.A(new_n14788), .B(new_n14787), .Y(new_n14789));
  AOI21xp33_ASAP7_75t_L     g14533(.A1(new_n14547), .A2(new_n14555), .B(new_n14559), .Y(new_n14790));
  AO21x2_ASAP7_75t_L        g14534(.A1(new_n14789), .A2(new_n14782), .B(new_n14790), .Y(new_n14791));
  NAND3xp33_ASAP7_75t_L     g14535(.A(new_n14782), .B(new_n14789), .C(new_n14790), .Y(new_n14792));
  NAND2xp33_ASAP7_75t_L     g14536(.A(new_n14792), .B(new_n14791), .Y(new_n14793));
  OAI21xp33_ASAP7_75t_L     g14537(.A1(new_n14683), .A2(new_n14685), .B(new_n14793), .Y(new_n14794));
  NOR2xp33_ASAP7_75t_L      g14538(.A(new_n14683), .B(new_n14685), .Y(new_n14795));
  AND2x2_ASAP7_75t_L        g14539(.A(new_n14792), .B(new_n14791), .Y(new_n14796));
  NAND2xp33_ASAP7_75t_L     g14540(.A(new_n14796), .B(new_n14795), .Y(new_n14797));
  NAND2xp33_ASAP7_75t_L     g14541(.A(new_n14794), .B(new_n14797), .Y(new_n14798));
  OA21x2_ASAP7_75t_L        g14542(.A1(new_n14675), .A2(new_n14677), .B(new_n14798), .Y(new_n14799));
  NOR3xp33_ASAP7_75t_L      g14543(.A(new_n14798), .B(new_n14677), .C(new_n14675), .Y(new_n14800));
  NOR2xp33_ASAP7_75t_L      g14544(.A(new_n14800), .B(new_n14799), .Y(new_n14801));
  XOR2x2_ASAP7_75t_L        g14545(.A(new_n14668), .B(new_n14801), .Y(new_n14802));
  OAI21xp33_ASAP7_75t_L     g14546(.A1(new_n14662), .A2(new_n14661), .B(new_n14802), .Y(new_n14803));
  OR3x1_ASAP7_75t_L         g14547(.A(new_n14572), .B(new_n14425), .C(new_n14659), .Y(new_n14804));
  AND2x2_ASAP7_75t_L        g14548(.A(new_n14801), .B(new_n14668), .Y(new_n14805));
  NOR2xp33_ASAP7_75t_L      g14549(.A(new_n14668), .B(new_n14801), .Y(new_n14806));
  OAI211xp5_ASAP7_75t_L     g14550(.A1(new_n14805), .A2(new_n14806), .B(new_n14804), .C(new_n14660), .Y(new_n14807));
  AND2x2_ASAP7_75t_L        g14551(.A(new_n14803), .B(new_n14807), .Y(new_n14808));
  AOI21xp33_ASAP7_75t_L     g14552(.A1(new_n14656), .A2(new_n14652), .B(new_n14808), .Y(new_n14809));
  INVx1_ASAP7_75t_L         g14553(.A(new_n14652), .Y(new_n14810));
  MAJx2_ASAP7_75t_L         g14554(.A(new_n14573), .B(new_n14582), .C(new_n14580), .Y(new_n14811));
  NOR2xp33_ASAP7_75t_L      g14555(.A(new_n14651), .B(new_n14811), .Y(new_n14812));
  NAND2xp33_ASAP7_75t_L     g14556(.A(new_n14803), .B(new_n14807), .Y(new_n14813));
  NOR3xp33_ASAP7_75t_L      g14557(.A(new_n14813), .B(new_n14810), .C(new_n14812), .Y(new_n14814));
  OR2x4_ASAP7_75t_L         g14558(.A(new_n14814), .B(new_n14809), .Y(new_n14815));
  NOR3xp33_ASAP7_75t_L      g14559(.A(new_n14815), .B(new_n14647), .C(new_n14646), .Y(new_n14816));
  INVx1_ASAP7_75t_L         g14560(.A(new_n14647), .Y(new_n14817));
  NOR2xp33_ASAP7_75t_L      g14561(.A(new_n14814), .B(new_n14809), .Y(new_n14818));
  AOI21xp33_ASAP7_75t_L     g14562(.A1(new_n14817), .A2(new_n14645), .B(new_n14818), .Y(new_n14819));
  NOR2xp33_ASAP7_75t_L      g14563(.A(new_n14819), .B(new_n14816), .Y(new_n14820));
  AOI21xp33_ASAP7_75t_L     g14564(.A1(new_n14639), .A2(new_n14637), .B(new_n14820), .Y(new_n14821));
  NAND3xp33_ASAP7_75t_L     g14565(.A(new_n14818), .B(new_n14817), .C(new_n14645), .Y(new_n14822));
  OAI21xp33_ASAP7_75t_L     g14566(.A1(new_n14646), .A2(new_n14647), .B(new_n14815), .Y(new_n14823));
  NAND2xp33_ASAP7_75t_L     g14567(.A(new_n14822), .B(new_n14823), .Y(new_n14824));
  NOR3xp33_ASAP7_75t_L      g14568(.A(new_n14824), .B(new_n14638), .C(new_n14636), .Y(new_n14825));
  OAI22xp33_ASAP7_75t_L     g14569(.A1(new_n14629), .A2(new_n14625), .B1(new_n14825), .B2(new_n14821), .Y(new_n14826));
  INVx1_ASAP7_75t_L         g14570(.A(new_n14625), .Y(new_n14827));
  NOR2xp33_ASAP7_75t_L      g14571(.A(new_n14825), .B(new_n14821), .Y(new_n14828));
  NAND3xp33_ASAP7_75t_L     g14572(.A(new_n14828), .B(new_n14628), .C(new_n14827), .Y(new_n14829));
  NAND3xp33_ASAP7_75t_L     g14573(.A(new_n14829), .B(new_n14826), .C(new_n14619), .Y(new_n14830));
  AO21x2_ASAP7_75t_L        g14574(.A1(new_n14826), .A2(new_n14829), .B(new_n14619), .Y(new_n14831));
  NAND2xp33_ASAP7_75t_L     g14575(.A(new_n14830), .B(new_n14831), .Y(new_n14832));
  INVx1_ASAP7_75t_L         g14576(.A(new_n14832), .Y(new_n14833));
  A2O1A1Ixp33_ASAP7_75t_L   g14577(.A1(new_n14616), .A2(new_n14613), .B(new_n14611), .C(new_n14833), .Y(new_n14834));
  A2O1A1O1Ixp25_ASAP7_75t_L g14578(.A1(new_n14395), .A2(new_n14398), .B(new_n14402), .C(new_n14613), .D(new_n14611), .Y(new_n14835));
  NAND2xp33_ASAP7_75t_L     g14579(.A(new_n14832), .B(new_n14835), .Y(new_n14836));
  AND2x2_ASAP7_75t_L        g14580(.A(new_n14836), .B(new_n14834), .Y(\f[72] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14581(.A1(new_n14593), .A2(new_n14413), .B(new_n14626), .C(new_n14624), .Y(new_n14838));
  A2O1A1Ixp33_ASAP7_75t_L   g14582(.A1(new_n14628), .A2(new_n14827), .B(new_n14828), .C(new_n14838), .Y(new_n14839));
  NAND2xp33_ASAP7_75t_L     g14583(.A(new_n14635), .B(new_n14630), .Y(new_n14840));
  A2O1A1Ixp33_ASAP7_75t_L   g14584(.A1(new_n14637), .A2(new_n14639), .B(new_n14824), .C(new_n14840), .Y(new_n14841));
  AOI22xp33_ASAP7_75t_L     g14585(.A1(new_n590), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n674), .Y(new_n14842));
  A2O1A1Ixp33_ASAP7_75t_L   g14586(.A1(new_n13506), .A2(new_n13507), .B(new_n675), .C(new_n14842), .Y(new_n14843));
  NOR2xp33_ASAP7_75t_L      g14587(.A(new_n594), .B(new_n14843), .Y(new_n14844));
  A2O1A1O1Ixp25_ASAP7_75t_L g14588(.A1(new_n13507), .A2(new_n13506), .B(new_n675), .C(new_n14842), .D(\a[11] ), .Y(new_n14845));
  NOR2xp33_ASAP7_75t_L      g14589(.A(new_n14845), .B(new_n14844), .Y(new_n14846));
  XNOR2x2_ASAP7_75t_L       g14590(.A(new_n14846), .B(new_n14841), .Y(new_n14847));
  NAND2xp33_ASAP7_75t_L     g14591(.A(\b[61] ), .B(new_n826), .Y(new_n14848));
  OAI221xp5_ASAP7_75t_L     g14592(.A1(new_n11226), .A2(new_n994), .B1(new_n911), .B2(new_n11920), .C(new_n14848), .Y(new_n14849));
  AOI211xp5_ASAP7_75t_L     g14593(.A1(\b[59] ), .A2(new_n908), .B(new_n813), .C(new_n14849), .Y(new_n14850));
  INVx1_ASAP7_75t_L         g14594(.A(new_n14850), .Y(new_n14851));
  A2O1A1Ixp33_ASAP7_75t_L   g14595(.A1(\b[59] ), .A2(new_n908), .B(new_n14849), .C(new_n813), .Y(new_n14852));
  NAND2xp33_ASAP7_75t_L     g14596(.A(new_n14852), .B(new_n14851), .Y(new_n14853));
  NAND3xp33_ASAP7_75t_L     g14597(.A(new_n14822), .B(new_n14817), .C(new_n14853), .Y(new_n14854));
  O2A1O1Ixp33_ASAP7_75t_L   g14598(.A1(new_n14646), .A2(new_n14815), .B(new_n14817), .C(new_n14853), .Y(new_n14855));
  INVx1_ASAP7_75t_L         g14599(.A(new_n14855), .Y(new_n14856));
  A2O1A1Ixp33_ASAP7_75t_L   g14600(.A1(new_n14580), .A2(new_n14582), .B(new_n14648), .C(new_n14655), .Y(new_n14857));
  AOI22xp33_ASAP7_75t_L     g14601(.A1(new_n1103), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n1113), .Y(new_n14858));
  OAI221xp5_ASAP7_75t_L     g14602(.A1(new_n1195), .A2(new_n10178), .B1(new_n1197), .B2(new_n10856), .C(new_n14858), .Y(new_n14859));
  XNOR2x2_ASAP7_75t_L       g14603(.A(\a[17] ), .B(new_n14859), .Y(new_n14860));
  INVx1_ASAP7_75t_L         g14604(.A(new_n14860), .Y(new_n14861));
  A2O1A1O1Ixp25_ASAP7_75t_L g14605(.A1(new_n14656), .A2(new_n14652), .B(new_n14808), .C(new_n14857), .D(new_n14861), .Y(new_n14862));
  INVx1_ASAP7_75t_L         g14606(.A(new_n14862), .Y(new_n14863));
  INVx1_ASAP7_75t_L         g14607(.A(new_n14857), .Y(new_n14864));
  O2A1O1Ixp33_ASAP7_75t_L   g14608(.A1(new_n14812), .A2(new_n14810), .B(new_n14813), .C(new_n14864), .Y(new_n14865));
  NAND2xp33_ASAP7_75t_L     g14609(.A(new_n14861), .B(new_n14865), .Y(new_n14866));
  NAND2xp33_ASAP7_75t_L     g14610(.A(new_n14866), .B(new_n14863), .Y(new_n14867));
  AOI22xp33_ASAP7_75t_L     g14611(.A1(new_n1406), .A2(\b[55] ), .B1(new_n1404), .B2(new_n9542), .Y(new_n14868));
  OAI221xp5_ASAP7_75t_L     g14612(.A1(new_n1398), .A2(new_n9199), .B1(new_n8882), .B2(new_n1549), .C(new_n14868), .Y(new_n14869));
  XNOR2x2_ASAP7_75t_L       g14613(.A(\a[20] ), .B(new_n14869), .Y(new_n14870));
  O2A1O1Ixp33_ASAP7_75t_L   g14614(.A1(new_n14806), .A2(new_n14805), .B(new_n14660), .C(new_n14662), .Y(new_n14871));
  XOR2x2_ASAP7_75t_L        g14615(.A(new_n14870), .B(new_n14871), .Y(new_n14872));
  NOR2xp33_ASAP7_75t_L      g14616(.A(new_n14665), .B(new_n14667), .Y(new_n14873));
  AOI22xp33_ASAP7_75t_L     g14617(.A1(new_n1766), .A2(\b[52] ), .B1(new_n1764), .B2(new_n8577), .Y(new_n14874));
  OAI221xp5_ASAP7_75t_L     g14618(.A1(new_n1758), .A2(new_n8249), .B1(new_n8228), .B2(new_n1911), .C(new_n14874), .Y(new_n14875));
  XNOR2x2_ASAP7_75t_L       g14619(.A(\a[23] ), .B(new_n14875), .Y(new_n14876));
  INVx1_ASAP7_75t_L         g14620(.A(new_n14876), .Y(new_n14877));
  OR3x1_ASAP7_75t_L         g14621(.A(new_n14805), .B(new_n14873), .C(new_n14877), .Y(new_n14878));
  A2O1A1Ixp33_ASAP7_75t_L   g14622(.A1(new_n14801), .A2(new_n14668), .B(new_n14873), .C(new_n14877), .Y(new_n14879));
  AOI22xp33_ASAP7_75t_L     g14623(.A1(new_n2228), .A2(\b[49] ), .B1(new_n2226), .B2(new_n7914), .Y(new_n14880));
  OAI221xp5_ASAP7_75t_L     g14624(.A1(new_n2220), .A2(new_n7333), .B1(new_n7316), .B2(new_n2387), .C(new_n14880), .Y(new_n14881));
  XNOR2x2_ASAP7_75t_L       g14625(.A(\a[26] ), .B(new_n14881), .Y(new_n14882));
  NOR2xp33_ASAP7_75t_L      g14626(.A(new_n14673), .B(new_n14670), .Y(new_n14883));
  O2A1O1Ixp33_ASAP7_75t_L   g14627(.A1(new_n14675), .A2(new_n14677), .B(new_n14798), .C(new_n14883), .Y(new_n14884));
  XNOR2x2_ASAP7_75t_L       g14628(.A(new_n14882), .B(new_n14884), .Y(new_n14885));
  O2A1O1Ixp33_ASAP7_75t_L   g14629(.A1(new_n14448), .A2(new_n14561), .B(new_n14678), .C(new_n14681), .Y(new_n14886));
  O2A1O1Ixp33_ASAP7_75t_L   g14630(.A1(new_n14683), .A2(new_n14685), .B(new_n14796), .C(new_n14886), .Y(new_n14887));
  AOI22xp33_ASAP7_75t_L     g14631(.A1(new_n2706), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n2702), .Y(new_n14888));
  OAI221xp5_ASAP7_75t_L     g14632(.A1(new_n2932), .A2(new_n6220), .B1(new_n2707), .B2(new_n7887), .C(new_n14888), .Y(new_n14889));
  XNOR2x2_ASAP7_75t_L       g14633(.A(\a[29] ), .B(new_n14889), .Y(new_n14890));
  XNOR2x2_ASAP7_75t_L       g14634(.A(new_n14890), .B(new_n14887), .Y(new_n14891));
  AOI22xp33_ASAP7_75t_L     g14635(.A1(new_n3256), .A2(\b[43] ), .B1(new_n3254), .B2(new_n6202), .Y(new_n14892));
  OAI221xp5_ASAP7_75t_L     g14636(.A1(new_n3248), .A2(new_n5680), .B1(new_n5666), .B2(new_n3492), .C(new_n14892), .Y(new_n14893));
  XNOR2x2_ASAP7_75t_L       g14637(.A(\a[32] ), .B(new_n14893), .Y(new_n14894));
  INVx1_ASAP7_75t_L         g14638(.A(new_n14894), .Y(new_n14895));
  NAND2xp33_ASAP7_75t_L     g14639(.A(new_n14788), .B(new_n14778), .Y(new_n14896));
  A2O1A1Ixp33_ASAP7_75t_L   g14640(.A1(new_n14782), .A2(new_n14789), .B(new_n14790), .C(new_n14896), .Y(new_n14897));
  NOR2xp33_ASAP7_75t_L      g14641(.A(new_n14895), .B(new_n14897), .Y(new_n14898));
  A2O1A1O1Ixp25_ASAP7_75t_L g14642(.A1(new_n14789), .A2(new_n14782), .B(new_n14790), .C(new_n14896), .D(new_n14894), .Y(new_n14899));
  NOR2xp33_ASAP7_75t_L      g14643(.A(new_n14899), .B(new_n14898), .Y(new_n14900));
  AOI22xp33_ASAP7_75t_L     g14644(.A1(new_n3884), .A2(\b[40] ), .B1(new_n3881), .B2(new_n5194), .Y(new_n14901));
  OAI221xp5_ASAP7_75t_L     g14645(.A1(new_n4312), .A2(new_n5166), .B1(new_n4915), .B2(new_n4986), .C(new_n14901), .Y(new_n14902));
  XNOR2x2_ASAP7_75t_L       g14646(.A(\a[35] ), .B(new_n14902), .Y(new_n14903));
  NAND2xp33_ASAP7_75t_L     g14647(.A(new_n14774), .B(new_n14786), .Y(new_n14904));
  AOI22xp33_ASAP7_75t_L     g14648(.A1(new_n4544), .A2(\b[37] ), .B1(new_n4542), .B2(new_n4709), .Y(new_n14905));
  OAI221xp5_ASAP7_75t_L     g14649(.A1(new_n4536), .A2(new_n4465), .B1(new_n4053), .B2(new_n4781), .C(new_n14905), .Y(new_n14906));
  XNOR2x2_ASAP7_75t_L       g14650(.A(\a[38] ), .B(new_n14906), .Y(new_n14907));
  INVx1_ASAP7_75t_L         g14651(.A(new_n14907), .Y(new_n14908));
  AOI22xp33_ASAP7_75t_L     g14652(.A1(new_n5249), .A2(\b[34] ), .B1(new_n5247), .B2(new_n3833), .Y(new_n14909));
  OAI221xp5_ASAP7_75t_L     g14653(.A1(new_n5241), .A2(new_n3807), .B1(new_n3443), .B2(new_n5521), .C(new_n14909), .Y(new_n14910));
  XNOR2x2_ASAP7_75t_L       g14654(.A(\a[41] ), .B(new_n14910), .Y(new_n14911));
  AOI22xp33_ASAP7_75t_L     g14655(.A1(new_n10594), .A2(\b[16] ), .B1(new_n10591), .B2(new_n1058), .Y(new_n14912));
  OAI221xp5_ASAP7_75t_L     g14656(.A1(new_n11335), .A2(new_n952), .B1(new_n871), .B2(new_n11330), .C(new_n14912), .Y(new_n14913));
  XNOR2x2_ASAP7_75t_L       g14657(.A(\a[59] ), .B(new_n14913), .Y(new_n14914));
  NAND2xp33_ASAP7_75t_L     g14658(.A(new_n11654), .B(new_n800), .Y(new_n14915));
  OAI221xp5_ASAP7_75t_L     g14659(.A1(new_n12023), .A2(new_n793), .B1(new_n763), .B2(new_n12364), .C(new_n14915), .Y(new_n14916));
  AOI21xp33_ASAP7_75t_L     g14660(.A1(new_n12021), .A2(\b[11] ), .B(new_n14916), .Y(new_n14917));
  NAND2xp33_ASAP7_75t_L     g14661(.A(\a[62] ), .B(new_n14917), .Y(new_n14918));
  A2O1A1Ixp33_ASAP7_75t_L   g14662(.A1(\b[11] ), .A2(new_n12021), .B(new_n14916), .C(new_n11651), .Y(new_n14919));
  NAND2xp33_ASAP7_75t_L     g14663(.A(new_n14919), .B(new_n14918), .Y(new_n14920));
  NOR2xp33_ASAP7_75t_L      g14664(.A(new_n559), .B(new_n12671), .Y(new_n14921));
  O2A1O1Ixp33_ASAP7_75t_L   g14665(.A1(new_n12353), .A2(new_n12355), .B(\b[10] ), .C(new_n14921), .Y(new_n14922));
  INVx1_ASAP7_75t_L         g14666(.A(new_n14711), .Y(new_n14923));
  O2A1O1Ixp33_ASAP7_75t_L   g14667(.A1(new_n503), .A2(new_n12356), .B(new_n14467), .C(\a[8] ), .Y(new_n14924));
  O2A1O1Ixp33_ASAP7_75t_L   g14668(.A1(new_n14707), .A2(new_n14706), .B(new_n14923), .C(new_n14924), .Y(new_n14925));
  NAND2xp33_ASAP7_75t_L     g14669(.A(new_n14922), .B(new_n14925), .Y(new_n14926));
  INVx1_ASAP7_75t_L         g14670(.A(new_n14922), .Y(new_n14927));
  A2O1A1Ixp33_ASAP7_75t_L   g14671(.A1(new_n14709), .A2(new_n14923), .B(new_n14924), .C(new_n14927), .Y(new_n14928));
  AND2x2_ASAP7_75t_L        g14672(.A(new_n14926), .B(new_n14928), .Y(new_n14929));
  XNOR2x2_ASAP7_75t_L       g14673(.A(new_n14929), .B(new_n14920), .Y(new_n14930));
  NAND3xp33_ASAP7_75t_L     g14674(.A(new_n14930), .B(new_n14718), .C(new_n14717), .Y(new_n14931));
  O2A1O1Ixp33_ASAP7_75t_L   g14675(.A1(new_n14719), .A2(new_n14720), .B(new_n14717), .C(new_n14930), .Y(new_n14932));
  INVx1_ASAP7_75t_L         g14676(.A(new_n14932), .Y(new_n14933));
  NAND3xp33_ASAP7_75t_L     g14677(.A(new_n14933), .B(new_n14931), .C(new_n14914), .Y(new_n14934));
  AO21x2_ASAP7_75t_L        g14678(.A1(new_n14931), .A2(new_n14933), .B(new_n14914), .Y(new_n14935));
  NAND4xp25_ASAP7_75t_L     g14679(.A(new_n14935), .B(new_n14727), .C(new_n14729), .D(new_n14934), .Y(new_n14936));
  NAND2xp33_ASAP7_75t_L     g14680(.A(new_n14934), .B(new_n14935), .Y(new_n14937));
  A2O1A1Ixp33_ASAP7_75t_L   g14681(.A1(new_n14726), .A2(new_n14722), .B(new_n14730), .C(new_n14937), .Y(new_n14938));
  NAND2xp33_ASAP7_75t_L     g14682(.A(\b[19] ), .B(new_n9623), .Y(new_n14939));
  OAI221xp5_ASAP7_75t_L     g14683(.A1(new_n1356), .A2(new_n10280), .B1(new_n9949), .B2(new_n2793), .C(new_n14939), .Y(new_n14940));
  AOI21xp33_ASAP7_75t_L     g14684(.A1(new_n9948), .A2(\b[17] ), .B(new_n14940), .Y(new_n14941));
  NAND2xp33_ASAP7_75t_L     g14685(.A(\a[56] ), .B(new_n14941), .Y(new_n14942));
  A2O1A1Ixp33_ASAP7_75t_L   g14686(.A1(\b[17] ), .A2(new_n9948), .B(new_n14940), .C(new_n9610), .Y(new_n14943));
  AND2x2_ASAP7_75t_L        g14687(.A(new_n14943), .B(new_n14942), .Y(new_n14944));
  NAND3xp33_ASAP7_75t_L     g14688(.A(new_n14938), .B(new_n14936), .C(new_n14944), .Y(new_n14945));
  AO21x2_ASAP7_75t_L        g14689(.A1(new_n14936), .A2(new_n14938), .B(new_n14944), .Y(new_n14946));
  NAND2xp33_ASAP7_75t_L     g14690(.A(new_n14945), .B(new_n14946), .Y(new_n14947));
  OAI31xp33_ASAP7_75t_L     g14691(.A1(new_n14730), .A2(new_n14735), .A3(new_n14731), .B(new_n14739), .Y(new_n14948));
  OR2x4_ASAP7_75t_L         g14692(.A(new_n14947), .B(new_n14948), .Y(new_n14949));
  NAND2xp33_ASAP7_75t_L     g14693(.A(new_n14947), .B(new_n14948), .Y(new_n14950));
  AOI22xp33_ASAP7_75t_L     g14694(.A1(new_n8645), .A2(\b[22] ), .B1(new_n8642), .B2(new_n1864), .Y(new_n14951));
  OAI221xp5_ASAP7_75t_L     g14695(.A1(new_n9322), .A2(new_n1709), .B1(new_n1594), .B2(new_n8965), .C(new_n14951), .Y(new_n14952));
  XNOR2x2_ASAP7_75t_L       g14696(.A(\a[53] ), .B(new_n14952), .Y(new_n14953));
  AND3x1_ASAP7_75t_L        g14697(.A(new_n14949), .B(new_n14953), .C(new_n14950), .Y(new_n14954));
  AOI21xp33_ASAP7_75t_L     g14698(.A1(new_n14949), .A2(new_n14950), .B(new_n14953), .Y(new_n14955));
  INVx1_ASAP7_75t_L         g14699(.A(new_n14743), .Y(new_n14956));
  NAND3xp33_ASAP7_75t_L     g14700(.A(new_n14738), .B(new_n14739), .C(new_n14956), .Y(new_n14957));
  A2O1A1Ixp33_ASAP7_75t_L   g14701(.A1(new_n14748), .A2(new_n14492), .B(new_n14744), .C(new_n14957), .Y(new_n14958));
  OR3x1_ASAP7_75t_L         g14702(.A(new_n14958), .B(new_n14954), .C(new_n14955), .Y(new_n14959));
  OAI21xp33_ASAP7_75t_L     g14703(.A1(new_n14954), .A2(new_n14955), .B(new_n14958), .Y(new_n14960));
  NAND2xp33_ASAP7_75t_L     g14704(.A(new_n14960), .B(new_n14959), .Y(new_n14961));
  INVx1_ASAP7_75t_L         g14705(.A(new_n14961), .Y(new_n14962));
  AOI22xp33_ASAP7_75t_L     g14706(.A1(new_n7659), .A2(\b[25] ), .B1(new_n7656), .B2(new_n2188), .Y(new_n14963));
  OAI221xp5_ASAP7_75t_L     g14707(.A1(new_n8326), .A2(new_n2019), .B1(new_n1995), .B2(new_n7994), .C(new_n14963), .Y(new_n14964));
  XNOR2x2_ASAP7_75t_L       g14708(.A(\a[50] ), .B(new_n14964), .Y(new_n14965));
  NAND2xp33_ASAP7_75t_L     g14709(.A(new_n14965), .B(new_n14962), .Y(new_n14966));
  INVx1_ASAP7_75t_L         g14710(.A(new_n14965), .Y(new_n14967));
  NAND2xp33_ASAP7_75t_L     g14711(.A(new_n14967), .B(new_n14961), .Y(new_n14968));
  NAND2xp33_ASAP7_75t_L     g14712(.A(new_n14968), .B(new_n14966), .Y(new_n14969));
  INVx1_ASAP7_75t_L         g14713(.A(new_n14699), .Y(new_n14970));
  MAJIxp5_ASAP7_75t_L       g14714(.A(new_n14696), .B(new_n14970), .C(new_n14750), .Y(new_n14971));
  XNOR2x2_ASAP7_75t_L       g14715(.A(new_n14971), .B(new_n14969), .Y(new_n14972));
  AOI22xp33_ASAP7_75t_L     g14716(.A1(new_n6822), .A2(\b[28] ), .B1(new_n6819), .B2(new_n2858), .Y(new_n14973));
  OAI221xp5_ASAP7_75t_L     g14717(.A1(new_n7392), .A2(new_n2650), .B1(new_n2477), .B2(new_n7115), .C(new_n14973), .Y(new_n14974));
  XNOR2x2_ASAP7_75t_L       g14718(.A(\a[47] ), .B(new_n14974), .Y(new_n14975));
  NAND2xp33_ASAP7_75t_L     g14719(.A(new_n14975), .B(new_n14972), .Y(new_n14976));
  INVx1_ASAP7_75t_L         g14720(.A(new_n14969), .Y(new_n14977));
  NAND2xp33_ASAP7_75t_L     g14721(.A(new_n14971), .B(new_n14977), .Y(new_n14978));
  AND2x2_ASAP7_75t_L        g14722(.A(new_n14970), .B(new_n14750), .Y(new_n14979));
  A2O1A1Ixp33_ASAP7_75t_L   g14723(.A1(new_n14696), .A2(new_n14751), .B(new_n14979), .C(new_n14969), .Y(new_n14980));
  AO21x2_ASAP7_75t_L        g14724(.A1(new_n14978), .A2(new_n14980), .B(new_n14975), .Y(new_n14981));
  MAJx2_ASAP7_75t_L         g14725(.A(new_n14752), .B(new_n14755), .C(new_n14757), .Y(new_n14982));
  NAND3xp33_ASAP7_75t_L     g14726(.A(new_n14981), .B(new_n14976), .C(new_n14982), .Y(new_n14983));
  AO21x2_ASAP7_75t_L        g14727(.A1(new_n14976), .A2(new_n14981), .B(new_n14982), .Y(new_n14984));
  NAND2xp33_ASAP7_75t_L     g14728(.A(new_n14983), .B(new_n14984), .Y(new_n14985));
  AOI22xp33_ASAP7_75t_L     g14729(.A1(new_n6002), .A2(\b[31] ), .B1(new_n5999), .B2(new_n3426), .Y(new_n14986));
  OAI221xp5_ASAP7_75t_L     g14730(.A1(new_n6544), .A2(new_n3212), .B1(new_n2871), .B2(new_n6309), .C(new_n14986), .Y(new_n14987));
  XNOR2x2_ASAP7_75t_L       g14731(.A(\a[44] ), .B(new_n14987), .Y(new_n14988));
  XOR2x2_ASAP7_75t_L        g14732(.A(new_n14988), .B(new_n14985), .Y(new_n14989));
  NAND2xp33_ASAP7_75t_L     g14733(.A(new_n14762), .B(new_n14764), .Y(new_n14990));
  NAND2xp33_ASAP7_75t_L     g14734(.A(new_n14989), .B(new_n14990), .Y(new_n14991));
  INVx1_ASAP7_75t_L         g14735(.A(new_n14991), .Y(new_n14992));
  NOR2xp33_ASAP7_75t_L      g14736(.A(new_n14989), .B(new_n14990), .Y(new_n14993));
  NOR3xp33_ASAP7_75t_L      g14737(.A(new_n14992), .B(new_n14993), .C(new_n14911), .Y(new_n14994));
  INVx1_ASAP7_75t_L         g14738(.A(new_n14911), .Y(new_n14995));
  XOR2x2_ASAP7_75t_L        g14739(.A(new_n14989), .B(new_n14990), .Y(new_n14996));
  NOR2xp33_ASAP7_75t_L      g14740(.A(new_n14995), .B(new_n14996), .Y(new_n14997));
  NOR2xp33_ASAP7_75t_L      g14741(.A(new_n14994), .B(new_n14997), .Y(new_n14998));
  A2O1A1Ixp33_ASAP7_75t_L   g14742(.A1(new_n14766), .A2(new_n14693), .B(new_n14768), .C(new_n14998), .Y(new_n14999));
  AOI21xp33_ASAP7_75t_L     g14743(.A1(new_n14766), .A2(new_n14693), .B(new_n14768), .Y(new_n15000));
  OAI21xp33_ASAP7_75t_L     g14744(.A1(new_n14994), .A2(new_n14997), .B(new_n15000), .Y(new_n15001));
  AND2x2_ASAP7_75t_L        g14745(.A(new_n14999), .B(new_n15001), .Y(new_n15002));
  XNOR2x2_ASAP7_75t_L       g14746(.A(new_n14908), .B(new_n15002), .Y(new_n15003));
  XNOR2x2_ASAP7_75t_L       g14747(.A(new_n14904), .B(new_n15003), .Y(new_n15004));
  NOR2xp33_ASAP7_75t_L      g14748(.A(new_n14903), .B(new_n15004), .Y(new_n15005));
  AND3x1_ASAP7_75t_L        g14749(.A(new_n15001), .B(new_n14999), .C(new_n14908), .Y(new_n15006));
  NOR2xp33_ASAP7_75t_L      g14750(.A(new_n14908), .B(new_n15002), .Y(new_n15007));
  NOR2xp33_ASAP7_75t_L      g14751(.A(new_n15006), .B(new_n15007), .Y(new_n15008));
  A2O1A1Ixp33_ASAP7_75t_L   g14752(.A1(new_n14770), .A2(new_n14773), .B(new_n14777), .C(new_n15008), .Y(new_n15009));
  NAND3xp33_ASAP7_75t_L     g14753(.A(new_n15003), .B(new_n14786), .C(new_n14774), .Y(new_n15010));
  AND3x1_ASAP7_75t_L        g14754(.A(new_n15009), .B(new_n15010), .C(new_n14903), .Y(new_n15011));
  NOR2xp33_ASAP7_75t_L      g14755(.A(new_n15011), .B(new_n15005), .Y(new_n15012));
  XOR2x2_ASAP7_75t_L        g14756(.A(new_n15012), .B(new_n14900), .Y(new_n15013));
  XNOR2x2_ASAP7_75t_L       g14757(.A(new_n15013), .B(new_n14891), .Y(new_n15014));
  XOR2x2_ASAP7_75t_L        g14758(.A(new_n15014), .B(new_n14885), .Y(new_n15015));
  NAND3xp33_ASAP7_75t_L     g14759(.A(new_n14878), .B(new_n15015), .C(new_n14879), .Y(new_n15016));
  AO21x2_ASAP7_75t_L        g14760(.A1(new_n14879), .A2(new_n14878), .B(new_n15015), .Y(new_n15017));
  NAND2xp33_ASAP7_75t_L     g14761(.A(new_n15016), .B(new_n15017), .Y(new_n15018));
  XOR2x2_ASAP7_75t_L        g14762(.A(new_n14872), .B(new_n15018), .Y(new_n15019));
  XNOR2x2_ASAP7_75t_L       g14763(.A(new_n15019), .B(new_n14867), .Y(new_n15020));
  AOI21xp33_ASAP7_75t_L     g14764(.A1(new_n14854), .A2(new_n14856), .B(new_n15020), .Y(new_n15021));
  INVx1_ASAP7_75t_L         g14765(.A(new_n14854), .Y(new_n15022));
  XNOR2x2_ASAP7_75t_L       g14766(.A(new_n14872), .B(new_n15018), .Y(new_n15023));
  XNOR2x2_ASAP7_75t_L       g14767(.A(new_n15023), .B(new_n14867), .Y(new_n15024));
  NOR3xp33_ASAP7_75t_L      g14768(.A(new_n15024), .B(new_n15022), .C(new_n14855), .Y(new_n15025));
  NOR2xp33_ASAP7_75t_L      g14769(.A(new_n15021), .B(new_n15025), .Y(new_n15026));
  NAND2xp33_ASAP7_75t_L     g14770(.A(new_n15026), .B(new_n14847), .Y(new_n15027));
  INVx1_ASAP7_75t_L         g14771(.A(new_n14846), .Y(new_n15028));
  A2O1A1O1Ixp25_ASAP7_75t_L g14772(.A1(new_n14639), .A2(new_n14637), .B(new_n14824), .C(new_n14840), .D(new_n15028), .Y(new_n15029));
  NOR2xp33_ASAP7_75t_L      g14773(.A(new_n14846), .B(new_n14841), .Y(new_n15030));
  OR3x1_ASAP7_75t_L         g14774(.A(new_n15026), .B(new_n15029), .C(new_n15030), .Y(new_n15031));
  AND3x1_ASAP7_75t_L        g14775(.A(new_n15031), .B(new_n15027), .C(new_n14839), .Y(new_n15032));
  AOI21xp33_ASAP7_75t_L     g14776(.A1(new_n15031), .A2(new_n15027), .B(new_n14839), .Y(new_n15033));
  NOR2xp33_ASAP7_75t_L      g14777(.A(new_n15033), .B(new_n15032), .Y(new_n15034));
  INVx1_ASAP7_75t_L         g14778(.A(new_n15034), .Y(new_n15035));
  O2A1O1Ixp33_ASAP7_75t_L   g14779(.A1(new_n14835), .A2(new_n14832), .B(new_n14830), .C(new_n15035), .Y(new_n15036));
  INVx1_ASAP7_75t_L         g14780(.A(new_n14611), .Y(new_n15037));
  A2O1A1Ixp33_ASAP7_75t_L   g14781(.A1(new_n14614), .A2(new_n15037), .B(new_n14832), .C(new_n14830), .Y(new_n15038));
  NOR2xp33_ASAP7_75t_L      g14782(.A(new_n15034), .B(new_n15038), .Y(new_n15039));
  NOR2xp33_ASAP7_75t_L      g14783(.A(new_n15039), .B(new_n15036), .Y(\f[73] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14784(.A1(new_n14639), .A2(new_n14637), .B(new_n14824), .C(new_n14840), .D(new_n14846), .Y(new_n15041));
  AO21x2_ASAP7_75t_L        g14785(.A1(new_n15026), .A2(new_n14847), .B(new_n15041), .Y(new_n15042));
  A2O1A1O1Ixp25_ASAP7_75t_L g14786(.A1(new_n14656), .A2(new_n14652), .B(new_n14808), .C(new_n14857), .D(new_n14860), .Y(new_n15043));
  AOI22xp33_ASAP7_75t_L     g14787(.A1(new_n817), .A2(\b[61] ), .B1(\b[62] ), .B2(new_n826), .Y(new_n15044));
  OAI221xp5_ASAP7_75t_L     g14788(.A1(new_n909), .A2(new_n11226), .B1(new_n911), .B2(new_n12281), .C(new_n15044), .Y(new_n15045));
  XNOR2x2_ASAP7_75t_L       g14789(.A(\a[14] ), .B(new_n15045), .Y(new_n15046));
  INVx1_ASAP7_75t_L         g14790(.A(new_n15046), .Y(new_n15047));
  A2O1A1Ixp33_ASAP7_75t_L   g14791(.A1(new_n14867), .A2(new_n15019), .B(new_n15043), .C(new_n15047), .Y(new_n15048));
  A2O1A1Ixp33_ASAP7_75t_L   g14792(.A1(new_n14656), .A2(new_n14652), .B(new_n14808), .C(new_n14857), .Y(new_n15049));
  NOR2xp33_ASAP7_75t_L      g14793(.A(new_n14860), .B(new_n15049), .Y(new_n15050));
  O2A1O1Ixp33_ASAP7_75t_L   g14794(.A1(new_n14862), .A2(new_n15050), .B(new_n15019), .C(new_n15043), .Y(new_n15051));
  NAND2xp33_ASAP7_75t_L     g14795(.A(new_n15046), .B(new_n15051), .Y(new_n15052));
  NAND2xp33_ASAP7_75t_L     g14796(.A(new_n15048), .B(new_n15052), .Y(new_n15053));
  AOI22xp33_ASAP7_75t_L     g14797(.A1(new_n1113), .A2(\b[59] ), .B1(new_n1110), .B2(new_n10887), .Y(new_n15054));
  OAI221xp5_ASAP7_75t_L     g14798(.A1(new_n1298), .A2(new_n10848), .B1(new_n10488), .B2(new_n1195), .C(new_n15054), .Y(new_n15055));
  XNOR2x2_ASAP7_75t_L       g14799(.A(\a[17] ), .B(new_n15055), .Y(new_n15056));
  OAI21xp33_ASAP7_75t_L     g14800(.A1(new_n14661), .A2(new_n14802), .B(new_n14804), .Y(new_n15057));
  MAJx2_ASAP7_75t_L         g14801(.A(new_n15018), .B(new_n15057), .C(new_n14870), .Y(new_n15058));
  NAND2xp33_ASAP7_75t_L     g14802(.A(new_n15056), .B(new_n15058), .Y(new_n15059));
  OR2x4_ASAP7_75t_L         g14803(.A(new_n15056), .B(new_n15058), .Y(new_n15060));
  AOI22xp33_ASAP7_75t_L     g14804(.A1(new_n1406), .A2(\b[56] ), .B1(new_n1404), .B2(new_n10185), .Y(new_n15061));
  OAI221xp5_ASAP7_75t_L     g14805(.A1(new_n1398), .A2(new_n9534), .B1(new_n9199), .B2(new_n1549), .C(new_n15061), .Y(new_n15062));
  XNOR2x2_ASAP7_75t_L       g14806(.A(\a[20] ), .B(new_n15062), .Y(new_n15063));
  INVx1_ASAP7_75t_L         g14807(.A(new_n15063), .Y(new_n15064));
  NAND2xp33_ASAP7_75t_L     g14808(.A(new_n14668), .B(new_n14801), .Y(new_n15065));
  O2A1O1Ixp33_ASAP7_75t_L   g14809(.A1(new_n14665), .A2(new_n14667), .B(new_n15065), .C(new_n14876), .Y(new_n15066));
  AOI21xp33_ASAP7_75t_L     g14810(.A1(new_n14878), .A2(new_n15015), .B(new_n15066), .Y(new_n15067));
  NAND2xp33_ASAP7_75t_L     g14811(.A(new_n15064), .B(new_n15067), .Y(new_n15068));
  A2O1A1Ixp33_ASAP7_75t_L   g14812(.A1(new_n14878), .A2(new_n15015), .B(new_n15066), .C(new_n15063), .Y(new_n15069));
  NAND2xp33_ASAP7_75t_L     g14813(.A(new_n15069), .B(new_n15068), .Y(new_n15070));
  INVx1_ASAP7_75t_L         g14814(.A(new_n14882), .Y(new_n15071));
  NAND2xp33_ASAP7_75t_L     g14815(.A(new_n15071), .B(new_n14884), .Y(new_n15072));
  A2O1A1Ixp33_ASAP7_75t_L   g14816(.A1(new_n14674), .A2(new_n14676), .B(new_n14799), .C(new_n14882), .Y(new_n15073));
  A2O1A1Ixp33_ASAP7_75t_L   g14817(.A1(new_n14674), .A2(new_n14676), .B(new_n14799), .C(new_n15071), .Y(new_n15074));
  A2O1A1Ixp33_ASAP7_75t_L   g14818(.A1(new_n15073), .A2(new_n15072), .B(new_n15014), .C(new_n15074), .Y(new_n15075));
  AOI22xp33_ASAP7_75t_L     g14819(.A1(new_n1770), .A2(\b[52] ), .B1(\b[53] ), .B2(new_n1766), .Y(new_n15076));
  OAI221xp5_ASAP7_75t_L     g14820(.A1(new_n1911), .A2(new_n8249), .B1(new_n1771), .B2(new_n8888), .C(new_n15076), .Y(new_n15077));
  XNOR2x2_ASAP7_75t_L       g14821(.A(\a[23] ), .B(new_n15077), .Y(new_n15078));
  XNOR2x2_ASAP7_75t_L       g14822(.A(new_n15078), .B(new_n15075), .Y(new_n15079));
  MAJIxp5_ASAP7_75t_L       g14823(.A(new_n15013), .B(new_n14887), .C(new_n14890), .Y(new_n15080));
  AOI22xp33_ASAP7_75t_L     g14824(.A1(new_n2232), .A2(\b[49] ), .B1(\b[50] ), .B2(new_n2228), .Y(new_n15081));
  OAI221xp5_ASAP7_75t_L     g14825(.A1(new_n2387), .A2(new_n7333), .B1(new_n2233), .B2(new_n8234), .C(new_n15081), .Y(new_n15082));
  XNOR2x2_ASAP7_75t_L       g14826(.A(\a[26] ), .B(new_n15082), .Y(new_n15083));
  INVx1_ASAP7_75t_L         g14827(.A(new_n15083), .Y(new_n15084));
  AND2x2_ASAP7_75t_L        g14828(.A(new_n15084), .B(new_n15080), .Y(new_n15085));
  NOR2xp33_ASAP7_75t_L      g14829(.A(new_n15084), .B(new_n15080), .Y(new_n15086));
  NOR2xp33_ASAP7_75t_L      g14830(.A(new_n15086), .B(new_n15085), .Y(new_n15087));
  INVx1_ASAP7_75t_L         g14831(.A(new_n14899), .Y(new_n15088));
  AOI22xp33_ASAP7_75t_L     g14832(.A1(new_n2702), .A2(\b[47] ), .B1(new_n2700), .B2(new_n7323), .Y(new_n15089));
  OAI221xp5_ASAP7_75t_L     g14833(.A1(new_n2694), .A2(new_n7033), .B1(new_n6756), .B2(new_n2932), .C(new_n15089), .Y(new_n15090));
  XNOR2x2_ASAP7_75t_L       g14834(.A(\a[29] ), .B(new_n15090), .Y(new_n15091));
  A2O1A1Ixp33_ASAP7_75t_L   g14835(.A1(new_n15012), .A2(new_n15088), .B(new_n14898), .C(new_n15091), .Y(new_n15092));
  AOI211xp5_ASAP7_75t_L     g14836(.A1(new_n15012), .A2(new_n15088), .B(new_n15091), .C(new_n14898), .Y(new_n15093));
  INVx1_ASAP7_75t_L         g14837(.A(new_n15093), .Y(new_n15094));
  NAND2xp33_ASAP7_75t_L     g14838(.A(new_n15092), .B(new_n15094), .Y(new_n15095));
  AOI22xp33_ASAP7_75t_L     g14839(.A1(new_n3260), .A2(\b[43] ), .B1(\b[44] ), .B2(new_n3256), .Y(new_n15096));
  OAI221xp5_ASAP7_75t_L     g14840(.A1(new_n3492), .A2(new_n5680), .B1(new_n3261), .B2(new_n6229), .C(new_n15096), .Y(new_n15097));
  XNOR2x2_ASAP7_75t_L       g14841(.A(\a[32] ), .B(new_n15097), .Y(new_n15098));
  INVx1_ASAP7_75t_L         g14842(.A(new_n15098), .Y(new_n15099));
  INVx1_ASAP7_75t_L         g14843(.A(new_n15010), .Y(new_n15100));
  NOR2xp33_ASAP7_75t_L      g14844(.A(new_n15100), .B(new_n15011), .Y(new_n15101));
  NAND2xp33_ASAP7_75t_L     g14845(.A(new_n15099), .B(new_n15101), .Y(new_n15102));
  A2O1A1Ixp33_ASAP7_75t_L   g14846(.A1(new_n15009), .A2(new_n14903), .B(new_n15100), .C(new_n15098), .Y(new_n15103));
  NAND2xp33_ASAP7_75t_L     g14847(.A(new_n15103), .B(new_n15102), .Y(new_n15104));
  AOI22xp33_ASAP7_75t_L     g14848(.A1(new_n3884), .A2(\b[41] ), .B1(new_n3881), .B2(new_n5669), .Y(new_n15105));
  OAI221xp5_ASAP7_75t_L     g14849(.A1(new_n4312), .A2(new_n5186), .B1(new_n5166), .B2(new_n4986), .C(new_n15105), .Y(new_n15106));
  XNOR2x2_ASAP7_75t_L       g14850(.A(\a[35] ), .B(new_n15106), .Y(new_n15107));
  A2O1A1O1Ixp25_ASAP7_75t_L g14851(.A1(new_n14766), .A2(new_n14693), .B(new_n14768), .C(new_n14998), .D(new_n15006), .Y(new_n15108));
  AOI22xp33_ASAP7_75t_L     g14852(.A1(new_n7659), .A2(\b[26] ), .B1(new_n7656), .B2(new_n2888), .Y(new_n15109));
  OAI221xp5_ASAP7_75t_L     g14853(.A1(new_n8326), .A2(new_n2180), .B1(new_n2019), .B2(new_n7994), .C(new_n15109), .Y(new_n15110));
  XNOR2x2_ASAP7_75t_L       g14854(.A(\a[50] ), .B(new_n15110), .Y(new_n15111));
  INVx1_ASAP7_75t_L         g14855(.A(new_n14954), .Y(new_n15112));
  AOI22xp33_ASAP7_75t_L     g14856(.A1(new_n8645), .A2(\b[23] ), .B1(new_n8642), .B2(new_n2002), .Y(new_n15113));
  OAI221xp5_ASAP7_75t_L     g14857(.A1(new_n9322), .A2(new_n1857), .B1(new_n1709), .B2(new_n8965), .C(new_n15113), .Y(new_n15114));
  XNOR2x2_ASAP7_75t_L       g14858(.A(\a[53] ), .B(new_n15114), .Y(new_n15115));
  AOI22xp33_ASAP7_75t_L     g14859(.A1(new_n10594), .A2(\b[17] ), .B1(new_n10591), .B2(new_n1252), .Y(new_n15116));
  OAI221xp5_ASAP7_75t_L     g14860(.A1(new_n11335), .A2(new_n1051), .B1(new_n952), .B2(new_n11330), .C(new_n15116), .Y(new_n15117));
  XNOR2x2_ASAP7_75t_L       g14861(.A(\a[59] ), .B(new_n15117), .Y(new_n15118));
  A2O1A1Ixp33_ASAP7_75t_L   g14862(.A1(new_n14709), .A2(new_n14923), .B(new_n14924), .C(new_n14922), .Y(new_n15119));
  NOR2xp33_ASAP7_75t_L      g14863(.A(new_n631), .B(new_n12671), .Y(new_n15120));
  O2A1O1Ixp33_ASAP7_75t_L   g14864(.A1(new_n12353), .A2(new_n12355), .B(\b[11] ), .C(new_n15120), .Y(new_n15121));
  NAND2xp33_ASAP7_75t_L     g14865(.A(new_n15121), .B(new_n14922), .Y(new_n15122));
  A2O1A1Ixp33_ASAP7_75t_L   g14866(.A1(\b[11] ), .A2(new_n12669), .B(new_n15120), .C(new_n14927), .Y(new_n15123));
  AND2x2_ASAP7_75t_L        g14867(.A(new_n15122), .B(new_n15123), .Y(new_n15124));
  INVx1_ASAP7_75t_L         g14868(.A(new_n15124), .Y(new_n15125));
  A2O1A1O1Ixp25_ASAP7_75t_L g14869(.A1(new_n14919), .A2(new_n14918), .B(new_n14929), .C(new_n15119), .D(new_n15125), .Y(new_n15126));
  A2O1A1Ixp33_ASAP7_75t_L   g14870(.A1(new_n14918), .A2(new_n14919), .B(new_n14929), .C(new_n15119), .Y(new_n15127));
  NOR2xp33_ASAP7_75t_L      g14871(.A(new_n15124), .B(new_n15127), .Y(new_n15128));
  AOI22xp33_ASAP7_75t_L     g14872(.A1(new_n11656), .A2(\b[14] ), .B1(new_n11654), .B2(new_n879), .Y(new_n15129));
  OAI221xp5_ASAP7_75t_L     g14873(.A1(new_n12364), .A2(new_n793), .B1(new_n763), .B2(new_n13003), .C(new_n15129), .Y(new_n15130));
  XNOR2x2_ASAP7_75t_L       g14874(.A(\a[62] ), .B(new_n15130), .Y(new_n15131));
  INVx1_ASAP7_75t_L         g14875(.A(new_n15131), .Y(new_n15132));
  OAI21xp33_ASAP7_75t_L     g14876(.A1(new_n15126), .A2(new_n15128), .B(new_n15132), .Y(new_n15133));
  NOR2xp33_ASAP7_75t_L      g14877(.A(new_n15126), .B(new_n15128), .Y(new_n15134));
  NAND2xp33_ASAP7_75t_L     g14878(.A(new_n15131), .B(new_n15134), .Y(new_n15135));
  AND3x1_ASAP7_75t_L        g14879(.A(new_n15118), .B(new_n15135), .C(new_n15133), .Y(new_n15136));
  AOI21xp33_ASAP7_75t_L     g14880(.A1(new_n15135), .A2(new_n15133), .B(new_n15118), .Y(new_n15137));
  NOR2xp33_ASAP7_75t_L      g14881(.A(new_n15137), .B(new_n15136), .Y(new_n15138));
  A2O1A1Ixp33_ASAP7_75t_L   g14882(.A1(new_n14931), .A2(new_n14914), .B(new_n14932), .C(new_n15138), .Y(new_n15139));
  A2O1A1Ixp33_ASAP7_75t_L   g14883(.A1(new_n14718), .A2(new_n14717), .B(new_n14930), .C(new_n14934), .Y(new_n15140));
  NOR2xp33_ASAP7_75t_L      g14884(.A(new_n15140), .B(new_n15138), .Y(new_n15141));
  INVx1_ASAP7_75t_L         g14885(.A(new_n15141), .Y(new_n15142));
  NAND2xp33_ASAP7_75t_L     g14886(.A(new_n15139), .B(new_n15142), .Y(new_n15143));
  AOI22xp33_ASAP7_75t_L     g14887(.A1(new_n9623), .A2(\b[20] ), .B1(new_n9620), .B2(new_n1600), .Y(new_n15144));
  OAI221xp5_ASAP7_75t_L     g14888(.A1(new_n10280), .A2(new_n1493), .B1(new_n1356), .B2(new_n12010), .C(new_n15144), .Y(new_n15145));
  XNOR2x2_ASAP7_75t_L       g14889(.A(\a[56] ), .B(new_n15145), .Y(new_n15146));
  NAND2xp33_ASAP7_75t_L     g14890(.A(new_n15146), .B(new_n15143), .Y(new_n15147));
  NOR2xp33_ASAP7_75t_L      g14891(.A(new_n15146), .B(new_n15143), .Y(new_n15148));
  INVx1_ASAP7_75t_L         g14892(.A(new_n15148), .Y(new_n15149));
  NAND2xp33_ASAP7_75t_L     g14893(.A(new_n15149), .B(new_n15147), .Y(new_n15150));
  NAND2xp33_ASAP7_75t_L     g14894(.A(new_n14936), .B(new_n14945), .Y(new_n15151));
  XOR2x2_ASAP7_75t_L        g14895(.A(new_n15151), .B(new_n15150), .Y(new_n15152));
  XNOR2x2_ASAP7_75t_L       g14896(.A(new_n15115), .B(new_n15152), .Y(new_n15153));
  OA211x2_ASAP7_75t_L       g14897(.A1(new_n14948), .A2(new_n14947), .B(new_n15153), .C(new_n15112), .Y(new_n15154));
  O2A1O1Ixp33_ASAP7_75t_L   g14898(.A1(new_n14947), .A2(new_n14948), .B(new_n15112), .C(new_n15153), .Y(new_n15155));
  NOR3xp33_ASAP7_75t_L      g14899(.A(new_n15154), .B(new_n15155), .C(new_n15111), .Y(new_n15156));
  INVx1_ASAP7_75t_L         g14900(.A(new_n15156), .Y(new_n15157));
  OAI21xp33_ASAP7_75t_L     g14901(.A1(new_n15155), .A2(new_n15154), .B(new_n15111), .Y(new_n15158));
  NAND2xp33_ASAP7_75t_L     g14902(.A(new_n15158), .B(new_n15157), .Y(new_n15159));
  NAND2xp33_ASAP7_75t_L     g14903(.A(new_n14959), .B(new_n14966), .Y(new_n15160));
  XNOR2x2_ASAP7_75t_L       g14904(.A(new_n15160), .B(new_n15159), .Y(new_n15161));
  AOI22xp33_ASAP7_75t_L     g14905(.A1(new_n6822), .A2(\b[29] ), .B1(new_n6819), .B2(new_n5472), .Y(new_n15162));
  OAI221xp5_ASAP7_75t_L     g14906(.A1(new_n7392), .A2(new_n2852), .B1(new_n2650), .B2(new_n7115), .C(new_n15162), .Y(new_n15163));
  XNOR2x2_ASAP7_75t_L       g14907(.A(\a[47] ), .B(new_n15163), .Y(new_n15164));
  INVx1_ASAP7_75t_L         g14908(.A(new_n15164), .Y(new_n15165));
  NOR2xp33_ASAP7_75t_L      g14909(.A(new_n15165), .B(new_n15161), .Y(new_n15166));
  AND2x2_ASAP7_75t_L        g14910(.A(new_n15165), .B(new_n15161), .Y(new_n15167));
  NOR2xp33_ASAP7_75t_L      g14911(.A(new_n15166), .B(new_n15167), .Y(new_n15168));
  NAND2xp33_ASAP7_75t_L     g14912(.A(new_n14978), .B(new_n14976), .Y(new_n15169));
  XOR2x2_ASAP7_75t_L        g14913(.A(new_n15169), .B(new_n15168), .Y(new_n15170));
  AOI22xp33_ASAP7_75t_L     g14914(.A1(new_n6002), .A2(\b[32] ), .B1(new_n5999), .B2(new_n3450), .Y(new_n15171));
  OAI221xp5_ASAP7_75t_L     g14915(.A1(new_n6544), .A2(new_n3419), .B1(new_n3212), .B2(new_n6309), .C(new_n15171), .Y(new_n15172));
  XNOR2x2_ASAP7_75t_L       g14916(.A(\a[44] ), .B(new_n15172), .Y(new_n15173));
  XNOR2x2_ASAP7_75t_L       g14917(.A(new_n15173), .B(new_n15170), .Y(new_n15174));
  OA21x2_ASAP7_75t_L        g14918(.A1(new_n14988), .A2(new_n14985), .B(new_n14984), .Y(new_n15175));
  XNOR2x2_ASAP7_75t_L       g14919(.A(new_n15175), .B(new_n15174), .Y(new_n15176));
  AOI22xp33_ASAP7_75t_L     g14920(.A1(new_n5249), .A2(\b[35] ), .B1(new_n5247), .B2(new_n5649), .Y(new_n15177));
  OAI221xp5_ASAP7_75t_L     g14921(.A1(new_n5241), .A2(new_n3827), .B1(new_n3807), .B2(new_n5521), .C(new_n15177), .Y(new_n15178));
  XNOR2x2_ASAP7_75t_L       g14922(.A(\a[41] ), .B(new_n15178), .Y(new_n15179));
  XOR2x2_ASAP7_75t_L        g14923(.A(new_n15179), .B(new_n15176), .Y(new_n15180));
  INVx1_ASAP7_75t_L         g14924(.A(new_n15180), .Y(new_n15181));
  OAI21xp33_ASAP7_75t_L     g14925(.A1(new_n14911), .A2(new_n14993), .B(new_n14991), .Y(new_n15182));
  NOR2xp33_ASAP7_75t_L      g14926(.A(new_n15182), .B(new_n15181), .Y(new_n15183));
  O2A1O1Ixp33_ASAP7_75t_L   g14927(.A1(new_n14911), .A2(new_n14993), .B(new_n14991), .C(new_n15180), .Y(new_n15184));
  AOI22xp33_ASAP7_75t_L     g14928(.A1(new_n4544), .A2(\b[38] ), .B1(new_n4542), .B2(new_n4923), .Y(new_n15185));
  OAI221xp5_ASAP7_75t_L     g14929(.A1(new_n4536), .A2(new_n4701), .B1(new_n4465), .B2(new_n4781), .C(new_n15185), .Y(new_n15186));
  XNOR2x2_ASAP7_75t_L       g14930(.A(\a[38] ), .B(new_n15186), .Y(new_n15187));
  OAI21xp33_ASAP7_75t_L     g14931(.A1(new_n15183), .A2(new_n15184), .B(new_n15187), .Y(new_n15188));
  OR3x1_ASAP7_75t_L         g14932(.A(new_n15183), .B(new_n15184), .C(new_n15187), .Y(new_n15189));
  NAND2xp33_ASAP7_75t_L     g14933(.A(new_n15188), .B(new_n15189), .Y(new_n15190));
  XOR2x2_ASAP7_75t_L        g14934(.A(new_n15108), .B(new_n15190), .Y(new_n15191));
  XNOR2x2_ASAP7_75t_L       g14935(.A(new_n15107), .B(new_n15191), .Y(new_n15192));
  XOR2x2_ASAP7_75t_L        g14936(.A(new_n15192), .B(new_n15104), .Y(new_n15193));
  NOR2xp33_ASAP7_75t_L      g14937(.A(new_n15095), .B(new_n15193), .Y(new_n15194));
  AND2x2_ASAP7_75t_L        g14938(.A(new_n15095), .B(new_n15193), .Y(new_n15195));
  NOR2xp33_ASAP7_75t_L      g14939(.A(new_n15194), .B(new_n15195), .Y(new_n15196));
  NAND2xp33_ASAP7_75t_L     g14940(.A(new_n15196), .B(new_n15087), .Y(new_n15197));
  OAI22xp33_ASAP7_75t_L     g14941(.A1(new_n15085), .A2(new_n15086), .B1(new_n15195), .B2(new_n15194), .Y(new_n15198));
  AND2x2_ASAP7_75t_L        g14942(.A(new_n15198), .B(new_n15197), .Y(new_n15199));
  XNOR2x2_ASAP7_75t_L       g14943(.A(new_n15079), .B(new_n15199), .Y(new_n15200));
  XNOR2x2_ASAP7_75t_L       g14944(.A(new_n15200), .B(new_n15070), .Y(new_n15201));
  NAND3xp33_ASAP7_75t_L     g14945(.A(new_n15060), .B(new_n15059), .C(new_n15201), .Y(new_n15202));
  AO21x2_ASAP7_75t_L        g14946(.A1(new_n15059), .A2(new_n15060), .B(new_n15201), .Y(new_n15203));
  AO21x2_ASAP7_75t_L        g14947(.A1(new_n15203), .A2(new_n15202), .B(new_n15053), .Y(new_n15204));
  NAND3xp33_ASAP7_75t_L     g14948(.A(new_n15053), .B(new_n15202), .C(new_n15203), .Y(new_n15205));
  NAND2xp33_ASAP7_75t_L     g14949(.A(new_n14854), .B(new_n14856), .Y(new_n15206));
  A2O1A1Ixp33_ASAP7_75t_L   g14950(.A1(new_n14818), .A2(new_n14645), .B(new_n14647), .C(new_n14853), .Y(new_n15207));
  INVx1_ASAP7_75t_L         g14951(.A(new_n15207), .Y(new_n15208));
  A2O1A1Ixp33_ASAP7_75t_L   g14952(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n597), .Y(new_n15209));
  A2O1A1Ixp33_ASAP7_75t_L   g14953(.A1(new_n15209), .A2(new_n1620), .B(new_n12599), .C(\a[11] ), .Y(new_n15210));
  O2A1O1Ixp33_ASAP7_75t_L   g14954(.A1(new_n675), .A2(new_n13934), .B(new_n1620), .C(new_n12599), .Y(new_n15211));
  NAND2xp33_ASAP7_75t_L     g14955(.A(new_n594), .B(new_n15211), .Y(new_n15212));
  AND2x2_ASAP7_75t_L        g14956(.A(new_n15212), .B(new_n15210), .Y(new_n15213));
  INVx1_ASAP7_75t_L         g14957(.A(new_n15213), .Y(new_n15214));
  A2O1A1Ixp33_ASAP7_75t_L   g14958(.A1(new_n15024), .A2(new_n15206), .B(new_n15208), .C(new_n15214), .Y(new_n15215));
  O2A1O1Ixp33_ASAP7_75t_L   g14959(.A1(new_n14855), .A2(new_n15022), .B(new_n15024), .C(new_n15208), .Y(new_n15216));
  NAND2xp33_ASAP7_75t_L     g14960(.A(new_n15213), .B(new_n15216), .Y(new_n15217));
  AND4x1_ASAP7_75t_L        g14961(.A(new_n15204), .B(new_n15217), .C(new_n15205), .D(new_n15215), .Y(new_n15218));
  AOI22xp33_ASAP7_75t_L     g14962(.A1(new_n15204), .A2(new_n15205), .B1(new_n15215), .B2(new_n15217), .Y(new_n15219));
  OA21x2_ASAP7_75t_L        g14963(.A1(new_n15219), .A2(new_n15218), .B(new_n15042), .Y(new_n15220));
  NOR3xp33_ASAP7_75t_L      g14964(.A(new_n15042), .B(new_n15218), .C(new_n15219), .Y(new_n15221));
  NOR2xp33_ASAP7_75t_L      g14965(.A(new_n15221), .B(new_n15220), .Y(new_n15222));
  A2O1A1Ixp33_ASAP7_75t_L   g14966(.A1(new_n15038), .A2(new_n15034), .B(new_n15032), .C(new_n15222), .Y(new_n15223));
  INVx1_ASAP7_75t_L         g14967(.A(new_n15223), .Y(new_n15224));
  INVx1_ASAP7_75t_L         g14968(.A(new_n15032), .Y(new_n15225));
  A2O1A1Ixp33_ASAP7_75t_L   g14969(.A1(new_n14834), .A2(new_n14830), .B(new_n15035), .C(new_n15225), .Y(new_n15226));
  NOR2xp33_ASAP7_75t_L      g14970(.A(new_n15222), .B(new_n15226), .Y(new_n15227));
  NOR2xp33_ASAP7_75t_L      g14971(.A(new_n15224), .B(new_n15227), .Y(\f[74] ));
  INVx1_ASAP7_75t_L         g14972(.A(new_n15060), .Y(new_n15229));
  AOI22xp33_ASAP7_75t_L     g14973(.A1(new_n1113), .A2(\b[60] ), .B1(new_n1110), .B2(new_n11234), .Y(new_n15230));
  OAI221xp5_ASAP7_75t_L     g14974(.A1(new_n1298), .A2(new_n10881), .B1(new_n10848), .B2(new_n1195), .C(new_n15230), .Y(new_n15231));
  XNOR2x2_ASAP7_75t_L       g14975(.A(\a[17] ), .B(new_n15231), .Y(new_n15232));
  A2O1A1Ixp33_ASAP7_75t_L   g14976(.A1(new_n15201), .A2(new_n15059), .B(new_n15229), .C(new_n15232), .Y(new_n15233));
  INVx1_ASAP7_75t_L         g14977(.A(new_n15233), .Y(new_n15234));
  AND3x1_ASAP7_75t_L        g14978(.A(new_n15060), .B(new_n15201), .C(new_n15059), .Y(new_n15235));
  NOR3xp33_ASAP7_75t_L      g14979(.A(new_n15235), .B(new_n15232), .C(new_n15229), .Y(new_n15236));
  AOI22xp33_ASAP7_75t_L     g14980(.A1(new_n1406), .A2(\b[57] ), .B1(new_n1404), .B2(new_n10495), .Y(new_n15237));
  OAI221xp5_ASAP7_75t_L     g14981(.A1(new_n1398), .A2(new_n10178), .B1(new_n9534), .B2(new_n1549), .C(new_n15237), .Y(new_n15238));
  XNOR2x2_ASAP7_75t_L       g14982(.A(\a[20] ), .B(new_n15238), .Y(new_n15239));
  INVx1_ASAP7_75t_L         g14983(.A(new_n15239), .Y(new_n15240));
  A2O1A1Ixp33_ASAP7_75t_L   g14984(.A1(new_n14878), .A2(new_n15015), .B(new_n15066), .C(new_n15064), .Y(new_n15241));
  A2O1A1Ixp33_ASAP7_75t_L   g14985(.A1(new_n15069), .A2(new_n15068), .B(new_n15200), .C(new_n15241), .Y(new_n15242));
  OR2x4_ASAP7_75t_L         g14986(.A(new_n15240), .B(new_n15242), .Y(new_n15243));
  NAND2xp33_ASAP7_75t_L     g14987(.A(new_n15240), .B(new_n15242), .Y(new_n15244));
  A2O1A1O1Ixp25_ASAP7_75t_L g14988(.A1(new_n15073), .A2(new_n15072), .B(new_n15014), .C(new_n15074), .D(new_n15078), .Y(new_n15245));
  AOI22xp33_ASAP7_75t_L     g14989(.A1(new_n1766), .A2(\b[54] ), .B1(new_n1764), .B2(new_n9208), .Y(new_n15246));
  OAI221xp5_ASAP7_75t_L     g14990(.A1(new_n1758), .A2(new_n8882), .B1(new_n8569), .B2(new_n1911), .C(new_n15246), .Y(new_n15247));
  XNOR2x2_ASAP7_75t_L       g14991(.A(\a[23] ), .B(new_n15247), .Y(new_n15248));
  A2O1A1Ixp33_ASAP7_75t_L   g14992(.A1(new_n15199), .A2(new_n15079), .B(new_n15245), .C(new_n15248), .Y(new_n15249));
  AOI21xp33_ASAP7_75t_L     g14993(.A1(new_n15199), .A2(new_n15079), .B(new_n15245), .Y(new_n15250));
  INVx1_ASAP7_75t_L         g14994(.A(new_n15248), .Y(new_n15251));
  NAND2xp33_ASAP7_75t_L     g14995(.A(new_n15251), .B(new_n15250), .Y(new_n15252));
  NAND2xp33_ASAP7_75t_L     g14996(.A(new_n15249), .B(new_n15252), .Y(new_n15253));
  AOI22xp33_ASAP7_75t_L     g14997(.A1(new_n2228), .A2(\b[51] ), .B1(new_n2226), .B2(new_n8257), .Y(new_n15254));
  OAI221xp5_ASAP7_75t_L     g14998(.A1(new_n2220), .A2(new_n8228), .B1(new_n7907), .B2(new_n2387), .C(new_n15254), .Y(new_n15255));
  XNOR2x2_ASAP7_75t_L       g14999(.A(\a[26] ), .B(new_n15255), .Y(new_n15256));
  INVx1_ASAP7_75t_L         g15000(.A(new_n15256), .Y(new_n15257));
  AOI211xp5_ASAP7_75t_L     g15001(.A1(new_n15087), .A2(new_n15196), .B(new_n15257), .C(new_n15085), .Y(new_n15258));
  A2O1A1Ixp33_ASAP7_75t_L   g15002(.A1(new_n15087), .A2(new_n15196), .B(new_n15085), .C(new_n15257), .Y(new_n15259));
  INVx1_ASAP7_75t_L         g15003(.A(new_n15259), .Y(new_n15260));
  NOR2xp33_ASAP7_75t_L      g15004(.A(new_n15258), .B(new_n15260), .Y(new_n15261));
  AOI22xp33_ASAP7_75t_L     g15005(.A1(new_n2702), .A2(\b[48] ), .B1(new_n2700), .B2(new_n7341), .Y(new_n15262));
  OAI221xp5_ASAP7_75t_L     g15006(.A1(new_n2694), .A2(new_n7316), .B1(new_n7033), .B2(new_n2932), .C(new_n15262), .Y(new_n15263));
  XNOR2x2_ASAP7_75t_L       g15007(.A(\a[29] ), .B(new_n15263), .Y(new_n15264));
  INVx1_ASAP7_75t_L         g15008(.A(new_n15264), .Y(new_n15265));
  O2A1O1Ixp33_ASAP7_75t_L   g15009(.A1(new_n15095), .A2(new_n15193), .B(new_n15094), .C(new_n15265), .Y(new_n15266));
  INVx1_ASAP7_75t_L         g15010(.A(new_n15266), .Y(new_n15267));
  OR2x4_ASAP7_75t_L         g15011(.A(new_n15095), .B(new_n15193), .Y(new_n15268));
  NAND3xp33_ASAP7_75t_L     g15012(.A(new_n15268), .B(new_n15094), .C(new_n15265), .Y(new_n15269));
  NAND2xp33_ASAP7_75t_L     g15013(.A(new_n15267), .B(new_n15269), .Y(new_n15270));
  AOI22xp33_ASAP7_75t_L     g15014(.A1(new_n3884), .A2(\b[42] ), .B1(new_n3881), .B2(new_n5688), .Y(new_n15271));
  OAI221xp5_ASAP7_75t_L     g15015(.A1(new_n4312), .A2(new_n5666), .B1(new_n5186), .B2(new_n4986), .C(new_n15271), .Y(new_n15272));
  XNOR2x2_ASAP7_75t_L       g15016(.A(\a[35] ), .B(new_n15272), .Y(new_n15273));
  INVx1_ASAP7_75t_L         g15017(.A(new_n15184), .Y(new_n15274));
  AOI22xp33_ASAP7_75t_L     g15018(.A1(new_n5249), .A2(\b[36] ), .B1(new_n5247), .B2(new_n4473), .Y(new_n15275));
  OAI221xp5_ASAP7_75t_L     g15019(.A1(new_n5241), .A2(new_n4053), .B1(new_n3827), .B2(new_n5521), .C(new_n15275), .Y(new_n15276));
  XNOR2x2_ASAP7_75t_L       g15020(.A(\a[41] ), .B(new_n15276), .Y(new_n15277));
  INVx1_ASAP7_75t_L         g15021(.A(new_n15277), .Y(new_n15278));
  MAJIxp5_ASAP7_75t_L       g15022(.A(new_n15168), .B(new_n15173), .C(new_n15169), .Y(new_n15279));
  AOI22xp33_ASAP7_75t_L     g15023(.A1(new_n6002), .A2(\b[33] ), .B1(new_n5999), .B2(new_n3813), .Y(new_n15280));
  OAI221xp5_ASAP7_75t_L     g15024(.A1(new_n6544), .A2(new_n3443), .B1(new_n3419), .B2(new_n6309), .C(new_n15280), .Y(new_n15281));
  XNOR2x2_ASAP7_75t_L       g15025(.A(\a[44] ), .B(new_n15281), .Y(new_n15282));
  NOR2xp33_ASAP7_75t_L      g15026(.A(new_n15154), .B(new_n15156), .Y(new_n15283));
  MAJIxp5_ASAP7_75t_L       g15027(.A(new_n15150), .B(new_n15115), .C(new_n15151), .Y(new_n15284));
  AOI22xp33_ASAP7_75t_L     g15028(.A1(new_n8645), .A2(\b[24] ), .B1(new_n8642), .B2(new_n2027), .Y(new_n15285));
  OAI221xp5_ASAP7_75t_L     g15029(.A1(new_n9322), .A2(new_n1995), .B1(new_n1857), .B2(new_n8965), .C(new_n15285), .Y(new_n15286));
  XNOR2x2_ASAP7_75t_L       g15030(.A(\a[53] ), .B(new_n15286), .Y(new_n15287));
  A2O1A1O1Ixp25_ASAP7_75t_L g15031(.A1(new_n14919), .A2(new_n14918), .B(new_n14929), .C(new_n15119), .D(new_n15124), .Y(new_n15288));
  A2O1A1O1Ixp25_ASAP7_75t_L g15032(.A1(new_n12669), .A2(\b[11] ), .B(new_n15120), .C(new_n14922), .D(new_n15288), .Y(new_n15289));
  AOI22xp33_ASAP7_75t_L     g15033(.A1(new_n11656), .A2(\b[15] ), .B1(new_n11654), .B2(new_n959), .Y(new_n15290));
  OAI221xp5_ASAP7_75t_L     g15034(.A1(new_n12364), .A2(new_n871), .B1(new_n793), .B2(new_n13003), .C(new_n15290), .Y(new_n15291));
  XNOR2x2_ASAP7_75t_L       g15035(.A(new_n11651), .B(new_n15291), .Y(new_n15292));
  NOR2xp33_ASAP7_75t_L      g15036(.A(new_n695), .B(new_n12671), .Y(new_n15293));
  O2A1O1Ixp33_ASAP7_75t_L   g15037(.A1(new_n12353), .A2(new_n12355), .B(\b[12] ), .C(new_n15293), .Y(new_n15294));
  A2O1A1Ixp33_ASAP7_75t_L   g15038(.A1(new_n12669), .A2(\b[10] ), .B(new_n14921), .C(\a[11] ), .Y(new_n15295));
  NOR2xp33_ASAP7_75t_L      g15039(.A(\a[11] ), .B(new_n14927), .Y(new_n15296));
  INVx1_ASAP7_75t_L         g15040(.A(new_n15296), .Y(new_n15297));
  AOI21xp33_ASAP7_75t_L     g15041(.A1(new_n15297), .A2(new_n15295), .B(new_n15294), .Y(new_n15298));
  AND3x1_ASAP7_75t_L        g15042(.A(new_n15297), .B(new_n15295), .C(new_n15294), .Y(new_n15299));
  NOR2xp33_ASAP7_75t_L      g15043(.A(new_n15298), .B(new_n15299), .Y(new_n15300));
  XNOR2x2_ASAP7_75t_L       g15044(.A(new_n15300), .B(new_n15292), .Y(new_n15301));
  XOR2x2_ASAP7_75t_L        g15045(.A(new_n15289), .B(new_n15301), .Y(new_n15302));
  AOI22xp33_ASAP7_75t_L     g15046(.A1(new_n10594), .A2(\b[18] ), .B1(new_n10591), .B2(new_n1363), .Y(new_n15303));
  OAI221xp5_ASAP7_75t_L     g15047(.A1(new_n11335), .A2(new_n1244), .B1(new_n1051), .B2(new_n11330), .C(new_n15303), .Y(new_n15304));
  XNOR2x2_ASAP7_75t_L       g15048(.A(\a[59] ), .B(new_n15304), .Y(new_n15305));
  INVx1_ASAP7_75t_L         g15049(.A(new_n15305), .Y(new_n15306));
  NAND2xp33_ASAP7_75t_L     g15050(.A(new_n15306), .B(new_n15302), .Y(new_n15307));
  INVx1_ASAP7_75t_L         g15051(.A(new_n15307), .Y(new_n15308));
  NOR2xp33_ASAP7_75t_L      g15052(.A(new_n15306), .B(new_n15302), .Y(new_n15309));
  OR2x4_ASAP7_75t_L         g15053(.A(new_n15309), .B(new_n15308), .Y(new_n15310));
  A2O1A1Ixp33_ASAP7_75t_L   g15054(.A1(new_n15131), .A2(new_n15134), .B(new_n15136), .C(new_n15310), .Y(new_n15311));
  INVx1_ASAP7_75t_L         g15055(.A(new_n15135), .Y(new_n15312));
  OR4x2_ASAP7_75t_L         g15056(.A(new_n15309), .B(new_n15308), .C(new_n15136), .D(new_n15312), .Y(new_n15313));
  NAND2xp33_ASAP7_75t_L     g15057(.A(new_n15313), .B(new_n15311), .Y(new_n15314));
  AOI22xp33_ASAP7_75t_L     g15058(.A1(new_n9623), .A2(\b[21] ), .B1(new_n9620), .B2(new_n1715), .Y(new_n15315));
  OAI221xp5_ASAP7_75t_L     g15059(.A1(new_n10280), .A2(new_n1594), .B1(new_n1493), .B2(new_n12010), .C(new_n15315), .Y(new_n15316));
  XNOR2x2_ASAP7_75t_L       g15060(.A(\a[56] ), .B(new_n15316), .Y(new_n15317));
  XNOR2x2_ASAP7_75t_L       g15061(.A(new_n15317), .B(new_n15314), .Y(new_n15318));
  INVx1_ASAP7_75t_L         g15062(.A(new_n15140), .Y(new_n15319));
  O2A1O1Ixp33_ASAP7_75t_L   g15063(.A1(new_n15136), .A2(new_n15137), .B(new_n15319), .C(new_n15148), .Y(new_n15320));
  XOR2x2_ASAP7_75t_L        g15064(.A(new_n15320), .B(new_n15318), .Y(new_n15321));
  XNOR2x2_ASAP7_75t_L       g15065(.A(new_n15287), .B(new_n15321), .Y(new_n15322));
  XNOR2x2_ASAP7_75t_L       g15066(.A(new_n15284), .B(new_n15322), .Y(new_n15323));
  AOI22xp33_ASAP7_75t_L     g15067(.A1(new_n7659), .A2(\b[27] ), .B1(new_n7656), .B2(new_n2657), .Y(new_n15324));
  OAI221xp5_ASAP7_75t_L     g15068(.A1(new_n8326), .A2(new_n2477), .B1(new_n2180), .B2(new_n7994), .C(new_n15324), .Y(new_n15325));
  XNOR2x2_ASAP7_75t_L       g15069(.A(\a[50] ), .B(new_n15325), .Y(new_n15326));
  XNOR2x2_ASAP7_75t_L       g15070(.A(new_n15326), .B(new_n15323), .Y(new_n15327));
  XOR2x2_ASAP7_75t_L        g15071(.A(new_n15283), .B(new_n15327), .Y(new_n15328));
  AOI22xp33_ASAP7_75t_L     g15072(.A1(new_n6822), .A2(\b[30] ), .B1(new_n6819), .B2(new_n3219), .Y(new_n15329));
  OAI221xp5_ASAP7_75t_L     g15073(.A1(new_n7392), .A2(new_n2871), .B1(new_n2852), .B2(new_n7115), .C(new_n15329), .Y(new_n15330));
  XNOR2x2_ASAP7_75t_L       g15074(.A(new_n6816), .B(new_n15330), .Y(new_n15331));
  XNOR2x2_ASAP7_75t_L       g15075(.A(new_n15331), .B(new_n15328), .Y(new_n15332));
  INVx1_ASAP7_75t_L         g15076(.A(new_n15158), .Y(new_n15333));
  O2A1O1Ixp33_ASAP7_75t_L   g15077(.A1(new_n15156), .A2(new_n15333), .B(new_n15160), .C(new_n15166), .Y(new_n15334));
  XNOR2x2_ASAP7_75t_L       g15078(.A(new_n15334), .B(new_n15332), .Y(new_n15335));
  XNOR2x2_ASAP7_75t_L       g15079(.A(new_n15282), .B(new_n15335), .Y(new_n15336));
  XOR2x2_ASAP7_75t_L        g15080(.A(new_n15279), .B(new_n15336), .Y(new_n15337));
  XNOR2x2_ASAP7_75t_L       g15081(.A(new_n15278), .B(new_n15337), .Y(new_n15338));
  INVx1_ASAP7_75t_L         g15082(.A(new_n15174), .Y(new_n15339));
  MAJx2_ASAP7_75t_L         g15083(.A(new_n15339), .B(new_n15175), .C(new_n15179), .Y(new_n15340));
  XNOR2x2_ASAP7_75t_L       g15084(.A(new_n15340), .B(new_n15338), .Y(new_n15341));
  AOI22xp33_ASAP7_75t_L     g15085(.A1(new_n4544), .A2(\b[39] ), .B1(new_n4542), .B2(new_n5174), .Y(new_n15342));
  OAI221xp5_ASAP7_75t_L     g15086(.A1(new_n4536), .A2(new_n4915), .B1(new_n4701), .B2(new_n4781), .C(new_n15342), .Y(new_n15343));
  XNOR2x2_ASAP7_75t_L       g15087(.A(\a[38] ), .B(new_n15343), .Y(new_n15344));
  XNOR2x2_ASAP7_75t_L       g15088(.A(new_n15344), .B(new_n15341), .Y(new_n15345));
  AO21x2_ASAP7_75t_L        g15089(.A1(new_n15274), .A2(new_n15189), .B(new_n15345), .Y(new_n15346));
  NAND3xp33_ASAP7_75t_L     g15090(.A(new_n15345), .B(new_n15189), .C(new_n15274), .Y(new_n15347));
  NAND2xp33_ASAP7_75t_L     g15091(.A(new_n15347), .B(new_n15346), .Y(new_n15348));
  XNOR2x2_ASAP7_75t_L       g15092(.A(new_n15273), .B(new_n15348), .Y(new_n15349));
  MAJx2_ASAP7_75t_L         g15093(.A(new_n15190), .B(new_n15108), .C(new_n15107), .Y(new_n15350));
  XNOR2x2_ASAP7_75t_L       g15094(.A(new_n15350), .B(new_n15349), .Y(new_n15351));
  AOI22xp33_ASAP7_75t_L     g15095(.A1(new_n3256), .A2(\b[45] ), .B1(new_n3254), .B2(new_n6764), .Y(new_n15352));
  OAI221xp5_ASAP7_75t_L     g15096(.A1(new_n3248), .A2(new_n6220), .B1(new_n6195), .B2(new_n3492), .C(new_n15352), .Y(new_n15353));
  XNOR2x2_ASAP7_75t_L       g15097(.A(\a[32] ), .B(new_n15353), .Y(new_n15354));
  MAJIxp5_ASAP7_75t_L       g15098(.A(new_n15192), .B(new_n15099), .C(new_n15101), .Y(new_n15355));
  XNOR2x2_ASAP7_75t_L       g15099(.A(new_n15354), .B(new_n15355), .Y(new_n15356));
  NOR2xp33_ASAP7_75t_L      g15100(.A(new_n15351), .B(new_n15356), .Y(new_n15357));
  AND2x2_ASAP7_75t_L        g15101(.A(new_n15351), .B(new_n15356), .Y(new_n15358));
  NOR2xp33_ASAP7_75t_L      g15102(.A(new_n15357), .B(new_n15358), .Y(new_n15359));
  XNOR2x2_ASAP7_75t_L       g15103(.A(new_n15359), .B(new_n15270), .Y(new_n15360));
  XNOR2x2_ASAP7_75t_L       g15104(.A(new_n15360), .B(new_n15261), .Y(new_n15361));
  XOR2x2_ASAP7_75t_L        g15105(.A(new_n15361), .B(new_n15253), .Y(new_n15362));
  NAND3xp33_ASAP7_75t_L     g15106(.A(new_n15362), .B(new_n15244), .C(new_n15243), .Y(new_n15363));
  AO21x2_ASAP7_75t_L        g15107(.A1(new_n15243), .A2(new_n15244), .B(new_n15362), .Y(new_n15364));
  AND2x2_ASAP7_75t_L        g15108(.A(new_n15363), .B(new_n15364), .Y(new_n15365));
  OAI21xp33_ASAP7_75t_L     g15109(.A1(new_n15236), .A2(new_n15234), .B(new_n15365), .Y(new_n15366));
  OR3x1_ASAP7_75t_L         g15110(.A(new_n15235), .B(new_n15229), .C(new_n15232), .Y(new_n15367));
  NAND2xp33_ASAP7_75t_L     g15111(.A(new_n15363), .B(new_n15364), .Y(new_n15368));
  NAND3xp33_ASAP7_75t_L     g15112(.A(new_n15367), .B(new_n15368), .C(new_n15233), .Y(new_n15369));
  AND2x2_ASAP7_75t_L        g15113(.A(new_n15369), .B(new_n15366), .Y(new_n15370));
  NAND2xp33_ASAP7_75t_L     g15114(.A(\b[63] ), .B(new_n826), .Y(new_n15371));
  A2O1A1Ixp33_ASAP7_75t_L   g15115(.A1(new_n12607), .A2(new_n12603), .B(new_n911), .C(new_n15371), .Y(new_n15372));
  AOI221xp5_ASAP7_75t_L     g15116(.A1(\b[61] ), .A2(new_n908), .B1(\b[62] ), .B2(new_n817), .C(new_n15372), .Y(new_n15373));
  XNOR2x2_ASAP7_75t_L       g15117(.A(new_n813), .B(new_n15373), .Y(new_n15374));
  INVx1_ASAP7_75t_L         g15118(.A(new_n15048), .Y(new_n15375));
  A2O1A1Ixp33_ASAP7_75t_L   g15119(.A1(new_n15203), .A2(new_n15202), .B(new_n15375), .C(new_n15052), .Y(new_n15376));
  NOR2xp33_ASAP7_75t_L      g15120(.A(new_n15374), .B(new_n15376), .Y(new_n15377));
  INVx1_ASAP7_75t_L         g15121(.A(new_n15377), .Y(new_n15378));
  INVx1_ASAP7_75t_L         g15122(.A(new_n15374), .Y(new_n15379));
  A2O1A1O1Ixp25_ASAP7_75t_L g15123(.A1(new_n15202), .A2(new_n15203), .B(new_n15375), .C(new_n15052), .D(new_n15379), .Y(new_n15380));
  INVx1_ASAP7_75t_L         g15124(.A(new_n15380), .Y(new_n15381));
  NAND3xp33_ASAP7_75t_L     g15125(.A(new_n15370), .B(new_n15378), .C(new_n15381), .Y(new_n15382));
  NAND2xp33_ASAP7_75t_L     g15126(.A(new_n15369), .B(new_n15366), .Y(new_n15383));
  OAI21xp33_ASAP7_75t_L     g15127(.A1(new_n15377), .A2(new_n15380), .B(new_n15383), .Y(new_n15384));
  INVx1_ASAP7_75t_L         g15128(.A(new_n15217), .Y(new_n15385));
  NOR2xp33_ASAP7_75t_L      g15129(.A(new_n15385), .B(new_n15218), .Y(new_n15386));
  NAND3xp33_ASAP7_75t_L     g15130(.A(new_n15382), .B(new_n15384), .C(new_n15386), .Y(new_n15387));
  NOR3xp33_ASAP7_75t_L      g15131(.A(new_n15383), .B(new_n15377), .C(new_n15380), .Y(new_n15388));
  AOI21xp33_ASAP7_75t_L     g15132(.A1(new_n15378), .A2(new_n15381), .B(new_n15370), .Y(new_n15389));
  OAI22xp33_ASAP7_75t_L     g15133(.A1(new_n15389), .A2(new_n15388), .B1(new_n15218), .B2(new_n15385), .Y(new_n15390));
  NAND2xp33_ASAP7_75t_L     g15134(.A(new_n15387), .B(new_n15390), .Y(new_n15391));
  INVx1_ASAP7_75t_L         g15135(.A(new_n15391), .Y(new_n15392));
  A2O1A1Ixp33_ASAP7_75t_L   g15136(.A1(new_n15226), .A2(new_n15222), .B(new_n15220), .C(new_n15392), .Y(new_n15393));
  A2O1A1O1Ixp25_ASAP7_75t_L g15137(.A1(new_n15034), .A2(new_n15038), .B(new_n15032), .C(new_n15222), .D(new_n15220), .Y(new_n15394));
  NAND2xp33_ASAP7_75t_L     g15138(.A(new_n15391), .B(new_n15394), .Y(new_n15395));
  AND2x2_ASAP7_75t_L        g15139(.A(new_n15395), .B(new_n15393), .Y(\f[75] ));
  NOR2xp33_ASAP7_75t_L      g15140(.A(new_n15377), .B(new_n15388), .Y(new_n15397));
  O2A1O1Ixp33_ASAP7_75t_L   g15141(.A1(new_n15056), .A2(new_n15058), .B(new_n15202), .C(new_n15232), .Y(new_n15398));
  INVx1_ASAP7_75t_L         g15142(.A(new_n15398), .Y(new_n15399));
  AOI22xp33_ASAP7_75t_L     g15143(.A1(new_n817), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n908), .Y(new_n15400));
  A2O1A1Ixp33_ASAP7_75t_L   g15144(.A1(new_n13506), .A2(new_n13507), .B(new_n911), .C(new_n15400), .Y(new_n15401));
  NOR2xp33_ASAP7_75t_L      g15145(.A(new_n813), .B(new_n15401), .Y(new_n15402));
  A2O1A1O1Ixp25_ASAP7_75t_L g15146(.A1(new_n13507), .A2(new_n13506), .B(new_n911), .C(new_n15400), .D(\a[14] ), .Y(new_n15403));
  NOR2xp33_ASAP7_75t_L      g15147(.A(new_n15403), .B(new_n15402), .Y(new_n15404));
  INVx1_ASAP7_75t_L         g15148(.A(new_n15404), .Y(new_n15405));
  A2O1A1O1Ixp25_ASAP7_75t_L g15149(.A1(new_n15233), .A2(new_n15367), .B(new_n15368), .C(new_n15399), .D(new_n15405), .Y(new_n15406));
  A2O1A1Ixp33_ASAP7_75t_L   g15150(.A1(new_n15367), .A2(new_n15233), .B(new_n15368), .C(new_n15399), .Y(new_n15407));
  NOR2xp33_ASAP7_75t_L      g15151(.A(new_n15404), .B(new_n15407), .Y(new_n15408));
  NOR2xp33_ASAP7_75t_L      g15152(.A(new_n15406), .B(new_n15408), .Y(new_n15409));
  AOI22xp33_ASAP7_75t_L     g15153(.A1(new_n1113), .A2(\b[61] ), .B1(new_n1110), .B2(new_n11919), .Y(new_n15410));
  OAI221xp5_ASAP7_75t_L     g15154(.A1(new_n1298), .A2(new_n11226), .B1(new_n10881), .B2(new_n1195), .C(new_n15410), .Y(new_n15411));
  XNOR2x2_ASAP7_75t_L       g15155(.A(\a[17] ), .B(new_n15411), .Y(new_n15412));
  NAND2xp33_ASAP7_75t_L     g15156(.A(new_n15244), .B(new_n15363), .Y(new_n15413));
  XNOR2x2_ASAP7_75t_L       g15157(.A(new_n15412), .B(new_n15413), .Y(new_n15414));
  NOR2xp33_ASAP7_75t_L      g15158(.A(new_n15248), .B(new_n15250), .Y(new_n15415));
  AOI22xp33_ASAP7_75t_L     g15159(.A1(new_n1410), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n1406), .Y(new_n15416));
  OAI221xp5_ASAP7_75t_L     g15160(.A1(new_n1549), .A2(new_n10178), .B1(new_n1411), .B2(new_n10856), .C(new_n15416), .Y(new_n15417));
  XNOR2x2_ASAP7_75t_L       g15161(.A(\a[20] ), .B(new_n15417), .Y(new_n15418));
  A2O1A1Ixp33_ASAP7_75t_L   g15162(.A1(new_n15253), .A2(new_n15361), .B(new_n15415), .C(new_n15418), .Y(new_n15419));
  A2O1A1Ixp33_ASAP7_75t_L   g15163(.A1(new_n15199), .A2(new_n15079), .B(new_n15245), .C(new_n15251), .Y(new_n15420));
  NAND2xp33_ASAP7_75t_L     g15164(.A(new_n15361), .B(new_n15253), .Y(new_n15421));
  INVx1_ASAP7_75t_L         g15165(.A(new_n15418), .Y(new_n15422));
  NAND3xp33_ASAP7_75t_L     g15166(.A(new_n15421), .B(new_n15420), .C(new_n15422), .Y(new_n15423));
  NAND2xp33_ASAP7_75t_L     g15167(.A(new_n15419), .B(new_n15423), .Y(new_n15424));
  AOI22xp33_ASAP7_75t_L     g15168(.A1(new_n1766), .A2(\b[55] ), .B1(new_n1764), .B2(new_n9542), .Y(new_n15425));
  OAI221xp5_ASAP7_75t_L     g15169(.A1(new_n1758), .A2(new_n9199), .B1(new_n8882), .B2(new_n1911), .C(new_n15425), .Y(new_n15426));
  XNOR2x2_ASAP7_75t_L       g15170(.A(\a[23] ), .B(new_n15426), .Y(new_n15427));
  OAI21xp33_ASAP7_75t_L     g15171(.A1(new_n15258), .A2(new_n15360), .B(new_n15259), .Y(new_n15428));
  XNOR2x2_ASAP7_75t_L       g15172(.A(new_n15427), .B(new_n15428), .Y(new_n15429));
  AOI22xp33_ASAP7_75t_L     g15173(.A1(new_n2702), .A2(\b[49] ), .B1(new_n2700), .B2(new_n7914), .Y(new_n15430));
  OAI221xp5_ASAP7_75t_L     g15174(.A1(new_n2694), .A2(new_n7333), .B1(new_n7316), .B2(new_n2932), .C(new_n15430), .Y(new_n15431));
  XNOR2x2_ASAP7_75t_L       g15175(.A(\a[29] ), .B(new_n15431), .Y(new_n15432));
  INVx1_ASAP7_75t_L         g15176(.A(new_n15432), .Y(new_n15433));
  MAJIxp5_ASAP7_75t_L       g15177(.A(new_n15351), .B(new_n15354), .C(new_n15355), .Y(new_n15434));
  XNOR2x2_ASAP7_75t_L       g15178(.A(new_n15433), .B(new_n15434), .Y(new_n15435));
  OR2x4_ASAP7_75t_L         g15179(.A(new_n15344), .B(new_n15341), .Y(new_n15436));
  A2O1A1Ixp33_ASAP7_75t_L   g15180(.A1(new_n15189), .A2(new_n15274), .B(new_n15345), .C(new_n15436), .Y(new_n15437));
  AOI22xp33_ASAP7_75t_L     g15181(.A1(new_n4544), .A2(\b[40] ), .B1(new_n4542), .B2(new_n5194), .Y(new_n15438));
  OAI221xp5_ASAP7_75t_L     g15182(.A1(new_n4536), .A2(new_n5166), .B1(new_n4915), .B2(new_n4781), .C(new_n15438), .Y(new_n15439));
  XNOR2x2_ASAP7_75t_L       g15183(.A(\a[38] ), .B(new_n15439), .Y(new_n15440));
  NOR2xp33_ASAP7_75t_L      g15184(.A(new_n15340), .B(new_n15338), .Y(new_n15441));
  AOI21xp33_ASAP7_75t_L     g15185(.A1(new_n15337), .A2(new_n15278), .B(new_n15441), .Y(new_n15442));
  AOI22xp33_ASAP7_75t_L     g15186(.A1(new_n5249), .A2(\b[37] ), .B1(new_n5247), .B2(new_n4709), .Y(new_n15443));
  OAI221xp5_ASAP7_75t_L     g15187(.A1(new_n5241), .A2(new_n4465), .B1(new_n4053), .B2(new_n5521), .C(new_n15443), .Y(new_n15444));
  XNOR2x2_ASAP7_75t_L       g15188(.A(\a[41] ), .B(new_n15444), .Y(new_n15445));
  INVx1_ASAP7_75t_L         g15189(.A(new_n15445), .Y(new_n15446));
  INVx1_ASAP7_75t_L         g15190(.A(new_n15335), .Y(new_n15447));
  NAND2xp33_ASAP7_75t_L     g15191(.A(new_n15279), .B(new_n15336), .Y(new_n15448));
  OAI21xp33_ASAP7_75t_L     g15192(.A1(new_n15282), .A2(new_n15447), .B(new_n15448), .Y(new_n15449));
  AOI22xp33_ASAP7_75t_L     g15193(.A1(new_n6002), .A2(\b[34] ), .B1(new_n5999), .B2(new_n3833), .Y(new_n15450));
  OAI221xp5_ASAP7_75t_L     g15194(.A1(new_n6544), .A2(new_n3807), .B1(new_n3443), .B2(new_n6309), .C(new_n15450), .Y(new_n15451));
  XNOR2x2_ASAP7_75t_L       g15195(.A(\a[44] ), .B(new_n15451), .Y(new_n15452));
  INVx1_ASAP7_75t_L         g15196(.A(new_n15452), .Y(new_n15453));
  AOI22xp33_ASAP7_75t_L     g15197(.A1(new_n6822), .A2(\b[31] ), .B1(new_n6819), .B2(new_n3426), .Y(new_n15454));
  OAI221xp5_ASAP7_75t_L     g15198(.A1(new_n7392), .A2(new_n3212), .B1(new_n2871), .B2(new_n7115), .C(new_n15454), .Y(new_n15455));
  XNOR2x2_ASAP7_75t_L       g15199(.A(\a[47] ), .B(new_n15455), .Y(new_n15456));
  NOR2xp33_ASAP7_75t_L      g15200(.A(new_n15326), .B(new_n15323), .Y(new_n15457));
  NAND2xp33_ASAP7_75t_L     g15201(.A(new_n15326), .B(new_n15323), .Y(new_n15458));
  O2A1O1Ixp33_ASAP7_75t_L   g15202(.A1(new_n15156), .A2(new_n15154), .B(new_n15458), .C(new_n15457), .Y(new_n15459));
  NOR2xp33_ASAP7_75t_L      g15203(.A(new_n763), .B(new_n12671), .Y(new_n15460));
  O2A1O1Ixp33_ASAP7_75t_L   g15204(.A1(new_n12353), .A2(new_n12355), .B(\b[13] ), .C(new_n15460), .Y(new_n15461));
  A2O1A1Ixp33_ASAP7_75t_L   g15205(.A1(new_n12669), .A2(\b[10] ), .B(new_n14921), .C(new_n594), .Y(new_n15462));
  A2O1A1Ixp33_ASAP7_75t_L   g15206(.A1(new_n15297), .A2(new_n15295), .B(new_n15294), .C(new_n15462), .Y(new_n15463));
  INVx1_ASAP7_75t_L         g15207(.A(new_n15463), .Y(new_n15464));
  NAND2xp33_ASAP7_75t_L     g15208(.A(new_n15461), .B(new_n15464), .Y(new_n15465));
  A2O1A1Ixp33_ASAP7_75t_L   g15209(.A1(new_n12669), .A2(\b[13] ), .B(new_n15460), .C(new_n15463), .Y(new_n15466));
  AND2x2_ASAP7_75t_L        g15210(.A(new_n15466), .B(new_n15465), .Y(new_n15467));
  AOI22xp33_ASAP7_75t_L     g15211(.A1(new_n11656), .A2(\b[16] ), .B1(new_n11654), .B2(new_n1058), .Y(new_n15468));
  OAI221xp5_ASAP7_75t_L     g15212(.A1(new_n12364), .A2(new_n952), .B1(new_n871), .B2(new_n13003), .C(new_n15468), .Y(new_n15469));
  XNOR2x2_ASAP7_75t_L       g15213(.A(\a[62] ), .B(new_n15469), .Y(new_n15470));
  XOR2x2_ASAP7_75t_L        g15214(.A(new_n15467), .B(new_n15470), .Y(new_n15471));
  A2O1A1Ixp33_ASAP7_75t_L   g15215(.A1(\b[11] ), .A2(new_n12669), .B(new_n15120), .C(new_n14922), .Y(new_n15472));
  INVx1_ASAP7_75t_L         g15216(.A(new_n15288), .Y(new_n15473));
  NAND2xp33_ASAP7_75t_L     g15217(.A(new_n15300), .B(new_n15292), .Y(new_n15474));
  A2O1A1Ixp33_ASAP7_75t_L   g15218(.A1(new_n15473), .A2(new_n15472), .B(new_n15301), .C(new_n15474), .Y(new_n15475));
  OR2x4_ASAP7_75t_L         g15219(.A(new_n15471), .B(new_n15475), .Y(new_n15476));
  O2A1O1Ixp33_ASAP7_75t_L   g15220(.A1(new_n14927), .A2(new_n15121), .B(new_n15473), .C(new_n15301), .Y(new_n15477));
  A2O1A1Ixp33_ASAP7_75t_L   g15221(.A1(new_n15292), .A2(new_n15300), .B(new_n15477), .C(new_n15471), .Y(new_n15478));
  NAND2xp33_ASAP7_75t_L     g15222(.A(new_n15478), .B(new_n15476), .Y(new_n15479));
  OAI22xp33_ASAP7_75t_L     g15223(.A1(new_n2793), .A2(new_n10974), .B1(new_n10975), .B2(new_n1493), .Y(new_n15480));
  AOI221xp5_ASAP7_75t_L     g15224(.A1(\b[17] ), .A2(new_n10973), .B1(\b[18] ), .B2(new_n10584), .C(new_n15480), .Y(new_n15481));
  XNOR2x2_ASAP7_75t_L       g15225(.A(\a[59] ), .B(new_n15481), .Y(new_n15482));
  OR2x4_ASAP7_75t_L         g15226(.A(new_n15482), .B(new_n15479), .Y(new_n15483));
  NAND2xp33_ASAP7_75t_L     g15227(.A(new_n15482), .B(new_n15479), .Y(new_n15484));
  NAND4xp25_ASAP7_75t_L     g15228(.A(new_n15313), .B(new_n15483), .C(new_n15484), .D(new_n15307), .Y(new_n15485));
  INVx1_ASAP7_75t_L         g15229(.A(new_n15313), .Y(new_n15486));
  NAND2xp33_ASAP7_75t_L     g15230(.A(new_n15484), .B(new_n15483), .Y(new_n15487));
  A2O1A1Ixp33_ASAP7_75t_L   g15231(.A1(new_n15306), .A2(new_n15302), .B(new_n15486), .C(new_n15487), .Y(new_n15488));
  AOI22xp33_ASAP7_75t_L     g15232(.A1(new_n9623), .A2(\b[22] ), .B1(new_n9620), .B2(new_n1864), .Y(new_n15489));
  OAI221xp5_ASAP7_75t_L     g15233(.A1(new_n10280), .A2(new_n1709), .B1(new_n1594), .B2(new_n12010), .C(new_n15489), .Y(new_n15490));
  XNOR2x2_ASAP7_75t_L       g15234(.A(\a[56] ), .B(new_n15490), .Y(new_n15491));
  NAND3xp33_ASAP7_75t_L     g15235(.A(new_n15488), .B(new_n15485), .C(new_n15491), .Y(new_n15492));
  NAND2xp33_ASAP7_75t_L     g15236(.A(new_n15485), .B(new_n15488), .Y(new_n15493));
  INVx1_ASAP7_75t_L         g15237(.A(new_n15491), .Y(new_n15494));
  NAND2xp33_ASAP7_75t_L     g15238(.A(new_n15494), .B(new_n15493), .Y(new_n15495));
  AND2x2_ASAP7_75t_L        g15239(.A(new_n15492), .B(new_n15495), .Y(new_n15496));
  O2A1O1Ixp33_ASAP7_75t_L   g15240(.A1(new_n15143), .A2(new_n15146), .B(new_n15142), .C(new_n15318), .Y(new_n15497));
  NOR2xp33_ASAP7_75t_L      g15241(.A(new_n15317), .B(new_n15314), .Y(new_n15498));
  NOR2xp33_ASAP7_75t_L      g15242(.A(new_n15498), .B(new_n15497), .Y(new_n15499));
  XOR2x2_ASAP7_75t_L        g15243(.A(new_n15496), .B(new_n15499), .Y(new_n15500));
  AOI22xp33_ASAP7_75t_L     g15244(.A1(new_n8645), .A2(\b[25] ), .B1(new_n8642), .B2(new_n2188), .Y(new_n15501));
  OAI221xp5_ASAP7_75t_L     g15245(.A1(new_n9322), .A2(new_n2019), .B1(new_n1995), .B2(new_n8965), .C(new_n15501), .Y(new_n15502));
  XNOR2x2_ASAP7_75t_L       g15246(.A(\a[53] ), .B(new_n15502), .Y(new_n15503));
  NAND2xp33_ASAP7_75t_L     g15247(.A(new_n15503), .B(new_n15500), .Y(new_n15504));
  NAND2xp33_ASAP7_75t_L     g15248(.A(new_n15496), .B(new_n15499), .Y(new_n15505));
  AO21x2_ASAP7_75t_L        g15249(.A1(new_n15492), .A2(new_n15495), .B(new_n15499), .Y(new_n15506));
  AO21x2_ASAP7_75t_L        g15250(.A1(new_n15505), .A2(new_n15506), .B(new_n15503), .Y(new_n15507));
  INVx1_ASAP7_75t_L         g15251(.A(new_n15287), .Y(new_n15508));
  MAJIxp5_ASAP7_75t_L       g15252(.A(new_n15321), .B(new_n15284), .C(new_n15508), .Y(new_n15509));
  NAND3xp33_ASAP7_75t_L     g15253(.A(new_n15504), .B(new_n15507), .C(new_n15509), .Y(new_n15510));
  NAND2xp33_ASAP7_75t_L     g15254(.A(new_n15507), .B(new_n15504), .Y(new_n15511));
  AND2x2_ASAP7_75t_L        g15255(.A(new_n15284), .B(new_n15322), .Y(new_n15512));
  A2O1A1Ixp33_ASAP7_75t_L   g15256(.A1(new_n15508), .A2(new_n15321), .B(new_n15512), .C(new_n15511), .Y(new_n15513));
  NAND2xp33_ASAP7_75t_L     g15257(.A(new_n15510), .B(new_n15513), .Y(new_n15514));
  AOI22xp33_ASAP7_75t_L     g15258(.A1(new_n7659), .A2(\b[28] ), .B1(new_n7656), .B2(new_n2858), .Y(new_n15515));
  OAI221xp5_ASAP7_75t_L     g15259(.A1(new_n8326), .A2(new_n2650), .B1(new_n2477), .B2(new_n7994), .C(new_n15515), .Y(new_n15516));
  XNOR2x2_ASAP7_75t_L       g15260(.A(\a[50] ), .B(new_n15516), .Y(new_n15517));
  NAND2xp33_ASAP7_75t_L     g15261(.A(new_n15517), .B(new_n15514), .Y(new_n15518));
  INVx1_ASAP7_75t_L         g15262(.A(new_n15517), .Y(new_n15519));
  NAND3xp33_ASAP7_75t_L     g15263(.A(new_n15510), .B(new_n15513), .C(new_n15519), .Y(new_n15520));
  NAND2xp33_ASAP7_75t_L     g15264(.A(new_n15520), .B(new_n15518), .Y(new_n15521));
  XNOR2x2_ASAP7_75t_L       g15265(.A(new_n15459), .B(new_n15521), .Y(new_n15522));
  XNOR2x2_ASAP7_75t_L       g15266(.A(new_n15456), .B(new_n15522), .Y(new_n15523));
  NAND2xp33_ASAP7_75t_L     g15267(.A(new_n15331), .B(new_n15328), .Y(new_n15524));
  OR2x4_ASAP7_75t_L         g15268(.A(new_n15331), .B(new_n15328), .Y(new_n15525));
  NAND3xp33_ASAP7_75t_L     g15269(.A(new_n15334), .B(new_n15525), .C(new_n15524), .Y(new_n15526));
  NAND2xp33_ASAP7_75t_L     g15270(.A(new_n15524), .B(new_n15526), .Y(new_n15527));
  XNOR2x2_ASAP7_75t_L       g15271(.A(new_n15527), .B(new_n15523), .Y(new_n15528));
  XNOR2x2_ASAP7_75t_L       g15272(.A(new_n15453), .B(new_n15528), .Y(new_n15529));
  XNOR2x2_ASAP7_75t_L       g15273(.A(new_n15449), .B(new_n15529), .Y(new_n15530));
  XNOR2x2_ASAP7_75t_L       g15274(.A(new_n15446), .B(new_n15530), .Y(new_n15531));
  XOR2x2_ASAP7_75t_L        g15275(.A(new_n15442), .B(new_n15531), .Y(new_n15532));
  XNOR2x2_ASAP7_75t_L       g15276(.A(new_n15440), .B(new_n15532), .Y(new_n15533));
  NAND2xp33_ASAP7_75t_L     g15277(.A(new_n15437), .B(new_n15533), .Y(new_n15534));
  INVx1_ASAP7_75t_L         g15278(.A(new_n15440), .Y(new_n15535));
  AND2x2_ASAP7_75t_L        g15279(.A(new_n15535), .B(new_n15532), .Y(new_n15536));
  NOR2xp33_ASAP7_75t_L      g15280(.A(new_n15535), .B(new_n15532), .Y(new_n15537));
  OAI211xp5_ASAP7_75t_L     g15281(.A1(new_n15537), .A2(new_n15536), .B(new_n15436), .C(new_n15346), .Y(new_n15538));
  NAND2xp33_ASAP7_75t_L     g15282(.A(new_n15538), .B(new_n15534), .Y(new_n15539));
  NAND2xp33_ASAP7_75t_L     g15283(.A(\b[43] ), .B(new_n3884), .Y(new_n15540));
  OAI221xp5_ASAP7_75t_L     g15284(.A1(new_n5680), .A2(new_n4312), .B1(new_n4114), .B2(new_n9799), .C(new_n15540), .Y(new_n15541));
  AOI21xp33_ASAP7_75t_L     g15285(.A1(new_n4111), .A2(\b[41] ), .B(new_n15541), .Y(new_n15542));
  NAND2xp33_ASAP7_75t_L     g15286(.A(\a[35] ), .B(new_n15542), .Y(new_n15543));
  A2O1A1Ixp33_ASAP7_75t_L   g15287(.A1(\b[41] ), .A2(new_n4111), .B(new_n15541), .C(new_n3878), .Y(new_n15544));
  NAND2xp33_ASAP7_75t_L     g15288(.A(new_n15544), .B(new_n15543), .Y(new_n15545));
  XOR2x2_ASAP7_75t_L        g15289(.A(new_n15545), .B(new_n15539), .Y(new_n15546));
  MAJx2_ASAP7_75t_L         g15290(.A(new_n15348), .B(new_n15273), .C(new_n15350), .Y(new_n15547));
  AOI22xp33_ASAP7_75t_L     g15291(.A1(new_n3260), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n3256), .Y(new_n15548));
  OAI221xp5_ASAP7_75t_L     g15292(.A1(new_n3492), .A2(new_n6220), .B1(new_n3261), .B2(new_n7887), .C(new_n15548), .Y(new_n15549));
  XNOR2x2_ASAP7_75t_L       g15293(.A(\a[32] ), .B(new_n15549), .Y(new_n15550));
  XNOR2x2_ASAP7_75t_L       g15294(.A(new_n15550), .B(new_n15547), .Y(new_n15551));
  XOR2x2_ASAP7_75t_L        g15295(.A(new_n15551), .B(new_n15546), .Y(new_n15552));
  XOR2x2_ASAP7_75t_L        g15296(.A(new_n15552), .B(new_n15435), .Y(new_n15553));
  O2A1O1Ixp33_ASAP7_75t_L   g15297(.A1(new_n15095), .A2(new_n15193), .B(new_n15094), .C(new_n15264), .Y(new_n15554));
  AOI22xp33_ASAP7_75t_L     g15298(.A1(new_n2232), .A2(\b[51] ), .B1(\b[52] ), .B2(new_n2228), .Y(new_n15555));
  OAI221xp5_ASAP7_75t_L     g15299(.A1(new_n2387), .A2(new_n8228), .B1(new_n2233), .B2(new_n10519), .C(new_n15555), .Y(new_n15556));
  XNOR2x2_ASAP7_75t_L       g15300(.A(\a[26] ), .B(new_n15556), .Y(new_n15557));
  INVx1_ASAP7_75t_L         g15301(.A(new_n15557), .Y(new_n15558));
  A2O1A1Ixp33_ASAP7_75t_L   g15302(.A1(new_n15270), .A2(new_n15359), .B(new_n15554), .C(new_n15558), .Y(new_n15559));
  INVx1_ASAP7_75t_L         g15303(.A(new_n15269), .Y(new_n15560));
  O2A1O1Ixp33_ASAP7_75t_L   g15304(.A1(new_n15266), .A2(new_n15560), .B(new_n15359), .C(new_n15554), .Y(new_n15561));
  NAND2xp33_ASAP7_75t_L     g15305(.A(new_n15557), .B(new_n15561), .Y(new_n15562));
  NAND2xp33_ASAP7_75t_L     g15306(.A(new_n15559), .B(new_n15562), .Y(new_n15563));
  XOR2x2_ASAP7_75t_L        g15307(.A(new_n15553), .B(new_n15563), .Y(new_n15564));
  XNOR2x2_ASAP7_75t_L       g15308(.A(new_n15429), .B(new_n15564), .Y(new_n15565));
  XOR2x2_ASAP7_75t_L        g15309(.A(new_n15565), .B(new_n15424), .Y(new_n15566));
  XOR2x2_ASAP7_75t_L        g15310(.A(new_n15566), .B(new_n15414), .Y(new_n15567));
  NOR2xp33_ASAP7_75t_L      g15311(.A(new_n15409), .B(new_n15567), .Y(new_n15568));
  XNOR2x2_ASAP7_75t_L       g15312(.A(new_n15404), .B(new_n15407), .Y(new_n15569));
  XNOR2x2_ASAP7_75t_L       g15313(.A(new_n15566), .B(new_n15414), .Y(new_n15570));
  NOR2xp33_ASAP7_75t_L      g15314(.A(new_n15569), .B(new_n15570), .Y(new_n15571));
  NOR3xp33_ASAP7_75t_L      g15315(.A(new_n15568), .B(new_n15571), .C(new_n15397), .Y(new_n15572));
  OA21x2_ASAP7_75t_L        g15316(.A1(new_n15571), .A2(new_n15568), .B(new_n15397), .Y(new_n15573));
  NOR2xp33_ASAP7_75t_L      g15317(.A(new_n15572), .B(new_n15573), .Y(new_n15574));
  INVx1_ASAP7_75t_L         g15318(.A(new_n15574), .Y(new_n15575));
  O2A1O1Ixp33_ASAP7_75t_L   g15319(.A1(new_n15394), .A2(new_n15391), .B(new_n15387), .C(new_n15575), .Y(new_n15576));
  INVx1_ASAP7_75t_L         g15320(.A(new_n15220), .Y(new_n15577));
  A2O1A1Ixp33_ASAP7_75t_L   g15321(.A1(new_n15223), .A2(new_n15577), .B(new_n15391), .C(new_n15387), .Y(new_n15578));
  NOR2xp33_ASAP7_75t_L      g15322(.A(new_n15574), .B(new_n15578), .Y(new_n15579));
  NOR2xp33_ASAP7_75t_L      g15323(.A(new_n15579), .B(new_n15576), .Y(\f[76] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g15324(.A1(new_n15233), .A2(new_n15367), .B(new_n15368), .C(new_n15399), .D(new_n15404), .Y(new_n15581));
  O2A1O1Ixp33_ASAP7_75t_L   g15325(.A1(new_n15406), .A2(new_n15408), .B(new_n15570), .C(new_n15581), .Y(new_n15582));
  A2O1A1Ixp33_ASAP7_75t_L   g15326(.A1(new_n15253), .A2(new_n15361), .B(new_n15415), .C(new_n15422), .Y(new_n15583));
  AOI22xp33_ASAP7_75t_L     g15327(.A1(new_n1103), .A2(\b[61] ), .B1(\b[62] ), .B2(new_n1113), .Y(new_n15584));
  OAI221xp5_ASAP7_75t_L     g15328(.A1(new_n1195), .A2(new_n11226), .B1(new_n1197), .B2(new_n12281), .C(new_n15584), .Y(new_n15585));
  NOR2xp33_ASAP7_75t_L      g15329(.A(new_n1107), .B(new_n15585), .Y(new_n15586));
  AND2x2_ASAP7_75t_L        g15330(.A(new_n1107), .B(new_n15585), .Y(new_n15587));
  NOR2xp33_ASAP7_75t_L      g15331(.A(new_n15586), .B(new_n15587), .Y(new_n15588));
  INVx1_ASAP7_75t_L         g15332(.A(new_n15588), .Y(new_n15589));
  A2O1A1O1Ixp25_ASAP7_75t_L g15333(.A1(new_n15423), .A2(new_n15419), .B(new_n15565), .C(new_n15583), .D(new_n15589), .Y(new_n15590));
  A2O1A1Ixp33_ASAP7_75t_L   g15334(.A1(new_n15423), .A2(new_n15419), .B(new_n15565), .C(new_n15583), .Y(new_n15591));
  NOR2xp33_ASAP7_75t_L      g15335(.A(new_n15588), .B(new_n15591), .Y(new_n15592));
  AOI22xp33_ASAP7_75t_L     g15336(.A1(new_n1406), .A2(\b[59] ), .B1(new_n1404), .B2(new_n10887), .Y(new_n15593));
  OAI221xp5_ASAP7_75t_L     g15337(.A1(new_n1398), .A2(new_n10848), .B1(new_n10488), .B2(new_n1549), .C(new_n15593), .Y(new_n15594));
  XNOR2x2_ASAP7_75t_L       g15338(.A(\a[20] ), .B(new_n15594), .Y(new_n15595));
  O2A1O1Ixp33_ASAP7_75t_L   g15339(.A1(new_n15258), .A2(new_n15360), .B(new_n15259), .C(new_n15427), .Y(new_n15596));
  AOI21xp33_ASAP7_75t_L     g15340(.A1(new_n15564), .A2(new_n15429), .B(new_n15596), .Y(new_n15597));
  AND2x2_ASAP7_75t_L        g15341(.A(new_n15595), .B(new_n15597), .Y(new_n15598));
  NOR2xp33_ASAP7_75t_L      g15342(.A(new_n15595), .B(new_n15597), .Y(new_n15599));
  NOR2xp33_ASAP7_75t_L      g15343(.A(new_n15599), .B(new_n15598), .Y(new_n15600));
  AOI22xp33_ASAP7_75t_L     g15344(.A1(new_n1766), .A2(\b[56] ), .B1(new_n1764), .B2(new_n10185), .Y(new_n15601));
  OAI221xp5_ASAP7_75t_L     g15345(.A1(new_n1758), .A2(new_n9534), .B1(new_n9199), .B2(new_n1911), .C(new_n15601), .Y(new_n15602));
  XNOR2x2_ASAP7_75t_L       g15346(.A(\a[23] ), .B(new_n15602), .Y(new_n15603));
  MAJx2_ASAP7_75t_L         g15347(.A(new_n15561), .B(new_n15553), .C(new_n15557), .Y(new_n15604));
  NAND2xp33_ASAP7_75t_L     g15348(.A(new_n15603), .B(new_n15604), .Y(new_n15605));
  NOR2xp33_ASAP7_75t_L      g15349(.A(new_n15603), .B(new_n15604), .Y(new_n15606));
  INVx1_ASAP7_75t_L         g15350(.A(new_n15606), .Y(new_n15607));
  NAND2xp33_ASAP7_75t_L     g15351(.A(\b[53] ), .B(new_n2228), .Y(new_n15608));
  OAI221xp5_ASAP7_75t_L     g15352(.A1(new_n8569), .A2(new_n2220), .B1(new_n2233), .B2(new_n8888), .C(new_n15608), .Y(new_n15609));
  AOI21xp33_ASAP7_75t_L     g15353(.A1(new_n2386), .A2(\b[51] ), .B(new_n15609), .Y(new_n15610));
  NAND2xp33_ASAP7_75t_L     g15354(.A(\a[26] ), .B(new_n15610), .Y(new_n15611));
  A2O1A1Ixp33_ASAP7_75t_L   g15355(.A1(\b[51] ), .A2(new_n2386), .B(new_n15609), .C(new_n2223), .Y(new_n15612));
  NAND2xp33_ASAP7_75t_L     g15356(.A(new_n15612), .B(new_n15611), .Y(new_n15613));
  MAJIxp5_ASAP7_75t_L       g15357(.A(new_n15552), .B(new_n15433), .C(new_n15434), .Y(new_n15614));
  INVx1_ASAP7_75t_L         g15358(.A(new_n15614), .Y(new_n15615));
  NOR2xp33_ASAP7_75t_L      g15359(.A(new_n15613), .B(new_n15615), .Y(new_n15616));
  INVx1_ASAP7_75t_L         g15360(.A(new_n15616), .Y(new_n15617));
  NAND2xp33_ASAP7_75t_L     g15361(.A(new_n15613), .B(new_n15615), .Y(new_n15618));
  NAND2xp33_ASAP7_75t_L     g15362(.A(new_n15618), .B(new_n15617), .Y(new_n15619));
  AOI22xp33_ASAP7_75t_L     g15363(.A1(new_n3260), .A2(\b[46] ), .B1(\b[47] ), .B2(new_n3256), .Y(new_n15620));
  OAI221xp5_ASAP7_75t_L     g15364(.A1(new_n3492), .A2(new_n6756), .B1(new_n3261), .B2(new_n7322), .C(new_n15620), .Y(new_n15621));
  XNOR2x2_ASAP7_75t_L       g15365(.A(\a[32] ), .B(new_n15621), .Y(new_n15622));
  INVx1_ASAP7_75t_L         g15366(.A(new_n15622), .Y(new_n15623));
  OAI211xp5_ASAP7_75t_L     g15367(.A1(new_n15545), .A2(new_n15539), .B(new_n15538), .C(new_n15623), .Y(new_n15624));
  INVx1_ASAP7_75t_L         g15368(.A(new_n15538), .Y(new_n15625));
  INVx1_ASAP7_75t_L         g15369(.A(new_n15545), .Y(new_n15626));
  A2O1A1Ixp33_ASAP7_75t_L   g15370(.A1(new_n15534), .A2(new_n15626), .B(new_n15625), .C(new_n15622), .Y(new_n15627));
  AOI22xp33_ASAP7_75t_L     g15371(.A1(new_n3884), .A2(\b[44] ), .B1(new_n3881), .B2(new_n7055), .Y(new_n15628));
  OAI221xp5_ASAP7_75t_L     g15372(.A1(new_n4312), .A2(new_n6195), .B1(new_n5680), .B2(new_n4986), .C(new_n15628), .Y(new_n15629));
  XNOR2x2_ASAP7_75t_L       g15373(.A(\a[35] ), .B(new_n15629), .Y(new_n15630));
  NOR2xp33_ASAP7_75t_L      g15374(.A(new_n15442), .B(new_n15531), .Y(new_n15631));
  NOR2xp33_ASAP7_75t_L      g15375(.A(new_n15631), .B(new_n15536), .Y(new_n15632));
  AOI22xp33_ASAP7_75t_L     g15376(.A1(new_n4544), .A2(\b[41] ), .B1(new_n4542), .B2(new_n5669), .Y(new_n15633));
  OAI221xp5_ASAP7_75t_L     g15377(.A1(new_n4536), .A2(new_n5186), .B1(new_n5166), .B2(new_n4781), .C(new_n15633), .Y(new_n15634));
  XNOR2x2_ASAP7_75t_L       g15378(.A(new_n4539), .B(new_n15634), .Y(new_n15635));
  O2A1O1Ixp33_ASAP7_75t_L   g15379(.A1(new_n15282), .A2(new_n15447), .B(new_n15448), .C(new_n15529), .Y(new_n15636));
  AO21x2_ASAP7_75t_L        g15380(.A1(new_n15446), .A2(new_n15530), .B(new_n15636), .Y(new_n15637));
  MAJIxp5_ASAP7_75t_L       g15381(.A(new_n15521), .B(new_n15456), .C(new_n15459), .Y(new_n15638));
  AOI22xp33_ASAP7_75t_L     g15382(.A1(new_n6822), .A2(\b[32] ), .B1(new_n6819), .B2(new_n3450), .Y(new_n15639));
  OAI221xp5_ASAP7_75t_L     g15383(.A1(new_n7392), .A2(new_n3419), .B1(new_n3212), .B2(new_n7115), .C(new_n15639), .Y(new_n15640));
  XNOR2x2_ASAP7_75t_L       g15384(.A(\a[47] ), .B(new_n15640), .Y(new_n15641));
  INVx1_ASAP7_75t_L         g15385(.A(new_n15641), .Y(new_n15642));
  AOI22xp33_ASAP7_75t_L     g15386(.A1(new_n8645), .A2(\b[26] ), .B1(new_n8642), .B2(new_n2888), .Y(new_n15643));
  OAI221xp5_ASAP7_75t_L     g15387(.A1(new_n9322), .A2(new_n2180), .B1(new_n2019), .B2(new_n8965), .C(new_n15643), .Y(new_n15644));
  XNOR2x2_ASAP7_75t_L       g15388(.A(\a[53] ), .B(new_n15644), .Y(new_n15645));
  INVx1_ASAP7_75t_L         g15389(.A(new_n15645), .Y(new_n15646));
  A2O1A1Ixp33_ASAP7_75t_L   g15390(.A1(new_n14927), .A2(new_n594), .B(new_n15298), .C(new_n15461), .Y(new_n15647));
  A2O1A1Ixp33_ASAP7_75t_L   g15391(.A1(new_n15466), .A2(new_n15465), .B(new_n15470), .C(new_n15647), .Y(new_n15648));
  NOR2xp33_ASAP7_75t_L      g15392(.A(new_n793), .B(new_n12671), .Y(new_n15649));
  A2O1A1Ixp33_ASAP7_75t_L   g15393(.A1(\b[14] ), .A2(new_n12669), .B(new_n15649), .C(new_n15461), .Y(new_n15650));
  O2A1O1Ixp33_ASAP7_75t_L   g15394(.A1(new_n12353), .A2(new_n12355), .B(\b[14] ), .C(new_n15649), .Y(new_n15651));
  A2O1A1Ixp33_ASAP7_75t_L   g15395(.A1(new_n12669), .A2(\b[13] ), .B(new_n15460), .C(new_n15651), .Y(new_n15652));
  NAND2xp33_ASAP7_75t_L     g15396(.A(new_n15652), .B(new_n15650), .Y(new_n15653));
  AOI22xp33_ASAP7_75t_L     g15397(.A1(new_n11647), .A2(\b[16] ), .B1(\b[17] ), .B2(new_n11656), .Y(new_n15654));
  OAI221xp5_ASAP7_75t_L     g15398(.A1(new_n13003), .A2(new_n952), .B1(new_n12022), .B2(new_n1251), .C(new_n15654), .Y(new_n15655));
  XNOR2x2_ASAP7_75t_L       g15399(.A(\a[62] ), .B(new_n15655), .Y(new_n15656));
  NOR2xp33_ASAP7_75t_L      g15400(.A(new_n15653), .B(new_n15656), .Y(new_n15657));
  AND2x2_ASAP7_75t_L        g15401(.A(new_n15653), .B(new_n15656), .Y(new_n15658));
  NOR2xp33_ASAP7_75t_L      g15402(.A(new_n15657), .B(new_n15658), .Y(new_n15659));
  NAND2xp33_ASAP7_75t_L     g15403(.A(new_n15648), .B(new_n15659), .Y(new_n15660));
  NOR2xp33_ASAP7_75t_L      g15404(.A(new_n15648), .B(new_n15659), .Y(new_n15661));
  INVx1_ASAP7_75t_L         g15405(.A(new_n15661), .Y(new_n15662));
  AOI22xp33_ASAP7_75t_L     g15406(.A1(new_n10594), .A2(\b[20] ), .B1(new_n10591), .B2(new_n1600), .Y(new_n15663));
  OAI221xp5_ASAP7_75t_L     g15407(.A1(new_n11335), .A2(new_n1493), .B1(new_n1356), .B2(new_n11330), .C(new_n15663), .Y(new_n15664));
  XNOR2x2_ASAP7_75t_L       g15408(.A(\a[59] ), .B(new_n15664), .Y(new_n15665));
  NAND3xp33_ASAP7_75t_L     g15409(.A(new_n15665), .B(new_n15662), .C(new_n15660), .Y(new_n15666));
  AO21x2_ASAP7_75t_L        g15410(.A1(new_n15660), .A2(new_n15662), .B(new_n15665), .Y(new_n15667));
  NAND2xp33_ASAP7_75t_L     g15411(.A(new_n15666), .B(new_n15667), .Y(new_n15668));
  O2A1O1Ixp33_ASAP7_75t_L   g15412(.A1(new_n15479), .A2(new_n15482), .B(new_n15476), .C(new_n15668), .Y(new_n15669));
  NAND2xp33_ASAP7_75t_L     g15413(.A(new_n15476), .B(new_n15483), .Y(new_n15670));
  AOI21xp33_ASAP7_75t_L     g15414(.A1(new_n15667), .A2(new_n15666), .B(new_n15670), .Y(new_n15671));
  NOR2xp33_ASAP7_75t_L      g15415(.A(new_n15669), .B(new_n15671), .Y(new_n15672));
  AOI22xp33_ASAP7_75t_L     g15416(.A1(new_n9623), .A2(\b[23] ), .B1(new_n9620), .B2(new_n2002), .Y(new_n15673));
  OAI221xp5_ASAP7_75t_L     g15417(.A1(new_n10280), .A2(new_n1857), .B1(new_n1709), .B2(new_n12010), .C(new_n15673), .Y(new_n15674));
  XNOR2x2_ASAP7_75t_L       g15418(.A(new_n9610), .B(new_n15674), .Y(new_n15675));
  XOR2x2_ASAP7_75t_L        g15419(.A(new_n15675), .B(new_n15672), .Y(new_n15676));
  INVx1_ASAP7_75t_L         g15420(.A(new_n15676), .Y(new_n15677));
  NAND2xp33_ASAP7_75t_L     g15421(.A(new_n15485), .B(new_n15492), .Y(new_n15678));
  NOR2xp33_ASAP7_75t_L      g15422(.A(new_n15678), .B(new_n15677), .Y(new_n15679));
  O2A1O1Ixp33_ASAP7_75t_L   g15423(.A1(new_n15493), .A2(new_n15494), .B(new_n15485), .C(new_n15676), .Y(new_n15680));
  NOR2xp33_ASAP7_75t_L      g15424(.A(new_n15680), .B(new_n15679), .Y(new_n15681));
  NAND2xp33_ASAP7_75t_L     g15425(.A(new_n15646), .B(new_n15681), .Y(new_n15682));
  NOR2xp33_ASAP7_75t_L      g15426(.A(new_n15646), .B(new_n15681), .Y(new_n15683));
  INVx1_ASAP7_75t_L         g15427(.A(new_n15683), .Y(new_n15684));
  NAND2xp33_ASAP7_75t_L     g15428(.A(new_n15682), .B(new_n15684), .Y(new_n15685));
  NAND2xp33_ASAP7_75t_L     g15429(.A(new_n15505), .B(new_n15504), .Y(new_n15686));
  XOR2x2_ASAP7_75t_L        g15430(.A(new_n15686), .B(new_n15685), .Y(new_n15687));
  AOI22xp33_ASAP7_75t_L     g15431(.A1(new_n7659), .A2(\b[29] ), .B1(new_n7656), .B2(new_n5472), .Y(new_n15688));
  OAI221xp5_ASAP7_75t_L     g15432(.A1(new_n8326), .A2(new_n2852), .B1(new_n2650), .B2(new_n7994), .C(new_n15688), .Y(new_n15689));
  XNOR2x2_ASAP7_75t_L       g15433(.A(\a[50] ), .B(new_n15689), .Y(new_n15690));
  NAND2xp33_ASAP7_75t_L     g15434(.A(new_n15690), .B(new_n15687), .Y(new_n15691));
  INVx1_ASAP7_75t_L         g15435(.A(new_n15691), .Y(new_n15692));
  NOR2xp33_ASAP7_75t_L      g15436(.A(new_n15690), .B(new_n15687), .Y(new_n15693));
  NOR2xp33_ASAP7_75t_L      g15437(.A(new_n15693), .B(new_n15692), .Y(new_n15694));
  O2A1O1Ixp33_ASAP7_75t_L   g15438(.A1(new_n15514), .A2(new_n15517), .B(new_n15513), .C(new_n15694), .Y(new_n15695));
  A2O1A1Ixp33_ASAP7_75t_L   g15439(.A1(new_n15507), .A2(new_n15504), .B(new_n15509), .C(new_n15520), .Y(new_n15696));
  NOR3xp33_ASAP7_75t_L      g15440(.A(new_n15696), .B(new_n15693), .C(new_n15692), .Y(new_n15697));
  NOR3xp33_ASAP7_75t_L      g15441(.A(new_n15695), .B(new_n15697), .C(new_n15642), .Y(new_n15698));
  INVx1_ASAP7_75t_L         g15442(.A(new_n15698), .Y(new_n15699));
  OAI21xp33_ASAP7_75t_L     g15443(.A1(new_n15697), .A2(new_n15695), .B(new_n15642), .Y(new_n15700));
  NAND2xp33_ASAP7_75t_L     g15444(.A(new_n15700), .B(new_n15699), .Y(new_n15701));
  NOR2xp33_ASAP7_75t_L      g15445(.A(new_n15638), .B(new_n15701), .Y(new_n15702));
  INVx1_ASAP7_75t_L         g15446(.A(new_n15638), .Y(new_n15703));
  AND2x2_ASAP7_75t_L        g15447(.A(new_n15700), .B(new_n15699), .Y(new_n15704));
  NOR2xp33_ASAP7_75t_L      g15448(.A(new_n15703), .B(new_n15704), .Y(new_n15705));
  NOR2xp33_ASAP7_75t_L      g15449(.A(new_n15702), .B(new_n15705), .Y(new_n15706));
  AOI22xp33_ASAP7_75t_L     g15450(.A1(new_n6002), .A2(\b[35] ), .B1(new_n5999), .B2(new_n5649), .Y(new_n15707));
  OAI221xp5_ASAP7_75t_L     g15451(.A1(new_n6544), .A2(new_n3827), .B1(new_n3807), .B2(new_n6309), .C(new_n15707), .Y(new_n15708));
  XNOR2x2_ASAP7_75t_L       g15452(.A(\a[44] ), .B(new_n15708), .Y(new_n15709));
  NAND2xp33_ASAP7_75t_L     g15453(.A(new_n15709), .B(new_n15706), .Y(new_n15710));
  INVx1_ASAP7_75t_L         g15454(.A(new_n15709), .Y(new_n15711));
  OAI21xp33_ASAP7_75t_L     g15455(.A1(new_n15702), .A2(new_n15705), .B(new_n15711), .Y(new_n15712));
  NAND2xp33_ASAP7_75t_L     g15456(.A(new_n15712), .B(new_n15710), .Y(new_n15713));
  NAND2xp33_ASAP7_75t_L     g15457(.A(new_n15453), .B(new_n15528), .Y(new_n15714));
  A2O1A1Ixp33_ASAP7_75t_L   g15458(.A1(new_n15526), .A2(new_n15524), .B(new_n15523), .C(new_n15714), .Y(new_n15715));
  NOR2xp33_ASAP7_75t_L      g15459(.A(new_n15715), .B(new_n15713), .Y(new_n15716));
  INVx1_ASAP7_75t_L         g15460(.A(new_n15713), .Y(new_n15717));
  A2O1A1O1Ixp25_ASAP7_75t_L g15461(.A1(new_n15526), .A2(new_n15524), .B(new_n15523), .C(new_n15714), .D(new_n15717), .Y(new_n15718));
  AOI22xp33_ASAP7_75t_L     g15462(.A1(new_n5249), .A2(\b[38] ), .B1(new_n5247), .B2(new_n4923), .Y(new_n15719));
  OAI221xp5_ASAP7_75t_L     g15463(.A1(new_n5241), .A2(new_n4701), .B1(new_n4465), .B2(new_n5521), .C(new_n15719), .Y(new_n15720));
  XNOR2x2_ASAP7_75t_L       g15464(.A(\a[41] ), .B(new_n15720), .Y(new_n15721));
  OAI21xp33_ASAP7_75t_L     g15465(.A1(new_n15716), .A2(new_n15718), .B(new_n15721), .Y(new_n15722));
  XOR2x2_ASAP7_75t_L        g15466(.A(new_n15715), .B(new_n15713), .Y(new_n15723));
  INVx1_ASAP7_75t_L         g15467(.A(new_n15721), .Y(new_n15724));
  NAND2xp33_ASAP7_75t_L     g15468(.A(new_n15724), .B(new_n15723), .Y(new_n15725));
  NAND3xp33_ASAP7_75t_L     g15469(.A(new_n15722), .B(new_n15637), .C(new_n15725), .Y(new_n15726));
  AO21x2_ASAP7_75t_L        g15470(.A1(new_n15725), .A2(new_n15722), .B(new_n15637), .Y(new_n15727));
  NAND3xp33_ASAP7_75t_L     g15471(.A(new_n15727), .B(new_n15726), .C(new_n15635), .Y(new_n15728));
  AO21x2_ASAP7_75t_L        g15472(.A1(new_n15726), .A2(new_n15727), .B(new_n15635), .Y(new_n15729));
  NAND2xp33_ASAP7_75t_L     g15473(.A(new_n15728), .B(new_n15729), .Y(new_n15730));
  XOR2x2_ASAP7_75t_L        g15474(.A(new_n15632), .B(new_n15730), .Y(new_n15731));
  XOR2x2_ASAP7_75t_L        g15475(.A(new_n15630), .B(new_n15731), .Y(new_n15732));
  NAND3xp33_ASAP7_75t_L     g15476(.A(new_n15732), .B(new_n15624), .C(new_n15627), .Y(new_n15733));
  AO21x2_ASAP7_75t_L        g15477(.A1(new_n15627), .A2(new_n15624), .B(new_n15732), .Y(new_n15734));
  NAND2xp33_ASAP7_75t_L     g15478(.A(new_n15733), .B(new_n15734), .Y(new_n15735));
  MAJIxp5_ASAP7_75t_L       g15479(.A(new_n15546), .B(new_n15547), .C(new_n15550), .Y(new_n15736));
  AOI22xp33_ASAP7_75t_L     g15480(.A1(new_n2706), .A2(\b[49] ), .B1(\b[50] ), .B2(new_n2702), .Y(new_n15737));
  OAI221xp5_ASAP7_75t_L     g15481(.A1(new_n2932), .A2(new_n7333), .B1(new_n2707), .B2(new_n8234), .C(new_n15737), .Y(new_n15738));
  XNOR2x2_ASAP7_75t_L       g15482(.A(new_n2697), .B(new_n15738), .Y(new_n15739));
  XNOR2x2_ASAP7_75t_L       g15483(.A(new_n15739), .B(new_n15736), .Y(new_n15740));
  AND2x2_ASAP7_75t_L        g15484(.A(new_n15735), .B(new_n15740), .Y(new_n15741));
  NOR2xp33_ASAP7_75t_L      g15485(.A(new_n15735), .B(new_n15740), .Y(new_n15742));
  NOR2xp33_ASAP7_75t_L      g15486(.A(new_n15742), .B(new_n15741), .Y(new_n15743));
  XOR2x2_ASAP7_75t_L        g15487(.A(new_n15743), .B(new_n15619), .Y(new_n15744));
  AND3x1_ASAP7_75t_L        g15488(.A(new_n15607), .B(new_n15744), .C(new_n15605), .Y(new_n15745));
  AOI21xp33_ASAP7_75t_L     g15489(.A1(new_n15607), .A2(new_n15605), .B(new_n15744), .Y(new_n15746));
  NOR2xp33_ASAP7_75t_L      g15490(.A(new_n15746), .B(new_n15745), .Y(new_n15747));
  NAND2xp33_ASAP7_75t_L     g15491(.A(new_n15747), .B(new_n15600), .Y(new_n15748));
  OAI22xp33_ASAP7_75t_L     g15492(.A1(new_n15598), .A2(new_n15599), .B1(new_n15746), .B2(new_n15745), .Y(new_n15749));
  OAI211xp5_ASAP7_75t_L     g15493(.A1(new_n15592), .A2(new_n15590), .B(new_n15748), .C(new_n15749), .Y(new_n15750));
  NOR2xp33_ASAP7_75t_L      g15494(.A(new_n15590), .B(new_n15592), .Y(new_n15751));
  NAND2xp33_ASAP7_75t_L     g15495(.A(new_n15749), .B(new_n15748), .Y(new_n15752));
  NAND2xp33_ASAP7_75t_L     g15496(.A(new_n15751), .B(new_n15752), .Y(new_n15753));
  NAND2xp33_ASAP7_75t_L     g15497(.A(new_n15750), .B(new_n15753), .Y(new_n15754));
  INVx1_ASAP7_75t_L         g15498(.A(new_n15413), .Y(new_n15755));
  MAJIxp5_ASAP7_75t_L       g15499(.A(new_n15566), .B(new_n15412), .C(new_n15755), .Y(new_n15756));
  O2A1O1Ixp33_ASAP7_75t_L   g15500(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n911), .Y(new_n15757));
  O2A1O1Ixp33_ASAP7_75t_L   g15501(.A1(new_n908), .A2(new_n15757), .B(\b[63] ), .C(new_n813), .Y(new_n15758));
  A2O1A1O1Ixp25_ASAP7_75t_L g15502(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n823), .D(new_n908), .Y(new_n15759));
  NOR3xp33_ASAP7_75t_L      g15503(.A(new_n15759), .B(new_n12599), .C(\a[14] ), .Y(new_n15760));
  NOR2xp33_ASAP7_75t_L      g15504(.A(new_n15758), .B(new_n15760), .Y(new_n15761));
  XOR2x2_ASAP7_75t_L        g15505(.A(new_n15761), .B(new_n15756), .Y(new_n15762));
  NOR2xp33_ASAP7_75t_L      g15506(.A(new_n15754), .B(new_n15762), .Y(new_n15763));
  XNOR2x2_ASAP7_75t_L       g15507(.A(new_n15761), .B(new_n15756), .Y(new_n15764));
  AOI21xp33_ASAP7_75t_L     g15508(.A1(new_n15753), .A2(new_n15750), .B(new_n15764), .Y(new_n15765));
  NOR3xp33_ASAP7_75t_L      g15509(.A(new_n15765), .B(new_n15763), .C(new_n15582), .Y(new_n15766));
  O2A1O1Ixp33_ASAP7_75t_L   g15510(.A1(new_n15234), .A2(new_n15236), .B(new_n15365), .C(new_n15398), .Y(new_n15767));
  MAJIxp5_ASAP7_75t_L       g15511(.A(new_n15567), .B(new_n15767), .C(new_n15404), .Y(new_n15768));
  NAND3xp33_ASAP7_75t_L     g15512(.A(new_n15764), .B(new_n15753), .C(new_n15750), .Y(new_n15769));
  NAND2xp33_ASAP7_75t_L     g15513(.A(new_n15754), .B(new_n15762), .Y(new_n15770));
  AOI21xp33_ASAP7_75t_L     g15514(.A1(new_n15769), .A2(new_n15770), .B(new_n15768), .Y(new_n15771));
  NOR2xp33_ASAP7_75t_L      g15515(.A(new_n15771), .B(new_n15766), .Y(new_n15772));
  A2O1A1Ixp33_ASAP7_75t_L   g15516(.A1(new_n15578), .A2(new_n15574), .B(new_n15572), .C(new_n15772), .Y(new_n15773));
  INVx1_ASAP7_75t_L         g15517(.A(new_n15773), .Y(new_n15774));
  INVx1_ASAP7_75t_L         g15518(.A(new_n15572), .Y(new_n15775));
  A2O1A1Ixp33_ASAP7_75t_L   g15519(.A1(new_n15393), .A2(new_n15387), .B(new_n15575), .C(new_n15775), .Y(new_n15776));
  NOR2xp33_ASAP7_75t_L      g15520(.A(new_n15772), .B(new_n15776), .Y(new_n15777));
  NOR2xp33_ASAP7_75t_L      g15521(.A(new_n15774), .B(new_n15777), .Y(\f[77] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15522(.A1(new_n15758), .A2(new_n15760), .B(new_n15756), .C(new_n15763), .Y(new_n15779));
  NAND2xp33_ASAP7_75t_L     g15523(.A(new_n15589), .B(new_n15591), .Y(new_n15780));
  NAND2xp33_ASAP7_75t_L     g15524(.A(new_n15780), .B(new_n15750), .Y(new_n15781));
  NAND2xp33_ASAP7_75t_L     g15525(.A(\b[63] ), .B(new_n1113), .Y(new_n15782));
  A2O1A1Ixp33_ASAP7_75t_L   g15526(.A1(new_n12607), .A2(new_n12603), .B(new_n1197), .C(new_n15782), .Y(new_n15783));
  AOI221xp5_ASAP7_75t_L     g15527(.A1(\b[61] ), .A2(new_n1194), .B1(\b[62] ), .B2(new_n1103), .C(new_n15783), .Y(new_n15784));
  XNOR2x2_ASAP7_75t_L       g15528(.A(new_n1107), .B(new_n15784), .Y(new_n15785));
  NAND2xp33_ASAP7_75t_L     g15529(.A(new_n15785), .B(new_n15781), .Y(new_n15786));
  INVx1_ASAP7_75t_L         g15530(.A(new_n15785), .Y(new_n15787));
  NAND3xp33_ASAP7_75t_L     g15531(.A(new_n15750), .B(new_n15780), .C(new_n15787), .Y(new_n15788));
  AND2x2_ASAP7_75t_L        g15532(.A(new_n15788), .B(new_n15786), .Y(new_n15789));
  AOI22xp33_ASAP7_75t_L     g15533(.A1(new_n1406), .A2(\b[60] ), .B1(new_n1404), .B2(new_n11234), .Y(new_n15790));
  OAI221xp5_ASAP7_75t_L     g15534(.A1(new_n1398), .A2(new_n10881), .B1(new_n10848), .B2(new_n1549), .C(new_n15790), .Y(new_n15791));
  XNOR2x2_ASAP7_75t_L       g15535(.A(\a[20] ), .B(new_n15791), .Y(new_n15792));
  INVx1_ASAP7_75t_L         g15536(.A(new_n15792), .Y(new_n15793));
  AOI211xp5_ASAP7_75t_L     g15537(.A1(new_n15600), .A2(new_n15747), .B(new_n15793), .C(new_n15599), .Y(new_n15794));
  O2A1O1Ixp33_ASAP7_75t_L   g15538(.A1(new_n15595), .A2(new_n15597), .B(new_n15748), .C(new_n15792), .Y(new_n15795));
  NOR2xp33_ASAP7_75t_L      g15539(.A(new_n15794), .B(new_n15795), .Y(new_n15796));
  AOI22xp33_ASAP7_75t_L     g15540(.A1(new_n1766), .A2(\b[57] ), .B1(new_n1764), .B2(new_n10495), .Y(new_n15797));
  OAI221xp5_ASAP7_75t_L     g15541(.A1(new_n1758), .A2(new_n10178), .B1(new_n9534), .B2(new_n1911), .C(new_n15797), .Y(new_n15798));
  XNOR2x2_ASAP7_75t_L       g15542(.A(\a[23] ), .B(new_n15798), .Y(new_n15799));
  A2O1A1Ixp33_ASAP7_75t_L   g15543(.A1(new_n15605), .A2(new_n15744), .B(new_n15606), .C(new_n15799), .Y(new_n15800));
  NOR2xp33_ASAP7_75t_L      g15544(.A(new_n15606), .B(new_n15745), .Y(new_n15801));
  INVx1_ASAP7_75t_L         g15545(.A(new_n15799), .Y(new_n15802));
  NAND2xp33_ASAP7_75t_L     g15546(.A(new_n15802), .B(new_n15801), .Y(new_n15803));
  AOI22xp33_ASAP7_75t_L     g15547(.A1(new_n2228), .A2(\b[54] ), .B1(new_n2226), .B2(new_n9208), .Y(new_n15804));
  OAI221xp5_ASAP7_75t_L     g15548(.A1(new_n2220), .A2(new_n8882), .B1(new_n8569), .B2(new_n2387), .C(new_n15804), .Y(new_n15805));
  XNOR2x2_ASAP7_75t_L       g15549(.A(\a[26] ), .B(new_n15805), .Y(new_n15806));
  INVx1_ASAP7_75t_L         g15550(.A(new_n15806), .Y(new_n15807));
  A2O1A1Ixp33_ASAP7_75t_L   g15551(.A1(new_n15612), .A2(new_n15611), .B(new_n15614), .C(new_n15743), .Y(new_n15808));
  O2A1O1Ixp33_ASAP7_75t_L   g15552(.A1(new_n15615), .A2(new_n15613), .B(new_n15808), .C(new_n15807), .Y(new_n15809));
  AOI21xp33_ASAP7_75t_L     g15553(.A1(new_n15743), .A2(new_n15618), .B(new_n15616), .Y(new_n15810));
  NAND2xp33_ASAP7_75t_L     g15554(.A(new_n15807), .B(new_n15810), .Y(new_n15811));
  INVx1_ASAP7_75t_L         g15555(.A(new_n15811), .Y(new_n15812));
  NOR2xp33_ASAP7_75t_L      g15556(.A(new_n15809), .B(new_n15812), .Y(new_n15813));
  AOI22xp33_ASAP7_75t_L     g15557(.A1(new_n2702), .A2(\b[51] ), .B1(new_n2700), .B2(new_n8257), .Y(new_n15814));
  OAI221xp5_ASAP7_75t_L     g15558(.A1(new_n2694), .A2(new_n8228), .B1(new_n7907), .B2(new_n2932), .C(new_n15814), .Y(new_n15815));
  XNOR2x2_ASAP7_75t_L       g15559(.A(\a[29] ), .B(new_n15815), .Y(new_n15816));
  INVx1_ASAP7_75t_L         g15560(.A(new_n15816), .Y(new_n15817));
  NOR2xp33_ASAP7_75t_L      g15561(.A(new_n15739), .B(new_n15736), .Y(new_n15818));
  NOR2xp33_ASAP7_75t_L      g15562(.A(new_n15818), .B(new_n15742), .Y(new_n15819));
  XNOR2x2_ASAP7_75t_L       g15563(.A(new_n15817), .B(new_n15819), .Y(new_n15820));
  NAND2xp33_ASAP7_75t_L     g15564(.A(new_n15726), .B(new_n15728), .Y(new_n15821));
  AOI22xp33_ASAP7_75t_L     g15565(.A1(new_n4544), .A2(\b[42] ), .B1(new_n4542), .B2(new_n5688), .Y(new_n15822));
  OAI221xp5_ASAP7_75t_L     g15566(.A1(new_n4536), .A2(new_n5666), .B1(new_n5186), .B2(new_n4781), .C(new_n15822), .Y(new_n15823));
  XNOR2x2_ASAP7_75t_L       g15567(.A(\a[38] ), .B(new_n15823), .Y(new_n15824));
  INVx1_ASAP7_75t_L         g15568(.A(new_n15824), .Y(new_n15825));
  AOI21xp33_ASAP7_75t_L     g15569(.A1(new_n15723), .A2(new_n15724), .B(new_n15718), .Y(new_n15826));
  AOI22xp33_ASAP7_75t_L     g15570(.A1(new_n6002), .A2(\b[36] ), .B1(new_n5999), .B2(new_n4473), .Y(new_n15827));
  OAI221xp5_ASAP7_75t_L     g15571(.A1(new_n6544), .A2(new_n4053), .B1(new_n3827), .B2(new_n6309), .C(new_n15827), .Y(new_n15828));
  XNOR2x2_ASAP7_75t_L       g15572(.A(new_n5996), .B(new_n15828), .Y(new_n15829));
  AOI22xp33_ASAP7_75t_L     g15573(.A1(new_n8645), .A2(\b[27] ), .B1(new_n8642), .B2(new_n2657), .Y(new_n15830));
  OAI221xp5_ASAP7_75t_L     g15574(.A1(new_n9322), .A2(new_n2477), .B1(new_n2180), .B2(new_n8965), .C(new_n15830), .Y(new_n15831));
  XNOR2x2_ASAP7_75t_L       g15575(.A(\a[53] ), .B(new_n15831), .Y(new_n15832));
  INVx1_ASAP7_75t_L         g15576(.A(new_n15832), .Y(new_n15833));
  NAND2xp33_ASAP7_75t_L     g15577(.A(new_n15675), .B(new_n15672), .Y(new_n15834));
  A2O1A1Ixp33_ASAP7_75t_L   g15578(.A1(new_n15667), .A2(new_n15666), .B(new_n15670), .C(new_n15834), .Y(new_n15835));
  AOI22xp33_ASAP7_75t_L     g15579(.A1(new_n11656), .A2(\b[18] ), .B1(new_n11654), .B2(new_n1363), .Y(new_n15836));
  OAI221xp5_ASAP7_75t_L     g15580(.A1(new_n12364), .A2(new_n1244), .B1(new_n1051), .B2(new_n13003), .C(new_n15836), .Y(new_n15837));
  XNOR2x2_ASAP7_75t_L       g15581(.A(new_n11651), .B(new_n15837), .Y(new_n15838));
  NOR2xp33_ASAP7_75t_L      g15582(.A(new_n871), .B(new_n12671), .Y(new_n15839));
  O2A1O1Ixp33_ASAP7_75t_L   g15583(.A1(new_n12353), .A2(new_n12355), .B(\b[15] ), .C(new_n15839), .Y(new_n15840));
  INVx1_ASAP7_75t_L         g15584(.A(new_n15840), .Y(new_n15841));
  NOR2xp33_ASAP7_75t_L      g15585(.A(\a[14] ), .B(new_n15841), .Y(new_n15842));
  INVx1_ASAP7_75t_L         g15586(.A(new_n15842), .Y(new_n15843));
  A2O1A1Ixp33_ASAP7_75t_L   g15587(.A1(new_n12669), .A2(\b[15] ), .B(new_n15839), .C(\a[14] ), .Y(new_n15844));
  NAND2xp33_ASAP7_75t_L     g15588(.A(new_n15844), .B(new_n15843), .Y(new_n15845));
  A2O1A1Ixp33_ASAP7_75t_L   g15589(.A1(new_n12669), .A2(\b[13] ), .B(new_n15460), .C(new_n15845), .Y(new_n15846));
  INVx1_ASAP7_75t_L         g15590(.A(new_n15846), .Y(new_n15847));
  AND3x1_ASAP7_75t_L        g15591(.A(new_n15843), .B(new_n15844), .C(new_n15461), .Y(new_n15848));
  NOR2xp33_ASAP7_75t_L      g15592(.A(new_n15848), .B(new_n15847), .Y(new_n15849));
  XNOR2x2_ASAP7_75t_L       g15593(.A(new_n15849), .B(new_n15838), .Y(new_n15850));
  A2O1A1O1Ixp25_ASAP7_75t_L g15594(.A1(new_n12669), .A2(\b[14] ), .B(new_n15649), .C(new_n15461), .D(new_n15657), .Y(new_n15851));
  XNOR2x2_ASAP7_75t_L       g15595(.A(new_n15851), .B(new_n15850), .Y(new_n15852));
  AOI22xp33_ASAP7_75t_L     g15596(.A1(new_n10594), .A2(\b[21] ), .B1(new_n10591), .B2(new_n1715), .Y(new_n15853));
  OAI221xp5_ASAP7_75t_L     g15597(.A1(new_n11335), .A2(new_n1594), .B1(new_n1493), .B2(new_n11330), .C(new_n15853), .Y(new_n15854));
  XNOR2x2_ASAP7_75t_L       g15598(.A(\a[59] ), .B(new_n15854), .Y(new_n15855));
  XNOR2x2_ASAP7_75t_L       g15599(.A(new_n15855), .B(new_n15852), .Y(new_n15856));
  AOI21xp33_ASAP7_75t_L     g15600(.A1(new_n15665), .A2(new_n15660), .B(new_n15661), .Y(new_n15857));
  XNOR2x2_ASAP7_75t_L       g15601(.A(new_n15857), .B(new_n15856), .Y(new_n15858));
  AOI22xp33_ASAP7_75t_L     g15602(.A1(new_n9623), .A2(\b[24] ), .B1(new_n9620), .B2(new_n2027), .Y(new_n15859));
  OAI221xp5_ASAP7_75t_L     g15603(.A1(new_n10280), .A2(new_n1995), .B1(new_n1857), .B2(new_n12010), .C(new_n15859), .Y(new_n15860));
  XNOR2x2_ASAP7_75t_L       g15604(.A(new_n9610), .B(new_n15860), .Y(new_n15861));
  XNOR2x2_ASAP7_75t_L       g15605(.A(new_n15861), .B(new_n15858), .Y(new_n15862));
  XNOR2x2_ASAP7_75t_L       g15606(.A(new_n15835), .B(new_n15862), .Y(new_n15863));
  XNOR2x2_ASAP7_75t_L       g15607(.A(new_n15833), .B(new_n15863), .Y(new_n15864));
  OAI211xp5_ASAP7_75t_L     g15608(.A1(new_n15677), .A2(new_n15678), .B(new_n15864), .C(new_n15682), .Y(new_n15865));
  O2A1O1Ixp33_ASAP7_75t_L   g15609(.A1(new_n15677), .A2(new_n15678), .B(new_n15682), .C(new_n15864), .Y(new_n15866));
  INVx1_ASAP7_75t_L         g15610(.A(new_n15866), .Y(new_n15867));
  NAND2xp33_ASAP7_75t_L     g15611(.A(new_n15865), .B(new_n15867), .Y(new_n15868));
  AOI22xp33_ASAP7_75t_L     g15612(.A1(new_n7659), .A2(\b[30] ), .B1(new_n7656), .B2(new_n3219), .Y(new_n15869));
  OAI221xp5_ASAP7_75t_L     g15613(.A1(new_n8326), .A2(new_n2871), .B1(new_n2852), .B2(new_n7994), .C(new_n15869), .Y(new_n15870));
  XNOR2x2_ASAP7_75t_L       g15614(.A(\a[50] ), .B(new_n15870), .Y(new_n15871));
  XNOR2x2_ASAP7_75t_L       g15615(.A(new_n15871), .B(new_n15868), .Y(new_n15872));
  A2O1A1Ixp33_ASAP7_75t_L   g15616(.A1(new_n15686), .A2(new_n15685), .B(new_n15692), .C(new_n15872), .Y(new_n15873));
  INVx1_ASAP7_75t_L         g15617(.A(new_n15872), .Y(new_n15874));
  INVx1_ASAP7_75t_L         g15618(.A(new_n15682), .Y(new_n15875));
  O2A1O1Ixp33_ASAP7_75t_L   g15619(.A1(new_n15875), .A2(new_n15683), .B(new_n15686), .C(new_n15692), .Y(new_n15876));
  NAND2xp33_ASAP7_75t_L     g15620(.A(new_n15874), .B(new_n15876), .Y(new_n15877));
  NAND2xp33_ASAP7_75t_L     g15621(.A(new_n15873), .B(new_n15877), .Y(new_n15878));
  AOI22xp33_ASAP7_75t_L     g15622(.A1(new_n6822), .A2(\b[33] ), .B1(new_n6819), .B2(new_n3813), .Y(new_n15879));
  OAI221xp5_ASAP7_75t_L     g15623(.A1(new_n7392), .A2(new_n3443), .B1(new_n3419), .B2(new_n7115), .C(new_n15879), .Y(new_n15880));
  XNOR2x2_ASAP7_75t_L       g15624(.A(\a[47] ), .B(new_n15880), .Y(new_n15881));
  XNOR2x2_ASAP7_75t_L       g15625(.A(new_n15881), .B(new_n15878), .Y(new_n15882));
  NOR3xp33_ASAP7_75t_L      g15626(.A(new_n15882), .B(new_n15698), .C(new_n15697), .Y(new_n15883));
  OA21x2_ASAP7_75t_L        g15627(.A1(new_n15697), .A2(new_n15698), .B(new_n15882), .Y(new_n15884));
  NOR2xp33_ASAP7_75t_L      g15628(.A(new_n15883), .B(new_n15884), .Y(new_n15885));
  NAND2xp33_ASAP7_75t_L     g15629(.A(new_n15829), .B(new_n15885), .Y(new_n15886));
  OR2x4_ASAP7_75t_L         g15630(.A(new_n15829), .B(new_n15885), .Y(new_n15887));
  NAND2xp33_ASAP7_75t_L     g15631(.A(new_n15886), .B(new_n15887), .Y(new_n15888));
  A2O1A1Ixp33_ASAP7_75t_L   g15632(.A1(new_n15706), .A2(new_n15709), .B(new_n15702), .C(new_n15888), .Y(new_n15889));
  INVx1_ASAP7_75t_L         g15633(.A(new_n15702), .Y(new_n15890));
  NAND4xp25_ASAP7_75t_L     g15634(.A(new_n15887), .B(new_n15890), .C(new_n15710), .D(new_n15886), .Y(new_n15891));
  NAND2xp33_ASAP7_75t_L     g15635(.A(new_n15891), .B(new_n15889), .Y(new_n15892));
  AOI22xp33_ASAP7_75t_L     g15636(.A1(new_n5249), .A2(\b[39] ), .B1(new_n5247), .B2(new_n5174), .Y(new_n15893));
  OAI221xp5_ASAP7_75t_L     g15637(.A1(new_n5241), .A2(new_n4915), .B1(new_n4701), .B2(new_n5521), .C(new_n15893), .Y(new_n15894));
  XNOR2x2_ASAP7_75t_L       g15638(.A(\a[41] ), .B(new_n15894), .Y(new_n15895));
  XOR2x2_ASAP7_75t_L        g15639(.A(new_n15895), .B(new_n15892), .Y(new_n15896));
  XNOR2x2_ASAP7_75t_L       g15640(.A(new_n15826), .B(new_n15896), .Y(new_n15897));
  AND2x2_ASAP7_75t_L        g15641(.A(new_n15825), .B(new_n15897), .Y(new_n15898));
  NOR2xp33_ASAP7_75t_L      g15642(.A(new_n15825), .B(new_n15897), .Y(new_n15899));
  NOR2xp33_ASAP7_75t_L      g15643(.A(new_n15899), .B(new_n15898), .Y(new_n15900));
  XNOR2x2_ASAP7_75t_L       g15644(.A(new_n15821), .B(new_n15900), .Y(new_n15901));
  AOI22xp33_ASAP7_75t_L     g15645(.A1(new_n3884), .A2(\b[45] ), .B1(new_n3881), .B2(new_n6764), .Y(new_n15902));
  OAI221xp5_ASAP7_75t_L     g15646(.A1(new_n4312), .A2(new_n6220), .B1(new_n6195), .B2(new_n4986), .C(new_n15902), .Y(new_n15903));
  XNOR2x2_ASAP7_75t_L       g15647(.A(\a[35] ), .B(new_n15903), .Y(new_n15904));
  XNOR2x2_ASAP7_75t_L       g15648(.A(new_n15904), .B(new_n15901), .Y(new_n15905));
  MAJx2_ASAP7_75t_L         g15649(.A(new_n15730), .B(new_n15630), .C(new_n15632), .Y(new_n15906));
  XNOR2x2_ASAP7_75t_L       g15650(.A(new_n15906), .B(new_n15905), .Y(new_n15907));
  AOI22xp33_ASAP7_75t_L     g15651(.A1(new_n3256), .A2(\b[48] ), .B1(new_n3254), .B2(new_n7341), .Y(new_n15908));
  OAI221xp5_ASAP7_75t_L     g15652(.A1(new_n3248), .A2(new_n7316), .B1(new_n7033), .B2(new_n3492), .C(new_n15908), .Y(new_n15909));
  XNOR2x2_ASAP7_75t_L       g15653(.A(\a[32] ), .B(new_n15909), .Y(new_n15910));
  NAND2xp33_ASAP7_75t_L     g15654(.A(new_n15627), .B(new_n15733), .Y(new_n15911));
  XNOR2x2_ASAP7_75t_L       g15655(.A(new_n15910), .B(new_n15911), .Y(new_n15912));
  NOR2xp33_ASAP7_75t_L      g15656(.A(new_n15907), .B(new_n15912), .Y(new_n15913));
  AND2x2_ASAP7_75t_L        g15657(.A(new_n15907), .B(new_n15912), .Y(new_n15914));
  NOR3xp33_ASAP7_75t_L      g15658(.A(new_n15820), .B(new_n15913), .C(new_n15914), .Y(new_n15915));
  OA21x2_ASAP7_75t_L        g15659(.A1(new_n15913), .A2(new_n15914), .B(new_n15820), .Y(new_n15916));
  NOR2xp33_ASAP7_75t_L      g15660(.A(new_n15915), .B(new_n15916), .Y(new_n15917));
  NAND2xp33_ASAP7_75t_L     g15661(.A(new_n15813), .B(new_n15917), .Y(new_n15918));
  OAI22xp33_ASAP7_75t_L     g15662(.A1(new_n15916), .A2(new_n15915), .B1(new_n15812), .B2(new_n15809), .Y(new_n15919));
  AOI22xp33_ASAP7_75t_L     g15663(.A1(new_n15918), .A2(new_n15919), .B1(new_n15800), .B2(new_n15803), .Y(new_n15920));
  AND4x1_ASAP7_75t_L        g15664(.A(new_n15803), .B(new_n15800), .C(new_n15919), .D(new_n15918), .Y(new_n15921));
  NOR2xp33_ASAP7_75t_L      g15665(.A(new_n15920), .B(new_n15921), .Y(new_n15922));
  XOR2x2_ASAP7_75t_L        g15666(.A(new_n15922), .B(new_n15796), .Y(new_n15923));
  NOR2xp33_ASAP7_75t_L      g15667(.A(new_n15923), .B(new_n15789), .Y(new_n15924));
  AND3x1_ASAP7_75t_L        g15668(.A(new_n15923), .B(new_n15788), .C(new_n15786), .Y(new_n15925));
  OAI21xp33_ASAP7_75t_L     g15669(.A1(new_n15924), .A2(new_n15925), .B(new_n15779), .Y(new_n15926));
  OA21x2_ASAP7_75t_L        g15670(.A1(new_n15758), .A2(new_n15760), .B(new_n15756), .Y(new_n15927));
  AO21x2_ASAP7_75t_L        g15671(.A1(new_n15788), .A2(new_n15786), .B(new_n15923), .Y(new_n15928));
  NAND2xp33_ASAP7_75t_L     g15672(.A(new_n15923), .B(new_n15789), .Y(new_n15929));
  OAI211xp5_ASAP7_75t_L     g15673(.A1(new_n15763), .A2(new_n15927), .B(new_n15928), .C(new_n15929), .Y(new_n15930));
  NAND2xp33_ASAP7_75t_L     g15674(.A(new_n15926), .B(new_n15930), .Y(new_n15931));
  INVx1_ASAP7_75t_L         g15675(.A(new_n15931), .Y(new_n15932));
  A2O1A1Ixp33_ASAP7_75t_L   g15676(.A1(new_n15776), .A2(new_n15772), .B(new_n15766), .C(new_n15932), .Y(new_n15933));
  A2O1A1O1Ixp25_ASAP7_75t_L g15677(.A1(new_n15574), .A2(new_n15578), .B(new_n15572), .C(new_n15772), .D(new_n15766), .Y(new_n15934));
  NAND2xp33_ASAP7_75t_L     g15678(.A(new_n15931), .B(new_n15934), .Y(new_n15935));
  AND2x2_ASAP7_75t_L        g15679(.A(new_n15935), .B(new_n15933), .Y(\f[78] ));
  INVx1_ASAP7_75t_L         g15680(.A(new_n15795), .Y(new_n15937));
  AOI22xp33_ASAP7_75t_L     g15681(.A1(new_n1103), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1194), .Y(new_n15938));
  A2O1A1Ixp33_ASAP7_75t_L   g15682(.A1(new_n13506), .A2(new_n13507), .B(new_n1197), .C(new_n15938), .Y(new_n15939));
  NOR2xp33_ASAP7_75t_L      g15683(.A(new_n1107), .B(new_n15939), .Y(new_n15940));
  A2O1A1O1Ixp25_ASAP7_75t_L g15684(.A1(new_n13507), .A2(new_n13506), .B(new_n1197), .C(new_n15938), .D(\a[17] ), .Y(new_n15941));
  NOR2xp33_ASAP7_75t_L      g15685(.A(new_n15941), .B(new_n15940), .Y(new_n15942));
  O2A1O1Ixp33_ASAP7_75t_L   g15686(.A1(new_n15922), .A2(new_n15794), .B(new_n15937), .C(new_n15942), .Y(new_n15943));
  INVx1_ASAP7_75t_L         g15687(.A(new_n15943), .Y(new_n15944));
  O2A1O1Ixp33_ASAP7_75t_L   g15688(.A1(new_n15920), .A2(new_n15921), .B(new_n15796), .C(new_n15795), .Y(new_n15945));
  NAND2xp33_ASAP7_75t_L     g15689(.A(new_n15942), .B(new_n15945), .Y(new_n15946));
  AOI22xp33_ASAP7_75t_L     g15690(.A1(new_n1406), .A2(\b[61] ), .B1(new_n1404), .B2(new_n11919), .Y(new_n15947));
  OAI221xp5_ASAP7_75t_L     g15691(.A1(new_n1398), .A2(new_n11226), .B1(new_n10881), .B2(new_n1549), .C(new_n15947), .Y(new_n15948));
  XNOR2x2_ASAP7_75t_L       g15692(.A(\a[20] ), .B(new_n15948), .Y(new_n15949));
  INVx1_ASAP7_75t_L         g15693(.A(new_n15949), .Y(new_n15950));
  NAND2xp33_ASAP7_75t_L     g15694(.A(new_n15919), .B(new_n15918), .Y(new_n15951));
  A2O1A1Ixp33_ASAP7_75t_L   g15695(.A1(new_n15605), .A2(new_n15744), .B(new_n15606), .C(new_n15802), .Y(new_n15952));
  A2O1A1Ixp33_ASAP7_75t_L   g15696(.A1(new_n15803), .A2(new_n15800), .B(new_n15951), .C(new_n15952), .Y(new_n15953));
  NOR2xp33_ASAP7_75t_L      g15697(.A(new_n15950), .B(new_n15953), .Y(new_n15954));
  A2O1A1O1Ixp25_ASAP7_75t_L g15698(.A1(new_n15800), .A2(new_n15803), .B(new_n15951), .C(new_n15952), .D(new_n15949), .Y(new_n15955));
  NOR2xp33_ASAP7_75t_L      g15699(.A(new_n15955), .B(new_n15954), .Y(new_n15956));
  AOI22xp33_ASAP7_75t_L     g15700(.A1(new_n1770), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n1766), .Y(new_n15957));
  OAI221xp5_ASAP7_75t_L     g15701(.A1(new_n1911), .A2(new_n10178), .B1(new_n1771), .B2(new_n10856), .C(new_n15957), .Y(new_n15958));
  XNOR2x2_ASAP7_75t_L       g15702(.A(\a[23] ), .B(new_n15958), .Y(new_n15959));
  INVx1_ASAP7_75t_L         g15703(.A(new_n15959), .Y(new_n15960));
  A2O1A1Ixp33_ASAP7_75t_L   g15704(.A1(new_n15917), .A2(new_n15813), .B(new_n15812), .C(new_n15960), .Y(new_n15961));
  NAND3xp33_ASAP7_75t_L     g15705(.A(new_n15918), .B(new_n15811), .C(new_n15959), .Y(new_n15962));
  NAND2xp33_ASAP7_75t_L     g15706(.A(new_n15961), .B(new_n15962), .Y(new_n15963));
  INVx1_ASAP7_75t_L         g15707(.A(new_n15963), .Y(new_n15964));
  AOI22xp33_ASAP7_75t_L     g15708(.A1(new_n2228), .A2(\b[55] ), .B1(new_n2226), .B2(new_n9542), .Y(new_n15965));
  OAI221xp5_ASAP7_75t_L     g15709(.A1(new_n2220), .A2(new_n9199), .B1(new_n8882), .B2(new_n2387), .C(new_n15965), .Y(new_n15966));
  XNOR2x2_ASAP7_75t_L       g15710(.A(\a[26] ), .B(new_n15966), .Y(new_n15967));
  AOI21xp33_ASAP7_75t_L     g15711(.A1(new_n15819), .A2(new_n15817), .B(new_n15915), .Y(new_n15968));
  XNOR2x2_ASAP7_75t_L       g15712(.A(new_n15967), .B(new_n15968), .Y(new_n15969));
  AOI22xp33_ASAP7_75t_L     g15713(.A1(new_n2702), .A2(\b[52] ), .B1(new_n2700), .B2(new_n8577), .Y(new_n15970));
  OAI221xp5_ASAP7_75t_L     g15714(.A1(new_n2694), .A2(new_n8249), .B1(new_n8228), .B2(new_n2932), .C(new_n15970), .Y(new_n15971));
  XNOR2x2_ASAP7_75t_L       g15715(.A(\a[29] ), .B(new_n15971), .Y(new_n15972));
  INVx1_ASAP7_75t_L         g15716(.A(new_n15972), .Y(new_n15973));
  MAJIxp5_ASAP7_75t_L       g15717(.A(new_n15907), .B(new_n15910), .C(new_n15911), .Y(new_n15974));
  XNOR2x2_ASAP7_75t_L       g15718(.A(new_n15973), .B(new_n15974), .Y(new_n15975));
  AOI22xp33_ASAP7_75t_L     g15719(.A1(new_n3256), .A2(\b[49] ), .B1(new_n3254), .B2(new_n7914), .Y(new_n15976));
  OAI221xp5_ASAP7_75t_L     g15720(.A1(new_n3248), .A2(new_n7333), .B1(new_n7316), .B2(new_n3492), .C(new_n15976), .Y(new_n15977));
  XNOR2x2_ASAP7_75t_L       g15721(.A(\a[32] ), .B(new_n15977), .Y(new_n15978));
  MAJIxp5_ASAP7_75t_L       g15722(.A(new_n15901), .B(new_n15904), .C(new_n15906), .Y(new_n15979));
  XNOR2x2_ASAP7_75t_L       g15723(.A(new_n15978), .B(new_n15979), .Y(new_n15980));
  INVx1_ASAP7_75t_L         g15724(.A(new_n15980), .Y(new_n15981));
  NOR2xp33_ASAP7_75t_L      g15725(.A(new_n15895), .B(new_n15892), .Y(new_n15982));
  A2O1A1O1Ixp25_ASAP7_75t_L g15726(.A1(new_n15723), .A2(new_n15724), .B(new_n15718), .C(new_n15896), .D(new_n15982), .Y(new_n15983));
  AOI22xp33_ASAP7_75t_L     g15727(.A1(new_n5249), .A2(\b[40] ), .B1(new_n5247), .B2(new_n5194), .Y(new_n15984));
  OAI221xp5_ASAP7_75t_L     g15728(.A1(new_n5241), .A2(new_n5166), .B1(new_n4915), .B2(new_n5521), .C(new_n15984), .Y(new_n15985));
  XNOR2x2_ASAP7_75t_L       g15729(.A(\a[41] ), .B(new_n15985), .Y(new_n15986));
  INVx1_ASAP7_75t_L         g15730(.A(new_n15986), .Y(new_n15987));
  NAND2xp33_ASAP7_75t_L     g15731(.A(new_n15886), .B(new_n15891), .Y(new_n15988));
  AOI22xp33_ASAP7_75t_L     g15732(.A1(new_n6002), .A2(\b[37] ), .B1(new_n5999), .B2(new_n4709), .Y(new_n15989));
  OAI221xp5_ASAP7_75t_L     g15733(.A1(new_n6544), .A2(new_n4465), .B1(new_n4053), .B2(new_n6309), .C(new_n15989), .Y(new_n15990));
  XNOR2x2_ASAP7_75t_L       g15734(.A(\a[44] ), .B(new_n15990), .Y(new_n15991));
  INVx1_ASAP7_75t_L         g15735(.A(new_n15991), .Y(new_n15992));
  INVx1_ASAP7_75t_L         g15736(.A(new_n15878), .Y(new_n15993));
  INVx1_ASAP7_75t_L         g15737(.A(new_n15881), .Y(new_n15994));
  O2A1O1Ixp33_ASAP7_75t_L   g15738(.A1(new_n15653), .A2(new_n15656), .B(new_n15650), .C(new_n15850), .Y(new_n15995));
  NOR2xp33_ASAP7_75t_L      g15739(.A(new_n952), .B(new_n12671), .Y(new_n15996));
  A2O1A1O1Ixp25_ASAP7_75t_L g15740(.A1(new_n12669), .A2(\b[15] ), .B(new_n15839), .C(new_n813), .D(new_n15847), .Y(new_n15997));
  A2O1A1Ixp33_ASAP7_75t_L   g15741(.A1(new_n12669), .A2(\b[16] ), .B(new_n15996), .C(new_n15997), .Y(new_n15998));
  O2A1O1Ixp33_ASAP7_75t_L   g15742(.A1(new_n12353), .A2(new_n12355), .B(\b[16] ), .C(new_n15996), .Y(new_n15999));
  INVx1_ASAP7_75t_L         g15743(.A(new_n15999), .Y(new_n16000));
  A2O1A1Ixp33_ASAP7_75t_L   g15744(.A1(new_n12669), .A2(\b[15] ), .B(new_n15839), .C(new_n813), .Y(new_n16001));
  A2O1A1O1Ixp25_ASAP7_75t_L g15745(.A1(new_n15844), .A2(new_n15843), .B(new_n15461), .C(new_n16001), .D(new_n16000), .Y(new_n16002));
  INVx1_ASAP7_75t_L         g15746(.A(new_n16002), .Y(new_n16003));
  NAND2xp33_ASAP7_75t_L     g15747(.A(new_n16003), .B(new_n15998), .Y(new_n16004));
  AOI22xp33_ASAP7_75t_L     g15748(.A1(new_n11647), .A2(\b[18] ), .B1(\b[19] ), .B2(new_n11656), .Y(new_n16005));
  OAI221xp5_ASAP7_75t_L     g15749(.A1(new_n13003), .A2(new_n1244), .B1(new_n12022), .B2(new_n2793), .C(new_n16005), .Y(new_n16006));
  XNOR2x2_ASAP7_75t_L       g15750(.A(\a[62] ), .B(new_n16006), .Y(new_n16007));
  NOR2xp33_ASAP7_75t_L      g15751(.A(new_n16004), .B(new_n16007), .Y(new_n16008));
  AND2x2_ASAP7_75t_L        g15752(.A(new_n16004), .B(new_n16007), .Y(new_n16009));
  NOR2xp33_ASAP7_75t_L      g15753(.A(new_n16008), .B(new_n16009), .Y(new_n16010));
  A2O1A1Ixp33_ASAP7_75t_L   g15754(.A1(new_n15849), .A2(new_n15838), .B(new_n15995), .C(new_n16010), .Y(new_n16011));
  INVx1_ASAP7_75t_L         g15755(.A(new_n15657), .Y(new_n16012));
  NAND2xp33_ASAP7_75t_L     g15756(.A(new_n15849), .B(new_n15838), .Y(new_n16013));
  A2O1A1Ixp33_ASAP7_75t_L   g15757(.A1(new_n16012), .A2(new_n15650), .B(new_n15850), .C(new_n16013), .Y(new_n16014));
  NOR2xp33_ASAP7_75t_L      g15758(.A(new_n16010), .B(new_n16014), .Y(new_n16015));
  INVx1_ASAP7_75t_L         g15759(.A(new_n16015), .Y(new_n16016));
  AOI22xp33_ASAP7_75t_L     g15760(.A1(new_n10594), .A2(\b[22] ), .B1(new_n10591), .B2(new_n1864), .Y(new_n16017));
  OAI221xp5_ASAP7_75t_L     g15761(.A1(new_n11335), .A2(new_n1709), .B1(new_n1594), .B2(new_n11330), .C(new_n16017), .Y(new_n16018));
  XNOR2x2_ASAP7_75t_L       g15762(.A(\a[59] ), .B(new_n16018), .Y(new_n16019));
  AND3x1_ASAP7_75t_L        g15763(.A(new_n16016), .B(new_n16019), .C(new_n16011), .Y(new_n16020));
  INVx1_ASAP7_75t_L         g15764(.A(new_n16020), .Y(new_n16021));
  AO21x2_ASAP7_75t_L        g15765(.A1(new_n16011), .A2(new_n16016), .B(new_n16019), .Y(new_n16022));
  AND2x2_ASAP7_75t_L        g15766(.A(new_n16022), .B(new_n16021), .Y(new_n16023));
  INVx1_ASAP7_75t_L         g15767(.A(new_n15857), .Y(new_n16024));
  MAJx2_ASAP7_75t_L         g15768(.A(new_n16024), .B(new_n15855), .C(new_n15852), .Y(new_n16025));
  NAND2xp33_ASAP7_75t_L     g15769(.A(new_n16025), .B(new_n16023), .Y(new_n16026));
  AO21x2_ASAP7_75t_L        g15770(.A1(new_n16022), .A2(new_n16021), .B(new_n16025), .Y(new_n16027));
  AOI22xp33_ASAP7_75t_L     g15771(.A1(new_n9623), .A2(\b[25] ), .B1(new_n9620), .B2(new_n2188), .Y(new_n16028));
  OAI221xp5_ASAP7_75t_L     g15772(.A1(new_n10280), .A2(new_n2019), .B1(new_n1995), .B2(new_n12010), .C(new_n16028), .Y(new_n16029));
  XNOR2x2_ASAP7_75t_L       g15773(.A(\a[56] ), .B(new_n16029), .Y(new_n16030));
  NAND3xp33_ASAP7_75t_L     g15774(.A(new_n16026), .B(new_n16027), .C(new_n16030), .Y(new_n16031));
  AO21x2_ASAP7_75t_L        g15775(.A1(new_n16027), .A2(new_n16026), .B(new_n16030), .Y(new_n16032));
  NAND2xp33_ASAP7_75t_L     g15776(.A(new_n16031), .B(new_n16032), .Y(new_n16033));
  A2O1A1O1Ixp25_ASAP7_75t_L g15777(.A1(new_n15667), .A2(new_n15666), .B(new_n15670), .C(new_n15834), .D(new_n15862), .Y(new_n16034));
  AOI21xp33_ASAP7_75t_L     g15778(.A1(new_n15861), .A2(new_n15858), .B(new_n16034), .Y(new_n16035));
  XOR2x2_ASAP7_75t_L        g15779(.A(new_n16033), .B(new_n16035), .Y(new_n16036));
  NAND2xp33_ASAP7_75t_L     g15780(.A(\b[28] ), .B(new_n8645), .Y(new_n16037));
  OAI221xp5_ASAP7_75t_L     g15781(.A1(new_n2650), .A2(new_n9322), .B1(new_n8967), .B2(new_n5212), .C(new_n16037), .Y(new_n16038));
  AOI21xp33_ASAP7_75t_L     g15782(.A1(new_n8964), .A2(\b[26] ), .B(new_n16038), .Y(new_n16039));
  NAND2xp33_ASAP7_75t_L     g15783(.A(\a[53] ), .B(new_n16039), .Y(new_n16040));
  A2O1A1Ixp33_ASAP7_75t_L   g15784(.A1(\b[26] ), .A2(new_n8964), .B(new_n16038), .C(new_n8639), .Y(new_n16041));
  AND3x1_ASAP7_75t_L        g15785(.A(new_n16036), .B(new_n16041), .C(new_n16040), .Y(new_n16042));
  AOI21xp33_ASAP7_75t_L     g15786(.A1(new_n16041), .A2(new_n16040), .B(new_n16036), .Y(new_n16043));
  NOR2xp33_ASAP7_75t_L      g15787(.A(new_n16043), .B(new_n16042), .Y(new_n16044));
  A2O1A1Ixp33_ASAP7_75t_L   g15788(.A1(new_n15863), .A2(new_n15833), .B(new_n15866), .C(new_n16044), .Y(new_n16045));
  NAND2xp33_ASAP7_75t_L     g15789(.A(new_n15833), .B(new_n15863), .Y(new_n16046));
  OAI211xp5_ASAP7_75t_L     g15790(.A1(new_n16043), .A2(new_n16042), .B(new_n15867), .C(new_n16046), .Y(new_n16047));
  NAND2xp33_ASAP7_75t_L     g15791(.A(new_n16047), .B(new_n16045), .Y(new_n16048));
  NAND2xp33_ASAP7_75t_L     g15792(.A(\b[31] ), .B(new_n7659), .Y(new_n16049));
  OAI221xp5_ASAP7_75t_L     g15793(.A1(new_n3212), .A2(new_n8326), .B1(new_n7996), .B2(new_n4030), .C(new_n16049), .Y(new_n16050));
  AOI21xp33_ASAP7_75t_L     g15794(.A1(new_n7993), .A2(\b[29] ), .B(new_n16050), .Y(new_n16051));
  NAND2xp33_ASAP7_75t_L     g15795(.A(\a[50] ), .B(new_n16051), .Y(new_n16052));
  A2O1A1Ixp33_ASAP7_75t_L   g15796(.A1(\b[29] ), .A2(new_n7993), .B(new_n16050), .C(new_n7653), .Y(new_n16053));
  NAND2xp33_ASAP7_75t_L     g15797(.A(new_n16053), .B(new_n16052), .Y(new_n16054));
  XNOR2x2_ASAP7_75t_L       g15798(.A(new_n16054), .B(new_n16048), .Y(new_n16055));
  INVx1_ASAP7_75t_L         g15799(.A(new_n16055), .Y(new_n16056));
  NOR2xp33_ASAP7_75t_L      g15800(.A(new_n15871), .B(new_n15868), .Y(new_n16057));
  AOI21xp33_ASAP7_75t_L     g15801(.A1(new_n15876), .A2(new_n15874), .B(new_n16057), .Y(new_n16058));
  NAND2xp33_ASAP7_75t_L     g15802(.A(new_n16058), .B(new_n16056), .Y(new_n16059));
  A2O1A1Ixp33_ASAP7_75t_L   g15803(.A1(new_n15874), .A2(new_n15876), .B(new_n16057), .C(new_n16055), .Y(new_n16060));
  AND2x2_ASAP7_75t_L        g15804(.A(new_n16060), .B(new_n16059), .Y(new_n16061));
  AOI22xp33_ASAP7_75t_L     g15805(.A1(new_n6822), .A2(\b[34] ), .B1(new_n6819), .B2(new_n3833), .Y(new_n16062));
  OAI221xp5_ASAP7_75t_L     g15806(.A1(new_n7392), .A2(new_n3807), .B1(new_n3443), .B2(new_n7115), .C(new_n16062), .Y(new_n16063));
  XNOR2x2_ASAP7_75t_L       g15807(.A(\a[47] ), .B(new_n16063), .Y(new_n16064));
  XNOR2x2_ASAP7_75t_L       g15808(.A(new_n16064), .B(new_n16061), .Y(new_n16065));
  A2O1A1Ixp33_ASAP7_75t_L   g15809(.A1(new_n15994), .A2(new_n15993), .B(new_n15883), .C(new_n16065), .Y(new_n16066));
  INVx1_ASAP7_75t_L         g15810(.A(new_n16066), .Y(new_n16067));
  AOI211xp5_ASAP7_75t_L     g15811(.A1(new_n15993), .A2(new_n15994), .B(new_n15883), .C(new_n16065), .Y(new_n16068));
  NOR2xp33_ASAP7_75t_L      g15812(.A(new_n16067), .B(new_n16068), .Y(new_n16069));
  XNOR2x2_ASAP7_75t_L       g15813(.A(new_n15992), .B(new_n16069), .Y(new_n16070));
  XNOR2x2_ASAP7_75t_L       g15814(.A(new_n15988), .B(new_n16070), .Y(new_n16071));
  AND2x2_ASAP7_75t_L        g15815(.A(new_n15987), .B(new_n16071), .Y(new_n16072));
  NOR2xp33_ASAP7_75t_L      g15816(.A(new_n15987), .B(new_n16071), .Y(new_n16073));
  OR3x1_ASAP7_75t_L         g15817(.A(new_n16072), .B(new_n15983), .C(new_n16073), .Y(new_n16074));
  OAI21xp33_ASAP7_75t_L     g15818(.A1(new_n16073), .A2(new_n16072), .B(new_n15983), .Y(new_n16075));
  NAND2xp33_ASAP7_75t_L     g15819(.A(new_n16075), .B(new_n16074), .Y(new_n16076));
  NAND2xp33_ASAP7_75t_L     g15820(.A(\b[43] ), .B(new_n4544), .Y(new_n16077));
  OAI221xp5_ASAP7_75t_L     g15821(.A1(new_n5680), .A2(new_n4536), .B1(new_n4549), .B2(new_n9799), .C(new_n16077), .Y(new_n16078));
  AOI21xp33_ASAP7_75t_L     g15822(.A1(new_n4780), .A2(\b[41] ), .B(new_n16078), .Y(new_n16079));
  NAND2xp33_ASAP7_75t_L     g15823(.A(\a[38] ), .B(new_n16079), .Y(new_n16080));
  A2O1A1Ixp33_ASAP7_75t_L   g15824(.A1(\b[41] ), .A2(new_n4780), .B(new_n16078), .C(new_n4539), .Y(new_n16081));
  NAND2xp33_ASAP7_75t_L     g15825(.A(new_n16081), .B(new_n16080), .Y(new_n16082));
  XNOR2x2_ASAP7_75t_L       g15826(.A(new_n16082), .B(new_n16076), .Y(new_n16083));
  NAND2xp33_ASAP7_75t_L     g15827(.A(new_n15825), .B(new_n15897), .Y(new_n16084));
  A2O1A1Ixp33_ASAP7_75t_L   g15828(.A1(new_n15728), .A2(new_n15726), .B(new_n15899), .C(new_n16084), .Y(new_n16085));
  XNOR2x2_ASAP7_75t_L       g15829(.A(new_n16085), .B(new_n16083), .Y(new_n16086));
  AOI22xp33_ASAP7_75t_L     g15830(.A1(new_n3884), .A2(\b[46] ), .B1(new_n3881), .B2(new_n7041), .Y(new_n16087));
  OAI221xp5_ASAP7_75t_L     g15831(.A1(new_n4312), .A2(new_n6756), .B1(new_n6220), .B2(new_n4986), .C(new_n16087), .Y(new_n16088));
  XNOR2x2_ASAP7_75t_L       g15832(.A(\a[35] ), .B(new_n16088), .Y(new_n16089));
  INVx1_ASAP7_75t_L         g15833(.A(new_n16089), .Y(new_n16090));
  OR2x4_ASAP7_75t_L         g15834(.A(new_n16090), .B(new_n16086), .Y(new_n16091));
  NAND2xp33_ASAP7_75t_L     g15835(.A(new_n16090), .B(new_n16086), .Y(new_n16092));
  NAND2xp33_ASAP7_75t_L     g15836(.A(new_n16092), .B(new_n16091), .Y(new_n16093));
  XNOR2x2_ASAP7_75t_L       g15837(.A(new_n15981), .B(new_n16093), .Y(new_n16094));
  XOR2x2_ASAP7_75t_L        g15838(.A(new_n16094), .B(new_n15975), .Y(new_n16095));
  NOR2xp33_ASAP7_75t_L      g15839(.A(new_n16095), .B(new_n15969), .Y(new_n16096));
  AND2x2_ASAP7_75t_L        g15840(.A(new_n16095), .B(new_n15969), .Y(new_n16097));
  NOR2xp33_ASAP7_75t_L      g15841(.A(new_n16096), .B(new_n16097), .Y(new_n16098));
  NAND2xp33_ASAP7_75t_L     g15842(.A(new_n15964), .B(new_n16098), .Y(new_n16099));
  OAI21xp33_ASAP7_75t_L     g15843(.A1(new_n16096), .A2(new_n16097), .B(new_n15963), .Y(new_n16100));
  NAND2xp33_ASAP7_75t_L     g15844(.A(new_n16100), .B(new_n16099), .Y(new_n16101));
  INVx1_ASAP7_75t_L         g15845(.A(new_n16101), .Y(new_n16102));
  NAND2xp33_ASAP7_75t_L     g15846(.A(new_n16102), .B(new_n15956), .Y(new_n16103));
  OAI21xp33_ASAP7_75t_L     g15847(.A1(new_n15955), .A2(new_n15954), .B(new_n16101), .Y(new_n16104));
  NAND2xp33_ASAP7_75t_L     g15848(.A(new_n16104), .B(new_n16103), .Y(new_n16105));
  NAND3xp33_ASAP7_75t_L     g15849(.A(new_n15946), .B(new_n15944), .C(new_n16105), .Y(new_n16106));
  AOI21xp33_ASAP7_75t_L     g15850(.A1(new_n15946), .A2(new_n15944), .B(new_n16105), .Y(new_n16107));
  INVx1_ASAP7_75t_L         g15851(.A(new_n16107), .Y(new_n16108));
  O2A1O1Ixp33_ASAP7_75t_L   g15852(.A1(new_n15751), .A2(new_n15752), .B(new_n15780), .C(new_n15785), .Y(new_n16109));
  NOR2xp33_ASAP7_75t_L      g15853(.A(new_n16109), .B(new_n15924), .Y(new_n16110));
  AND3x1_ASAP7_75t_L        g15854(.A(new_n16110), .B(new_n16108), .C(new_n16106), .Y(new_n16111));
  AOI21xp33_ASAP7_75t_L     g15855(.A1(new_n16108), .A2(new_n16106), .B(new_n16110), .Y(new_n16112));
  NOR2xp33_ASAP7_75t_L      g15856(.A(new_n16112), .B(new_n16111), .Y(new_n16113));
  INVx1_ASAP7_75t_L         g15857(.A(new_n16113), .Y(new_n16114));
  O2A1O1Ixp33_ASAP7_75t_L   g15858(.A1(new_n15931), .A2(new_n15934), .B(new_n15930), .C(new_n16114), .Y(new_n16115));
  INVx1_ASAP7_75t_L         g15859(.A(new_n15766), .Y(new_n16116));
  A2O1A1Ixp33_ASAP7_75t_L   g15860(.A1(new_n15773), .A2(new_n16116), .B(new_n15931), .C(new_n15930), .Y(new_n16117));
  NOR2xp33_ASAP7_75t_L      g15861(.A(new_n16113), .B(new_n16117), .Y(new_n16118));
  NOR2xp33_ASAP7_75t_L      g15862(.A(new_n16118), .B(new_n16115), .Y(\f[79] ));
  AOI22xp33_ASAP7_75t_L     g15863(.A1(new_n1406), .A2(\b[62] ), .B1(new_n1404), .B2(new_n12280), .Y(new_n16120));
  OAI221xp5_ASAP7_75t_L     g15864(.A1(new_n1398), .A2(new_n11911), .B1(new_n11226), .B2(new_n1549), .C(new_n16120), .Y(new_n16121));
  XNOR2x2_ASAP7_75t_L       g15865(.A(\a[20] ), .B(new_n16121), .Y(new_n16122));
  INVx1_ASAP7_75t_L         g15866(.A(new_n16122), .Y(new_n16123));
  A2O1A1Ixp33_ASAP7_75t_L   g15867(.A1(new_n15918), .A2(new_n15811), .B(new_n15959), .C(new_n16099), .Y(new_n16124));
  NOR2xp33_ASAP7_75t_L      g15868(.A(new_n16123), .B(new_n16124), .Y(new_n16125));
  A2O1A1O1Ixp25_ASAP7_75t_L g15869(.A1(new_n15918), .A2(new_n15811), .B(new_n15959), .C(new_n16099), .D(new_n16122), .Y(new_n16126));
  NOR2xp33_ASAP7_75t_L      g15870(.A(new_n16126), .B(new_n16125), .Y(new_n16127));
  AOI22xp33_ASAP7_75t_L     g15871(.A1(new_n1766), .A2(\b[59] ), .B1(new_n1764), .B2(new_n10887), .Y(new_n16128));
  OAI221xp5_ASAP7_75t_L     g15872(.A1(new_n1758), .A2(new_n10848), .B1(new_n10488), .B2(new_n1911), .C(new_n16128), .Y(new_n16129));
  XNOR2x2_ASAP7_75t_L       g15873(.A(\a[23] ), .B(new_n16129), .Y(new_n16130));
  MAJIxp5_ASAP7_75t_L       g15874(.A(new_n16095), .B(new_n15967), .C(new_n15968), .Y(new_n16131));
  XNOR2x2_ASAP7_75t_L       g15875(.A(new_n16130), .B(new_n16131), .Y(new_n16132));
  AOI22xp33_ASAP7_75t_L     g15876(.A1(new_n2228), .A2(\b[56] ), .B1(new_n2226), .B2(new_n10185), .Y(new_n16133));
  OAI221xp5_ASAP7_75t_L     g15877(.A1(new_n2220), .A2(new_n9534), .B1(new_n9199), .B2(new_n2387), .C(new_n16133), .Y(new_n16134));
  XNOR2x2_ASAP7_75t_L       g15878(.A(\a[26] ), .B(new_n16134), .Y(new_n16135));
  MAJIxp5_ASAP7_75t_L       g15879(.A(new_n16094), .B(new_n15973), .C(new_n15974), .Y(new_n16136));
  AND2x2_ASAP7_75t_L        g15880(.A(new_n16135), .B(new_n16136), .Y(new_n16137));
  NOR2xp33_ASAP7_75t_L      g15881(.A(new_n16135), .B(new_n16136), .Y(new_n16138));
  NOR2xp33_ASAP7_75t_L      g15882(.A(new_n16138), .B(new_n16137), .Y(new_n16139));
  AOI22xp33_ASAP7_75t_L     g15883(.A1(new_n2702), .A2(\b[53] ), .B1(new_n2700), .B2(new_n8889), .Y(new_n16140));
  OAI221xp5_ASAP7_75t_L     g15884(.A1(new_n2694), .A2(new_n8569), .B1(new_n8249), .B2(new_n2932), .C(new_n16140), .Y(new_n16141));
  NOR2xp33_ASAP7_75t_L      g15885(.A(new_n2697), .B(new_n16141), .Y(new_n16142));
  AND2x2_ASAP7_75t_L        g15886(.A(new_n2697), .B(new_n16141), .Y(new_n16143));
  NOR2xp33_ASAP7_75t_L      g15887(.A(new_n16142), .B(new_n16143), .Y(new_n16144));
  INVx1_ASAP7_75t_L         g15888(.A(new_n15978), .Y(new_n16145));
  NAND2xp33_ASAP7_75t_L     g15889(.A(new_n16145), .B(new_n15979), .Y(new_n16146));
  A2O1A1Ixp33_ASAP7_75t_L   g15890(.A1(new_n16091), .A2(new_n16092), .B(new_n15981), .C(new_n16146), .Y(new_n16147));
  NOR2xp33_ASAP7_75t_L      g15891(.A(new_n16144), .B(new_n16147), .Y(new_n16148));
  INVx1_ASAP7_75t_L         g15892(.A(new_n16144), .Y(new_n16149));
  A2O1A1O1Ixp25_ASAP7_75t_L g15893(.A1(new_n16092), .A2(new_n16091), .B(new_n15981), .C(new_n16146), .D(new_n16149), .Y(new_n16150));
  NOR2xp33_ASAP7_75t_L      g15894(.A(new_n16150), .B(new_n16148), .Y(new_n16151));
  AOI22xp33_ASAP7_75t_L     g15895(.A1(new_n3256), .A2(\b[50] ), .B1(new_n3254), .B2(new_n8235), .Y(new_n16152));
  OAI221xp5_ASAP7_75t_L     g15896(.A1(new_n3248), .A2(new_n7907), .B1(new_n7333), .B2(new_n3492), .C(new_n16152), .Y(new_n16153));
  XNOR2x2_ASAP7_75t_L       g15897(.A(\a[32] ), .B(new_n16153), .Y(new_n16154));
  MAJx2_ASAP7_75t_L         g15898(.A(new_n16083), .B(new_n16085), .C(new_n16090), .Y(new_n16155));
  INVx1_ASAP7_75t_L         g15899(.A(new_n16155), .Y(new_n16156));
  AND2x2_ASAP7_75t_L        g15900(.A(new_n16154), .B(new_n16156), .Y(new_n16157));
  NOR2xp33_ASAP7_75t_L      g15901(.A(new_n16154), .B(new_n16156), .Y(new_n16158));
  NOR2xp33_ASAP7_75t_L      g15902(.A(new_n16158), .B(new_n16157), .Y(new_n16159));
  AOI22xp33_ASAP7_75t_L     g15903(.A1(new_n4544), .A2(\b[44] ), .B1(new_n4542), .B2(new_n7055), .Y(new_n16160));
  OAI221xp5_ASAP7_75t_L     g15904(.A1(new_n4536), .A2(new_n6195), .B1(new_n5680), .B2(new_n4781), .C(new_n16160), .Y(new_n16161));
  XNOR2x2_ASAP7_75t_L       g15905(.A(\a[38] ), .B(new_n16161), .Y(new_n16162));
  INVx1_ASAP7_75t_L         g15906(.A(new_n16072), .Y(new_n16163));
  AOI22xp33_ASAP7_75t_L     g15907(.A1(new_n5249), .A2(\b[41] ), .B1(new_n5247), .B2(new_n5669), .Y(new_n16164));
  OAI221xp5_ASAP7_75t_L     g15908(.A1(new_n5241), .A2(new_n5186), .B1(new_n5166), .B2(new_n5521), .C(new_n16164), .Y(new_n16165));
  XNOR2x2_ASAP7_75t_L       g15909(.A(\a[41] ), .B(new_n16165), .Y(new_n16166));
  INVx1_ASAP7_75t_L         g15910(.A(new_n16166), .Y(new_n16167));
  AOI21xp33_ASAP7_75t_L     g15911(.A1(new_n16069), .A2(new_n15992), .B(new_n16067), .Y(new_n16168));
  AOI22xp33_ASAP7_75t_L     g15912(.A1(new_n6002), .A2(\b[38] ), .B1(new_n5999), .B2(new_n4923), .Y(new_n16169));
  OAI221xp5_ASAP7_75t_L     g15913(.A1(new_n6544), .A2(new_n4701), .B1(new_n4465), .B2(new_n6309), .C(new_n16169), .Y(new_n16170));
  XNOR2x2_ASAP7_75t_L       g15914(.A(\a[44] ), .B(new_n16170), .Y(new_n16171));
  INVx1_ASAP7_75t_L         g15915(.A(new_n16061), .Y(new_n16172));
  AOI22xp33_ASAP7_75t_L     g15916(.A1(new_n7659), .A2(\b[32] ), .B1(new_n7656), .B2(new_n3450), .Y(new_n16173));
  OAI221xp5_ASAP7_75t_L     g15917(.A1(new_n8326), .A2(new_n3419), .B1(new_n3212), .B2(new_n7994), .C(new_n16173), .Y(new_n16174));
  XNOR2x2_ASAP7_75t_L       g15918(.A(\a[50] ), .B(new_n16174), .Y(new_n16175));
  INVx1_ASAP7_75t_L         g15919(.A(new_n16035), .Y(new_n16176));
  AOI22xp33_ASAP7_75t_L     g15920(.A1(new_n9623), .A2(\b[26] ), .B1(new_n9620), .B2(new_n2888), .Y(new_n16177));
  OAI221xp5_ASAP7_75t_L     g15921(.A1(new_n10280), .A2(new_n2180), .B1(new_n2019), .B2(new_n12010), .C(new_n16177), .Y(new_n16178));
  XNOR2x2_ASAP7_75t_L       g15922(.A(\a[56] ), .B(new_n16178), .Y(new_n16179));
  INVx1_ASAP7_75t_L         g15923(.A(new_n16179), .Y(new_n16180));
  A2O1A1O1Ixp25_ASAP7_75t_L g15924(.A1(new_n15841), .A2(new_n813), .B(new_n15847), .C(new_n15999), .D(new_n16008), .Y(new_n16181));
  AOI22xp33_ASAP7_75t_L     g15925(.A1(new_n11656), .A2(\b[20] ), .B1(new_n11654), .B2(new_n1600), .Y(new_n16182));
  OAI221xp5_ASAP7_75t_L     g15926(.A1(new_n12364), .A2(new_n1493), .B1(new_n1356), .B2(new_n13003), .C(new_n16182), .Y(new_n16183));
  XNOR2x2_ASAP7_75t_L       g15927(.A(new_n11651), .B(new_n16183), .Y(new_n16184));
  NOR2xp33_ASAP7_75t_L      g15928(.A(new_n1051), .B(new_n12671), .Y(new_n16185));
  A2O1A1Ixp33_ASAP7_75t_L   g15929(.A1(\b[17] ), .A2(new_n12669), .B(new_n16185), .C(new_n15999), .Y(new_n16186));
  O2A1O1Ixp33_ASAP7_75t_L   g15930(.A1(new_n12353), .A2(new_n12355), .B(\b[17] ), .C(new_n16185), .Y(new_n16187));
  A2O1A1Ixp33_ASAP7_75t_L   g15931(.A1(new_n12669), .A2(\b[16] ), .B(new_n15996), .C(new_n16187), .Y(new_n16188));
  AND2x2_ASAP7_75t_L        g15932(.A(new_n16186), .B(new_n16188), .Y(new_n16189));
  XNOR2x2_ASAP7_75t_L       g15933(.A(new_n16189), .B(new_n16184), .Y(new_n16190));
  NAND2xp33_ASAP7_75t_L     g15934(.A(new_n16181), .B(new_n16190), .Y(new_n16191));
  O2A1O1Ixp33_ASAP7_75t_L   g15935(.A1(new_n16004), .A2(new_n16007), .B(new_n16003), .C(new_n16190), .Y(new_n16192));
  INVx1_ASAP7_75t_L         g15936(.A(new_n16192), .Y(new_n16193));
  NAND2xp33_ASAP7_75t_L     g15937(.A(new_n16191), .B(new_n16193), .Y(new_n16194));
  AOI22xp33_ASAP7_75t_L     g15938(.A1(new_n10594), .A2(\b[23] ), .B1(new_n10591), .B2(new_n2002), .Y(new_n16195));
  OAI221xp5_ASAP7_75t_L     g15939(.A1(new_n11335), .A2(new_n1857), .B1(new_n1709), .B2(new_n11330), .C(new_n16195), .Y(new_n16196));
  XNOR2x2_ASAP7_75t_L       g15940(.A(\a[59] ), .B(new_n16196), .Y(new_n16197));
  NAND2xp33_ASAP7_75t_L     g15941(.A(new_n16197), .B(new_n16194), .Y(new_n16198));
  NOR2xp33_ASAP7_75t_L      g15942(.A(new_n16197), .B(new_n16194), .Y(new_n16199));
  INVx1_ASAP7_75t_L         g15943(.A(new_n16199), .Y(new_n16200));
  NAND2xp33_ASAP7_75t_L     g15944(.A(new_n16198), .B(new_n16200), .Y(new_n16201));
  INVx1_ASAP7_75t_L         g15945(.A(new_n16014), .Y(new_n16202));
  O2A1O1Ixp33_ASAP7_75t_L   g15946(.A1(new_n16008), .A2(new_n16009), .B(new_n16202), .C(new_n16020), .Y(new_n16203));
  XNOR2x2_ASAP7_75t_L       g15947(.A(new_n16203), .B(new_n16201), .Y(new_n16204));
  NAND2xp33_ASAP7_75t_L     g15948(.A(new_n16180), .B(new_n16204), .Y(new_n16205));
  INVx1_ASAP7_75t_L         g15949(.A(new_n16201), .Y(new_n16206));
  NAND2xp33_ASAP7_75t_L     g15950(.A(new_n16203), .B(new_n16206), .Y(new_n16207));
  INVx1_ASAP7_75t_L         g15951(.A(new_n16207), .Y(new_n16208));
  O2A1O1Ixp33_ASAP7_75t_L   g15952(.A1(new_n16014), .A2(new_n16010), .B(new_n16021), .C(new_n16206), .Y(new_n16209));
  OAI21xp33_ASAP7_75t_L     g15953(.A1(new_n16209), .A2(new_n16208), .B(new_n16179), .Y(new_n16210));
  NAND2xp33_ASAP7_75t_L     g15954(.A(new_n16205), .B(new_n16210), .Y(new_n16211));
  NAND2xp33_ASAP7_75t_L     g15955(.A(new_n16026), .B(new_n16031), .Y(new_n16212));
  INVx1_ASAP7_75t_L         g15956(.A(new_n16212), .Y(new_n16213));
  XNOR2x2_ASAP7_75t_L       g15957(.A(new_n16213), .B(new_n16211), .Y(new_n16214));
  AOI22xp33_ASAP7_75t_L     g15958(.A1(new_n8645), .A2(\b[29] ), .B1(new_n8642), .B2(new_n5472), .Y(new_n16215));
  OAI221xp5_ASAP7_75t_L     g15959(.A1(new_n9322), .A2(new_n2852), .B1(new_n2650), .B2(new_n8965), .C(new_n16215), .Y(new_n16216));
  XNOR2x2_ASAP7_75t_L       g15960(.A(\a[53] ), .B(new_n16216), .Y(new_n16217));
  NAND2xp33_ASAP7_75t_L     g15961(.A(new_n16217), .B(new_n16214), .Y(new_n16218));
  INVx1_ASAP7_75t_L         g15962(.A(new_n16211), .Y(new_n16219));
  NAND2xp33_ASAP7_75t_L     g15963(.A(new_n16213), .B(new_n16219), .Y(new_n16220));
  INVx1_ASAP7_75t_L         g15964(.A(new_n16026), .Y(new_n16221));
  A2O1A1Ixp33_ASAP7_75t_L   g15965(.A1(new_n16027), .A2(new_n16030), .B(new_n16221), .C(new_n16211), .Y(new_n16222));
  AO21x2_ASAP7_75t_L        g15966(.A1(new_n16222), .A2(new_n16220), .B(new_n16217), .Y(new_n16223));
  NAND2xp33_ASAP7_75t_L     g15967(.A(new_n16218), .B(new_n16223), .Y(new_n16224));
  A2O1A1Ixp33_ASAP7_75t_L   g15968(.A1(new_n16176), .A2(new_n16033), .B(new_n16043), .C(new_n16224), .Y(new_n16225));
  A2O1A1O1Ixp25_ASAP7_75t_L g15969(.A1(new_n15861), .A2(new_n15858), .B(new_n16034), .C(new_n16033), .D(new_n16043), .Y(new_n16226));
  NAND3xp33_ASAP7_75t_L     g15970(.A(new_n16223), .B(new_n16218), .C(new_n16226), .Y(new_n16227));
  NAND3xp33_ASAP7_75t_L     g15971(.A(new_n16225), .B(new_n16175), .C(new_n16227), .Y(new_n16228));
  AO21x2_ASAP7_75t_L        g15972(.A1(new_n16227), .A2(new_n16225), .B(new_n16175), .Y(new_n16229));
  NAND2xp33_ASAP7_75t_L     g15973(.A(new_n16228), .B(new_n16229), .Y(new_n16230));
  O2A1O1Ixp33_ASAP7_75t_L   g15974(.A1(new_n16048), .A2(new_n16054), .B(new_n16047), .C(new_n16230), .Y(new_n16231));
  INVx1_ASAP7_75t_L         g15975(.A(new_n16231), .Y(new_n16232));
  OA21x2_ASAP7_75t_L        g15976(.A1(new_n16054), .A2(new_n16048), .B(new_n16047), .Y(new_n16233));
  NAND2xp33_ASAP7_75t_L     g15977(.A(new_n16233), .B(new_n16230), .Y(new_n16234));
  AOI22xp33_ASAP7_75t_L     g15978(.A1(new_n6822), .A2(\b[35] ), .B1(new_n6819), .B2(new_n5649), .Y(new_n16235));
  OAI221xp5_ASAP7_75t_L     g15979(.A1(new_n7392), .A2(new_n3827), .B1(new_n3807), .B2(new_n7115), .C(new_n16235), .Y(new_n16236));
  XNOR2x2_ASAP7_75t_L       g15980(.A(\a[47] ), .B(new_n16236), .Y(new_n16237));
  AND3x1_ASAP7_75t_L        g15981(.A(new_n16232), .B(new_n16237), .C(new_n16234), .Y(new_n16238));
  AND2x2_ASAP7_75t_L        g15982(.A(new_n16234), .B(new_n16232), .Y(new_n16239));
  NOR2xp33_ASAP7_75t_L      g15983(.A(new_n16237), .B(new_n16239), .Y(new_n16240));
  NOR2xp33_ASAP7_75t_L      g15984(.A(new_n16238), .B(new_n16240), .Y(new_n16241));
  O2A1O1Ixp33_ASAP7_75t_L   g15985(.A1(new_n16172), .A2(new_n16064), .B(new_n16060), .C(new_n16241), .Y(new_n16242));
  NOR2xp33_ASAP7_75t_L      g15986(.A(new_n16064), .B(new_n16172), .Y(new_n16243));
  A2O1A1O1Ixp25_ASAP7_75t_L g15987(.A1(new_n15876), .A2(new_n15874), .B(new_n16057), .C(new_n16055), .D(new_n16243), .Y(new_n16244));
  AND2x2_ASAP7_75t_L        g15988(.A(new_n16244), .B(new_n16241), .Y(new_n16245));
  NOR2xp33_ASAP7_75t_L      g15989(.A(new_n16242), .B(new_n16245), .Y(new_n16246));
  XNOR2x2_ASAP7_75t_L       g15990(.A(new_n16171), .B(new_n16246), .Y(new_n16247));
  XNOR2x2_ASAP7_75t_L       g15991(.A(new_n16168), .B(new_n16247), .Y(new_n16248));
  XNOR2x2_ASAP7_75t_L       g15992(.A(new_n16167), .B(new_n16248), .Y(new_n16249));
  A2O1A1O1Ixp25_ASAP7_75t_L g15993(.A1(new_n15891), .A2(new_n15886), .B(new_n16070), .C(new_n16163), .D(new_n16249), .Y(new_n16250));
  A2O1A1Ixp33_ASAP7_75t_L   g15994(.A1(new_n15891), .A2(new_n15886), .B(new_n16070), .C(new_n16163), .Y(new_n16251));
  INVx1_ASAP7_75t_L         g15995(.A(new_n16249), .Y(new_n16252));
  NOR2xp33_ASAP7_75t_L      g15996(.A(new_n16251), .B(new_n16252), .Y(new_n16253));
  NOR2xp33_ASAP7_75t_L      g15997(.A(new_n16250), .B(new_n16253), .Y(new_n16254));
  XNOR2x2_ASAP7_75t_L       g15998(.A(new_n16162), .B(new_n16254), .Y(new_n16255));
  NOR2xp33_ASAP7_75t_L      g15999(.A(new_n16082), .B(new_n16076), .Y(new_n16256));
  O2A1O1Ixp33_ASAP7_75t_L   g16000(.A1(new_n16072), .A2(new_n16073), .B(new_n15983), .C(new_n16256), .Y(new_n16257));
  XOR2x2_ASAP7_75t_L        g16001(.A(new_n16257), .B(new_n16255), .Y(new_n16258));
  AOI22xp33_ASAP7_75t_L     g16002(.A1(new_n3884), .A2(\b[47] ), .B1(new_n3881), .B2(new_n7323), .Y(new_n16259));
  OAI221xp5_ASAP7_75t_L     g16003(.A1(new_n4312), .A2(new_n7033), .B1(new_n6756), .B2(new_n4986), .C(new_n16259), .Y(new_n16260));
  XNOR2x2_ASAP7_75t_L       g16004(.A(\a[35] ), .B(new_n16260), .Y(new_n16261));
  XNOR2x2_ASAP7_75t_L       g16005(.A(new_n16261), .B(new_n16258), .Y(new_n16262));
  XNOR2x2_ASAP7_75t_L       g16006(.A(new_n16159), .B(new_n16262), .Y(new_n16263));
  NOR2xp33_ASAP7_75t_L      g16007(.A(new_n16151), .B(new_n16263), .Y(new_n16264));
  AND2x2_ASAP7_75t_L        g16008(.A(new_n16151), .B(new_n16263), .Y(new_n16265));
  NOR2xp33_ASAP7_75t_L      g16009(.A(new_n16264), .B(new_n16265), .Y(new_n16266));
  NAND2xp33_ASAP7_75t_L     g16010(.A(new_n16266), .B(new_n16139), .Y(new_n16267));
  OAI22xp33_ASAP7_75t_L     g16011(.A1(new_n16137), .A2(new_n16138), .B1(new_n16265), .B2(new_n16264), .Y(new_n16268));
  NAND2xp33_ASAP7_75t_L     g16012(.A(new_n16268), .B(new_n16267), .Y(new_n16269));
  XOR2x2_ASAP7_75t_L        g16013(.A(new_n16269), .B(new_n16132), .Y(new_n16270));
  INVx1_ASAP7_75t_L         g16014(.A(new_n16270), .Y(new_n16271));
  NOR2xp33_ASAP7_75t_L      g16015(.A(new_n16271), .B(new_n16127), .Y(new_n16272));
  NOR3xp33_ASAP7_75t_L      g16016(.A(new_n16125), .B(new_n16126), .C(new_n16270), .Y(new_n16273));
  A2O1A1Ixp33_ASAP7_75t_L   g16017(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n1110), .Y(new_n16274));
  A2O1A1Ixp33_ASAP7_75t_L   g16018(.A1(new_n16274), .A2(new_n1195), .B(new_n12599), .C(\a[17] ), .Y(new_n16275));
  O2A1O1Ixp33_ASAP7_75t_L   g16019(.A1(new_n1197), .A2(new_n13934), .B(new_n1195), .C(new_n12599), .Y(new_n16276));
  NAND2xp33_ASAP7_75t_L     g16020(.A(new_n1107), .B(new_n16276), .Y(new_n16277));
  AND2x2_ASAP7_75t_L        g16021(.A(new_n16277), .B(new_n16275), .Y(new_n16278));
  INVx1_ASAP7_75t_L         g16022(.A(new_n16278), .Y(new_n16279));
  A2O1A1Ixp33_ASAP7_75t_L   g16023(.A1(new_n15956), .A2(new_n16102), .B(new_n15955), .C(new_n16279), .Y(new_n16280));
  INVx1_ASAP7_75t_L         g16024(.A(new_n15955), .Y(new_n16281));
  NAND3xp33_ASAP7_75t_L     g16025(.A(new_n16103), .B(new_n16281), .C(new_n16278), .Y(new_n16282));
  NAND2xp33_ASAP7_75t_L     g16026(.A(new_n16280), .B(new_n16282), .Y(new_n16283));
  OR3x1_ASAP7_75t_L         g16027(.A(new_n16283), .B(new_n16272), .C(new_n16273), .Y(new_n16284));
  OR2x4_ASAP7_75t_L         g16028(.A(new_n16273), .B(new_n16272), .Y(new_n16285));
  NAND2xp33_ASAP7_75t_L     g16029(.A(new_n16283), .B(new_n16285), .Y(new_n16286));
  AND2x2_ASAP7_75t_L        g16030(.A(new_n15946), .B(new_n16106), .Y(new_n16287));
  AND3x1_ASAP7_75t_L        g16031(.A(new_n16287), .B(new_n16286), .C(new_n16284), .Y(new_n16288));
  AOI21xp33_ASAP7_75t_L     g16032(.A1(new_n16284), .A2(new_n16286), .B(new_n16287), .Y(new_n16289));
  NOR2xp33_ASAP7_75t_L      g16033(.A(new_n16289), .B(new_n16288), .Y(new_n16290));
  A2O1A1Ixp33_ASAP7_75t_L   g16034(.A1(new_n16117), .A2(new_n16113), .B(new_n16112), .C(new_n16290), .Y(new_n16291));
  INVx1_ASAP7_75t_L         g16035(.A(new_n16291), .Y(new_n16292));
  INVx1_ASAP7_75t_L         g16036(.A(new_n16112), .Y(new_n16293));
  A2O1A1Ixp33_ASAP7_75t_L   g16037(.A1(new_n15933), .A2(new_n15930), .B(new_n16114), .C(new_n16293), .Y(new_n16294));
  NOR2xp33_ASAP7_75t_L      g16038(.A(new_n16290), .B(new_n16294), .Y(new_n16295));
  NOR2xp33_ASAP7_75t_L      g16039(.A(new_n16292), .B(new_n16295), .Y(\f[80] ));
  NOR2xp33_ASAP7_75t_L      g16040(.A(new_n16283), .B(new_n16285), .Y(new_n16297));
  A2O1A1O1Ixp25_ASAP7_75t_L g16041(.A1(new_n15956), .A2(new_n16102), .B(new_n15955), .C(new_n16279), .D(new_n16297), .Y(new_n16298));
  INVx1_ASAP7_75t_L         g16042(.A(new_n16126), .Y(new_n16299));
  NAND2xp33_ASAP7_75t_L     g16043(.A(\b[63] ), .B(new_n1406), .Y(new_n16300));
  A2O1A1Ixp33_ASAP7_75t_L   g16044(.A1(new_n12607), .A2(new_n12603), .B(new_n1411), .C(new_n16300), .Y(new_n16301));
  AOI221xp5_ASAP7_75t_L     g16045(.A1(\b[61] ), .A2(new_n1548), .B1(\b[62] ), .B2(new_n1410), .C(new_n16301), .Y(new_n16302));
  XNOR2x2_ASAP7_75t_L       g16046(.A(new_n1401), .B(new_n16302), .Y(new_n16303));
  INVx1_ASAP7_75t_L         g16047(.A(new_n16303), .Y(new_n16304));
  O2A1O1Ixp33_ASAP7_75t_L   g16048(.A1(new_n16270), .A2(new_n16125), .B(new_n16299), .C(new_n16304), .Y(new_n16305));
  INVx1_ASAP7_75t_L         g16049(.A(new_n16305), .Y(new_n16306));
  INVx1_ASAP7_75t_L         g16050(.A(new_n15961), .Y(new_n16307));
  A2O1A1O1Ixp25_ASAP7_75t_L g16051(.A1(new_n15962), .A2(new_n16098), .B(new_n16307), .C(new_n16123), .D(new_n16273), .Y(new_n16308));
  NAND2xp33_ASAP7_75t_L     g16052(.A(new_n16304), .B(new_n16308), .Y(new_n16309));
  AOI22xp33_ASAP7_75t_L     g16053(.A1(new_n1766), .A2(\b[60] ), .B1(new_n1764), .B2(new_n11234), .Y(new_n16310));
  OAI221xp5_ASAP7_75t_L     g16054(.A1(new_n1758), .A2(new_n10881), .B1(new_n10848), .B2(new_n1911), .C(new_n16310), .Y(new_n16311));
  XNOR2x2_ASAP7_75t_L       g16055(.A(new_n1761), .B(new_n16311), .Y(new_n16312));
  INVx1_ASAP7_75t_L         g16056(.A(new_n16131), .Y(new_n16313));
  MAJIxp5_ASAP7_75t_L       g16057(.A(new_n16269), .B(new_n16130), .C(new_n16313), .Y(new_n16314));
  NOR2xp33_ASAP7_75t_L      g16058(.A(new_n16312), .B(new_n16314), .Y(new_n16315));
  AND2x2_ASAP7_75t_L        g16059(.A(new_n16312), .B(new_n16314), .Y(new_n16316));
  NOR2xp33_ASAP7_75t_L      g16060(.A(new_n16315), .B(new_n16316), .Y(new_n16317));
  AOI22xp33_ASAP7_75t_L     g16061(.A1(new_n2702), .A2(\b[54] ), .B1(new_n2700), .B2(new_n9208), .Y(new_n16318));
  OAI221xp5_ASAP7_75t_L     g16062(.A1(new_n2694), .A2(new_n8882), .B1(new_n8569), .B2(new_n2932), .C(new_n16318), .Y(new_n16319));
  XNOR2x2_ASAP7_75t_L       g16063(.A(\a[29] ), .B(new_n16319), .Y(new_n16320));
  INVx1_ASAP7_75t_L         g16064(.A(new_n16320), .Y(new_n16321));
  A2O1A1O1Ixp25_ASAP7_75t_L g16065(.A1(new_n16092), .A2(new_n16091), .B(new_n15981), .C(new_n16146), .D(new_n16144), .Y(new_n16322));
  OR3x1_ASAP7_75t_L         g16066(.A(new_n16264), .B(new_n16321), .C(new_n16322), .Y(new_n16323));
  A2O1A1Ixp33_ASAP7_75t_L   g16067(.A1(new_n16147), .A2(new_n16149), .B(new_n16264), .C(new_n16321), .Y(new_n16324));
  O2A1O1Ixp33_ASAP7_75t_L   g16068(.A1(new_n16076), .A2(new_n16082), .B(new_n16075), .C(new_n16255), .Y(new_n16325));
  A2O1A1Ixp33_ASAP7_75t_L   g16069(.A1(new_n16069), .A2(new_n15992), .B(new_n16067), .C(new_n16247), .Y(new_n16326));
  NAND2xp33_ASAP7_75t_L     g16070(.A(new_n16167), .B(new_n16248), .Y(new_n16327));
  AND2x2_ASAP7_75t_L        g16071(.A(new_n16326), .B(new_n16327), .Y(new_n16328));
  AOI22xp33_ASAP7_75t_L     g16072(.A1(new_n5249), .A2(\b[42] ), .B1(new_n5247), .B2(new_n5688), .Y(new_n16329));
  OAI221xp5_ASAP7_75t_L     g16073(.A1(new_n5241), .A2(new_n5666), .B1(new_n5186), .B2(new_n5521), .C(new_n16329), .Y(new_n16330));
  XNOR2x2_ASAP7_75t_L       g16074(.A(new_n5244), .B(new_n16330), .Y(new_n16331));
  MAJIxp5_ASAP7_75t_L       g16075(.A(new_n16241), .B(new_n16171), .C(new_n16244), .Y(new_n16332));
  INVx1_ASAP7_75t_L         g16076(.A(new_n16218), .Y(new_n16333));
  INVx1_ASAP7_75t_L         g16077(.A(new_n16181), .Y(new_n16334));
  INVx1_ASAP7_75t_L         g16078(.A(new_n16190), .Y(new_n16335));
  AOI22xp33_ASAP7_75t_L     g16079(.A1(new_n10594), .A2(\b[24] ), .B1(new_n10591), .B2(new_n2027), .Y(new_n16336));
  OAI221xp5_ASAP7_75t_L     g16080(.A1(new_n11335), .A2(new_n1995), .B1(new_n1857), .B2(new_n11330), .C(new_n16336), .Y(new_n16337));
  XNOR2x2_ASAP7_75t_L       g16081(.A(\a[59] ), .B(new_n16337), .Y(new_n16338));
  INVx1_ASAP7_75t_L         g16082(.A(new_n16338), .Y(new_n16339));
  AOI22xp33_ASAP7_75t_L     g16083(.A1(new_n11656), .A2(\b[21] ), .B1(new_n11654), .B2(new_n1715), .Y(new_n16340));
  OAI221xp5_ASAP7_75t_L     g16084(.A1(new_n12364), .A2(new_n1594), .B1(new_n1493), .B2(new_n13003), .C(new_n16340), .Y(new_n16341));
  XNOR2x2_ASAP7_75t_L       g16085(.A(\a[62] ), .B(new_n16341), .Y(new_n16342));
  INVx1_ASAP7_75t_L         g16086(.A(new_n16187), .Y(new_n16343));
  NOR2xp33_ASAP7_75t_L      g16087(.A(new_n1244), .B(new_n12671), .Y(new_n16344));
  A2O1A1Ixp33_ASAP7_75t_L   g16088(.A1(new_n12669), .A2(\b[18] ), .B(new_n16344), .C(new_n1107), .Y(new_n16345));
  O2A1O1Ixp33_ASAP7_75t_L   g16089(.A1(new_n12353), .A2(new_n12355), .B(\b[18] ), .C(new_n16344), .Y(new_n16346));
  NAND2xp33_ASAP7_75t_L     g16090(.A(\a[17] ), .B(new_n16346), .Y(new_n16347));
  NAND2xp33_ASAP7_75t_L     g16091(.A(new_n16345), .B(new_n16347), .Y(new_n16348));
  XNOR2x2_ASAP7_75t_L       g16092(.A(new_n16343), .B(new_n16348), .Y(new_n16349));
  INVx1_ASAP7_75t_L         g16093(.A(new_n16349), .Y(new_n16350));
  XNOR2x2_ASAP7_75t_L       g16094(.A(new_n16350), .B(new_n16342), .Y(new_n16351));
  INVx1_ASAP7_75t_L         g16095(.A(new_n16351), .Y(new_n16352));
  A2O1A1O1Ixp25_ASAP7_75t_L g16096(.A1(new_n12669), .A2(\b[16] ), .B(new_n15996), .C(new_n16187), .D(new_n16184), .Y(new_n16353));
  A2O1A1O1Ixp25_ASAP7_75t_L g16097(.A1(new_n12669), .A2(\b[17] ), .B(new_n16185), .C(new_n15999), .D(new_n16353), .Y(new_n16354));
  NAND2xp33_ASAP7_75t_L     g16098(.A(new_n16354), .B(new_n16352), .Y(new_n16355));
  A2O1A1Ixp33_ASAP7_75t_L   g16099(.A1(new_n15999), .A2(new_n16343), .B(new_n16353), .C(new_n16351), .Y(new_n16356));
  AO21x2_ASAP7_75t_L        g16100(.A1(new_n16356), .A2(new_n16355), .B(new_n16339), .Y(new_n16357));
  AND2x2_ASAP7_75t_L        g16101(.A(new_n16356), .B(new_n16355), .Y(new_n16358));
  NAND2xp33_ASAP7_75t_L     g16102(.A(new_n16339), .B(new_n16358), .Y(new_n16359));
  AND2x2_ASAP7_75t_L        g16103(.A(new_n16357), .B(new_n16359), .Y(new_n16360));
  A2O1A1Ixp33_ASAP7_75t_L   g16104(.A1(new_n16335), .A2(new_n16334), .B(new_n16199), .C(new_n16360), .Y(new_n16361));
  INVx1_ASAP7_75t_L         g16105(.A(new_n16361), .Y(new_n16362));
  NOR3xp33_ASAP7_75t_L      g16106(.A(new_n16360), .B(new_n16199), .C(new_n16192), .Y(new_n16363));
  NOR2xp33_ASAP7_75t_L      g16107(.A(new_n16363), .B(new_n16362), .Y(new_n16364));
  AOI22xp33_ASAP7_75t_L     g16108(.A1(new_n9623), .A2(\b[27] ), .B1(new_n9620), .B2(new_n2657), .Y(new_n16365));
  OAI221xp5_ASAP7_75t_L     g16109(.A1(new_n10280), .A2(new_n2477), .B1(new_n2180), .B2(new_n12010), .C(new_n16365), .Y(new_n16366));
  XNOR2x2_ASAP7_75t_L       g16110(.A(\a[56] ), .B(new_n16366), .Y(new_n16367));
  INVx1_ASAP7_75t_L         g16111(.A(new_n16367), .Y(new_n16368));
  XNOR2x2_ASAP7_75t_L       g16112(.A(new_n16368), .B(new_n16364), .Y(new_n16369));
  AND3x1_ASAP7_75t_L        g16113(.A(new_n16369), .B(new_n16205), .C(new_n16207), .Y(new_n16370));
  O2A1O1Ixp33_ASAP7_75t_L   g16114(.A1(new_n16179), .A2(new_n16209), .B(new_n16207), .C(new_n16369), .Y(new_n16371));
  NOR2xp33_ASAP7_75t_L      g16115(.A(new_n16371), .B(new_n16370), .Y(new_n16372));
  AOI22xp33_ASAP7_75t_L     g16116(.A1(new_n8645), .A2(\b[30] ), .B1(new_n8642), .B2(new_n3219), .Y(new_n16373));
  OAI221xp5_ASAP7_75t_L     g16117(.A1(new_n9322), .A2(new_n2871), .B1(new_n2852), .B2(new_n8965), .C(new_n16373), .Y(new_n16374));
  XNOR2x2_ASAP7_75t_L       g16118(.A(\a[53] ), .B(new_n16374), .Y(new_n16375));
  INVx1_ASAP7_75t_L         g16119(.A(new_n16375), .Y(new_n16376));
  XNOR2x2_ASAP7_75t_L       g16120(.A(new_n16376), .B(new_n16372), .Y(new_n16377));
  A2O1A1Ixp33_ASAP7_75t_L   g16121(.A1(new_n16212), .A2(new_n16211), .B(new_n16333), .C(new_n16377), .Y(new_n16378));
  A2O1A1Ixp33_ASAP7_75t_L   g16122(.A1(new_n16031), .A2(new_n16026), .B(new_n16219), .C(new_n16218), .Y(new_n16379));
  OR2x4_ASAP7_75t_L         g16123(.A(new_n16379), .B(new_n16377), .Y(new_n16380));
  NAND2xp33_ASAP7_75t_L     g16124(.A(new_n16378), .B(new_n16380), .Y(new_n16381));
  AOI22xp33_ASAP7_75t_L     g16125(.A1(new_n7659), .A2(\b[33] ), .B1(new_n7656), .B2(new_n3813), .Y(new_n16382));
  OAI221xp5_ASAP7_75t_L     g16126(.A1(new_n8326), .A2(new_n3443), .B1(new_n3419), .B2(new_n7994), .C(new_n16382), .Y(new_n16383));
  XNOR2x2_ASAP7_75t_L       g16127(.A(\a[50] ), .B(new_n16383), .Y(new_n16384));
  INVx1_ASAP7_75t_L         g16128(.A(new_n16384), .Y(new_n16385));
  NAND3xp33_ASAP7_75t_L     g16129(.A(new_n16228), .B(new_n16227), .C(new_n16385), .Y(new_n16386));
  INVx1_ASAP7_75t_L         g16130(.A(new_n16226), .Y(new_n16387));
  O2A1O1Ixp33_ASAP7_75t_L   g16131(.A1(new_n16224), .A2(new_n16387), .B(new_n16228), .C(new_n16385), .Y(new_n16388));
  INVx1_ASAP7_75t_L         g16132(.A(new_n16388), .Y(new_n16389));
  AND2x2_ASAP7_75t_L        g16133(.A(new_n16386), .B(new_n16389), .Y(new_n16390));
  NAND2xp33_ASAP7_75t_L     g16134(.A(new_n16381), .B(new_n16390), .Y(new_n16391));
  AO21x2_ASAP7_75t_L        g16135(.A1(new_n16386), .A2(new_n16389), .B(new_n16381), .Y(new_n16392));
  AOI22xp33_ASAP7_75t_L     g16136(.A1(new_n6822), .A2(\b[36] ), .B1(new_n6819), .B2(new_n4473), .Y(new_n16393));
  OAI221xp5_ASAP7_75t_L     g16137(.A1(new_n7392), .A2(new_n4053), .B1(new_n3827), .B2(new_n7115), .C(new_n16393), .Y(new_n16394));
  XNOR2x2_ASAP7_75t_L       g16138(.A(\a[47] ), .B(new_n16394), .Y(new_n16395));
  AO21x2_ASAP7_75t_L        g16139(.A1(new_n16392), .A2(new_n16391), .B(new_n16395), .Y(new_n16396));
  NAND3xp33_ASAP7_75t_L     g16140(.A(new_n16391), .B(new_n16392), .C(new_n16395), .Y(new_n16397));
  AND2x2_ASAP7_75t_L        g16141(.A(new_n16397), .B(new_n16396), .Y(new_n16398));
  INVx1_ASAP7_75t_L         g16142(.A(new_n16398), .Y(new_n16399));
  A2O1A1Ixp33_ASAP7_75t_L   g16143(.A1(new_n16234), .A2(new_n16237), .B(new_n16231), .C(new_n16399), .Y(new_n16400));
  NOR2xp33_ASAP7_75t_L      g16144(.A(new_n16231), .B(new_n16238), .Y(new_n16401));
  NAND2xp33_ASAP7_75t_L     g16145(.A(new_n16401), .B(new_n16398), .Y(new_n16402));
  NAND2xp33_ASAP7_75t_L     g16146(.A(new_n16402), .B(new_n16400), .Y(new_n16403));
  AOI22xp33_ASAP7_75t_L     g16147(.A1(new_n6002), .A2(\b[39] ), .B1(new_n5999), .B2(new_n5174), .Y(new_n16404));
  OAI221xp5_ASAP7_75t_L     g16148(.A1(new_n6544), .A2(new_n4915), .B1(new_n4701), .B2(new_n6309), .C(new_n16404), .Y(new_n16405));
  XNOR2x2_ASAP7_75t_L       g16149(.A(\a[44] ), .B(new_n16405), .Y(new_n16406));
  XNOR2x2_ASAP7_75t_L       g16150(.A(new_n16406), .B(new_n16403), .Y(new_n16407));
  XNOR2x2_ASAP7_75t_L       g16151(.A(new_n16332), .B(new_n16407), .Y(new_n16408));
  NAND2xp33_ASAP7_75t_L     g16152(.A(new_n16331), .B(new_n16408), .Y(new_n16409));
  INVx1_ASAP7_75t_L         g16153(.A(new_n16409), .Y(new_n16410));
  NOR2xp33_ASAP7_75t_L      g16154(.A(new_n16331), .B(new_n16408), .Y(new_n16411));
  OAI21xp33_ASAP7_75t_L     g16155(.A1(new_n16411), .A2(new_n16410), .B(new_n16328), .Y(new_n16412));
  OR3x1_ASAP7_75t_L         g16156(.A(new_n16410), .B(new_n16328), .C(new_n16411), .Y(new_n16413));
  NAND2xp33_ASAP7_75t_L     g16157(.A(new_n16412), .B(new_n16413), .Y(new_n16414));
  AOI22xp33_ASAP7_75t_L     g16158(.A1(new_n4544), .A2(\b[45] ), .B1(new_n4542), .B2(new_n6764), .Y(new_n16415));
  OAI221xp5_ASAP7_75t_L     g16159(.A1(new_n4536), .A2(new_n6220), .B1(new_n6195), .B2(new_n4781), .C(new_n16415), .Y(new_n16416));
  XNOR2x2_ASAP7_75t_L       g16160(.A(\a[38] ), .B(new_n16416), .Y(new_n16417));
  XNOR2x2_ASAP7_75t_L       g16161(.A(new_n16417), .B(new_n16414), .Y(new_n16418));
  INVx1_ASAP7_75t_L         g16162(.A(new_n16162), .Y(new_n16419));
  AOI21xp33_ASAP7_75t_L     g16163(.A1(new_n16254), .A2(new_n16419), .B(new_n16250), .Y(new_n16420));
  XOR2x2_ASAP7_75t_L        g16164(.A(new_n16420), .B(new_n16418), .Y(new_n16421));
  AOI22xp33_ASAP7_75t_L     g16165(.A1(new_n3884), .A2(\b[48] ), .B1(new_n3881), .B2(new_n7341), .Y(new_n16422));
  OAI221xp5_ASAP7_75t_L     g16166(.A1(new_n4312), .A2(new_n7316), .B1(new_n7033), .B2(new_n4986), .C(new_n16422), .Y(new_n16423));
  XNOR2x2_ASAP7_75t_L       g16167(.A(\a[35] ), .B(new_n16423), .Y(new_n16424));
  XNOR2x2_ASAP7_75t_L       g16168(.A(new_n16424), .B(new_n16421), .Y(new_n16425));
  INVx1_ASAP7_75t_L         g16169(.A(new_n16425), .Y(new_n16426));
  A2O1A1Ixp33_ASAP7_75t_L   g16170(.A1(new_n16258), .A2(new_n16261), .B(new_n16325), .C(new_n16426), .Y(new_n16427));
  AOI21xp33_ASAP7_75t_L     g16171(.A1(new_n16258), .A2(new_n16261), .B(new_n16325), .Y(new_n16428));
  NAND2xp33_ASAP7_75t_L     g16172(.A(new_n16428), .B(new_n16425), .Y(new_n16429));
  NAND2xp33_ASAP7_75t_L     g16173(.A(new_n16429), .B(new_n16427), .Y(new_n16430));
  AOI22xp33_ASAP7_75t_L     g16174(.A1(new_n3256), .A2(\b[51] ), .B1(new_n3254), .B2(new_n8257), .Y(new_n16431));
  OAI221xp5_ASAP7_75t_L     g16175(.A1(new_n3248), .A2(new_n8228), .B1(new_n7907), .B2(new_n3492), .C(new_n16431), .Y(new_n16432));
  XNOR2x2_ASAP7_75t_L       g16176(.A(\a[32] ), .B(new_n16432), .Y(new_n16433));
  INVx1_ASAP7_75t_L         g16177(.A(new_n16433), .Y(new_n16434));
  A2O1A1Ixp33_ASAP7_75t_L   g16178(.A1(new_n16262), .A2(new_n16159), .B(new_n16158), .C(new_n16434), .Y(new_n16435));
  AOI21xp33_ASAP7_75t_L     g16179(.A1(new_n16262), .A2(new_n16159), .B(new_n16158), .Y(new_n16436));
  NAND2xp33_ASAP7_75t_L     g16180(.A(new_n16433), .B(new_n16436), .Y(new_n16437));
  NAND2xp33_ASAP7_75t_L     g16181(.A(new_n16435), .B(new_n16437), .Y(new_n16438));
  XNOR2x2_ASAP7_75t_L       g16182(.A(new_n16438), .B(new_n16430), .Y(new_n16439));
  NAND3xp33_ASAP7_75t_L     g16183(.A(new_n16439), .B(new_n16324), .C(new_n16323), .Y(new_n16440));
  AO21x2_ASAP7_75t_L        g16184(.A1(new_n16323), .A2(new_n16324), .B(new_n16439), .Y(new_n16441));
  AOI22xp33_ASAP7_75t_L     g16185(.A1(new_n2228), .A2(\b[57] ), .B1(new_n2226), .B2(new_n10495), .Y(new_n16442));
  OAI221xp5_ASAP7_75t_L     g16186(.A1(new_n2220), .A2(new_n10178), .B1(new_n9534), .B2(new_n2387), .C(new_n16442), .Y(new_n16443));
  XNOR2x2_ASAP7_75t_L       g16187(.A(\a[26] ), .B(new_n16443), .Y(new_n16444));
  O2A1O1Ixp33_ASAP7_75t_L   g16188(.A1(new_n16135), .A2(new_n16136), .B(new_n16267), .C(new_n16444), .Y(new_n16445));
  INVx1_ASAP7_75t_L         g16189(.A(new_n16444), .Y(new_n16446));
  OAI21xp33_ASAP7_75t_L     g16190(.A1(new_n16135), .A2(new_n16136), .B(new_n16267), .Y(new_n16447));
  NOR2xp33_ASAP7_75t_L      g16191(.A(new_n16446), .B(new_n16447), .Y(new_n16448));
  NOR2xp33_ASAP7_75t_L      g16192(.A(new_n16445), .B(new_n16448), .Y(new_n16449));
  AO21x2_ASAP7_75t_L        g16193(.A1(new_n16440), .A2(new_n16441), .B(new_n16449), .Y(new_n16450));
  AND2x2_ASAP7_75t_L        g16194(.A(new_n16440), .B(new_n16441), .Y(new_n16451));
  NAND2xp33_ASAP7_75t_L     g16195(.A(new_n16451), .B(new_n16449), .Y(new_n16452));
  AND2x2_ASAP7_75t_L        g16196(.A(new_n16452), .B(new_n16450), .Y(new_n16453));
  NAND2xp33_ASAP7_75t_L     g16197(.A(new_n16317), .B(new_n16453), .Y(new_n16454));
  AO21x2_ASAP7_75t_L        g16198(.A1(new_n16452), .A2(new_n16450), .B(new_n16317), .Y(new_n16455));
  AND2x2_ASAP7_75t_L        g16199(.A(new_n16455), .B(new_n16454), .Y(new_n16456));
  AOI21xp33_ASAP7_75t_L     g16200(.A1(new_n16309), .A2(new_n16306), .B(new_n16456), .Y(new_n16457));
  AND3x1_ASAP7_75t_L        g16201(.A(new_n16309), .B(new_n16456), .C(new_n16306), .Y(new_n16458));
  OR3x1_ASAP7_75t_L         g16202(.A(new_n16298), .B(new_n16458), .C(new_n16457), .Y(new_n16459));
  OAI21xp33_ASAP7_75t_L     g16203(.A1(new_n16457), .A2(new_n16458), .B(new_n16298), .Y(new_n16460));
  NAND2xp33_ASAP7_75t_L     g16204(.A(new_n16460), .B(new_n16459), .Y(new_n16461));
  INVx1_ASAP7_75t_L         g16205(.A(new_n16461), .Y(new_n16462));
  A2O1A1Ixp33_ASAP7_75t_L   g16206(.A1(new_n16294), .A2(new_n16290), .B(new_n16288), .C(new_n16462), .Y(new_n16463));
  A2O1A1O1Ixp25_ASAP7_75t_L g16207(.A1(new_n16113), .A2(new_n16117), .B(new_n16112), .C(new_n16290), .D(new_n16288), .Y(new_n16464));
  NAND2xp33_ASAP7_75t_L     g16208(.A(new_n16461), .B(new_n16464), .Y(new_n16465));
  AND2x2_ASAP7_75t_L        g16209(.A(new_n16465), .B(new_n16463), .Y(\f[81] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16210(.A1(new_n16127), .A2(new_n16271), .B(new_n16126), .C(new_n16304), .Y(new_n16467));
  AOI22xp33_ASAP7_75t_L     g16211(.A1(new_n1766), .A2(\b[61] ), .B1(new_n1764), .B2(new_n11919), .Y(new_n16468));
  OAI221xp5_ASAP7_75t_L     g16212(.A1(new_n1758), .A2(new_n11226), .B1(new_n10881), .B2(new_n1911), .C(new_n16468), .Y(new_n16469));
  XNOR2x2_ASAP7_75t_L       g16213(.A(\a[23] ), .B(new_n16469), .Y(new_n16470));
  INVx1_ASAP7_75t_L         g16214(.A(new_n16470), .Y(new_n16471));
  O2A1O1Ixp33_ASAP7_75t_L   g16215(.A1(new_n16446), .A2(new_n16447), .B(new_n16452), .C(new_n16471), .Y(new_n16472));
  INVx1_ASAP7_75t_L         g16216(.A(new_n16472), .Y(new_n16473));
  AOI21xp33_ASAP7_75t_L     g16217(.A1(new_n16449), .A2(new_n16451), .B(new_n16448), .Y(new_n16474));
  NAND2xp33_ASAP7_75t_L     g16218(.A(new_n16471), .B(new_n16474), .Y(new_n16475));
  NAND2xp33_ASAP7_75t_L     g16219(.A(new_n16475), .B(new_n16473), .Y(new_n16476));
  AOI22xp33_ASAP7_75t_L     g16220(.A1(new_n2228), .A2(\b[58] ), .B1(new_n2226), .B2(new_n10857), .Y(new_n16477));
  OAI221xp5_ASAP7_75t_L     g16221(.A1(new_n2220), .A2(new_n10488), .B1(new_n10178), .B2(new_n2387), .C(new_n16477), .Y(new_n16478));
  XNOR2x2_ASAP7_75t_L       g16222(.A(\a[26] ), .B(new_n16478), .Y(new_n16479));
  NAND2xp33_ASAP7_75t_L     g16223(.A(new_n16323), .B(new_n16440), .Y(new_n16480));
  XNOR2x2_ASAP7_75t_L       g16224(.A(new_n16479), .B(new_n16480), .Y(new_n16481));
  AOI22xp33_ASAP7_75t_L     g16225(.A1(new_n2702), .A2(\b[55] ), .B1(new_n2700), .B2(new_n9542), .Y(new_n16482));
  OAI221xp5_ASAP7_75t_L     g16226(.A1(new_n2694), .A2(new_n9199), .B1(new_n8882), .B2(new_n2932), .C(new_n16482), .Y(new_n16483));
  XNOR2x2_ASAP7_75t_L       g16227(.A(\a[29] ), .B(new_n16483), .Y(new_n16484));
  A2O1A1Ixp33_ASAP7_75t_L   g16228(.A1(new_n16427), .A2(new_n16429), .B(new_n16438), .C(new_n16437), .Y(new_n16485));
  XNOR2x2_ASAP7_75t_L       g16229(.A(new_n16484), .B(new_n16485), .Y(new_n16486));
  AOI22xp33_ASAP7_75t_L     g16230(.A1(new_n3256), .A2(\b[52] ), .B1(new_n3254), .B2(new_n8577), .Y(new_n16487));
  OAI221xp5_ASAP7_75t_L     g16231(.A1(new_n3248), .A2(new_n8249), .B1(new_n8228), .B2(new_n3492), .C(new_n16487), .Y(new_n16488));
  XNOR2x2_ASAP7_75t_L       g16232(.A(\a[32] ), .B(new_n16488), .Y(new_n16489));
  INVx1_ASAP7_75t_L         g16233(.A(new_n16424), .Y(new_n16490));
  NAND2xp33_ASAP7_75t_L     g16234(.A(new_n16490), .B(new_n16421), .Y(new_n16491));
  AND3x1_ASAP7_75t_L        g16235(.A(new_n16429), .B(new_n16491), .C(new_n16489), .Y(new_n16492));
  INVx1_ASAP7_75t_L         g16236(.A(new_n16428), .Y(new_n16493));
  O2A1O1Ixp33_ASAP7_75t_L   g16237(.A1(new_n16493), .A2(new_n16426), .B(new_n16491), .C(new_n16489), .Y(new_n16494));
  INVx1_ASAP7_75t_L         g16238(.A(new_n16332), .Y(new_n16495));
  MAJIxp5_ASAP7_75t_L       g16239(.A(new_n16403), .B(new_n16495), .C(new_n16406), .Y(new_n16496));
  INVx1_ASAP7_75t_L         g16240(.A(new_n16496), .Y(new_n16497));
  AOI22xp33_ASAP7_75t_L     g16241(.A1(new_n6002), .A2(\b[40] ), .B1(new_n5999), .B2(new_n5194), .Y(new_n16498));
  OAI221xp5_ASAP7_75t_L     g16242(.A1(new_n6544), .A2(new_n5166), .B1(new_n4915), .B2(new_n6309), .C(new_n16498), .Y(new_n16499));
  XNOR2x2_ASAP7_75t_L       g16243(.A(\a[44] ), .B(new_n16499), .Y(new_n16500));
  INVx1_ASAP7_75t_L         g16244(.A(new_n16500), .Y(new_n16501));
  A2O1A1Ixp33_ASAP7_75t_L   g16245(.A1(new_n16392), .A2(new_n16391), .B(new_n16395), .C(new_n16402), .Y(new_n16502));
  AOI22xp33_ASAP7_75t_L     g16246(.A1(new_n9623), .A2(\b[28] ), .B1(new_n9620), .B2(new_n2858), .Y(new_n16503));
  OAI221xp5_ASAP7_75t_L     g16247(.A1(new_n10280), .A2(new_n2650), .B1(new_n2477), .B2(new_n12010), .C(new_n16503), .Y(new_n16504));
  XNOR2x2_ASAP7_75t_L       g16248(.A(\a[56] ), .B(new_n16504), .Y(new_n16505));
  INVx1_ASAP7_75t_L         g16249(.A(new_n16359), .Y(new_n16506));
  O2A1O1Ixp33_ASAP7_75t_L   g16250(.A1(new_n16192), .A2(new_n16199), .B(new_n16357), .C(new_n16506), .Y(new_n16507));
  NOR2xp33_ASAP7_75t_L      g16251(.A(new_n1356), .B(new_n12671), .Y(new_n16508));
  INVx1_ASAP7_75t_L         g16252(.A(new_n16345), .Y(new_n16509));
  A2O1A1O1Ixp25_ASAP7_75t_L g16253(.A1(new_n12669), .A2(\b[17] ), .B(new_n16185), .C(new_n16347), .D(new_n16509), .Y(new_n16510));
  A2O1A1Ixp33_ASAP7_75t_L   g16254(.A1(new_n12669), .A2(\b[19] ), .B(new_n16508), .C(new_n16510), .Y(new_n16511));
  O2A1O1Ixp33_ASAP7_75t_L   g16255(.A1(new_n12353), .A2(new_n12355), .B(\b[19] ), .C(new_n16508), .Y(new_n16512));
  INVx1_ASAP7_75t_L         g16256(.A(new_n16512), .Y(new_n16513));
  O2A1O1Ixp33_ASAP7_75t_L   g16257(.A1(new_n16187), .A2(new_n16348), .B(new_n16345), .C(new_n16513), .Y(new_n16514));
  INVx1_ASAP7_75t_L         g16258(.A(new_n16514), .Y(new_n16515));
  NAND2xp33_ASAP7_75t_L     g16259(.A(new_n16511), .B(new_n16515), .Y(new_n16516));
  AOI22xp33_ASAP7_75t_L     g16260(.A1(new_n11656), .A2(\b[22] ), .B1(new_n11654), .B2(new_n1864), .Y(new_n16517));
  OAI221xp5_ASAP7_75t_L     g16261(.A1(new_n12364), .A2(new_n1709), .B1(new_n1594), .B2(new_n13003), .C(new_n16517), .Y(new_n16518));
  XNOR2x2_ASAP7_75t_L       g16262(.A(\a[62] ), .B(new_n16518), .Y(new_n16519));
  NAND2xp33_ASAP7_75t_L     g16263(.A(new_n16516), .B(new_n16519), .Y(new_n16520));
  NOR2xp33_ASAP7_75t_L      g16264(.A(new_n16516), .B(new_n16519), .Y(new_n16521));
  INVx1_ASAP7_75t_L         g16265(.A(new_n16521), .Y(new_n16522));
  AND2x2_ASAP7_75t_L        g16266(.A(new_n16520), .B(new_n16522), .Y(new_n16523));
  OAI21xp33_ASAP7_75t_L     g16267(.A1(new_n16342), .A2(new_n16350), .B(new_n16355), .Y(new_n16524));
  NAND2xp33_ASAP7_75t_L     g16268(.A(new_n16524), .B(new_n16523), .Y(new_n16525));
  NOR2xp33_ASAP7_75t_L      g16269(.A(new_n16524), .B(new_n16523), .Y(new_n16526));
  INVx1_ASAP7_75t_L         g16270(.A(new_n16526), .Y(new_n16527));
  AOI22xp33_ASAP7_75t_L     g16271(.A1(new_n10594), .A2(\b[25] ), .B1(new_n10591), .B2(new_n2188), .Y(new_n16528));
  OAI221xp5_ASAP7_75t_L     g16272(.A1(new_n11335), .A2(new_n2019), .B1(new_n1995), .B2(new_n11330), .C(new_n16528), .Y(new_n16529));
  XNOR2x2_ASAP7_75t_L       g16273(.A(\a[59] ), .B(new_n16529), .Y(new_n16530));
  NAND3xp33_ASAP7_75t_L     g16274(.A(new_n16527), .B(new_n16525), .C(new_n16530), .Y(new_n16531));
  AO21x2_ASAP7_75t_L        g16275(.A1(new_n16525), .A2(new_n16527), .B(new_n16530), .Y(new_n16532));
  AND2x2_ASAP7_75t_L        g16276(.A(new_n16531), .B(new_n16532), .Y(new_n16533));
  XOR2x2_ASAP7_75t_L        g16277(.A(new_n16507), .B(new_n16533), .Y(new_n16534));
  INVx1_ASAP7_75t_L         g16278(.A(new_n16534), .Y(new_n16535));
  NAND2xp33_ASAP7_75t_L     g16279(.A(new_n16505), .B(new_n16535), .Y(new_n16536));
  INVx1_ASAP7_75t_L         g16280(.A(new_n16505), .Y(new_n16537));
  NAND2xp33_ASAP7_75t_L     g16281(.A(new_n16537), .B(new_n16534), .Y(new_n16538));
  NAND2xp33_ASAP7_75t_L     g16282(.A(new_n16368), .B(new_n16364), .Y(new_n16539));
  A2O1A1Ixp33_ASAP7_75t_L   g16283(.A1(new_n16205), .A2(new_n16207), .B(new_n16369), .C(new_n16539), .Y(new_n16540));
  NAND3xp33_ASAP7_75t_L     g16284(.A(new_n16540), .B(new_n16538), .C(new_n16536), .Y(new_n16541));
  AO21x2_ASAP7_75t_L        g16285(.A1(new_n16538), .A2(new_n16536), .B(new_n16540), .Y(new_n16542));
  NAND2xp33_ASAP7_75t_L     g16286(.A(new_n16541), .B(new_n16542), .Y(new_n16543));
  NAND2xp33_ASAP7_75t_L     g16287(.A(\b[31] ), .B(new_n8645), .Y(new_n16544));
  OAI221xp5_ASAP7_75t_L     g16288(.A1(new_n3212), .A2(new_n9322), .B1(new_n8967), .B2(new_n4030), .C(new_n16544), .Y(new_n16545));
  AOI21xp33_ASAP7_75t_L     g16289(.A1(new_n8964), .A2(\b[29] ), .B(new_n16545), .Y(new_n16546));
  NAND2xp33_ASAP7_75t_L     g16290(.A(\a[53] ), .B(new_n16546), .Y(new_n16547));
  A2O1A1Ixp33_ASAP7_75t_L   g16291(.A1(\b[29] ), .A2(new_n8964), .B(new_n16545), .C(new_n8639), .Y(new_n16548));
  NAND2xp33_ASAP7_75t_L     g16292(.A(new_n16548), .B(new_n16547), .Y(new_n16549));
  NOR2xp33_ASAP7_75t_L      g16293(.A(new_n16549), .B(new_n16543), .Y(new_n16550));
  INVx1_ASAP7_75t_L         g16294(.A(new_n16550), .Y(new_n16551));
  NAND2xp33_ASAP7_75t_L     g16295(.A(new_n16549), .B(new_n16543), .Y(new_n16552));
  NAND2xp33_ASAP7_75t_L     g16296(.A(new_n16552), .B(new_n16551), .Y(new_n16553));
  OAI31xp33_ASAP7_75t_L     g16297(.A1(new_n16370), .A2(new_n16375), .A3(new_n16371), .B(new_n16380), .Y(new_n16554));
  XNOR2x2_ASAP7_75t_L       g16298(.A(new_n16553), .B(new_n16554), .Y(new_n16555));
  AOI22xp33_ASAP7_75t_L     g16299(.A1(new_n7659), .A2(\b[34] ), .B1(new_n7656), .B2(new_n3833), .Y(new_n16556));
  OAI221xp5_ASAP7_75t_L     g16300(.A1(new_n8326), .A2(new_n3807), .B1(new_n3443), .B2(new_n7994), .C(new_n16556), .Y(new_n16557));
  XNOR2x2_ASAP7_75t_L       g16301(.A(\a[50] ), .B(new_n16557), .Y(new_n16558));
  INVx1_ASAP7_75t_L         g16302(.A(new_n16558), .Y(new_n16559));
  OR2x4_ASAP7_75t_L         g16303(.A(new_n16559), .B(new_n16555), .Y(new_n16560));
  NAND2xp33_ASAP7_75t_L     g16304(.A(new_n16559), .B(new_n16555), .Y(new_n16561));
  NAND2xp33_ASAP7_75t_L     g16305(.A(new_n16561), .B(new_n16560), .Y(new_n16562));
  A2O1A1Ixp33_ASAP7_75t_L   g16306(.A1(new_n16228), .A2(new_n16227), .B(new_n16385), .C(new_n16391), .Y(new_n16563));
  XNOR2x2_ASAP7_75t_L       g16307(.A(new_n16563), .B(new_n16562), .Y(new_n16564));
  AOI22xp33_ASAP7_75t_L     g16308(.A1(new_n6822), .A2(\b[37] ), .B1(new_n6819), .B2(new_n4709), .Y(new_n16565));
  OAI221xp5_ASAP7_75t_L     g16309(.A1(new_n7392), .A2(new_n4465), .B1(new_n4053), .B2(new_n7115), .C(new_n16565), .Y(new_n16566));
  XNOR2x2_ASAP7_75t_L       g16310(.A(\a[47] ), .B(new_n16566), .Y(new_n16567));
  XNOR2x2_ASAP7_75t_L       g16311(.A(new_n16567), .B(new_n16564), .Y(new_n16568));
  XOR2x2_ASAP7_75t_L        g16312(.A(new_n16502), .B(new_n16568), .Y(new_n16569));
  NAND2xp33_ASAP7_75t_L     g16313(.A(new_n16501), .B(new_n16569), .Y(new_n16570));
  INVx1_ASAP7_75t_L         g16314(.A(new_n16570), .Y(new_n16571));
  NOR2xp33_ASAP7_75t_L      g16315(.A(new_n16501), .B(new_n16569), .Y(new_n16572));
  OR3x1_ASAP7_75t_L         g16316(.A(new_n16571), .B(new_n16497), .C(new_n16572), .Y(new_n16573));
  OAI21xp33_ASAP7_75t_L     g16317(.A1(new_n16572), .A2(new_n16571), .B(new_n16497), .Y(new_n16574));
  NAND2xp33_ASAP7_75t_L     g16318(.A(new_n16574), .B(new_n16573), .Y(new_n16575));
  NAND2xp33_ASAP7_75t_L     g16319(.A(\b[43] ), .B(new_n5249), .Y(new_n16576));
  OAI221xp5_ASAP7_75t_L     g16320(.A1(new_n5680), .A2(new_n5241), .B1(new_n5252), .B2(new_n9799), .C(new_n16576), .Y(new_n16577));
  AOI21xp33_ASAP7_75t_L     g16321(.A1(new_n5526), .A2(\b[41] ), .B(new_n16577), .Y(new_n16578));
  NAND2xp33_ASAP7_75t_L     g16322(.A(\a[41] ), .B(new_n16578), .Y(new_n16579));
  A2O1A1Ixp33_ASAP7_75t_L   g16323(.A1(\b[41] ), .A2(new_n5526), .B(new_n16577), .C(new_n5244), .Y(new_n16580));
  NAND2xp33_ASAP7_75t_L     g16324(.A(new_n16580), .B(new_n16579), .Y(new_n16581));
  XNOR2x2_ASAP7_75t_L       g16325(.A(new_n16581), .B(new_n16575), .Y(new_n16582));
  A2O1A1Ixp33_ASAP7_75t_L   g16326(.A1(new_n16326), .A2(new_n16327), .B(new_n16411), .C(new_n16409), .Y(new_n16583));
  XNOR2x2_ASAP7_75t_L       g16327(.A(new_n16583), .B(new_n16582), .Y(new_n16584));
  AOI22xp33_ASAP7_75t_L     g16328(.A1(new_n4544), .A2(\b[46] ), .B1(new_n4542), .B2(new_n7041), .Y(new_n16585));
  OAI221xp5_ASAP7_75t_L     g16329(.A1(new_n4536), .A2(new_n6756), .B1(new_n6220), .B2(new_n4781), .C(new_n16585), .Y(new_n16586));
  XNOR2x2_ASAP7_75t_L       g16330(.A(\a[38] ), .B(new_n16586), .Y(new_n16587));
  INVx1_ASAP7_75t_L         g16331(.A(new_n16587), .Y(new_n16588));
  XNOR2x2_ASAP7_75t_L       g16332(.A(new_n16588), .B(new_n16584), .Y(new_n16589));
  MAJIxp5_ASAP7_75t_L       g16333(.A(new_n16420), .B(new_n16417), .C(new_n16414), .Y(new_n16590));
  NOR2xp33_ASAP7_75t_L      g16334(.A(new_n16590), .B(new_n16589), .Y(new_n16591));
  AND2x2_ASAP7_75t_L        g16335(.A(new_n16590), .B(new_n16589), .Y(new_n16592));
  NOR2xp33_ASAP7_75t_L      g16336(.A(new_n16591), .B(new_n16592), .Y(new_n16593));
  AOI22xp33_ASAP7_75t_L     g16337(.A1(new_n3884), .A2(\b[49] ), .B1(new_n3881), .B2(new_n7914), .Y(new_n16594));
  OAI221xp5_ASAP7_75t_L     g16338(.A1(new_n4312), .A2(new_n7333), .B1(new_n7316), .B2(new_n4986), .C(new_n16594), .Y(new_n16595));
  XNOR2x2_ASAP7_75t_L       g16339(.A(\a[35] ), .B(new_n16595), .Y(new_n16596));
  NAND2xp33_ASAP7_75t_L     g16340(.A(new_n16596), .B(new_n16593), .Y(new_n16597));
  INVx1_ASAP7_75t_L         g16341(.A(new_n16596), .Y(new_n16598));
  OAI21xp33_ASAP7_75t_L     g16342(.A1(new_n16591), .A2(new_n16592), .B(new_n16598), .Y(new_n16599));
  AND2x2_ASAP7_75t_L        g16343(.A(new_n16599), .B(new_n16597), .Y(new_n16600));
  OR3x1_ASAP7_75t_L         g16344(.A(new_n16600), .B(new_n16492), .C(new_n16494), .Y(new_n16601));
  OAI21xp33_ASAP7_75t_L     g16345(.A1(new_n16494), .A2(new_n16492), .B(new_n16600), .Y(new_n16602));
  NAND2xp33_ASAP7_75t_L     g16346(.A(new_n16602), .B(new_n16601), .Y(new_n16603));
  XNOR2x2_ASAP7_75t_L       g16347(.A(new_n16603), .B(new_n16486), .Y(new_n16604));
  NOR2xp33_ASAP7_75t_L      g16348(.A(new_n16604), .B(new_n16481), .Y(new_n16605));
  AND2x2_ASAP7_75t_L        g16349(.A(new_n16604), .B(new_n16481), .Y(new_n16606));
  NOR2xp33_ASAP7_75t_L      g16350(.A(new_n16605), .B(new_n16606), .Y(new_n16607));
  NOR2xp33_ASAP7_75t_L      g16351(.A(new_n16607), .B(new_n16476), .Y(new_n16608));
  INVx1_ASAP7_75t_L         g16352(.A(new_n16607), .Y(new_n16609));
  AOI21xp33_ASAP7_75t_L     g16353(.A1(new_n16475), .A2(new_n16473), .B(new_n16609), .Y(new_n16610));
  NOR2xp33_ASAP7_75t_L      g16354(.A(new_n16608), .B(new_n16610), .Y(new_n16611));
  A2O1A1Ixp33_ASAP7_75t_L   g16355(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n1404), .Y(new_n16612));
  AOI22xp33_ASAP7_75t_L     g16356(.A1(new_n1410), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1548), .Y(new_n16613));
  NAND3xp33_ASAP7_75t_L     g16357(.A(new_n16612), .B(\a[20] ), .C(new_n16613), .Y(new_n16614));
  INVx1_ASAP7_75t_L         g16358(.A(new_n16614), .Y(new_n16615));
  A2O1A1O1Ixp25_ASAP7_75t_L g16359(.A1(new_n13507), .A2(new_n13506), .B(new_n1411), .C(new_n16613), .D(\a[20] ), .Y(new_n16616));
  NOR2xp33_ASAP7_75t_L      g16360(.A(new_n16616), .B(new_n16615), .Y(new_n16617));
  OAI21xp33_ASAP7_75t_L     g16361(.A1(new_n16312), .A2(new_n16314), .B(new_n16454), .Y(new_n16618));
  NOR2xp33_ASAP7_75t_L      g16362(.A(new_n16617), .B(new_n16618), .Y(new_n16619));
  A2O1A1Ixp33_ASAP7_75t_L   g16363(.A1(new_n16453), .A2(new_n16317), .B(new_n16315), .C(new_n16617), .Y(new_n16620));
  INVx1_ASAP7_75t_L         g16364(.A(new_n16620), .Y(new_n16621));
  NOR3xp33_ASAP7_75t_L      g16365(.A(new_n16611), .B(new_n16619), .C(new_n16621), .Y(new_n16622));
  INVx1_ASAP7_75t_L         g16366(.A(new_n16622), .Y(new_n16623));
  OAI21xp33_ASAP7_75t_L     g16367(.A1(new_n16621), .A2(new_n16619), .B(new_n16611), .Y(new_n16624));
  NAND2xp33_ASAP7_75t_L     g16368(.A(new_n16624), .B(new_n16623), .Y(new_n16625));
  A2O1A1O1Ixp25_ASAP7_75t_L g16369(.A1(new_n16309), .A2(new_n16306), .B(new_n16456), .C(new_n16467), .D(new_n16625), .Y(new_n16626));
  A2O1A1Ixp33_ASAP7_75t_L   g16370(.A1(new_n16309), .A2(new_n16306), .B(new_n16456), .C(new_n16467), .Y(new_n16627));
  AOI21xp33_ASAP7_75t_L     g16371(.A1(new_n16623), .A2(new_n16624), .B(new_n16627), .Y(new_n16628));
  NOR2xp33_ASAP7_75t_L      g16372(.A(new_n16628), .B(new_n16626), .Y(new_n16629));
  INVx1_ASAP7_75t_L         g16373(.A(new_n16629), .Y(new_n16630));
  O2A1O1Ixp33_ASAP7_75t_L   g16374(.A1(new_n16461), .A2(new_n16464), .B(new_n16459), .C(new_n16630), .Y(new_n16631));
  INVx1_ASAP7_75t_L         g16375(.A(new_n16288), .Y(new_n16632));
  A2O1A1Ixp33_ASAP7_75t_L   g16376(.A1(new_n16291), .A2(new_n16632), .B(new_n16461), .C(new_n16459), .Y(new_n16633));
  NOR2xp33_ASAP7_75t_L      g16377(.A(new_n16629), .B(new_n16633), .Y(new_n16634));
  NOR2xp33_ASAP7_75t_L      g16378(.A(new_n16631), .B(new_n16634), .Y(\f[82] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16379(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n1404), .Y(new_n16636));
  A2O1A1Ixp33_ASAP7_75t_L   g16380(.A1(new_n16636), .A2(new_n1549), .B(new_n12599), .C(\a[20] ), .Y(new_n16637));
  O2A1O1Ixp33_ASAP7_75t_L   g16381(.A1(new_n1411), .A2(new_n13934), .B(new_n1549), .C(new_n12599), .Y(new_n16638));
  NAND2xp33_ASAP7_75t_L     g16382(.A(new_n1401), .B(new_n16638), .Y(new_n16639));
  AND2x2_ASAP7_75t_L        g16383(.A(new_n16639), .B(new_n16637), .Y(new_n16640));
  NOR3xp33_ASAP7_75t_L      g16384(.A(new_n16608), .B(new_n16640), .C(new_n16472), .Y(new_n16641));
  INVx1_ASAP7_75t_L         g16385(.A(new_n16641), .Y(new_n16642));
  A2O1A1Ixp33_ASAP7_75t_L   g16386(.A1(new_n16609), .A2(new_n16475), .B(new_n16472), .C(new_n16640), .Y(new_n16643));
  NAND2xp33_ASAP7_75t_L     g16387(.A(new_n16643), .B(new_n16642), .Y(new_n16644));
  AOI22xp33_ASAP7_75t_L     g16388(.A1(new_n1766), .A2(\b[62] ), .B1(new_n1764), .B2(new_n12280), .Y(new_n16645));
  OAI221xp5_ASAP7_75t_L     g16389(.A1(new_n1758), .A2(new_n11911), .B1(new_n11226), .B2(new_n1911), .C(new_n16645), .Y(new_n16646));
  XNOR2x2_ASAP7_75t_L       g16390(.A(\a[23] ), .B(new_n16646), .Y(new_n16647));
  INVx1_ASAP7_75t_L         g16391(.A(new_n16647), .Y(new_n16648));
  MAJIxp5_ASAP7_75t_L       g16392(.A(new_n16604), .B(new_n16479), .C(new_n16480), .Y(new_n16649));
  XNOR2x2_ASAP7_75t_L       g16393(.A(new_n16648), .B(new_n16649), .Y(new_n16650));
  INVx1_ASAP7_75t_L         g16394(.A(new_n16650), .Y(new_n16651));
  AOI22xp33_ASAP7_75t_L     g16395(.A1(new_n2228), .A2(\b[59] ), .B1(new_n2226), .B2(new_n10887), .Y(new_n16652));
  OAI221xp5_ASAP7_75t_L     g16396(.A1(new_n2220), .A2(new_n10848), .B1(new_n10488), .B2(new_n2387), .C(new_n16652), .Y(new_n16653));
  XNOR2x2_ASAP7_75t_L       g16397(.A(new_n2223), .B(new_n16653), .Y(new_n16654));
  MAJIxp5_ASAP7_75t_L       g16398(.A(new_n16603), .B(new_n16484), .C(new_n16485), .Y(new_n16655));
  OR2x4_ASAP7_75t_L         g16399(.A(new_n16654), .B(new_n16655), .Y(new_n16656));
  NAND2xp33_ASAP7_75t_L     g16400(.A(new_n16654), .B(new_n16655), .Y(new_n16657));
  NAND2xp33_ASAP7_75t_L     g16401(.A(new_n16657), .B(new_n16656), .Y(new_n16658));
  AOI22xp33_ASAP7_75t_L     g16402(.A1(new_n2702), .A2(\b[56] ), .B1(new_n2700), .B2(new_n10185), .Y(new_n16659));
  OAI221xp5_ASAP7_75t_L     g16403(.A1(new_n2694), .A2(new_n9534), .B1(new_n9199), .B2(new_n2932), .C(new_n16659), .Y(new_n16660));
  XNOR2x2_ASAP7_75t_L       g16404(.A(\a[29] ), .B(new_n16660), .Y(new_n16661));
  A2O1A1Ixp33_ASAP7_75t_L   g16405(.A1(new_n16491), .A2(new_n16429), .B(new_n16489), .C(new_n16601), .Y(new_n16662));
  XNOR2x2_ASAP7_75t_L       g16406(.A(new_n16661), .B(new_n16662), .Y(new_n16663));
  AOI22xp33_ASAP7_75t_L     g16407(.A1(new_n3256), .A2(\b[53] ), .B1(new_n3254), .B2(new_n8889), .Y(new_n16664));
  OAI221xp5_ASAP7_75t_L     g16408(.A1(new_n3248), .A2(new_n8569), .B1(new_n8249), .B2(new_n3492), .C(new_n16664), .Y(new_n16665));
  XNOR2x2_ASAP7_75t_L       g16409(.A(\a[32] ), .B(new_n16665), .Y(new_n16666));
  AOI21xp33_ASAP7_75t_L     g16410(.A1(new_n16593), .A2(new_n16596), .B(new_n16591), .Y(new_n16667));
  XNOR2x2_ASAP7_75t_L       g16411(.A(new_n16666), .B(new_n16667), .Y(new_n16668));
  AOI22xp33_ASAP7_75t_L     g16412(.A1(new_n5249), .A2(\b[44] ), .B1(new_n5247), .B2(new_n7055), .Y(new_n16669));
  OAI221xp5_ASAP7_75t_L     g16413(.A1(new_n5241), .A2(new_n6195), .B1(new_n5680), .B2(new_n5521), .C(new_n16669), .Y(new_n16670));
  XNOR2x2_ASAP7_75t_L       g16414(.A(\a[41] ), .B(new_n16670), .Y(new_n16671));
  INVx1_ASAP7_75t_L         g16415(.A(new_n16568), .Y(new_n16672));
  AOI22xp33_ASAP7_75t_L     g16416(.A1(new_n6002), .A2(\b[41] ), .B1(new_n5999), .B2(new_n5669), .Y(new_n16673));
  OAI221xp5_ASAP7_75t_L     g16417(.A1(new_n6544), .A2(new_n5186), .B1(new_n5166), .B2(new_n6309), .C(new_n16673), .Y(new_n16674));
  XNOR2x2_ASAP7_75t_L       g16418(.A(\a[44] ), .B(new_n16674), .Y(new_n16675));
  A2O1A1O1Ixp25_ASAP7_75t_L g16419(.A1(new_n16228), .A2(new_n16227), .B(new_n16385), .C(new_n16391), .D(new_n16562), .Y(new_n16676));
  INVx1_ASAP7_75t_L         g16420(.A(new_n16562), .Y(new_n16677));
  NOR2xp33_ASAP7_75t_L      g16421(.A(new_n16563), .B(new_n16677), .Y(new_n16678));
  INVx1_ASAP7_75t_L         g16422(.A(new_n16678), .Y(new_n16679));
  AOI22xp33_ASAP7_75t_L     g16423(.A1(new_n6822), .A2(\b[38] ), .B1(new_n6819), .B2(new_n4923), .Y(new_n16680));
  OAI221xp5_ASAP7_75t_L     g16424(.A1(new_n7392), .A2(new_n4701), .B1(new_n4465), .B2(new_n7115), .C(new_n16680), .Y(new_n16681));
  XNOR2x2_ASAP7_75t_L       g16425(.A(\a[47] ), .B(new_n16681), .Y(new_n16682));
  AOI22xp33_ASAP7_75t_L     g16426(.A1(new_n7659), .A2(\b[35] ), .B1(new_n7656), .B2(new_n5649), .Y(new_n16683));
  OAI221xp5_ASAP7_75t_L     g16427(.A1(new_n8326), .A2(new_n3827), .B1(new_n3807), .B2(new_n7994), .C(new_n16683), .Y(new_n16684));
  XNOR2x2_ASAP7_75t_L       g16428(.A(\a[50] ), .B(new_n16684), .Y(new_n16685));
  INVx1_ASAP7_75t_L         g16429(.A(new_n16685), .Y(new_n16686));
  AOI22xp33_ASAP7_75t_L     g16430(.A1(new_n8645), .A2(\b[32] ), .B1(new_n8642), .B2(new_n3450), .Y(new_n16687));
  OAI221xp5_ASAP7_75t_L     g16431(.A1(new_n9322), .A2(new_n3419), .B1(new_n3212), .B2(new_n8965), .C(new_n16687), .Y(new_n16688));
  XNOR2x2_ASAP7_75t_L       g16432(.A(\a[53] ), .B(new_n16688), .Y(new_n16689));
  AOI22xp33_ASAP7_75t_L     g16433(.A1(new_n10594), .A2(\b[26] ), .B1(new_n10591), .B2(new_n2888), .Y(new_n16690));
  OAI221xp5_ASAP7_75t_L     g16434(.A1(new_n11335), .A2(new_n2180), .B1(new_n2019), .B2(new_n11330), .C(new_n16690), .Y(new_n16691));
  XNOR2x2_ASAP7_75t_L       g16435(.A(\a[59] ), .B(new_n16691), .Y(new_n16692));
  INVx1_ASAP7_75t_L         g16436(.A(new_n16692), .Y(new_n16693));
  NOR2xp33_ASAP7_75t_L      g16437(.A(new_n1493), .B(new_n12671), .Y(new_n16694));
  O2A1O1Ixp33_ASAP7_75t_L   g16438(.A1(new_n12353), .A2(new_n12355), .B(\b[20] ), .C(new_n16694), .Y(new_n16695));
  A2O1A1Ixp33_ASAP7_75t_L   g16439(.A1(new_n12669), .A2(\b[19] ), .B(new_n16508), .C(new_n16695), .Y(new_n16696));
  A2O1A1Ixp33_ASAP7_75t_L   g16440(.A1(\b[20] ), .A2(new_n12669), .B(new_n16694), .C(new_n16512), .Y(new_n16697));
  NAND2xp33_ASAP7_75t_L     g16441(.A(new_n16697), .B(new_n16696), .Y(new_n16698));
  AOI22xp33_ASAP7_75t_L     g16442(.A1(new_n11647), .A2(\b[22] ), .B1(\b[23] ), .B2(new_n11656), .Y(new_n16699));
  OAI221xp5_ASAP7_75t_L     g16443(.A1(new_n13003), .A2(new_n1709), .B1(new_n12022), .B2(new_n4860), .C(new_n16699), .Y(new_n16700));
  XNOR2x2_ASAP7_75t_L       g16444(.A(\a[62] ), .B(new_n16700), .Y(new_n16701));
  NOR2xp33_ASAP7_75t_L      g16445(.A(new_n16698), .B(new_n16701), .Y(new_n16702));
  AND2x2_ASAP7_75t_L        g16446(.A(new_n16698), .B(new_n16701), .Y(new_n16703));
  NOR2xp33_ASAP7_75t_L      g16447(.A(new_n16702), .B(new_n16703), .Y(new_n16704));
  INVx1_ASAP7_75t_L         g16448(.A(new_n16704), .Y(new_n16705));
  O2A1O1Ixp33_ASAP7_75t_L   g16449(.A1(new_n16516), .A2(new_n16519), .B(new_n16515), .C(new_n16705), .Y(new_n16706));
  INVx1_ASAP7_75t_L         g16450(.A(new_n16706), .Y(new_n16707));
  A2O1A1O1Ixp25_ASAP7_75t_L g16451(.A1(new_n16343), .A2(new_n16347), .B(new_n16509), .C(new_n16512), .D(new_n16521), .Y(new_n16708));
  NAND2xp33_ASAP7_75t_L     g16452(.A(new_n16708), .B(new_n16705), .Y(new_n16709));
  NAND3xp33_ASAP7_75t_L     g16453(.A(new_n16707), .B(new_n16693), .C(new_n16709), .Y(new_n16710));
  AO21x2_ASAP7_75t_L        g16454(.A1(new_n16709), .A2(new_n16707), .B(new_n16693), .Y(new_n16711));
  AND2x2_ASAP7_75t_L        g16455(.A(new_n16710), .B(new_n16711), .Y(new_n16712));
  NAND3xp33_ASAP7_75t_L     g16456(.A(new_n16712), .B(new_n16531), .C(new_n16527), .Y(new_n16713));
  O2A1O1Ixp33_ASAP7_75t_L   g16457(.A1(new_n16523), .A2(new_n16524), .B(new_n16531), .C(new_n16712), .Y(new_n16714));
  INVx1_ASAP7_75t_L         g16458(.A(new_n16714), .Y(new_n16715));
  AOI22xp33_ASAP7_75t_L     g16459(.A1(new_n9623), .A2(\b[29] ), .B1(new_n9620), .B2(new_n5472), .Y(new_n16716));
  OAI221xp5_ASAP7_75t_L     g16460(.A1(new_n10280), .A2(new_n2852), .B1(new_n2650), .B2(new_n12010), .C(new_n16716), .Y(new_n16717));
  XNOR2x2_ASAP7_75t_L       g16461(.A(\a[56] ), .B(new_n16717), .Y(new_n16718));
  NAND3xp33_ASAP7_75t_L     g16462(.A(new_n16715), .B(new_n16713), .C(new_n16718), .Y(new_n16719));
  INVx1_ASAP7_75t_L         g16463(.A(new_n16719), .Y(new_n16720));
  AOI21xp33_ASAP7_75t_L     g16464(.A1(new_n16715), .A2(new_n16713), .B(new_n16718), .Y(new_n16721));
  NOR2xp33_ASAP7_75t_L      g16465(.A(new_n16721), .B(new_n16720), .Y(new_n16722));
  O2A1O1Ixp33_ASAP7_75t_L   g16466(.A1(new_n16507), .A2(new_n16533), .B(new_n16538), .C(new_n16722), .Y(new_n16723));
  A2O1A1Ixp33_ASAP7_75t_L   g16467(.A1(new_n16531), .A2(new_n16532), .B(new_n16507), .C(new_n16538), .Y(new_n16724));
  NOR3xp33_ASAP7_75t_L      g16468(.A(new_n16724), .B(new_n16721), .C(new_n16720), .Y(new_n16725));
  NOR2xp33_ASAP7_75t_L      g16469(.A(new_n16725), .B(new_n16723), .Y(new_n16726));
  NAND2xp33_ASAP7_75t_L     g16470(.A(new_n16689), .B(new_n16726), .Y(new_n16727));
  INVx1_ASAP7_75t_L         g16471(.A(new_n16689), .Y(new_n16728));
  OAI21xp33_ASAP7_75t_L     g16472(.A1(new_n16725), .A2(new_n16723), .B(new_n16728), .Y(new_n16729));
  AND2x2_ASAP7_75t_L        g16473(.A(new_n16729), .B(new_n16727), .Y(new_n16730));
  INVx1_ASAP7_75t_L         g16474(.A(new_n16730), .Y(new_n16731));
  AND2x2_ASAP7_75t_L        g16475(.A(new_n16542), .B(new_n16551), .Y(new_n16732));
  NAND2xp33_ASAP7_75t_L     g16476(.A(new_n16732), .B(new_n16731), .Y(new_n16733));
  INVx1_ASAP7_75t_L         g16477(.A(new_n16733), .Y(new_n16734));
  O2A1O1Ixp33_ASAP7_75t_L   g16478(.A1(new_n16543), .A2(new_n16549), .B(new_n16542), .C(new_n16731), .Y(new_n16735));
  NOR2xp33_ASAP7_75t_L      g16479(.A(new_n16735), .B(new_n16734), .Y(new_n16736));
  NAND2xp33_ASAP7_75t_L     g16480(.A(new_n16686), .B(new_n16736), .Y(new_n16737));
  OAI21xp33_ASAP7_75t_L     g16481(.A1(new_n16735), .A2(new_n16734), .B(new_n16685), .Y(new_n16738));
  NAND2xp33_ASAP7_75t_L     g16482(.A(new_n16738), .B(new_n16737), .Y(new_n16739));
  OAI21xp33_ASAP7_75t_L     g16483(.A1(new_n16553), .A2(new_n16554), .B(new_n16560), .Y(new_n16740));
  XNOR2x2_ASAP7_75t_L       g16484(.A(new_n16739), .B(new_n16740), .Y(new_n16741));
  XNOR2x2_ASAP7_75t_L       g16485(.A(new_n16682), .B(new_n16741), .Y(new_n16742));
  O2A1O1Ixp33_ASAP7_75t_L   g16486(.A1(new_n16676), .A2(new_n16567), .B(new_n16679), .C(new_n16742), .Y(new_n16743));
  OA21x2_ASAP7_75t_L        g16487(.A1(new_n16567), .A2(new_n16676), .B(new_n16679), .Y(new_n16744));
  AND2x2_ASAP7_75t_L        g16488(.A(new_n16744), .B(new_n16742), .Y(new_n16745));
  NOR3xp33_ASAP7_75t_L      g16489(.A(new_n16745), .B(new_n16743), .C(new_n16675), .Y(new_n16746));
  INVx1_ASAP7_75t_L         g16490(.A(new_n16746), .Y(new_n16747));
  OAI21xp33_ASAP7_75t_L     g16491(.A1(new_n16743), .A2(new_n16745), .B(new_n16675), .Y(new_n16748));
  NAND2xp33_ASAP7_75t_L     g16492(.A(new_n16748), .B(new_n16747), .Y(new_n16749));
  A2O1A1O1Ixp25_ASAP7_75t_L g16493(.A1(new_n16402), .A2(new_n16396), .B(new_n16672), .C(new_n16570), .D(new_n16749), .Y(new_n16750));
  A2O1A1Ixp33_ASAP7_75t_L   g16494(.A1(new_n16402), .A2(new_n16396), .B(new_n16672), .C(new_n16570), .Y(new_n16751));
  AOI21xp33_ASAP7_75t_L     g16495(.A1(new_n16748), .A2(new_n16747), .B(new_n16751), .Y(new_n16752));
  NOR3xp33_ASAP7_75t_L      g16496(.A(new_n16750), .B(new_n16752), .C(new_n16671), .Y(new_n16753));
  INVx1_ASAP7_75t_L         g16497(.A(new_n16671), .Y(new_n16754));
  NOR2xp33_ASAP7_75t_L      g16498(.A(new_n16752), .B(new_n16750), .Y(new_n16755));
  NOR2xp33_ASAP7_75t_L      g16499(.A(new_n16754), .B(new_n16755), .Y(new_n16756));
  NOR2xp33_ASAP7_75t_L      g16500(.A(new_n16581), .B(new_n16575), .Y(new_n16757));
  O2A1O1Ixp33_ASAP7_75t_L   g16501(.A1(new_n16571), .A2(new_n16572), .B(new_n16497), .C(new_n16757), .Y(new_n16758));
  INVx1_ASAP7_75t_L         g16502(.A(new_n16758), .Y(new_n16759));
  NOR3xp33_ASAP7_75t_L      g16503(.A(new_n16759), .B(new_n16756), .C(new_n16753), .Y(new_n16760));
  NOR2xp33_ASAP7_75t_L      g16504(.A(new_n16753), .B(new_n16756), .Y(new_n16761));
  O2A1O1Ixp33_ASAP7_75t_L   g16505(.A1(new_n16575), .A2(new_n16581), .B(new_n16574), .C(new_n16761), .Y(new_n16762));
  NOR2xp33_ASAP7_75t_L      g16506(.A(new_n16762), .B(new_n16760), .Y(new_n16763));
  AOI22xp33_ASAP7_75t_L     g16507(.A1(new_n4544), .A2(\b[47] ), .B1(new_n4542), .B2(new_n7323), .Y(new_n16764));
  OAI221xp5_ASAP7_75t_L     g16508(.A1(new_n4536), .A2(new_n7033), .B1(new_n6756), .B2(new_n4781), .C(new_n16764), .Y(new_n16765));
  XNOR2x2_ASAP7_75t_L       g16509(.A(\a[38] ), .B(new_n16765), .Y(new_n16766));
  XNOR2x2_ASAP7_75t_L       g16510(.A(new_n16766), .B(new_n16763), .Y(new_n16767));
  MAJx2_ASAP7_75t_L         g16511(.A(new_n16582), .B(new_n16583), .C(new_n16588), .Y(new_n16768));
  XNOR2x2_ASAP7_75t_L       g16512(.A(new_n16768), .B(new_n16767), .Y(new_n16769));
  AOI22xp33_ASAP7_75t_L     g16513(.A1(new_n3884), .A2(\b[50] ), .B1(new_n3881), .B2(new_n8235), .Y(new_n16770));
  OAI221xp5_ASAP7_75t_L     g16514(.A1(new_n4312), .A2(new_n7907), .B1(new_n7333), .B2(new_n4986), .C(new_n16770), .Y(new_n16771));
  XNOR2x2_ASAP7_75t_L       g16515(.A(\a[35] ), .B(new_n16771), .Y(new_n16772));
  INVx1_ASAP7_75t_L         g16516(.A(new_n16772), .Y(new_n16773));
  XNOR2x2_ASAP7_75t_L       g16517(.A(new_n16773), .B(new_n16769), .Y(new_n16774));
  XNOR2x2_ASAP7_75t_L       g16518(.A(new_n16774), .B(new_n16668), .Y(new_n16775));
  XNOR2x2_ASAP7_75t_L       g16519(.A(new_n16775), .B(new_n16663), .Y(new_n16776));
  XNOR2x2_ASAP7_75t_L       g16520(.A(new_n16658), .B(new_n16776), .Y(new_n16777));
  NAND2xp33_ASAP7_75t_L     g16521(.A(new_n16777), .B(new_n16651), .Y(new_n16778));
  INVx1_ASAP7_75t_L         g16522(.A(new_n16777), .Y(new_n16779));
  NAND2xp33_ASAP7_75t_L     g16523(.A(new_n16650), .B(new_n16779), .Y(new_n16780));
  NAND2xp33_ASAP7_75t_L     g16524(.A(new_n16778), .B(new_n16780), .Y(new_n16781));
  NOR2xp33_ASAP7_75t_L      g16525(.A(new_n16781), .B(new_n16644), .Y(new_n16782));
  INVx1_ASAP7_75t_L         g16526(.A(new_n16782), .Y(new_n16783));
  NAND2xp33_ASAP7_75t_L     g16527(.A(new_n16781), .B(new_n16644), .Y(new_n16784));
  NAND2xp33_ASAP7_75t_L     g16528(.A(new_n16784), .B(new_n16783), .Y(new_n16785));
  O2A1O1Ixp33_ASAP7_75t_L   g16529(.A1(new_n16617), .A2(new_n16618), .B(new_n16623), .C(new_n16785), .Y(new_n16786));
  AOI211xp5_ASAP7_75t_L     g16530(.A1(new_n16783), .A2(new_n16784), .B(new_n16622), .C(new_n16619), .Y(new_n16787));
  NOR2xp33_ASAP7_75t_L      g16531(.A(new_n16787), .B(new_n16786), .Y(new_n16788));
  A2O1A1Ixp33_ASAP7_75t_L   g16532(.A1(new_n16633), .A2(new_n16629), .B(new_n16626), .C(new_n16788), .Y(new_n16789));
  INVx1_ASAP7_75t_L         g16533(.A(new_n16789), .Y(new_n16790));
  INVx1_ASAP7_75t_L         g16534(.A(new_n16626), .Y(new_n16791));
  A2O1A1Ixp33_ASAP7_75t_L   g16535(.A1(new_n16463), .A2(new_n16459), .B(new_n16630), .C(new_n16791), .Y(new_n16792));
  NOR2xp33_ASAP7_75t_L      g16536(.A(new_n16788), .B(new_n16792), .Y(new_n16793));
  NOR2xp33_ASAP7_75t_L      g16537(.A(new_n16790), .B(new_n16793), .Y(\f[83] ));
  NOR2xp33_ASAP7_75t_L      g16538(.A(new_n16641), .B(new_n16782), .Y(new_n16795));
  INVx1_ASAP7_75t_L         g16539(.A(new_n16795), .Y(new_n16796));
  INVx1_ASAP7_75t_L         g16540(.A(new_n16778), .Y(new_n16797));
  NAND2xp33_ASAP7_75t_L     g16541(.A(\b[63] ), .B(new_n1766), .Y(new_n16798));
  A2O1A1Ixp33_ASAP7_75t_L   g16542(.A1(new_n12607), .A2(new_n12603), .B(new_n1771), .C(new_n16798), .Y(new_n16799));
  AOI221xp5_ASAP7_75t_L     g16543(.A1(\b[61] ), .A2(new_n1910), .B1(\b[62] ), .B2(new_n1770), .C(new_n16799), .Y(new_n16800));
  XNOR2x2_ASAP7_75t_L       g16544(.A(new_n1761), .B(new_n16800), .Y(new_n16801));
  A2O1A1Ixp33_ASAP7_75t_L   g16545(.A1(new_n16649), .A2(new_n16648), .B(new_n16797), .C(new_n16801), .Y(new_n16802));
  NAND2xp33_ASAP7_75t_L     g16546(.A(new_n16648), .B(new_n16649), .Y(new_n16803));
  INVx1_ASAP7_75t_L         g16547(.A(new_n16801), .Y(new_n16804));
  NAND3xp33_ASAP7_75t_L     g16548(.A(new_n16778), .B(new_n16803), .C(new_n16804), .Y(new_n16805));
  NAND2xp33_ASAP7_75t_L     g16549(.A(new_n16805), .B(new_n16802), .Y(new_n16806));
  AOI22xp33_ASAP7_75t_L     g16550(.A1(new_n2228), .A2(\b[60] ), .B1(new_n2226), .B2(new_n11234), .Y(new_n16807));
  OAI221xp5_ASAP7_75t_L     g16551(.A1(new_n2220), .A2(new_n10881), .B1(new_n10848), .B2(new_n2387), .C(new_n16807), .Y(new_n16808));
  XNOR2x2_ASAP7_75t_L       g16552(.A(\a[26] ), .B(new_n16808), .Y(new_n16809));
  INVx1_ASAP7_75t_L         g16553(.A(new_n16809), .Y(new_n16810));
  O2A1O1Ixp33_ASAP7_75t_L   g16554(.A1(new_n16658), .A2(new_n16776), .B(new_n16656), .C(new_n16810), .Y(new_n16811));
  OA211x2_ASAP7_75t_L       g16555(.A1(new_n16658), .A2(new_n16776), .B(new_n16810), .C(new_n16656), .Y(new_n16812));
  NOR2xp33_ASAP7_75t_L      g16556(.A(new_n16811), .B(new_n16812), .Y(new_n16813));
  INVx1_ASAP7_75t_L         g16557(.A(new_n16662), .Y(new_n16814));
  MAJIxp5_ASAP7_75t_L       g16558(.A(new_n16814), .B(new_n16661), .C(new_n16775), .Y(new_n16815));
  AOI22xp33_ASAP7_75t_L     g16559(.A1(new_n2702), .A2(\b[57] ), .B1(new_n2700), .B2(new_n10495), .Y(new_n16816));
  OAI221xp5_ASAP7_75t_L     g16560(.A1(new_n2694), .A2(new_n10178), .B1(new_n9534), .B2(new_n2932), .C(new_n16816), .Y(new_n16817));
  XNOR2x2_ASAP7_75t_L       g16561(.A(new_n2697), .B(new_n16817), .Y(new_n16818));
  XNOR2x2_ASAP7_75t_L       g16562(.A(new_n16818), .B(new_n16815), .Y(new_n16819));
  AOI22xp33_ASAP7_75t_L     g16563(.A1(new_n3256), .A2(\b[54] ), .B1(new_n3254), .B2(new_n9208), .Y(new_n16820));
  OAI221xp5_ASAP7_75t_L     g16564(.A1(new_n3248), .A2(new_n8882), .B1(new_n8569), .B2(new_n3492), .C(new_n16820), .Y(new_n16821));
  XNOR2x2_ASAP7_75t_L       g16565(.A(\a[32] ), .B(new_n16821), .Y(new_n16822));
  A2O1A1Ixp33_ASAP7_75t_L   g16566(.A1(new_n16593), .A2(new_n16596), .B(new_n16591), .C(new_n16666), .Y(new_n16823));
  AOI211xp5_ASAP7_75t_L     g16567(.A1(new_n16593), .A2(new_n16596), .B(new_n16666), .C(new_n16591), .Y(new_n16824));
  AOI21xp33_ASAP7_75t_L     g16568(.A1(new_n16774), .A2(new_n16823), .B(new_n16824), .Y(new_n16825));
  XNOR2x2_ASAP7_75t_L       g16569(.A(new_n16822), .B(new_n16825), .Y(new_n16826));
  MAJx2_ASAP7_75t_L         g16570(.A(new_n16767), .B(new_n16768), .C(new_n16773), .Y(new_n16827));
  AND2x2_ASAP7_75t_L        g16571(.A(new_n16766), .B(new_n16763), .Y(new_n16828));
  AOI22xp33_ASAP7_75t_L     g16572(.A1(new_n10594), .A2(\b[27] ), .B1(new_n10591), .B2(new_n2657), .Y(new_n16829));
  OAI221xp5_ASAP7_75t_L     g16573(.A1(new_n11335), .A2(new_n2477), .B1(new_n2180), .B2(new_n11330), .C(new_n16829), .Y(new_n16830));
  XNOR2x2_ASAP7_75t_L       g16574(.A(\a[59] ), .B(new_n16830), .Y(new_n16831));
  INVx1_ASAP7_75t_L         g16575(.A(new_n16831), .Y(new_n16832));
  NOR2xp33_ASAP7_75t_L      g16576(.A(new_n1594), .B(new_n12671), .Y(new_n16833));
  A2O1A1Ixp33_ASAP7_75t_L   g16577(.A1(new_n12669), .A2(\b[21] ), .B(new_n16833), .C(new_n1401), .Y(new_n16834));
  INVx1_ASAP7_75t_L         g16578(.A(new_n16834), .Y(new_n16835));
  O2A1O1Ixp33_ASAP7_75t_L   g16579(.A1(new_n12353), .A2(new_n12355), .B(\b[21] ), .C(new_n16833), .Y(new_n16836));
  NAND2xp33_ASAP7_75t_L     g16580(.A(\a[20] ), .B(new_n16836), .Y(new_n16837));
  INVx1_ASAP7_75t_L         g16581(.A(new_n16837), .Y(new_n16838));
  NOR2xp33_ASAP7_75t_L      g16582(.A(new_n16835), .B(new_n16838), .Y(new_n16839));
  XNOR2x2_ASAP7_75t_L       g16583(.A(new_n16695), .B(new_n16839), .Y(new_n16840));
  INVx1_ASAP7_75t_L         g16584(.A(new_n16840), .Y(new_n16841));
  AOI22xp33_ASAP7_75t_L     g16585(.A1(new_n11656), .A2(\b[24] ), .B1(new_n11654), .B2(new_n2027), .Y(new_n16842));
  OAI221xp5_ASAP7_75t_L     g16586(.A1(new_n12364), .A2(new_n1995), .B1(new_n1857), .B2(new_n13003), .C(new_n16842), .Y(new_n16843));
  XNOR2x2_ASAP7_75t_L       g16587(.A(\a[62] ), .B(new_n16843), .Y(new_n16844));
  XNOR2x2_ASAP7_75t_L       g16588(.A(new_n16841), .B(new_n16844), .Y(new_n16845));
  O2A1O1Ixp33_ASAP7_75t_L   g16589(.A1(new_n16698), .A2(new_n16701), .B(new_n16696), .C(new_n16845), .Y(new_n16846));
  A2O1A1O1Ixp25_ASAP7_75t_L g16590(.A1(new_n12669), .A2(\b[19] ), .B(new_n16508), .C(new_n16695), .D(new_n16702), .Y(new_n16847));
  AND2x2_ASAP7_75t_L        g16591(.A(new_n16847), .B(new_n16845), .Y(new_n16848));
  NOR2xp33_ASAP7_75t_L      g16592(.A(new_n16846), .B(new_n16848), .Y(new_n16849));
  XNOR2x2_ASAP7_75t_L       g16593(.A(new_n16832), .B(new_n16849), .Y(new_n16850));
  INVx1_ASAP7_75t_L         g16594(.A(new_n16850), .Y(new_n16851));
  A2O1A1Ixp33_ASAP7_75t_L   g16595(.A1(new_n16522), .A2(new_n16515), .B(new_n16705), .C(new_n16710), .Y(new_n16852));
  NOR2xp33_ASAP7_75t_L      g16596(.A(new_n16852), .B(new_n16851), .Y(new_n16853));
  O2A1O1Ixp33_ASAP7_75t_L   g16597(.A1(new_n16708), .A2(new_n16705), .B(new_n16710), .C(new_n16850), .Y(new_n16854));
  NOR2xp33_ASAP7_75t_L      g16598(.A(new_n16854), .B(new_n16853), .Y(new_n16855));
  AOI22xp33_ASAP7_75t_L     g16599(.A1(new_n9623), .A2(\b[30] ), .B1(new_n9620), .B2(new_n3219), .Y(new_n16856));
  OAI221xp5_ASAP7_75t_L     g16600(.A1(new_n10280), .A2(new_n2871), .B1(new_n2852), .B2(new_n12010), .C(new_n16856), .Y(new_n16857));
  XNOR2x2_ASAP7_75t_L       g16601(.A(\a[56] ), .B(new_n16857), .Y(new_n16858));
  INVx1_ASAP7_75t_L         g16602(.A(new_n16858), .Y(new_n16859));
  XNOR2x2_ASAP7_75t_L       g16603(.A(new_n16859), .B(new_n16855), .Y(new_n16860));
  A2O1A1Ixp33_ASAP7_75t_L   g16604(.A1(new_n16718), .A2(new_n16713), .B(new_n16714), .C(new_n16860), .Y(new_n16861));
  A2O1A1Ixp33_ASAP7_75t_L   g16605(.A1(new_n16531), .A2(new_n16527), .B(new_n16712), .C(new_n16719), .Y(new_n16862));
  OR2x4_ASAP7_75t_L         g16606(.A(new_n16862), .B(new_n16860), .Y(new_n16863));
  AND2x2_ASAP7_75t_L        g16607(.A(new_n16861), .B(new_n16863), .Y(new_n16864));
  AOI22xp33_ASAP7_75t_L     g16608(.A1(new_n8645), .A2(\b[33] ), .B1(new_n8642), .B2(new_n3813), .Y(new_n16865));
  OAI221xp5_ASAP7_75t_L     g16609(.A1(new_n9322), .A2(new_n3443), .B1(new_n3419), .B2(new_n8965), .C(new_n16865), .Y(new_n16866));
  XNOR2x2_ASAP7_75t_L       g16610(.A(\a[53] ), .B(new_n16866), .Y(new_n16867));
  INVx1_ASAP7_75t_L         g16611(.A(new_n16867), .Y(new_n16868));
  OAI311xp33_ASAP7_75t_L    g16612(.A1(new_n16724), .A2(new_n16721), .A3(new_n16720), .B1(new_n16868), .C1(new_n16727), .Y(new_n16869));
  A2O1A1Ixp33_ASAP7_75t_L   g16613(.A1(new_n16726), .A2(new_n16689), .B(new_n16725), .C(new_n16867), .Y(new_n16870));
  NAND2xp33_ASAP7_75t_L     g16614(.A(new_n16870), .B(new_n16869), .Y(new_n16871));
  XOR2x2_ASAP7_75t_L        g16615(.A(new_n16864), .B(new_n16871), .Y(new_n16872));
  AOI22xp33_ASAP7_75t_L     g16616(.A1(new_n7659), .A2(\b[36] ), .B1(new_n7656), .B2(new_n4473), .Y(new_n16873));
  OAI221xp5_ASAP7_75t_L     g16617(.A1(new_n8326), .A2(new_n4053), .B1(new_n3827), .B2(new_n7994), .C(new_n16873), .Y(new_n16874));
  XNOR2x2_ASAP7_75t_L       g16618(.A(\a[50] ), .B(new_n16874), .Y(new_n16875));
  NOR2xp33_ASAP7_75t_L      g16619(.A(new_n16875), .B(new_n16872), .Y(new_n16876));
  INVx1_ASAP7_75t_L         g16620(.A(new_n16876), .Y(new_n16877));
  NAND2xp33_ASAP7_75t_L     g16621(.A(new_n16875), .B(new_n16872), .Y(new_n16878));
  AND2x2_ASAP7_75t_L        g16622(.A(new_n16878), .B(new_n16877), .Y(new_n16879));
  INVx1_ASAP7_75t_L         g16623(.A(new_n16879), .Y(new_n16880));
  NAND3xp33_ASAP7_75t_L     g16624(.A(new_n16880), .B(new_n16737), .C(new_n16733), .Y(new_n16881));
  O2A1O1Ixp33_ASAP7_75t_L   g16625(.A1(new_n16685), .A2(new_n16735), .B(new_n16733), .C(new_n16880), .Y(new_n16882));
  INVx1_ASAP7_75t_L         g16626(.A(new_n16882), .Y(new_n16883));
  NAND2xp33_ASAP7_75t_L     g16627(.A(new_n16881), .B(new_n16883), .Y(new_n16884));
  AOI22xp33_ASAP7_75t_L     g16628(.A1(new_n6822), .A2(\b[39] ), .B1(new_n6819), .B2(new_n5174), .Y(new_n16885));
  OAI221xp5_ASAP7_75t_L     g16629(.A1(new_n7392), .A2(new_n4915), .B1(new_n4701), .B2(new_n7115), .C(new_n16885), .Y(new_n16886));
  XNOR2x2_ASAP7_75t_L       g16630(.A(\a[47] ), .B(new_n16886), .Y(new_n16887));
  XNOR2x2_ASAP7_75t_L       g16631(.A(new_n16887), .B(new_n16884), .Y(new_n16888));
  MAJIxp5_ASAP7_75t_L       g16632(.A(new_n16740), .B(new_n16682), .C(new_n16739), .Y(new_n16889));
  INVx1_ASAP7_75t_L         g16633(.A(new_n16889), .Y(new_n16890));
  NAND2xp33_ASAP7_75t_L     g16634(.A(new_n16890), .B(new_n16888), .Y(new_n16891));
  INVx1_ASAP7_75t_L         g16635(.A(new_n16888), .Y(new_n16892));
  NAND2xp33_ASAP7_75t_L     g16636(.A(new_n16889), .B(new_n16892), .Y(new_n16893));
  NAND2xp33_ASAP7_75t_L     g16637(.A(new_n16891), .B(new_n16893), .Y(new_n16894));
  AOI22xp33_ASAP7_75t_L     g16638(.A1(new_n6002), .A2(\b[42] ), .B1(new_n5999), .B2(new_n5688), .Y(new_n16895));
  OAI221xp5_ASAP7_75t_L     g16639(.A1(new_n6544), .A2(new_n5666), .B1(new_n5186), .B2(new_n6309), .C(new_n16895), .Y(new_n16896));
  XNOR2x2_ASAP7_75t_L       g16640(.A(\a[44] ), .B(new_n16896), .Y(new_n16897));
  XNOR2x2_ASAP7_75t_L       g16641(.A(new_n16897), .B(new_n16894), .Y(new_n16898));
  NOR2xp33_ASAP7_75t_L      g16642(.A(new_n16743), .B(new_n16746), .Y(new_n16899));
  NAND2xp33_ASAP7_75t_L     g16643(.A(new_n16899), .B(new_n16898), .Y(new_n16900));
  O2A1O1Ixp33_ASAP7_75t_L   g16644(.A1(new_n16744), .A2(new_n16742), .B(new_n16747), .C(new_n16898), .Y(new_n16901));
  INVx1_ASAP7_75t_L         g16645(.A(new_n16901), .Y(new_n16902));
  NAND2xp33_ASAP7_75t_L     g16646(.A(new_n16902), .B(new_n16900), .Y(new_n16903));
  AOI22xp33_ASAP7_75t_L     g16647(.A1(new_n5249), .A2(\b[45] ), .B1(new_n5247), .B2(new_n6764), .Y(new_n16904));
  OAI221xp5_ASAP7_75t_L     g16648(.A1(new_n5241), .A2(new_n6220), .B1(new_n6195), .B2(new_n5521), .C(new_n16904), .Y(new_n16905));
  XNOR2x2_ASAP7_75t_L       g16649(.A(\a[41] ), .B(new_n16905), .Y(new_n16906));
  XOR2x2_ASAP7_75t_L        g16650(.A(new_n16906), .B(new_n16903), .Y(new_n16907));
  OR3x1_ASAP7_75t_L         g16651(.A(new_n16907), .B(new_n16750), .C(new_n16753), .Y(new_n16908));
  A2O1A1Ixp33_ASAP7_75t_L   g16652(.A1(new_n16755), .A2(new_n16754), .B(new_n16750), .C(new_n16907), .Y(new_n16909));
  NAND2xp33_ASAP7_75t_L     g16653(.A(new_n16909), .B(new_n16908), .Y(new_n16910));
  AOI22xp33_ASAP7_75t_L     g16654(.A1(new_n4544), .A2(\b[48] ), .B1(new_n4542), .B2(new_n7341), .Y(new_n16911));
  OAI221xp5_ASAP7_75t_L     g16655(.A1(new_n4536), .A2(new_n7316), .B1(new_n7033), .B2(new_n4781), .C(new_n16911), .Y(new_n16912));
  XNOR2x2_ASAP7_75t_L       g16656(.A(\a[38] ), .B(new_n16912), .Y(new_n16913));
  XNOR2x2_ASAP7_75t_L       g16657(.A(new_n16913), .B(new_n16910), .Y(new_n16914));
  OA21x2_ASAP7_75t_L        g16658(.A1(new_n16762), .A2(new_n16828), .B(new_n16914), .Y(new_n16915));
  NOR3xp33_ASAP7_75t_L      g16659(.A(new_n16914), .B(new_n16828), .C(new_n16762), .Y(new_n16916));
  NOR2xp33_ASAP7_75t_L      g16660(.A(new_n16916), .B(new_n16915), .Y(new_n16917));
  AOI22xp33_ASAP7_75t_L     g16661(.A1(new_n3884), .A2(\b[51] ), .B1(new_n3881), .B2(new_n8257), .Y(new_n16918));
  OAI221xp5_ASAP7_75t_L     g16662(.A1(new_n4312), .A2(new_n8228), .B1(new_n7907), .B2(new_n4986), .C(new_n16918), .Y(new_n16919));
  XNOR2x2_ASAP7_75t_L       g16663(.A(new_n3878), .B(new_n16919), .Y(new_n16920));
  NAND2xp33_ASAP7_75t_L     g16664(.A(new_n16920), .B(new_n16917), .Y(new_n16921));
  OR2x4_ASAP7_75t_L         g16665(.A(new_n16920), .B(new_n16917), .Y(new_n16922));
  AO21x2_ASAP7_75t_L        g16666(.A1(new_n16921), .A2(new_n16922), .B(new_n16827), .Y(new_n16923));
  NAND3xp33_ASAP7_75t_L     g16667(.A(new_n16922), .B(new_n16921), .C(new_n16827), .Y(new_n16924));
  NAND2xp33_ASAP7_75t_L     g16668(.A(new_n16924), .B(new_n16923), .Y(new_n16925));
  NOR2xp33_ASAP7_75t_L      g16669(.A(new_n16826), .B(new_n16925), .Y(new_n16926));
  AND2x2_ASAP7_75t_L        g16670(.A(new_n16826), .B(new_n16925), .Y(new_n16927));
  NOR2xp33_ASAP7_75t_L      g16671(.A(new_n16926), .B(new_n16927), .Y(new_n16928));
  XNOR2x2_ASAP7_75t_L       g16672(.A(new_n16819), .B(new_n16928), .Y(new_n16929));
  AND2x2_ASAP7_75t_L        g16673(.A(new_n16813), .B(new_n16929), .Y(new_n16930));
  NOR2xp33_ASAP7_75t_L      g16674(.A(new_n16813), .B(new_n16929), .Y(new_n16931));
  NOR2xp33_ASAP7_75t_L      g16675(.A(new_n16931), .B(new_n16930), .Y(new_n16932));
  INVx1_ASAP7_75t_L         g16676(.A(new_n16932), .Y(new_n16933));
  XNOR2x2_ASAP7_75t_L       g16677(.A(new_n16933), .B(new_n16806), .Y(new_n16934));
  NOR2xp33_ASAP7_75t_L      g16678(.A(new_n16934), .B(new_n16796), .Y(new_n16935));
  INVx1_ASAP7_75t_L         g16679(.A(new_n16640), .Y(new_n16936));
  O2A1O1Ixp33_ASAP7_75t_L   g16680(.A1(new_n16605), .A2(new_n16606), .B(new_n16475), .C(new_n16472), .Y(new_n16937));
  A2O1A1Ixp33_ASAP7_75t_L   g16681(.A1(new_n16937), .A2(new_n16936), .B(new_n16782), .C(new_n16934), .Y(new_n16938));
  INVx1_ASAP7_75t_L         g16682(.A(new_n16938), .Y(new_n16939));
  NOR2xp33_ASAP7_75t_L      g16683(.A(new_n16935), .B(new_n16939), .Y(new_n16940));
  A2O1A1Ixp33_ASAP7_75t_L   g16684(.A1(new_n16792), .A2(new_n16788), .B(new_n16786), .C(new_n16940), .Y(new_n16941));
  INVx1_ASAP7_75t_L         g16685(.A(new_n16941), .Y(new_n16942));
  NOR3xp33_ASAP7_75t_L      g16686(.A(new_n16790), .B(new_n16940), .C(new_n16786), .Y(new_n16943));
  NOR2xp33_ASAP7_75t_L      g16687(.A(new_n16943), .B(new_n16942), .Y(\f[84] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g16688(.A1(new_n16629), .A2(new_n16633), .B(new_n16626), .C(new_n16788), .D(new_n16786), .Y(new_n16945));
  AOI22xp33_ASAP7_75t_L     g16689(.A1(new_n1770), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1910), .Y(new_n16946));
  A2O1A1Ixp33_ASAP7_75t_L   g16690(.A1(new_n13506), .A2(new_n13507), .B(new_n1771), .C(new_n16946), .Y(new_n16947));
  NOR2xp33_ASAP7_75t_L      g16691(.A(new_n1761), .B(new_n16947), .Y(new_n16948));
  A2O1A1O1Ixp25_ASAP7_75t_L g16692(.A1(new_n13507), .A2(new_n13506), .B(new_n1771), .C(new_n16946), .D(\a[23] ), .Y(new_n16949));
  NOR2xp33_ASAP7_75t_L      g16693(.A(new_n16949), .B(new_n16948), .Y(new_n16950));
  INVx1_ASAP7_75t_L         g16694(.A(new_n16950), .Y(new_n16951));
  A2O1A1Ixp33_ASAP7_75t_L   g16695(.A1(new_n16929), .A2(new_n16813), .B(new_n16812), .C(new_n16951), .Y(new_n16952));
  NOR2xp33_ASAP7_75t_L      g16696(.A(new_n16812), .B(new_n16930), .Y(new_n16953));
  NAND2xp33_ASAP7_75t_L     g16697(.A(new_n16950), .B(new_n16953), .Y(new_n16954));
  AND2x2_ASAP7_75t_L        g16698(.A(new_n16952), .B(new_n16954), .Y(new_n16955));
  INVx1_ASAP7_75t_L         g16699(.A(new_n16955), .Y(new_n16956));
  AOI22xp33_ASAP7_75t_L     g16700(.A1(new_n2228), .A2(\b[61] ), .B1(new_n2226), .B2(new_n11919), .Y(new_n16957));
  OAI221xp5_ASAP7_75t_L     g16701(.A1(new_n2220), .A2(new_n11226), .B1(new_n10881), .B2(new_n2387), .C(new_n16957), .Y(new_n16958));
  XNOR2x2_ASAP7_75t_L       g16702(.A(\a[26] ), .B(new_n16958), .Y(new_n16959));
  INVx1_ASAP7_75t_L         g16703(.A(new_n16959), .Y(new_n16960));
  MAJx2_ASAP7_75t_L         g16704(.A(new_n16928), .B(new_n16818), .C(new_n16815), .Y(new_n16961));
  NOR2xp33_ASAP7_75t_L      g16705(.A(new_n16960), .B(new_n16961), .Y(new_n16962));
  AND2x2_ASAP7_75t_L        g16706(.A(new_n16960), .B(new_n16961), .Y(new_n16963));
  NOR2xp33_ASAP7_75t_L      g16707(.A(new_n16962), .B(new_n16963), .Y(new_n16964));
  INVx1_ASAP7_75t_L         g16708(.A(new_n16964), .Y(new_n16965));
  NOR2xp33_ASAP7_75t_L      g16709(.A(new_n16822), .B(new_n16825), .Y(new_n16966));
  NOR2xp33_ASAP7_75t_L      g16710(.A(new_n16966), .B(new_n16926), .Y(new_n16967));
  AOI22xp33_ASAP7_75t_L     g16711(.A1(new_n2706), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n2702), .Y(new_n16968));
  OAI221xp5_ASAP7_75t_L     g16712(.A1(new_n2932), .A2(new_n10178), .B1(new_n2707), .B2(new_n10856), .C(new_n16968), .Y(new_n16969));
  XNOR2x2_ASAP7_75t_L       g16713(.A(\a[29] ), .B(new_n16969), .Y(new_n16970));
  XNOR2x2_ASAP7_75t_L       g16714(.A(new_n16970), .B(new_n16967), .Y(new_n16971));
  AOI22xp33_ASAP7_75t_L     g16715(.A1(new_n3256), .A2(\b[55] ), .B1(new_n3254), .B2(new_n9542), .Y(new_n16972));
  OAI221xp5_ASAP7_75t_L     g16716(.A1(new_n3248), .A2(new_n9199), .B1(new_n8882), .B2(new_n3492), .C(new_n16972), .Y(new_n16973));
  XNOR2x2_ASAP7_75t_L       g16717(.A(\a[32] ), .B(new_n16973), .Y(new_n16974));
  INVx1_ASAP7_75t_L         g16718(.A(new_n16974), .Y(new_n16975));
  NAND2xp33_ASAP7_75t_L     g16719(.A(new_n16921), .B(new_n16924), .Y(new_n16976));
  XNOR2x2_ASAP7_75t_L       g16720(.A(new_n16975), .B(new_n16976), .Y(new_n16977));
  OAI21xp33_ASAP7_75t_L     g16721(.A1(new_n16884), .A2(new_n16887), .B(new_n16893), .Y(new_n16978));
  AOI22xp33_ASAP7_75t_L     g16722(.A1(new_n6822), .A2(\b[40] ), .B1(new_n6819), .B2(new_n5194), .Y(new_n16979));
  OAI221xp5_ASAP7_75t_L     g16723(.A1(new_n7392), .A2(new_n5166), .B1(new_n4915), .B2(new_n7115), .C(new_n16979), .Y(new_n16980));
  XNOR2x2_ASAP7_75t_L       g16724(.A(\a[47] ), .B(new_n16980), .Y(new_n16981));
  INVx1_ASAP7_75t_L         g16725(.A(new_n16981), .Y(new_n16982));
  AOI22xp33_ASAP7_75t_L     g16726(.A1(new_n10594), .A2(\b[28] ), .B1(new_n10591), .B2(new_n2858), .Y(new_n16983));
  OAI221xp5_ASAP7_75t_L     g16727(.A1(new_n11335), .A2(new_n2650), .B1(new_n2477), .B2(new_n11330), .C(new_n16983), .Y(new_n16984));
  XNOR2x2_ASAP7_75t_L       g16728(.A(\a[59] ), .B(new_n16984), .Y(new_n16985));
  INVx1_ASAP7_75t_L         g16729(.A(new_n16985), .Y(new_n16986));
  INVx1_ASAP7_75t_L         g16730(.A(new_n16845), .Y(new_n16987));
  A2O1A1Ixp33_ASAP7_75t_L   g16731(.A1(new_n16695), .A2(new_n16513), .B(new_n16702), .C(new_n16987), .Y(new_n16988));
  NOR2xp33_ASAP7_75t_L      g16732(.A(new_n1709), .B(new_n12671), .Y(new_n16989));
  A2O1A1O1Ixp25_ASAP7_75t_L g16733(.A1(new_n12669), .A2(\b[20] ), .B(new_n16694), .C(new_n16837), .D(new_n16835), .Y(new_n16990));
  A2O1A1Ixp33_ASAP7_75t_L   g16734(.A1(new_n12669), .A2(\b[22] ), .B(new_n16989), .C(new_n16990), .Y(new_n16991));
  O2A1O1Ixp33_ASAP7_75t_L   g16735(.A1(new_n12353), .A2(new_n12355), .B(\b[22] ), .C(new_n16989), .Y(new_n16992));
  INVx1_ASAP7_75t_L         g16736(.A(new_n16992), .Y(new_n16993));
  O2A1O1Ixp33_ASAP7_75t_L   g16737(.A1(new_n16695), .A2(new_n16838), .B(new_n16834), .C(new_n16993), .Y(new_n16994));
  INVx1_ASAP7_75t_L         g16738(.A(new_n16994), .Y(new_n16995));
  NAND2xp33_ASAP7_75t_L     g16739(.A(new_n16991), .B(new_n16995), .Y(new_n16996));
  AOI22xp33_ASAP7_75t_L     g16740(.A1(new_n11647), .A2(\b[24] ), .B1(\b[25] ), .B2(new_n11656), .Y(new_n16997));
  OAI221xp5_ASAP7_75t_L     g16741(.A1(new_n13003), .A2(new_n1995), .B1(new_n12022), .B2(new_n2187), .C(new_n16997), .Y(new_n16998));
  XNOR2x2_ASAP7_75t_L       g16742(.A(\a[62] ), .B(new_n16998), .Y(new_n16999));
  NOR2xp33_ASAP7_75t_L      g16743(.A(new_n16996), .B(new_n16999), .Y(new_n17000));
  INVx1_ASAP7_75t_L         g16744(.A(new_n17000), .Y(new_n17001));
  NAND2xp33_ASAP7_75t_L     g16745(.A(new_n16996), .B(new_n16999), .Y(new_n17002));
  AND2x2_ASAP7_75t_L        g16746(.A(new_n17002), .B(new_n17001), .Y(new_n17003));
  INVx1_ASAP7_75t_L         g16747(.A(new_n17003), .Y(new_n17004));
  O2A1O1Ixp33_ASAP7_75t_L   g16748(.A1(new_n16841), .A2(new_n16844), .B(new_n16988), .C(new_n17004), .Y(new_n17005));
  OA211x2_ASAP7_75t_L       g16749(.A1(new_n16841), .A2(new_n16844), .B(new_n16988), .C(new_n17004), .Y(new_n17006));
  NOR2xp33_ASAP7_75t_L      g16750(.A(new_n17005), .B(new_n17006), .Y(new_n17007));
  NAND2xp33_ASAP7_75t_L     g16751(.A(new_n16986), .B(new_n17007), .Y(new_n17008));
  OAI21xp33_ASAP7_75t_L     g16752(.A1(new_n17005), .A2(new_n17006), .B(new_n16985), .Y(new_n17009));
  AND2x2_ASAP7_75t_L        g16753(.A(new_n17009), .B(new_n17008), .Y(new_n17010));
  A2O1A1Ixp33_ASAP7_75t_L   g16754(.A1(new_n16849), .A2(new_n16832), .B(new_n16854), .C(new_n17010), .Y(new_n17011));
  NAND2xp33_ASAP7_75t_L     g16755(.A(new_n16832), .B(new_n16849), .Y(new_n17012));
  A2O1A1Ixp33_ASAP7_75t_L   g16756(.A1(new_n16710), .A2(new_n16707), .B(new_n16850), .C(new_n17012), .Y(new_n17013));
  NOR2xp33_ASAP7_75t_L      g16757(.A(new_n17013), .B(new_n17010), .Y(new_n17014));
  INVx1_ASAP7_75t_L         g16758(.A(new_n17014), .Y(new_n17015));
  AOI22xp33_ASAP7_75t_L     g16759(.A1(new_n9623), .A2(\b[31] ), .B1(new_n9620), .B2(new_n3426), .Y(new_n17016));
  OAI221xp5_ASAP7_75t_L     g16760(.A1(new_n10280), .A2(new_n3212), .B1(new_n2871), .B2(new_n12010), .C(new_n17016), .Y(new_n17017));
  XNOR2x2_ASAP7_75t_L       g16761(.A(\a[56] ), .B(new_n17017), .Y(new_n17018));
  NAND3xp33_ASAP7_75t_L     g16762(.A(new_n17015), .B(new_n17011), .C(new_n17018), .Y(new_n17019));
  INVx1_ASAP7_75t_L         g16763(.A(new_n17019), .Y(new_n17020));
  AOI21xp33_ASAP7_75t_L     g16764(.A1(new_n17015), .A2(new_n17011), .B(new_n17018), .Y(new_n17021));
  NOR2xp33_ASAP7_75t_L      g16765(.A(new_n17021), .B(new_n17020), .Y(new_n17022));
  NAND2xp33_ASAP7_75t_L     g16766(.A(new_n16859), .B(new_n16855), .Y(new_n17023));
  AND2x2_ASAP7_75t_L        g16767(.A(new_n17023), .B(new_n16863), .Y(new_n17024));
  NAND2xp33_ASAP7_75t_L     g16768(.A(new_n17022), .B(new_n17024), .Y(new_n17025));
  INVx1_ASAP7_75t_L         g16769(.A(new_n17025), .Y(new_n17026));
  O2A1O1Ixp33_ASAP7_75t_L   g16770(.A1(new_n16862), .A2(new_n16860), .B(new_n17023), .C(new_n17022), .Y(new_n17027));
  NOR2xp33_ASAP7_75t_L      g16771(.A(new_n17027), .B(new_n17026), .Y(new_n17028));
  AOI22xp33_ASAP7_75t_L     g16772(.A1(new_n8645), .A2(\b[34] ), .B1(new_n8642), .B2(new_n3833), .Y(new_n17029));
  OAI221xp5_ASAP7_75t_L     g16773(.A1(new_n9322), .A2(new_n3807), .B1(new_n3443), .B2(new_n8965), .C(new_n17029), .Y(new_n17030));
  XNOR2x2_ASAP7_75t_L       g16774(.A(\a[53] ), .B(new_n17030), .Y(new_n17031));
  NAND2xp33_ASAP7_75t_L     g16775(.A(new_n17031), .B(new_n17028), .Y(new_n17032));
  INVx1_ASAP7_75t_L         g16776(.A(new_n17031), .Y(new_n17033));
  OAI21xp33_ASAP7_75t_L     g16777(.A1(new_n17027), .A2(new_n17026), .B(new_n17033), .Y(new_n17034));
  AND2x2_ASAP7_75t_L        g16778(.A(new_n17034), .B(new_n17032), .Y(new_n17035));
  INVx1_ASAP7_75t_L         g16779(.A(new_n17035), .Y(new_n17036));
  O2A1O1Ixp33_ASAP7_75t_L   g16780(.A1(new_n16864), .A2(new_n16871), .B(new_n16870), .C(new_n17036), .Y(new_n17037));
  A2O1A1Ixp33_ASAP7_75t_L   g16781(.A1(new_n16861), .A2(new_n16863), .B(new_n16871), .C(new_n16870), .Y(new_n17038));
  NOR2xp33_ASAP7_75t_L      g16782(.A(new_n17038), .B(new_n17035), .Y(new_n17039));
  NOR2xp33_ASAP7_75t_L      g16783(.A(new_n17039), .B(new_n17037), .Y(new_n17040));
  INVx1_ASAP7_75t_L         g16784(.A(new_n17040), .Y(new_n17041));
  AOI22xp33_ASAP7_75t_L     g16785(.A1(new_n7659), .A2(\b[37] ), .B1(new_n7656), .B2(new_n4709), .Y(new_n17042));
  OAI221xp5_ASAP7_75t_L     g16786(.A1(new_n8326), .A2(new_n4465), .B1(new_n4053), .B2(new_n7994), .C(new_n17042), .Y(new_n17043));
  XNOR2x2_ASAP7_75t_L       g16787(.A(\a[50] ), .B(new_n17043), .Y(new_n17044));
  AND2x2_ASAP7_75t_L        g16788(.A(new_n17044), .B(new_n17041), .Y(new_n17045));
  NOR2xp33_ASAP7_75t_L      g16789(.A(new_n17044), .B(new_n17041), .Y(new_n17046));
  NOR2xp33_ASAP7_75t_L      g16790(.A(new_n17046), .B(new_n17045), .Y(new_n17047));
  INVx1_ASAP7_75t_L         g16791(.A(new_n17047), .Y(new_n17048));
  O2A1O1Ixp33_ASAP7_75t_L   g16792(.A1(new_n16872), .A2(new_n16875), .B(new_n16883), .C(new_n17048), .Y(new_n17049));
  NOR3xp33_ASAP7_75t_L      g16793(.A(new_n17047), .B(new_n16882), .C(new_n16876), .Y(new_n17050));
  NOR2xp33_ASAP7_75t_L      g16794(.A(new_n17050), .B(new_n17049), .Y(new_n17051));
  NAND2xp33_ASAP7_75t_L     g16795(.A(new_n16982), .B(new_n17051), .Y(new_n17052));
  INVx1_ASAP7_75t_L         g16796(.A(new_n17052), .Y(new_n17053));
  NOR2xp33_ASAP7_75t_L      g16797(.A(new_n16982), .B(new_n17051), .Y(new_n17054));
  NOR2xp33_ASAP7_75t_L      g16798(.A(new_n17053), .B(new_n17054), .Y(new_n17055));
  XNOR2x2_ASAP7_75t_L       g16799(.A(new_n16978), .B(new_n17055), .Y(new_n17056));
  NAND2xp33_ASAP7_75t_L     g16800(.A(\b[43] ), .B(new_n6002), .Y(new_n17057));
  OAI221xp5_ASAP7_75t_L     g16801(.A1(new_n5680), .A2(new_n6544), .B1(new_n6311), .B2(new_n9799), .C(new_n17057), .Y(new_n17058));
  AOI21xp33_ASAP7_75t_L     g16802(.A1(new_n6308), .A2(\b[41] ), .B(new_n17058), .Y(new_n17059));
  NAND2xp33_ASAP7_75t_L     g16803(.A(\a[44] ), .B(new_n17059), .Y(new_n17060));
  A2O1A1Ixp33_ASAP7_75t_L   g16804(.A1(\b[41] ), .A2(new_n6308), .B(new_n17058), .C(new_n5996), .Y(new_n17061));
  NAND2xp33_ASAP7_75t_L     g16805(.A(new_n17061), .B(new_n17060), .Y(new_n17062));
  XOR2x2_ASAP7_75t_L        g16806(.A(new_n17062), .B(new_n17056), .Y(new_n17063));
  OA21x2_ASAP7_75t_L        g16807(.A1(new_n16894), .A2(new_n16897), .B(new_n16902), .Y(new_n17064));
  NAND2xp33_ASAP7_75t_L     g16808(.A(new_n17064), .B(new_n17063), .Y(new_n17065));
  OR2x4_ASAP7_75t_L         g16809(.A(new_n17064), .B(new_n17063), .Y(new_n17066));
  AOI22xp33_ASAP7_75t_L     g16810(.A1(new_n5249), .A2(\b[46] ), .B1(new_n5247), .B2(new_n7041), .Y(new_n17067));
  OAI221xp5_ASAP7_75t_L     g16811(.A1(new_n5241), .A2(new_n6756), .B1(new_n6220), .B2(new_n5521), .C(new_n17067), .Y(new_n17068));
  XNOR2x2_ASAP7_75t_L       g16812(.A(\a[41] ), .B(new_n17068), .Y(new_n17069));
  NAND3xp33_ASAP7_75t_L     g16813(.A(new_n17066), .B(new_n17065), .C(new_n17069), .Y(new_n17070));
  INVx1_ASAP7_75t_L         g16814(.A(new_n17070), .Y(new_n17071));
  AOI21xp33_ASAP7_75t_L     g16815(.A1(new_n17066), .A2(new_n17065), .B(new_n17069), .Y(new_n17072));
  NOR2xp33_ASAP7_75t_L      g16816(.A(new_n17071), .B(new_n17072), .Y(new_n17073));
  NOR2xp33_ASAP7_75t_L      g16817(.A(new_n16906), .B(new_n16903), .Y(new_n17074));
  O2A1O1Ixp33_ASAP7_75t_L   g16818(.A1(new_n16750), .A2(new_n16753), .B(new_n16907), .C(new_n17074), .Y(new_n17075));
  NAND2xp33_ASAP7_75t_L     g16819(.A(new_n17075), .B(new_n17073), .Y(new_n17076));
  INVx1_ASAP7_75t_L         g16820(.A(new_n17076), .Y(new_n17077));
  O2A1O1Ixp33_ASAP7_75t_L   g16821(.A1(new_n16903), .A2(new_n16906), .B(new_n16909), .C(new_n17073), .Y(new_n17078));
  NOR2xp33_ASAP7_75t_L      g16822(.A(new_n17077), .B(new_n17078), .Y(new_n17079));
  AOI22xp33_ASAP7_75t_L     g16823(.A1(new_n4544), .A2(\b[49] ), .B1(new_n4542), .B2(new_n7914), .Y(new_n17080));
  OAI221xp5_ASAP7_75t_L     g16824(.A1(new_n4536), .A2(new_n7333), .B1(new_n7316), .B2(new_n4781), .C(new_n17080), .Y(new_n17081));
  XNOR2x2_ASAP7_75t_L       g16825(.A(\a[38] ), .B(new_n17081), .Y(new_n17082));
  NAND2xp33_ASAP7_75t_L     g16826(.A(new_n17082), .B(new_n17079), .Y(new_n17083));
  INVx1_ASAP7_75t_L         g16827(.A(new_n17082), .Y(new_n17084));
  OAI21xp33_ASAP7_75t_L     g16828(.A1(new_n17078), .A2(new_n17077), .B(new_n17084), .Y(new_n17085));
  INVx1_ASAP7_75t_L         g16829(.A(new_n16910), .Y(new_n17086));
  INVx1_ASAP7_75t_L         g16830(.A(new_n16913), .Y(new_n17087));
  AOI21xp33_ASAP7_75t_L     g16831(.A1(new_n17087), .A2(new_n17086), .B(new_n16916), .Y(new_n17088));
  NAND3xp33_ASAP7_75t_L     g16832(.A(new_n17088), .B(new_n17085), .C(new_n17083), .Y(new_n17089));
  NAND2xp33_ASAP7_75t_L     g16833(.A(new_n17085), .B(new_n17083), .Y(new_n17090));
  A2O1A1Ixp33_ASAP7_75t_L   g16834(.A1(new_n17087), .A2(new_n17086), .B(new_n16916), .C(new_n17090), .Y(new_n17091));
  AOI22xp33_ASAP7_75t_L     g16835(.A1(new_n3884), .A2(\b[52] ), .B1(new_n3881), .B2(new_n8577), .Y(new_n17092));
  OAI221xp5_ASAP7_75t_L     g16836(.A1(new_n4312), .A2(new_n8249), .B1(new_n8228), .B2(new_n4986), .C(new_n17092), .Y(new_n17093));
  XNOR2x2_ASAP7_75t_L       g16837(.A(\a[35] ), .B(new_n17093), .Y(new_n17094));
  AND3x1_ASAP7_75t_L        g16838(.A(new_n17091), .B(new_n17094), .C(new_n17089), .Y(new_n17095));
  AOI21xp33_ASAP7_75t_L     g16839(.A1(new_n17091), .A2(new_n17089), .B(new_n17094), .Y(new_n17096));
  NOR2xp33_ASAP7_75t_L      g16840(.A(new_n17096), .B(new_n17095), .Y(new_n17097));
  NOR2xp33_ASAP7_75t_L      g16841(.A(new_n17097), .B(new_n16977), .Y(new_n17098));
  AND2x2_ASAP7_75t_L        g16842(.A(new_n17097), .B(new_n16977), .Y(new_n17099));
  NOR2xp33_ASAP7_75t_L      g16843(.A(new_n17098), .B(new_n17099), .Y(new_n17100));
  XOR2x2_ASAP7_75t_L        g16844(.A(new_n16971), .B(new_n17100), .Y(new_n17101));
  NOR2xp33_ASAP7_75t_L      g16845(.A(new_n17101), .B(new_n16965), .Y(new_n17102));
  INVx1_ASAP7_75t_L         g16846(.A(new_n17102), .Y(new_n17103));
  NAND2xp33_ASAP7_75t_L     g16847(.A(new_n17101), .B(new_n16965), .Y(new_n17104));
  AOI21xp33_ASAP7_75t_L     g16848(.A1(new_n17104), .A2(new_n17103), .B(new_n16956), .Y(new_n17105));
  AND3x1_ASAP7_75t_L        g16849(.A(new_n16956), .B(new_n17104), .C(new_n17103), .Y(new_n17106));
  A2O1A1Ixp33_ASAP7_75t_L   g16850(.A1(new_n16649), .A2(new_n16648), .B(new_n16797), .C(new_n16804), .Y(new_n17107));
  A2O1A1Ixp33_ASAP7_75t_L   g16851(.A1(new_n16805), .A2(new_n16802), .B(new_n16933), .C(new_n17107), .Y(new_n17108));
  NOR3xp33_ASAP7_75t_L      g16852(.A(new_n17106), .B(new_n17108), .C(new_n17105), .Y(new_n17109));
  INVx1_ASAP7_75t_L         g16853(.A(new_n16806), .Y(new_n17110));
  NOR2xp33_ASAP7_75t_L      g16854(.A(new_n17105), .B(new_n17106), .Y(new_n17111));
  O2A1O1Ixp33_ASAP7_75t_L   g16855(.A1(new_n16933), .A2(new_n17110), .B(new_n17107), .C(new_n17111), .Y(new_n17112));
  NOR2xp33_ASAP7_75t_L      g16856(.A(new_n17109), .B(new_n17112), .Y(new_n17113));
  INVx1_ASAP7_75t_L         g16857(.A(new_n17113), .Y(new_n17114));
  O2A1O1Ixp33_ASAP7_75t_L   g16858(.A1(new_n16935), .A2(new_n16945), .B(new_n16938), .C(new_n17114), .Y(new_n17115));
  INVx1_ASAP7_75t_L         g16859(.A(new_n16786), .Y(new_n17116));
  A2O1A1Ixp33_ASAP7_75t_L   g16860(.A1(new_n16789), .A2(new_n17116), .B(new_n16935), .C(new_n16938), .Y(new_n17117));
  NOR2xp33_ASAP7_75t_L      g16861(.A(new_n17113), .B(new_n17117), .Y(new_n17118));
  NOR2xp33_ASAP7_75t_L      g16862(.A(new_n17118), .B(new_n17115), .Y(\f[85] ));
  INVx1_ASAP7_75t_L         g16863(.A(new_n16963), .Y(new_n17120));
  A2O1A1Ixp33_ASAP7_75t_L   g16864(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n1764), .Y(new_n17121));
  A2O1A1Ixp33_ASAP7_75t_L   g16865(.A1(new_n17121), .A2(new_n1911), .B(new_n12599), .C(\a[23] ), .Y(new_n17122));
  O2A1O1Ixp33_ASAP7_75t_L   g16866(.A1(new_n1771), .A2(new_n13934), .B(new_n1911), .C(new_n12599), .Y(new_n17123));
  NAND2xp33_ASAP7_75t_L     g16867(.A(new_n1761), .B(new_n17123), .Y(new_n17124));
  AND2x2_ASAP7_75t_L        g16868(.A(new_n17124), .B(new_n17122), .Y(new_n17125));
  O2A1O1Ixp33_ASAP7_75t_L   g16869(.A1(new_n16962), .A2(new_n17101), .B(new_n17120), .C(new_n17125), .Y(new_n17126));
  INVx1_ASAP7_75t_L         g16870(.A(new_n17126), .Y(new_n17127));
  NAND3xp33_ASAP7_75t_L     g16871(.A(new_n17103), .B(new_n17120), .C(new_n17125), .Y(new_n17128));
  NAND2xp33_ASAP7_75t_L     g16872(.A(new_n17127), .B(new_n17128), .Y(new_n17129));
  AOI22xp33_ASAP7_75t_L     g16873(.A1(new_n2228), .A2(\b[62] ), .B1(new_n2226), .B2(new_n12280), .Y(new_n17130));
  OAI221xp5_ASAP7_75t_L     g16874(.A1(new_n2220), .A2(new_n11911), .B1(new_n11226), .B2(new_n2387), .C(new_n17130), .Y(new_n17131));
  XNOR2x2_ASAP7_75t_L       g16875(.A(\a[26] ), .B(new_n17131), .Y(new_n17132));
  INVx1_ASAP7_75t_L         g16876(.A(new_n16970), .Y(new_n17133));
  NOR3xp33_ASAP7_75t_L      g16877(.A(new_n16971), .B(new_n17098), .C(new_n17099), .Y(new_n17134));
  O2A1O1Ixp33_ASAP7_75t_L   g16878(.A1(new_n16966), .A2(new_n16926), .B(new_n17133), .C(new_n17134), .Y(new_n17135));
  AND2x2_ASAP7_75t_L        g16879(.A(new_n17132), .B(new_n17135), .Y(new_n17136));
  NOR2xp33_ASAP7_75t_L      g16880(.A(new_n17132), .B(new_n17135), .Y(new_n17137));
  AOI22xp33_ASAP7_75t_L     g16881(.A1(new_n2702), .A2(\b[59] ), .B1(new_n2700), .B2(new_n10887), .Y(new_n17138));
  OAI221xp5_ASAP7_75t_L     g16882(.A1(new_n2694), .A2(new_n10848), .B1(new_n10488), .B2(new_n2932), .C(new_n17138), .Y(new_n17139));
  XNOR2x2_ASAP7_75t_L       g16883(.A(\a[29] ), .B(new_n17139), .Y(new_n17140));
  AOI21xp33_ASAP7_75t_L     g16884(.A1(new_n16976), .A2(new_n16975), .B(new_n17098), .Y(new_n17141));
  XNOR2x2_ASAP7_75t_L       g16885(.A(new_n17140), .B(new_n17141), .Y(new_n17142));
  AOI22xp33_ASAP7_75t_L     g16886(.A1(new_n3256), .A2(\b[56] ), .B1(new_n3254), .B2(new_n10185), .Y(new_n17143));
  OAI221xp5_ASAP7_75t_L     g16887(.A1(new_n3248), .A2(new_n9534), .B1(new_n9199), .B2(new_n3492), .C(new_n17143), .Y(new_n17144));
  XNOR2x2_ASAP7_75t_L       g16888(.A(new_n3251), .B(new_n17144), .Y(new_n17145));
  AOI31xp33_ASAP7_75t_L     g16889(.A1(new_n17085), .A2(new_n17083), .A3(new_n17088), .B(new_n17095), .Y(new_n17146));
  NOR2xp33_ASAP7_75t_L      g16890(.A(new_n17145), .B(new_n17146), .Y(new_n17147));
  AND2x2_ASAP7_75t_L        g16891(.A(new_n17145), .B(new_n17146), .Y(new_n17148));
  NOR2xp33_ASAP7_75t_L      g16892(.A(new_n17147), .B(new_n17148), .Y(new_n17149));
  AOI22xp33_ASAP7_75t_L     g16893(.A1(new_n3884), .A2(\b[53] ), .B1(new_n3881), .B2(new_n8889), .Y(new_n17150));
  OAI221xp5_ASAP7_75t_L     g16894(.A1(new_n4312), .A2(new_n8569), .B1(new_n8249), .B2(new_n4986), .C(new_n17150), .Y(new_n17151));
  XNOR2x2_ASAP7_75t_L       g16895(.A(\a[35] ), .B(new_n17151), .Y(new_n17152));
  INVx1_ASAP7_75t_L         g16896(.A(new_n17152), .Y(new_n17153));
  AOI22xp33_ASAP7_75t_L     g16897(.A1(new_n6002), .A2(\b[44] ), .B1(new_n5999), .B2(new_n7055), .Y(new_n17154));
  OAI221xp5_ASAP7_75t_L     g16898(.A1(new_n6544), .A2(new_n6195), .B1(new_n5680), .B2(new_n6309), .C(new_n17154), .Y(new_n17155));
  XNOR2x2_ASAP7_75t_L       g16899(.A(\a[44] ), .B(new_n17155), .Y(new_n17156));
  INVx1_ASAP7_75t_L         g16900(.A(new_n17156), .Y(new_n17157));
  INVx1_ASAP7_75t_L         g16901(.A(new_n17049), .Y(new_n17158));
  AOI22xp33_ASAP7_75t_L     g16902(.A1(new_n6822), .A2(\b[41] ), .B1(new_n6819), .B2(new_n5669), .Y(new_n17159));
  OAI221xp5_ASAP7_75t_L     g16903(.A1(new_n7392), .A2(new_n5186), .B1(new_n5166), .B2(new_n7115), .C(new_n17159), .Y(new_n17160));
  XNOR2x2_ASAP7_75t_L       g16904(.A(\a[47] ), .B(new_n17160), .Y(new_n17161));
  AOI22xp33_ASAP7_75t_L     g16905(.A1(new_n8645), .A2(\b[35] ), .B1(new_n8642), .B2(new_n5649), .Y(new_n17162));
  OAI221xp5_ASAP7_75t_L     g16906(.A1(new_n9322), .A2(new_n3827), .B1(new_n3807), .B2(new_n8965), .C(new_n17162), .Y(new_n17163));
  XNOR2x2_ASAP7_75t_L       g16907(.A(\a[53] ), .B(new_n17163), .Y(new_n17164));
  INVx1_ASAP7_75t_L         g16908(.A(new_n17164), .Y(new_n17165));
  INVx1_ASAP7_75t_L         g16909(.A(new_n16999), .Y(new_n17166));
  NOR2xp33_ASAP7_75t_L      g16910(.A(new_n1857), .B(new_n12671), .Y(new_n17167));
  O2A1O1Ixp33_ASAP7_75t_L   g16911(.A1(new_n12353), .A2(new_n12355), .B(\b[23] ), .C(new_n17167), .Y(new_n17168));
  A2O1A1Ixp33_ASAP7_75t_L   g16912(.A1(new_n12669), .A2(\b[22] ), .B(new_n16989), .C(new_n17168), .Y(new_n17169));
  A2O1A1Ixp33_ASAP7_75t_L   g16913(.A1(\b[23] ), .A2(new_n12669), .B(new_n17167), .C(new_n16992), .Y(new_n17170));
  NAND2xp33_ASAP7_75t_L     g16914(.A(new_n17170), .B(new_n17169), .Y(new_n17171));
  AOI22xp33_ASAP7_75t_L     g16915(.A1(new_n11647), .A2(\b[25] ), .B1(\b[26] ), .B2(new_n11656), .Y(new_n17172));
  OAI221xp5_ASAP7_75t_L     g16916(.A1(new_n13003), .A2(new_n2019), .B1(new_n12022), .B2(new_n2487), .C(new_n17172), .Y(new_n17173));
  XNOR2x2_ASAP7_75t_L       g16917(.A(\a[62] ), .B(new_n17173), .Y(new_n17174));
  NOR2xp33_ASAP7_75t_L      g16918(.A(new_n17171), .B(new_n17174), .Y(new_n17175));
  INVx1_ASAP7_75t_L         g16919(.A(new_n17175), .Y(new_n17176));
  NAND2xp33_ASAP7_75t_L     g16920(.A(new_n17171), .B(new_n17174), .Y(new_n17177));
  AND2x2_ASAP7_75t_L        g16921(.A(new_n17177), .B(new_n17176), .Y(new_n17178));
  A2O1A1Ixp33_ASAP7_75t_L   g16922(.A1(new_n17166), .A2(new_n16991), .B(new_n16994), .C(new_n17178), .Y(new_n17179));
  A2O1A1Ixp33_ASAP7_75t_L   g16923(.A1(new_n12669), .A2(\b[20] ), .B(new_n16694), .C(new_n16839), .Y(new_n17180));
  A2O1A1Ixp33_ASAP7_75t_L   g16924(.A1(new_n17180), .A2(new_n16834), .B(new_n16993), .C(new_n17001), .Y(new_n17181));
  NOR2xp33_ASAP7_75t_L      g16925(.A(new_n17181), .B(new_n17178), .Y(new_n17182));
  INVx1_ASAP7_75t_L         g16926(.A(new_n17182), .Y(new_n17183));
  AOI22xp33_ASAP7_75t_L     g16927(.A1(new_n10594), .A2(\b[29] ), .B1(new_n10591), .B2(new_n5472), .Y(new_n17184));
  OAI221xp5_ASAP7_75t_L     g16928(.A1(new_n11335), .A2(new_n2852), .B1(new_n2650), .B2(new_n11330), .C(new_n17184), .Y(new_n17185));
  XNOR2x2_ASAP7_75t_L       g16929(.A(\a[59] ), .B(new_n17185), .Y(new_n17186));
  NAND3xp33_ASAP7_75t_L     g16930(.A(new_n17183), .B(new_n17179), .C(new_n17186), .Y(new_n17187));
  INVx1_ASAP7_75t_L         g16931(.A(new_n17187), .Y(new_n17188));
  AOI21xp33_ASAP7_75t_L     g16932(.A1(new_n17183), .A2(new_n17179), .B(new_n17186), .Y(new_n17189));
  INVx1_ASAP7_75t_L         g16933(.A(new_n17005), .Y(new_n17190));
  NAND2xp33_ASAP7_75t_L     g16934(.A(new_n17190), .B(new_n17008), .Y(new_n17191));
  NOR3xp33_ASAP7_75t_L      g16935(.A(new_n17191), .B(new_n17189), .C(new_n17188), .Y(new_n17192));
  NOR2xp33_ASAP7_75t_L      g16936(.A(new_n17189), .B(new_n17188), .Y(new_n17193));
  O2A1O1Ixp33_ASAP7_75t_L   g16937(.A1(new_n16985), .A2(new_n17006), .B(new_n17190), .C(new_n17193), .Y(new_n17194));
  AOI22xp33_ASAP7_75t_L     g16938(.A1(new_n9623), .A2(\b[32] ), .B1(new_n9620), .B2(new_n3450), .Y(new_n17195));
  OAI221xp5_ASAP7_75t_L     g16939(.A1(new_n10280), .A2(new_n3419), .B1(new_n3212), .B2(new_n12010), .C(new_n17195), .Y(new_n17196));
  XNOR2x2_ASAP7_75t_L       g16940(.A(\a[56] ), .B(new_n17196), .Y(new_n17197));
  OAI21xp33_ASAP7_75t_L     g16941(.A1(new_n17194), .A2(new_n17192), .B(new_n17197), .Y(new_n17198));
  NOR2xp33_ASAP7_75t_L      g16942(.A(new_n17194), .B(new_n17192), .Y(new_n17199));
  INVx1_ASAP7_75t_L         g16943(.A(new_n17197), .Y(new_n17200));
  NAND2xp33_ASAP7_75t_L     g16944(.A(new_n17200), .B(new_n17199), .Y(new_n17201));
  AND2x2_ASAP7_75t_L        g16945(.A(new_n17198), .B(new_n17201), .Y(new_n17202));
  INVx1_ASAP7_75t_L         g16946(.A(new_n17202), .Y(new_n17203));
  A2O1A1Ixp33_ASAP7_75t_L   g16947(.A1(new_n17008), .A2(new_n17009), .B(new_n17013), .C(new_n17019), .Y(new_n17204));
  NOR2xp33_ASAP7_75t_L      g16948(.A(new_n17204), .B(new_n17203), .Y(new_n17205));
  O2A1O1Ixp33_ASAP7_75t_L   g16949(.A1(new_n17013), .A2(new_n17010), .B(new_n17019), .C(new_n17202), .Y(new_n17206));
  NOR2xp33_ASAP7_75t_L      g16950(.A(new_n17206), .B(new_n17205), .Y(new_n17207));
  NAND2xp33_ASAP7_75t_L     g16951(.A(new_n17165), .B(new_n17207), .Y(new_n17208));
  INVx1_ASAP7_75t_L         g16952(.A(new_n17208), .Y(new_n17209));
  NOR2xp33_ASAP7_75t_L      g16953(.A(new_n17165), .B(new_n17207), .Y(new_n17210));
  NOR2xp33_ASAP7_75t_L      g16954(.A(new_n17210), .B(new_n17209), .Y(new_n17211));
  NAND3xp33_ASAP7_75t_L     g16955(.A(new_n17211), .B(new_n17032), .C(new_n17025), .Y(new_n17212));
  O2A1O1Ixp33_ASAP7_75t_L   g16956(.A1(new_n17027), .A2(new_n17033), .B(new_n17025), .C(new_n17211), .Y(new_n17213));
  INVx1_ASAP7_75t_L         g16957(.A(new_n17213), .Y(new_n17214));
  AOI22xp33_ASAP7_75t_L     g16958(.A1(new_n7659), .A2(\b[38] ), .B1(new_n7656), .B2(new_n4923), .Y(new_n17215));
  OAI221xp5_ASAP7_75t_L     g16959(.A1(new_n8326), .A2(new_n4701), .B1(new_n4465), .B2(new_n7994), .C(new_n17215), .Y(new_n17216));
  XNOR2x2_ASAP7_75t_L       g16960(.A(\a[50] ), .B(new_n17216), .Y(new_n17217));
  NAND3xp33_ASAP7_75t_L     g16961(.A(new_n17214), .B(new_n17212), .C(new_n17217), .Y(new_n17218));
  INVx1_ASAP7_75t_L         g16962(.A(new_n17218), .Y(new_n17219));
  AOI21xp33_ASAP7_75t_L     g16963(.A1(new_n17214), .A2(new_n17212), .B(new_n17217), .Y(new_n17220));
  NOR2xp33_ASAP7_75t_L      g16964(.A(new_n17220), .B(new_n17219), .Y(new_n17221));
  NOR2xp33_ASAP7_75t_L      g16965(.A(new_n17039), .B(new_n17046), .Y(new_n17222));
  XNOR2x2_ASAP7_75t_L       g16966(.A(new_n17221), .B(new_n17222), .Y(new_n17223));
  XNOR2x2_ASAP7_75t_L       g16967(.A(new_n17161), .B(new_n17223), .Y(new_n17224));
  O2A1O1Ixp33_ASAP7_75t_L   g16968(.A1(new_n16981), .A2(new_n17050), .B(new_n17158), .C(new_n17224), .Y(new_n17225));
  INVx1_ASAP7_75t_L         g16969(.A(new_n17225), .Y(new_n17226));
  NAND3xp33_ASAP7_75t_L     g16970(.A(new_n17052), .B(new_n17158), .C(new_n17224), .Y(new_n17227));
  NAND3xp33_ASAP7_75t_L     g16971(.A(new_n17226), .B(new_n17157), .C(new_n17227), .Y(new_n17228));
  AO21x2_ASAP7_75t_L        g16972(.A1(new_n17227), .A2(new_n17226), .B(new_n17157), .Y(new_n17229));
  MAJx2_ASAP7_75t_L         g16973(.A(new_n17055), .B(new_n16978), .C(new_n17062), .Y(new_n17230));
  AND3x1_ASAP7_75t_L        g16974(.A(new_n17230), .B(new_n17229), .C(new_n17228), .Y(new_n17231));
  AOI21xp33_ASAP7_75t_L     g16975(.A1(new_n17229), .A2(new_n17228), .B(new_n17230), .Y(new_n17232));
  NOR2xp33_ASAP7_75t_L      g16976(.A(new_n17232), .B(new_n17231), .Y(new_n17233));
  AOI22xp33_ASAP7_75t_L     g16977(.A1(new_n5249), .A2(\b[47] ), .B1(new_n5247), .B2(new_n7323), .Y(new_n17234));
  OAI221xp5_ASAP7_75t_L     g16978(.A1(new_n5241), .A2(new_n7033), .B1(new_n6756), .B2(new_n5521), .C(new_n17234), .Y(new_n17235));
  XNOR2x2_ASAP7_75t_L       g16979(.A(\a[41] ), .B(new_n17235), .Y(new_n17236));
  AND2x2_ASAP7_75t_L        g16980(.A(new_n17236), .B(new_n17233), .Y(new_n17237));
  NOR2xp33_ASAP7_75t_L      g16981(.A(new_n17236), .B(new_n17233), .Y(new_n17238));
  NOR2xp33_ASAP7_75t_L      g16982(.A(new_n17238), .B(new_n17237), .Y(new_n17239));
  A2O1A1Ixp33_ASAP7_75t_L   g16983(.A1(new_n17064), .A2(new_n17063), .B(new_n17071), .C(new_n17239), .Y(new_n17240));
  NAND2xp33_ASAP7_75t_L     g16984(.A(new_n17065), .B(new_n17070), .Y(new_n17241));
  NOR2xp33_ASAP7_75t_L      g16985(.A(new_n17239), .B(new_n17241), .Y(new_n17242));
  INVx1_ASAP7_75t_L         g16986(.A(new_n17242), .Y(new_n17243));
  NAND2xp33_ASAP7_75t_L     g16987(.A(new_n17240), .B(new_n17243), .Y(new_n17244));
  AOI22xp33_ASAP7_75t_L     g16988(.A1(new_n4544), .A2(\b[50] ), .B1(new_n4542), .B2(new_n8235), .Y(new_n17245));
  OAI221xp5_ASAP7_75t_L     g16989(.A1(new_n4536), .A2(new_n7907), .B1(new_n7333), .B2(new_n4781), .C(new_n17245), .Y(new_n17246));
  XNOR2x2_ASAP7_75t_L       g16990(.A(\a[38] ), .B(new_n17246), .Y(new_n17247));
  NAND2xp33_ASAP7_75t_L     g16991(.A(new_n17247), .B(new_n17244), .Y(new_n17248));
  NOR2xp33_ASAP7_75t_L      g16992(.A(new_n17247), .B(new_n17244), .Y(new_n17249));
  INVx1_ASAP7_75t_L         g16993(.A(new_n17249), .Y(new_n17250));
  AND2x2_ASAP7_75t_L        g16994(.A(new_n17248), .B(new_n17250), .Y(new_n17251));
  INVx1_ASAP7_75t_L         g16995(.A(new_n17251), .Y(new_n17252));
  NAND2xp33_ASAP7_75t_L     g16996(.A(new_n17076), .B(new_n17083), .Y(new_n17253));
  NOR2xp33_ASAP7_75t_L      g16997(.A(new_n17253), .B(new_n17252), .Y(new_n17254));
  O2A1O1Ixp33_ASAP7_75t_L   g16998(.A1(new_n17078), .A2(new_n17084), .B(new_n17076), .C(new_n17251), .Y(new_n17255));
  OA21x2_ASAP7_75t_L        g16999(.A1(new_n17255), .A2(new_n17254), .B(new_n17153), .Y(new_n17256));
  NOR3xp33_ASAP7_75t_L      g17000(.A(new_n17254), .B(new_n17255), .C(new_n17153), .Y(new_n17257));
  NOR2xp33_ASAP7_75t_L      g17001(.A(new_n17257), .B(new_n17256), .Y(new_n17258));
  XOR2x2_ASAP7_75t_L        g17002(.A(new_n17258), .B(new_n17149), .Y(new_n17259));
  XNOR2x2_ASAP7_75t_L       g17003(.A(new_n17259), .B(new_n17142), .Y(new_n17260));
  OR3x1_ASAP7_75t_L         g17004(.A(new_n17260), .B(new_n17136), .C(new_n17137), .Y(new_n17261));
  OAI21xp33_ASAP7_75t_L     g17005(.A1(new_n17137), .A2(new_n17136), .B(new_n17260), .Y(new_n17262));
  AND2x2_ASAP7_75t_L        g17006(.A(new_n17262), .B(new_n17261), .Y(new_n17263));
  XNOR2x2_ASAP7_75t_L       g17007(.A(new_n17263), .B(new_n17129), .Y(new_n17264));
  AOI21xp33_ASAP7_75t_L     g17008(.A1(new_n16950), .A2(new_n16953), .B(new_n17105), .Y(new_n17265));
  XOR2x2_ASAP7_75t_L        g17009(.A(new_n17265), .B(new_n17264), .Y(new_n17266));
  A2O1A1Ixp33_ASAP7_75t_L   g17010(.A1(new_n17117), .A2(new_n17113), .B(new_n17112), .C(new_n17266), .Y(new_n17267));
  INVx1_ASAP7_75t_L         g17011(.A(new_n17267), .Y(new_n17268));
  INVx1_ASAP7_75t_L         g17012(.A(new_n17112), .Y(new_n17269));
  A2O1A1Ixp33_ASAP7_75t_L   g17013(.A1(new_n16941), .A2(new_n16938), .B(new_n17114), .C(new_n17269), .Y(new_n17270));
  NOR2xp33_ASAP7_75t_L      g17014(.A(new_n17266), .B(new_n17270), .Y(new_n17271));
  NOR2xp33_ASAP7_75t_L      g17015(.A(new_n17268), .B(new_n17271), .Y(\f[86] ));
  NAND2xp33_ASAP7_75t_L     g17016(.A(\b[63] ), .B(new_n2228), .Y(new_n17273));
  A2O1A1Ixp33_ASAP7_75t_L   g17017(.A1(new_n12607), .A2(new_n12603), .B(new_n2233), .C(new_n17273), .Y(new_n17274));
  AOI221xp5_ASAP7_75t_L     g17018(.A1(\b[61] ), .A2(new_n2386), .B1(\b[62] ), .B2(new_n2232), .C(new_n17274), .Y(new_n17275));
  XNOR2x2_ASAP7_75t_L       g17019(.A(new_n2223), .B(new_n17275), .Y(new_n17276));
  INVx1_ASAP7_75t_L         g17020(.A(new_n17276), .Y(new_n17277));
  O2A1O1Ixp33_ASAP7_75t_L   g17021(.A1(new_n17132), .A2(new_n17135), .B(new_n17261), .C(new_n17277), .Y(new_n17278));
  INVx1_ASAP7_75t_L         g17022(.A(new_n17261), .Y(new_n17279));
  NOR3xp33_ASAP7_75t_L      g17023(.A(new_n17279), .B(new_n17276), .C(new_n17137), .Y(new_n17280));
  NOR2xp33_ASAP7_75t_L      g17024(.A(new_n17278), .B(new_n17280), .Y(new_n17281));
  MAJIxp5_ASAP7_75t_L       g17025(.A(new_n17259), .B(new_n17140), .C(new_n17141), .Y(new_n17282));
  AOI22xp33_ASAP7_75t_L     g17026(.A1(new_n2702), .A2(\b[60] ), .B1(new_n2700), .B2(new_n11234), .Y(new_n17283));
  OAI221xp5_ASAP7_75t_L     g17027(.A1(new_n2694), .A2(new_n10881), .B1(new_n10848), .B2(new_n2932), .C(new_n17283), .Y(new_n17284));
  XNOR2x2_ASAP7_75t_L       g17028(.A(\a[29] ), .B(new_n17284), .Y(new_n17285));
  XNOR2x2_ASAP7_75t_L       g17029(.A(new_n17285), .B(new_n17282), .Y(new_n17286));
  AOI22xp33_ASAP7_75t_L     g17030(.A1(new_n3256), .A2(\b[57] ), .B1(new_n3254), .B2(new_n10495), .Y(new_n17287));
  OAI221xp5_ASAP7_75t_L     g17031(.A1(new_n3248), .A2(new_n10178), .B1(new_n9534), .B2(new_n3492), .C(new_n17287), .Y(new_n17288));
  XNOR2x2_ASAP7_75t_L       g17032(.A(\a[32] ), .B(new_n17288), .Y(new_n17289));
  NOR2xp33_ASAP7_75t_L      g17033(.A(new_n17258), .B(new_n17147), .Y(new_n17290));
  NOR2xp33_ASAP7_75t_L      g17034(.A(new_n17148), .B(new_n17290), .Y(new_n17291));
  XNOR2x2_ASAP7_75t_L       g17035(.A(new_n17289), .B(new_n17291), .Y(new_n17292));
  AOI22xp33_ASAP7_75t_L     g17036(.A1(new_n3884), .A2(\b[54] ), .B1(new_n3881), .B2(new_n9208), .Y(new_n17293));
  OAI221xp5_ASAP7_75t_L     g17037(.A1(new_n4312), .A2(new_n8882), .B1(new_n8569), .B2(new_n4986), .C(new_n17293), .Y(new_n17294));
  XNOR2x2_ASAP7_75t_L       g17038(.A(\a[35] ), .B(new_n17294), .Y(new_n17295));
  INVx1_ASAP7_75t_L         g17039(.A(new_n17241), .Y(new_n17296));
  O2A1O1Ixp33_ASAP7_75t_L   g17040(.A1(new_n17237), .A2(new_n17238), .B(new_n17296), .C(new_n17249), .Y(new_n17297));
  AOI22xp33_ASAP7_75t_L     g17041(.A1(new_n6002), .A2(\b[45] ), .B1(new_n5999), .B2(new_n6764), .Y(new_n17298));
  OAI221xp5_ASAP7_75t_L     g17042(.A1(new_n6544), .A2(new_n6220), .B1(new_n6195), .B2(new_n6309), .C(new_n17298), .Y(new_n17299));
  XNOR2x2_ASAP7_75t_L       g17043(.A(new_n5996), .B(new_n17299), .Y(new_n17300));
  AOI22xp33_ASAP7_75t_L     g17044(.A1(new_n10594), .A2(\b[30] ), .B1(new_n10591), .B2(new_n3219), .Y(new_n17301));
  OAI221xp5_ASAP7_75t_L     g17045(.A1(new_n11335), .A2(new_n2871), .B1(new_n2852), .B2(new_n11330), .C(new_n17301), .Y(new_n17302));
  XNOR2x2_ASAP7_75t_L       g17046(.A(\a[59] ), .B(new_n17302), .Y(new_n17303));
  INVx1_ASAP7_75t_L         g17047(.A(new_n17303), .Y(new_n17304));
  NOR2xp33_ASAP7_75t_L      g17048(.A(new_n1995), .B(new_n12671), .Y(new_n17305));
  A2O1A1Ixp33_ASAP7_75t_L   g17049(.A1(new_n12669), .A2(\b[24] ), .B(new_n17305), .C(new_n1761), .Y(new_n17306));
  INVx1_ASAP7_75t_L         g17050(.A(new_n17306), .Y(new_n17307));
  O2A1O1Ixp33_ASAP7_75t_L   g17051(.A1(new_n12353), .A2(new_n12355), .B(\b[24] ), .C(new_n17305), .Y(new_n17308));
  NAND2xp33_ASAP7_75t_L     g17052(.A(\a[23] ), .B(new_n17308), .Y(new_n17309));
  INVx1_ASAP7_75t_L         g17053(.A(new_n17309), .Y(new_n17310));
  NOR2xp33_ASAP7_75t_L      g17054(.A(new_n17307), .B(new_n17310), .Y(new_n17311));
  XNOR2x2_ASAP7_75t_L       g17055(.A(new_n17168), .B(new_n17311), .Y(new_n17312));
  INVx1_ASAP7_75t_L         g17056(.A(new_n17312), .Y(new_n17313));
  AOI22xp33_ASAP7_75t_L     g17057(.A1(new_n11656), .A2(\b[27] ), .B1(new_n11654), .B2(new_n2657), .Y(new_n17314));
  OAI221xp5_ASAP7_75t_L     g17058(.A1(new_n12364), .A2(new_n2477), .B1(new_n2180), .B2(new_n13003), .C(new_n17314), .Y(new_n17315));
  XNOR2x2_ASAP7_75t_L       g17059(.A(\a[62] ), .B(new_n17315), .Y(new_n17316));
  XNOR2x2_ASAP7_75t_L       g17060(.A(new_n17313), .B(new_n17316), .Y(new_n17317));
  INVx1_ASAP7_75t_L         g17061(.A(new_n17317), .Y(new_n17318));
  A2O1A1Ixp33_ASAP7_75t_L   g17062(.A1(new_n17168), .A2(new_n16993), .B(new_n17175), .C(new_n17318), .Y(new_n17319));
  A2O1A1O1Ixp25_ASAP7_75t_L g17063(.A1(new_n12669), .A2(\b[22] ), .B(new_n16989), .C(new_n17168), .D(new_n17175), .Y(new_n17320));
  NAND2xp33_ASAP7_75t_L     g17064(.A(new_n17320), .B(new_n17317), .Y(new_n17321));
  AND2x2_ASAP7_75t_L        g17065(.A(new_n17321), .B(new_n17319), .Y(new_n17322));
  NAND2xp33_ASAP7_75t_L     g17066(.A(new_n17304), .B(new_n17322), .Y(new_n17323));
  AO21x2_ASAP7_75t_L        g17067(.A1(new_n17321), .A2(new_n17319), .B(new_n17304), .Y(new_n17324));
  AND2x2_ASAP7_75t_L        g17068(.A(new_n17324), .B(new_n17323), .Y(new_n17325));
  O2A1O1Ixp33_ASAP7_75t_L   g17069(.A1(new_n17181), .A2(new_n17178), .B(new_n17187), .C(new_n17325), .Y(new_n17326));
  INVx1_ASAP7_75t_L         g17070(.A(new_n17325), .Y(new_n17327));
  A2O1A1Ixp33_ASAP7_75t_L   g17071(.A1(new_n17176), .A2(new_n17177), .B(new_n17181), .C(new_n17187), .Y(new_n17328));
  NOR2xp33_ASAP7_75t_L      g17072(.A(new_n17328), .B(new_n17327), .Y(new_n17329));
  NOR2xp33_ASAP7_75t_L      g17073(.A(new_n17326), .B(new_n17329), .Y(new_n17330));
  AOI22xp33_ASAP7_75t_L     g17074(.A1(new_n9623), .A2(\b[33] ), .B1(new_n9620), .B2(new_n3813), .Y(new_n17331));
  OAI221xp5_ASAP7_75t_L     g17075(.A1(new_n10280), .A2(new_n3443), .B1(new_n3419), .B2(new_n12010), .C(new_n17331), .Y(new_n17332));
  XNOR2x2_ASAP7_75t_L       g17076(.A(\a[56] ), .B(new_n17332), .Y(new_n17333));
  A2O1A1O1Ixp25_ASAP7_75t_L g17077(.A1(new_n17008), .A2(new_n17190), .B(new_n17193), .C(new_n17201), .D(new_n17333), .Y(new_n17334));
  INVx1_ASAP7_75t_L         g17078(.A(new_n17333), .Y(new_n17335));
  A2O1A1Ixp33_ASAP7_75t_L   g17079(.A1(new_n17008), .A2(new_n17190), .B(new_n17193), .C(new_n17201), .Y(new_n17336));
  NOR2xp33_ASAP7_75t_L      g17080(.A(new_n17335), .B(new_n17336), .Y(new_n17337));
  NOR2xp33_ASAP7_75t_L      g17081(.A(new_n17334), .B(new_n17337), .Y(new_n17338));
  NAND2xp33_ASAP7_75t_L     g17082(.A(new_n17330), .B(new_n17338), .Y(new_n17339));
  INVx1_ASAP7_75t_L         g17083(.A(new_n17339), .Y(new_n17340));
  NOR2xp33_ASAP7_75t_L      g17084(.A(new_n17330), .B(new_n17338), .Y(new_n17341));
  NOR2xp33_ASAP7_75t_L      g17085(.A(new_n17341), .B(new_n17340), .Y(new_n17342));
  AOI22xp33_ASAP7_75t_L     g17086(.A1(new_n8645), .A2(\b[36] ), .B1(new_n8642), .B2(new_n4473), .Y(new_n17343));
  OAI221xp5_ASAP7_75t_L     g17087(.A1(new_n9322), .A2(new_n4053), .B1(new_n3827), .B2(new_n8965), .C(new_n17343), .Y(new_n17344));
  XNOR2x2_ASAP7_75t_L       g17088(.A(\a[53] ), .B(new_n17344), .Y(new_n17345));
  INVx1_ASAP7_75t_L         g17089(.A(new_n17345), .Y(new_n17346));
  XNOR2x2_ASAP7_75t_L       g17090(.A(new_n17346), .B(new_n17342), .Y(new_n17347));
  INVx1_ASAP7_75t_L         g17091(.A(new_n17347), .Y(new_n17348));
  NOR3xp33_ASAP7_75t_L      g17092(.A(new_n17348), .B(new_n17209), .C(new_n17205), .Y(new_n17349));
  O2A1O1Ixp33_ASAP7_75t_L   g17093(.A1(new_n17203), .A2(new_n17204), .B(new_n17208), .C(new_n17347), .Y(new_n17350));
  NOR2xp33_ASAP7_75t_L      g17094(.A(new_n17350), .B(new_n17349), .Y(new_n17351));
  AOI22xp33_ASAP7_75t_L     g17095(.A1(new_n7659), .A2(\b[39] ), .B1(new_n7656), .B2(new_n5174), .Y(new_n17352));
  OAI221xp5_ASAP7_75t_L     g17096(.A1(new_n8326), .A2(new_n4915), .B1(new_n4701), .B2(new_n7994), .C(new_n17352), .Y(new_n17353));
  XNOR2x2_ASAP7_75t_L       g17097(.A(\a[50] ), .B(new_n17353), .Y(new_n17354));
  INVx1_ASAP7_75t_L         g17098(.A(new_n17354), .Y(new_n17355));
  XNOR2x2_ASAP7_75t_L       g17099(.A(new_n17355), .B(new_n17351), .Y(new_n17356));
  A2O1A1Ixp33_ASAP7_75t_L   g17100(.A1(new_n17217), .A2(new_n17212), .B(new_n17213), .C(new_n17356), .Y(new_n17357));
  A2O1A1Ixp33_ASAP7_75t_L   g17101(.A1(new_n17032), .A2(new_n17025), .B(new_n17211), .C(new_n17218), .Y(new_n17358));
  NOR2xp33_ASAP7_75t_L      g17102(.A(new_n17358), .B(new_n17356), .Y(new_n17359));
  INVx1_ASAP7_75t_L         g17103(.A(new_n17359), .Y(new_n17360));
  NAND2xp33_ASAP7_75t_L     g17104(.A(new_n17357), .B(new_n17360), .Y(new_n17361));
  AOI22xp33_ASAP7_75t_L     g17105(.A1(new_n6822), .A2(\b[42] ), .B1(new_n6819), .B2(new_n5688), .Y(new_n17362));
  OAI221xp5_ASAP7_75t_L     g17106(.A1(new_n7392), .A2(new_n5666), .B1(new_n5186), .B2(new_n7115), .C(new_n17362), .Y(new_n17363));
  XNOR2x2_ASAP7_75t_L       g17107(.A(\a[47] ), .B(new_n17363), .Y(new_n17364));
  XNOR2x2_ASAP7_75t_L       g17108(.A(new_n17364), .B(new_n17361), .Y(new_n17365));
  MAJx2_ASAP7_75t_L         g17109(.A(new_n17222), .B(new_n17221), .C(new_n17161), .Y(new_n17366));
  XOR2x2_ASAP7_75t_L        g17110(.A(new_n17366), .B(new_n17365), .Y(new_n17367));
  XOR2x2_ASAP7_75t_L        g17111(.A(new_n17300), .B(new_n17367), .Y(new_n17368));
  INVx1_ASAP7_75t_L         g17112(.A(new_n17368), .Y(new_n17369));
  NAND3xp33_ASAP7_75t_L     g17113(.A(new_n17369), .B(new_n17228), .C(new_n17226), .Y(new_n17370));
  A2O1A1O1Ixp25_ASAP7_75t_L g17114(.A1(new_n17052), .A2(new_n17158), .B(new_n17224), .C(new_n17228), .D(new_n17369), .Y(new_n17371));
  INVx1_ASAP7_75t_L         g17115(.A(new_n17371), .Y(new_n17372));
  NAND2xp33_ASAP7_75t_L     g17116(.A(new_n17370), .B(new_n17372), .Y(new_n17373));
  AOI22xp33_ASAP7_75t_L     g17117(.A1(new_n5249), .A2(\b[48] ), .B1(new_n5247), .B2(new_n7341), .Y(new_n17374));
  OAI221xp5_ASAP7_75t_L     g17118(.A1(new_n5241), .A2(new_n7316), .B1(new_n7033), .B2(new_n5521), .C(new_n17374), .Y(new_n17375));
  XNOR2x2_ASAP7_75t_L       g17119(.A(\a[41] ), .B(new_n17375), .Y(new_n17376));
  XNOR2x2_ASAP7_75t_L       g17120(.A(new_n17376), .B(new_n17373), .Y(new_n17377));
  A2O1A1Ixp33_ASAP7_75t_L   g17121(.A1(new_n17233), .A2(new_n17236), .B(new_n17232), .C(new_n17377), .Y(new_n17378));
  OR3x1_ASAP7_75t_L         g17122(.A(new_n17377), .B(new_n17232), .C(new_n17237), .Y(new_n17379));
  AND2x2_ASAP7_75t_L        g17123(.A(new_n17378), .B(new_n17379), .Y(new_n17380));
  AOI22xp33_ASAP7_75t_L     g17124(.A1(new_n4544), .A2(\b[51] ), .B1(new_n4542), .B2(new_n8257), .Y(new_n17381));
  OAI221xp5_ASAP7_75t_L     g17125(.A1(new_n4536), .A2(new_n8228), .B1(new_n7907), .B2(new_n4781), .C(new_n17381), .Y(new_n17382));
  XNOR2x2_ASAP7_75t_L       g17126(.A(\a[38] ), .B(new_n17382), .Y(new_n17383));
  INVx1_ASAP7_75t_L         g17127(.A(new_n17383), .Y(new_n17384));
  NAND2xp33_ASAP7_75t_L     g17128(.A(new_n17384), .B(new_n17380), .Y(new_n17385));
  AO21x2_ASAP7_75t_L        g17129(.A1(new_n17378), .A2(new_n17379), .B(new_n17384), .Y(new_n17386));
  AND2x2_ASAP7_75t_L        g17130(.A(new_n17386), .B(new_n17385), .Y(new_n17387));
  XNOR2x2_ASAP7_75t_L       g17131(.A(new_n17297), .B(new_n17387), .Y(new_n17388));
  INVx1_ASAP7_75t_L         g17132(.A(new_n17388), .Y(new_n17389));
  NAND2xp33_ASAP7_75t_L     g17133(.A(new_n17295), .B(new_n17389), .Y(new_n17390));
  INVx1_ASAP7_75t_L         g17134(.A(new_n17295), .Y(new_n17391));
  NAND2xp33_ASAP7_75t_L     g17135(.A(new_n17391), .B(new_n17388), .Y(new_n17392));
  A2O1A1O1Ixp25_ASAP7_75t_L g17136(.A1(new_n17079), .A2(new_n17082), .B(new_n17077), .C(new_n17252), .D(new_n17257), .Y(new_n17393));
  NAND3xp33_ASAP7_75t_L     g17137(.A(new_n17393), .B(new_n17392), .C(new_n17390), .Y(new_n17394));
  NAND2xp33_ASAP7_75t_L     g17138(.A(new_n17392), .B(new_n17390), .Y(new_n17395));
  A2O1A1Ixp33_ASAP7_75t_L   g17139(.A1(new_n17253), .A2(new_n17252), .B(new_n17257), .C(new_n17395), .Y(new_n17396));
  NAND2xp33_ASAP7_75t_L     g17140(.A(new_n17394), .B(new_n17396), .Y(new_n17397));
  XOR2x2_ASAP7_75t_L        g17141(.A(new_n17397), .B(new_n17292), .Y(new_n17398));
  XNOR2x2_ASAP7_75t_L       g17142(.A(new_n17398), .B(new_n17286), .Y(new_n17399));
  INVx1_ASAP7_75t_L         g17143(.A(new_n17399), .Y(new_n17400));
  XNOR2x2_ASAP7_75t_L       g17144(.A(new_n17400), .B(new_n17281), .Y(new_n17401));
  A2O1A1Ixp33_ASAP7_75t_L   g17145(.A1(new_n17128), .A2(new_n17263), .B(new_n17126), .C(new_n17401), .Y(new_n17402));
  INVx1_ASAP7_75t_L         g17146(.A(new_n17402), .Y(new_n17403));
  AOI211xp5_ASAP7_75t_L     g17147(.A1(new_n17128), .A2(new_n17263), .B(new_n17126), .C(new_n17401), .Y(new_n17404));
  NOR2xp33_ASAP7_75t_L      g17148(.A(new_n17404), .B(new_n17403), .Y(new_n17405));
  A2O1A1Ixp33_ASAP7_75t_L   g17149(.A1(new_n17265), .A2(new_n17264), .B(new_n17268), .C(new_n17405), .Y(new_n17406));
  NAND2xp33_ASAP7_75t_L     g17150(.A(new_n17265), .B(new_n17264), .Y(new_n17407));
  INVx1_ASAP7_75t_L         g17151(.A(new_n17407), .Y(new_n17408));
  A2O1A1O1Ixp25_ASAP7_75t_L g17152(.A1(new_n17113), .A2(new_n17117), .B(new_n17112), .C(new_n17266), .D(new_n17408), .Y(new_n17409));
  OAI21xp33_ASAP7_75t_L     g17153(.A1(new_n17403), .A2(new_n17404), .B(new_n17409), .Y(new_n17410));
  AND2x2_ASAP7_75t_L        g17154(.A(new_n17410), .B(new_n17406), .Y(\f[87] ));
  O2A1O1Ixp33_ASAP7_75t_L   g17155(.A1(new_n17132), .A2(new_n17135), .B(new_n17261), .C(new_n17276), .Y(new_n17412));
  O2A1O1Ixp33_ASAP7_75t_L   g17156(.A1(new_n17278), .A2(new_n17280), .B(new_n17400), .C(new_n17412), .Y(new_n17413));
  AOI22xp33_ASAP7_75t_L     g17157(.A1(new_n2702), .A2(\b[61] ), .B1(new_n2700), .B2(new_n11919), .Y(new_n17414));
  OAI221xp5_ASAP7_75t_L     g17158(.A1(new_n2694), .A2(new_n11226), .B1(new_n10881), .B2(new_n2932), .C(new_n17414), .Y(new_n17415));
  XNOR2x2_ASAP7_75t_L       g17159(.A(\a[29] ), .B(new_n17415), .Y(new_n17416));
  MAJIxp5_ASAP7_75t_L       g17160(.A(new_n17397), .B(new_n17289), .C(new_n17291), .Y(new_n17417));
  XNOR2x2_ASAP7_75t_L       g17161(.A(new_n17416), .B(new_n17417), .Y(new_n17418));
  INVx1_ASAP7_75t_L         g17162(.A(new_n17392), .Y(new_n17419));
  AOI22xp33_ASAP7_75t_L     g17163(.A1(new_n3260), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n3256), .Y(new_n17420));
  OAI221xp5_ASAP7_75t_L     g17164(.A1(new_n3492), .A2(new_n10178), .B1(new_n3261), .B2(new_n10856), .C(new_n17420), .Y(new_n17421));
  XNOR2x2_ASAP7_75t_L       g17165(.A(\a[32] ), .B(new_n17421), .Y(new_n17422));
  INVx1_ASAP7_75t_L         g17166(.A(new_n17422), .Y(new_n17423));
  A2O1A1Ixp33_ASAP7_75t_L   g17167(.A1(new_n17393), .A2(new_n17390), .B(new_n17419), .C(new_n17423), .Y(new_n17424));
  NAND3xp33_ASAP7_75t_L     g17168(.A(new_n17394), .B(new_n17392), .C(new_n17422), .Y(new_n17425));
  AND2x2_ASAP7_75t_L        g17169(.A(new_n17424), .B(new_n17425), .Y(new_n17426));
  INVx1_ASAP7_75t_L         g17170(.A(new_n17297), .Y(new_n17427));
  INVx1_ASAP7_75t_L         g17171(.A(new_n17385), .Y(new_n17428));
  NAND2xp33_ASAP7_75t_L     g17172(.A(new_n17300), .B(new_n17367), .Y(new_n17429));
  AOI22xp33_ASAP7_75t_L     g17173(.A1(new_n7659), .A2(\b[40] ), .B1(new_n7656), .B2(new_n5194), .Y(new_n17430));
  OAI221xp5_ASAP7_75t_L     g17174(.A1(new_n8326), .A2(new_n5166), .B1(new_n4915), .B2(new_n7994), .C(new_n17430), .Y(new_n17431));
  XNOR2x2_ASAP7_75t_L       g17175(.A(\a[50] ), .B(new_n17431), .Y(new_n17432));
  INVx1_ASAP7_75t_L         g17176(.A(new_n17432), .Y(new_n17433));
  INVx1_ASAP7_75t_L         g17177(.A(new_n17320), .Y(new_n17434));
  NOR2xp33_ASAP7_75t_L      g17178(.A(new_n17313), .B(new_n17316), .Y(new_n17435));
  NOR2xp33_ASAP7_75t_L      g17179(.A(new_n2019), .B(new_n12671), .Y(new_n17436));
  A2O1A1O1Ixp25_ASAP7_75t_L g17180(.A1(new_n12669), .A2(\b[23] ), .B(new_n17167), .C(new_n17309), .D(new_n17307), .Y(new_n17437));
  A2O1A1Ixp33_ASAP7_75t_L   g17181(.A1(new_n12669), .A2(\b[25] ), .B(new_n17436), .C(new_n17437), .Y(new_n17438));
  O2A1O1Ixp33_ASAP7_75t_L   g17182(.A1(new_n12353), .A2(new_n12355), .B(\b[25] ), .C(new_n17436), .Y(new_n17439));
  INVx1_ASAP7_75t_L         g17183(.A(new_n17439), .Y(new_n17440));
  O2A1O1Ixp33_ASAP7_75t_L   g17184(.A1(new_n17168), .A2(new_n17310), .B(new_n17306), .C(new_n17440), .Y(new_n17441));
  INVx1_ASAP7_75t_L         g17185(.A(new_n17441), .Y(new_n17442));
  NAND2xp33_ASAP7_75t_L     g17186(.A(new_n17438), .B(new_n17442), .Y(new_n17443));
  AOI22xp33_ASAP7_75t_L     g17187(.A1(new_n11647), .A2(\b[27] ), .B1(\b[28] ), .B2(new_n11656), .Y(new_n17444));
  OAI221xp5_ASAP7_75t_L     g17188(.A1(new_n13003), .A2(new_n2477), .B1(new_n12022), .B2(new_n5212), .C(new_n17444), .Y(new_n17445));
  XNOR2x2_ASAP7_75t_L       g17189(.A(\a[62] ), .B(new_n17445), .Y(new_n17446));
  NOR2xp33_ASAP7_75t_L      g17190(.A(new_n17443), .B(new_n17446), .Y(new_n17447));
  INVx1_ASAP7_75t_L         g17191(.A(new_n17447), .Y(new_n17448));
  NAND2xp33_ASAP7_75t_L     g17192(.A(new_n17443), .B(new_n17446), .Y(new_n17449));
  AND2x2_ASAP7_75t_L        g17193(.A(new_n17449), .B(new_n17448), .Y(new_n17450));
  A2O1A1Ixp33_ASAP7_75t_L   g17194(.A1(new_n17318), .A2(new_n17434), .B(new_n17435), .C(new_n17450), .Y(new_n17451));
  A2O1A1O1Ixp25_ASAP7_75t_L g17195(.A1(new_n17168), .A2(new_n16993), .B(new_n17175), .C(new_n17318), .D(new_n17435), .Y(new_n17452));
  INVx1_ASAP7_75t_L         g17196(.A(new_n17452), .Y(new_n17453));
  NOR2xp33_ASAP7_75t_L      g17197(.A(new_n17450), .B(new_n17453), .Y(new_n17454));
  INVx1_ASAP7_75t_L         g17198(.A(new_n17454), .Y(new_n17455));
  AOI22xp33_ASAP7_75t_L     g17199(.A1(new_n10594), .A2(\b[31] ), .B1(new_n10591), .B2(new_n3426), .Y(new_n17456));
  OAI221xp5_ASAP7_75t_L     g17200(.A1(new_n11335), .A2(new_n3212), .B1(new_n2871), .B2(new_n11330), .C(new_n17456), .Y(new_n17457));
  XNOR2x2_ASAP7_75t_L       g17201(.A(\a[59] ), .B(new_n17457), .Y(new_n17458));
  NAND3xp33_ASAP7_75t_L     g17202(.A(new_n17455), .B(new_n17451), .C(new_n17458), .Y(new_n17459));
  INVx1_ASAP7_75t_L         g17203(.A(new_n17459), .Y(new_n17460));
  AOI21xp33_ASAP7_75t_L     g17204(.A1(new_n17455), .A2(new_n17451), .B(new_n17458), .Y(new_n17461));
  NOR2xp33_ASAP7_75t_L      g17205(.A(new_n17461), .B(new_n17460), .Y(new_n17462));
  AOI21xp33_ASAP7_75t_L     g17206(.A1(new_n17322), .A2(new_n17304), .B(new_n17329), .Y(new_n17463));
  NAND2xp33_ASAP7_75t_L     g17207(.A(new_n17462), .B(new_n17463), .Y(new_n17464));
  INVx1_ASAP7_75t_L         g17208(.A(new_n17464), .Y(new_n17465));
  O2A1O1Ixp33_ASAP7_75t_L   g17209(.A1(new_n17327), .A2(new_n17328), .B(new_n17323), .C(new_n17462), .Y(new_n17466));
  NOR2xp33_ASAP7_75t_L      g17210(.A(new_n17466), .B(new_n17465), .Y(new_n17467));
  AOI22xp33_ASAP7_75t_L     g17211(.A1(new_n9623), .A2(\b[34] ), .B1(new_n9620), .B2(new_n3833), .Y(new_n17468));
  OAI221xp5_ASAP7_75t_L     g17212(.A1(new_n10280), .A2(new_n3807), .B1(new_n3443), .B2(new_n12010), .C(new_n17468), .Y(new_n17469));
  XNOR2x2_ASAP7_75t_L       g17213(.A(\a[56] ), .B(new_n17469), .Y(new_n17470));
  NAND2xp33_ASAP7_75t_L     g17214(.A(new_n17470), .B(new_n17467), .Y(new_n17471));
  INVx1_ASAP7_75t_L         g17215(.A(new_n17470), .Y(new_n17472));
  OAI21xp33_ASAP7_75t_L     g17216(.A1(new_n17466), .A2(new_n17465), .B(new_n17472), .Y(new_n17473));
  AND2x2_ASAP7_75t_L        g17217(.A(new_n17473), .B(new_n17471), .Y(new_n17474));
  A2O1A1O1Ixp25_ASAP7_75t_L g17218(.A1(new_n17199), .A2(new_n17200), .B(new_n17194), .C(new_n17335), .D(new_n17340), .Y(new_n17475));
  NAND2xp33_ASAP7_75t_L     g17219(.A(new_n17474), .B(new_n17475), .Y(new_n17476));
  INVx1_ASAP7_75t_L         g17220(.A(new_n17474), .Y(new_n17477));
  A2O1A1Ixp33_ASAP7_75t_L   g17221(.A1(new_n17338), .A2(new_n17330), .B(new_n17334), .C(new_n17477), .Y(new_n17478));
  AND2x2_ASAP7_75t_L        g17222(.A(new_n17476), .B(new_n17478), .Y(new_n17479));
  INVx1_ASAP7_75t_L         g17223(.A(new_n17479), .Y(new_n17480));
  AOI22xp33_ASAP7_75t_L     g17224(.A1(new_n8645), .A2(\b[37] ), .B1(new_n8642), .B2(new_n4709), .Y(new_n17481));
  OAI221xp5_ASAP7_75t_L     g17225(.A1(new_n9322), .A2(new_n4465), .B1(new_n4053), .B2(new_n8965), .C(new_n17481), .Y(new_n17482));
  XNOR2x2_ASAP7_75t_L       g17226(.A(\a[53] ), .B(new_n17482), .Y(new_n17483));
  AND2x2_ASAP7_75t_L        g17227(.A(new_n17483), .B(new_n17480), .Y(new_n17484));
  NOR2xp33_ASAP7_75t_L      g17228(.A(new_n17483), .B(new_n17480), .Y(new_n17485));
  NOR2xp33_ASAP7_75t_L      g17229(.A(new_n17485), .B(new_n17484), .Y(new_n17486));
  A2O1A1Ixp33_ASAP7_75t_L   g17230(.A1(new_n17346), .A2(new_n17342), .B(new_n17350), .C(new_n17486), .Y(new_n17487));
  INVx1_ASAP7_75t_L         g17231(.A(new_n17487), .Y(new_n17488));
  AOI211xp5_ASAP7_75t_L     g17232(.A1(new_n17342), .A2(new_n17346), .B(new_n17350), .C(new_n17486), .Y(new_n17489));
  NOR2xp33_ASAP7_75t_L      g17233(.A(new_n17489), .B(new_n17488), .Y(new_n17490));
  NAND2xp33_ASAP7_75t_L     g17234(.A(new_n17433), .B(new_n17490), .Y(new_n17491));
  OAI21xp33_ASAP7_75t_L     g17235(.A1(new_n17489), .A2(new_n17488), .B(new_n17432), .Y(new_n17492));
  AND2x2_ASAP7_75t_L        g17236(.A(new_n17492), .B(new_n17491), .Y(new_n17493));
  A2O1A1Ixp33_ASAP7_75t_L   g17237(.A1(new_n17355), .A2(new_n17351), .B(new_n17359), .C(new_n17493), .Y(new_n17494));
  AOI21xp33_ASAP7_75t_L     g17238(.A1(new_n17355), .A2(new_n17351), .B(new_n17359), .Y(new_n17495));
  INVx1_ASAP7_75t_L         g17239(.A(new_n17495), .Y(new_n17496));
  NOR2xp33_ASAP7_75t_L      g17240(.A(new_n17496), .B(new_n17493), .Y(new_n17497));
  INVx1_ASAP7_75t_L         g17241(.A(new_n17497), .Y(new_n17498));
  AOI22xp33_ASAP7_75t_L     g17242(.A1(new_n6822), .A2(\b[43] ), .B1(new_n6819), .B2(new_n6202), .Y(new_n17499));
  OAI221xp5_ASAP7_75t_L     g17243(.A1(new_n7392), .A2(new_n5680), .B1(new_n5666), .B2(new_n7115), .C(new_n17499), .Y(new_n17500));
  XNOR2x2_ASAP7_75t_L       g17244(.A(\a[47] ), .B(new_n17500), .Y(new_n17501));
  NAND3xp33_ASAP7_75t_L     g17245(.A(new_n17498), .B(new_n17494), .C(new_n17501), .Y(new_n17502));
  AO21x2_ASAP7_75t_L        g17246(.A1(new_n17494), .A2(new_n17498), .B(new_n17501), .Y(new_n17503));
  NAND2xp33_ASAP7_75t_L     g17247(.A(new_n17502), .B(new_n17503), .Y(new_n17504));
  MAJIxp5_ASAP7_75t_L       g17248(.A(new_n17361), .B(new_n17364), .C(new_n17366), .Y(new_n17505));
  NOR2xp33_ASAP7_75t_L      g17249(.A(new_n17505), .B(new_n17504), .Y(new_n17506));
  INVx1_ASAP7_75t_L         g17250(.A(new_n17506), .Y(new_n17507));
  NAND2xp33_ASAP7_75t_L     g17251(.A(new_n17505), .B(new_n17504), .Y(new_n17508));
  AOI22xp33_ASAP7_75t_L     g17252(.A1(new_n6002), .A2(\b[46] ), .B1(new_n5999), .B2(new_n7041), .Y(new_n17509));
  OAI221xp5_ASAP7_75t_L     g17253(.A1(new_n6544), .A2(new_n6756), .B1(new_n6220), .B2(new_n6309), .C(new_n17509), .Y(new_n17510));
  XNOR2x2_ASAP7_75t_L       g17254(.A(\a[44] ), .B(new_n17510), .Y(new_n17511));
  NAND3xp33_ASAP7_75t_L     g17255(.A(new_n17507), .B(new_n17508), .C(new_n17511), .Y(new_n17512));
  AO21x2_ASAP7_75t_L        g17256(.A1(new_n17508), .A2(new_n17507), .B(new_n17511), .Y(new_n17513));
  NAND4xp25_ASAP7_75t_L     g17257(.A(new_n17513), .B(new_n17429), .C(new_n17372), .D(new_n17512), .Y(new_n17514));
  NAND2xp33_ASAP7_75t_L     g17258(.A(new_n17512), .B(new_n17513), .Y(new_n17515));
  A2O1A1Ixp33_ASAP7_75t_L   g17259(.A1(new_n17367), .A2(new_n17300), .B(new_n17371), .C(new_n17515), .Y(new_n17516));
  NAND2xp33_ASAP7_75t_L     g17260(.A(new_n5247), .B(new_n7914), .Y(new_n17517));
  OAI221xp5_ASAP7_75t_L     g17261(.A1(new_n5253), .A2(new_n7907), .B1(new_n7333), .B2(new_n5241), .C(new_n17517), .Y(new_n17518));
  AOI21xp33_ASAP7_75t_L     g17262(.A1(new_n5526), .A2(\b[47] ), .B(new_n17518), .Y(new_n17519));
  NAND2xp33_ASAP7_75t_L     g17263(.A(\a[41] ), .B(new_n17519), .Y(new_n17520));
  A2O1A1Ixp33_ASAP7_75t_L   g17264(.A1(\b[47] ), .A2(new_n5526), .B(new_n17518), .C(new_n5244), .Y(new_n17521));
  AND2x2_ASAP7_75t_L        g17265(.A(new_n17521), .B(new_n17520), .Y(new_n17522));
  NAND3xp33_ASAP7_75t_L     g17266(.A(new_n17516), .B(new_n17514), .C(new_n17522), .Y(new_n17523));
  AO21x2_ASAP7_75t_L        g17267(.A1(new_n17514), .A2(new_n17516), .B(new_n17522), .Y(new_n17524));
  NAND2xp33_ASAP7_75t_L     g17268(.A(new_n17523), .B(new_n17524), .Y(new_n17525));
  OAI21xp33_ASAP7_75t_L     g17269(.A1(new_n17373), .A2(new_n17376), .B(new_n17379), .Y(new_n17526));
  NOR2xp33_ASAP7_75t_L      g17270(.A(new_n17525), .B(new_n17526), .Y(new_n17527));
  INVx1_ASAP7_75t_L         g17271(.A(new_n17527), .Y(new_n17528));
  NAND2xp33_ASAP7_75t_L     g17272(.A(new_n17525), .B(new_n17526), .Y(new_n17529));
  NAND2xp33_ASAP7_75t_L     g17273(.A(new_n17529), .B(new_n17528), .Y(new_n17530));
  AOI22xp33_ASAP7_75t_L     g17274(.A1(new_n4544), .A2(\b[52] ), .B1(new_n4542), .B2(new_n8577), .Y(new_n17531));
  OAI221xp5_ASAP7_75t_L     g17275(.A1(new_n4536), .A2(new_n8249), .B1(new_n8228), .B2(new_n4781), .C(new_n17531), .Y(new_n17532));
  XNOR2x2_ASAP7_75t_L       g17276(.A(\a[38] ), .B(new_n17532), .Y(new_n17533));
  INVx1_ASAP7_75t_L         g17277(.A(new_n17533), .Y(new_n17534));
  NOR2xp33_ASAP7_75t_L      g17278(.A(new_n17534), .B(new_n17530), .Y(new_n17535));
  AOI21xp33_ASAP7_75t_L     g17279(.A1(new_n17528), .A2(new_n17529), .B(new_n17533), .Y(new_n17536));
  NOR2xp33_ASAP7_75t_L      g17280(.A(new_n17536), .B(new_n17535), .Y(new_n17537));
  A2O1A1Ixp33_ASAP7_75t_L   g17281(.A1(new_n17386), .A2(new_n17427), .B(new_n17428), .C(new_n17537), .Y(new_n17538));
  INVx1_ASAP7_75t_L         g17282(.A(new_n17537), .Y(new_n17539));
  O2A1O1Ixp33_ASAP7_75t_L   g17283(.A1(new_n17249), .A2(new_n17242), .B(new_n17386), .C(new_n17428), .Y(new_n17540));
  NAND2xp33_ASAP7_75t_L     g17284(.A(new_n17540), .B(new_n17539), .Y(new_n17541));
  NAND2xp33_ASAP7_75t_L     g17285(.A(new_n17538), .B(new_n17541), .Y(new_n17542));
  NAND2xp33_ASAP7_75t_L     g17286(.A(new_n3881), .B(new_n9542), .Y(new_n17543));
  OAI221xp5_ASAP7_75t_L     g17287(.A1(new_n4115), .A2(new_n9534), .B1(new_n9199), .B2(new_n4312), .C(new_n17543), .Y(new_n17544));
  AOI21xp33_ASAP7_75t_L     g17288(.A1(new_n4111), .A2(\b[53] ), .B(new_n17544), .Y(new_n17545));
  NAND2xp33_ASAP7_75t_L     g17289(.A(\a[35] ), .B(new_n17545), .Y(new_n17546));
  A2O1A1Ixp33_ASAP7_75t_L   g17290(.A1(\b[53] ), .A2(new_n4111), .B(new_n17544), .C(new_n3878), .Y(new_n17547));
  AND2x2_ASAP7_75t_L        g17291(.A(new_n17547), .B(new_n17546), .Y(new_n17548));
  INVx1_ASAP7_75t_L         g17292(.A(new_n17548), .Y(new_n17549));
  NAND2xp33_ASAP7_75t_L     g17293(.A(new_n17549), .B(new_n17542), .Y(new_n17550));
  INVx1_ASAP7_75t_L         g17294(.A(new_n17542), .Y(new_n17551));
  NAND2xp33_ASAP7_75t_L     g17295(.A(new_n17548), .B(new_n17551), .Y(new_n17552));
  AND2x2_ASAP7_75t_L        g17296(.A(new_n17550), .B(new_n17552), .Y(new_n17553));
  NAND2xp33_ASAP7_75t_L     g17297(.A(new_n17426), .B(new_n17553), .Y(new_n17554));
  AO21x2_ASAP7_75t_L        g17298(.A1(new_n17552), .A2(new_n17550), .B(new_n17426), .Y(new_n17555));
  NAND2xp33_ASAP7_75t_L     g17299(.A(new_n17554), .B(new_n17555), .Y(new_n17556));
  XNOR2x2_ASAP7_75t_L       g17300(.A(new_n17556), .B(new_n17418), .Y(new_n17557));
  INVx1_ASAP7_75t_L         g17301(.A(new_n17285), .Y(new_n17558));
  MAJIxp5_ASAP7_75t_L       g17302(.A(new_n17398), .B(new_n17282), .C(new_n17558), .Y(new_n17559));
  AOI22xp33_ASAP7_75t_L     g17303(.A1(new_n2232), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2386), .Y(new_n17560));
  A2O1A1Ixp33_ASAP7_75t_L   g17304(.A1(new_n13506), .A2(new_n13507), .B(new_n2233), .C(new_n17560), .Y(new_n17561));
  NOR2xp33_ASAP7_75t_L      g17305(.A(new_n2223), .B(new_n17561), .Y(new_n17562));
  A2O1A1O1Ixp25_ASAP7_75t_L g17306(.A1(new_n13507), .A2(new_n13506), .B(new_n2233), .C(new_n17560), .D(\a[26] ), .Y(new_n17563));
  NOR2xp33_ASAP7_75t_L      g17307(.A(new_n17563), .B(new_n17562), .Y(new_n17564));
  INVx1_ASAP7_75t_L         g17308(.A(new_n17564), .Y(new_n17565));
  XNOR2x2_ASAP7_75t_L       g17309(.A(new_n17565), .B(new_n17559), .Y(new_n17566));
  XNOR2x2_ASAP7_75t_L       g17310(.A(new_n17557), .B(new_n17566), .Y(new_n17567));
  NOR2xp33_ASAP7_75t_L      g17311(.A(new_n17567), .B(new_n17413), .Y(new_n17568));
  INVx1_ASAP7_75t_L         g17312(.A(new_n17568), .Y(new_n17569));
  NAND2xp33_ASAP7_75t_L     g17313(.A(new_n17567), .B(new_n17413), .Y(new_n17570));
  NAND2xp33_ASAP7_75t_L     g17314(.A(new_n17570), .B(new_n17569), .Y(new_n17571));
  A2O1A1O1Ixp25_ASAP7_75t_L g17315(.A1(new_n17407), .A2(new_n17267), .B(new_n17404), .C(new_n17402), .D(new_n17571), .Y(new_n17572));
  A2O1A1Ixp33_ASAP7_75t_L   g17316(.A1(new_n17267), .A2(new_n17407), .B(new_n17404), .C(new_n17402), .Y(new_n17573));
  INVx1_ASAP7_75t_L         g17317(.A(new_n17571), .Y(new_n17574));
  NOR2xp33_ASAP7_75t_L      g17318(.A(new_n17574), .B(new_n17573), .Y(new_n17575));
  NOR2xp33_ASAP7_75t_L      g17319(.A(new_n17572), .B(new_n17575), .Y(\f[88] ));
  NAND2xp33_ASAP7_75t_L     g17320(.A(new_n17557), .B(new_n17566), .Y(new_n17577));
  OAI21xp33_ASAP7_75t_L     g17321(.A1(new_n17559), .A2(new_n17564), .B(new_n17577), .Y(new_n17578));
  AOI22xp33_ASAP7_75t_L     g17322(.A1(new_n2702), .A2(\b[62] ), .B1(new_n2700), .B2(new_n12280), .Y(new_n17579));
  OAI221xp5_ASAP7_75t_L     g17323(.A1(new_n2694), .A2(new_n11911), .B1(new_n11226), .B2(new_n2932), .C(new_n17579), .Y(new_n17580));
  XNOR2x2_ASAP7_75t_L       g17324(.A(\a[29] ), .B(new_n17580), .Y(new_n17581));
  INVx1_ASAP7_75t_L         g17325(.A(new_n17581), .Y(new_n17582));
  A2O1A1Ixp33_ASAP7_75t_L   g17326(.A1(new_n17394), .A2(new_n17392), .B(new_n17422), .C(new_n17554), .Y(new_n17583));
  NOR2xp33_ASAP7_75t_L      g17327(.A(new_n17582), .B(new_n17583), .Y(new_n17584));
  A2O1A1O1Ixp25_ASAP7_75t_L g17328(.A1(new_n17394), .A2(new_n17392), .B(new_n17422), .C(new_n17554), .D(new_n17581), .Y(new_n17585));
  NOR2xp33_ASAP7_75t_L      g17329(.A(new_n17585), .B(new_n17584), .Y(new_n17586));
  AOI22xp33_ASAP7_75t_L     g17330(.A1(new_n3256), .A2(\b[59] ), .B1(new_n3254), .B2(new_n10887), .Y(new_n17587));
  OAI221xp5_ASAP7_75t_L     g17331(.A1(new_n3248), .A2(new_n10848), .B1(new_n10488), .B2(new_n3492), .C(new_n17587), .Y(new_n17588));
  XNOR2x2_ASAP7_75t_L       g17332(.A(\a[32] ), .B(new_n17588), .Y(new_n17589));
  INVx1_ASAP7_75t_L         g17333(.A(new_n17589), .Y(new_n17590));
  A2O1A1Ixp33_ASAP7_75t_L   g17334(.A1(new_n17386), .A2(new_n17427), .B(new_n17428), .C(new_n17539), .Y(new_n17591));
  A2O1A1Ixp33_ASAP7_75t_L   g17335(.A1(new_n17541), .A2(new_n17538), .B(new_n17548), .C(new_n17591), .Y(new_n17592));
  NOR2xp33_ASAP7_75t_L      g17336(.A(new_n17590), .B(new_n17592), .Y(new_n17593));
  A2O1A1O1Ixp25_ASAP7_75t_L g17337(.A1(new_n17538), .A2(new_n17541), .B(new_n17548), .C(new_n17591), .D(new_n17589), .Y(new_n17594));
  AOI22xp33_ASAP7_75t_L     g17338(.A1(new_n3884), .A2(\b[56] ), .B1(new_n3881), .B2(new_n10185), .Y(new_n17595));
  OAI221xp5_ASAP7_75t_L     g17339(.A1(new_n4312), .A2(new_n9534), .B1(new_n9199), .B2(new_n4986), .C(new_n17595), .Y(new_n17596));
  XNOR2x2_ASAP7_75t_L       g17340(.A(\a[35] ), .B(new_n17596), .Y(new_n17597));
  AOI22xp33_ASAP7_75t_L     g17341(.A1(new_n4544), .A2(\b[53] ), .B1(new_n4542), .B2(new_n8889), .Y(new_n17598));
  OAI221xp5_ASAP7_75t_L     g17342(.A1(new_n4536), .A2(new_n8569), .B1(new_n8249), .B2(new_n4781), .C(new_n17598), .Y(new_n17599));
  XNOR2x2_ASAP7_75t_L       g17343(.A(\a[38] ), .B(new_n17599), .Y(new_n17600));
  INVx1_ASAP7_75t_L         g17344(.A(new_n17600), .Y(new_n17601));
  AOI22xp33_ASAP7_75t_L     g17345(.A1(new_n6822), .A2(\b[44] ), .B1(new_n6819), .B2(new_n7055), .Y(new_n17602));
  OAI221xp5_ASAP7_75t_L     g17346(.A1(new_n7392), .A2(new_n6195), .B1(new_n5680), .B2(new_n7115), .C(new_n17602), .Y(new_n17603));
  XNOR2x2_ASAP7_75t_L       g17347(.A(\a[47] ), .B(new_n17603), .Y(new_n17604));
  INVx1_ASAP7_75t_L         g17348(.A(new_n17604), .Y(new_n17605));
  AOI22xp33_ASAP7_75t_L     g17349(.A1(new_n7659), .A2(\b[41] ), .B1(new_n7656), .B2(new_n5669), .Y(new_n17606));
  OAI221xp5_ASAP7_75t_L     g17350(.A1(new_n8326), .A2(new_n5186), .B1(new_n5166), .B2(new_n7994), .C(new_n17606), .Y(new_n17607));
  XNOR2x2_ASAP7_75t_L       g17351(.A(\a[50] ), .B(new_n17607), .Y(new_n17608));
  AOI22xp33_ASAP7_75t_L     g17352(.A1(new_n9623), .A2(\b[35] ), .B1(new_n9620), .B2(new_n5649), .Y(new_n17609));
  OAI221xp5_ASAP7_75t_L     g17353(.A1(new_n10280), .A2(new_n3827), .B1(new_n3807), .B2(new_n12010), .C(new_n17609), .Y(new_n17610));
  XNOR2x2_ASAP7_75t_L       g17354(.A(\a[56] ), .B(new_n17610), .Y(new_n17611));
  INVx1_ASAP7_75t_L         g17355(.A(new_n17611), .Y(new_n17612));
  AOI22xp33_ASAP7_75t_L     g17356(.A1(new_n10594), .A2(\b[32] ), .B1(new_n10591), .B2(new_n3450), .Y(new_n17613));
  OAI221xp5_ASAP7_75t_L     g17357(.A1(new_n11335), .A2(new_n3419), .B1(new_n3212), .B2(new_n11330), .C(new_n17613), .Y(new_n17614));
  XNOR2x2_ASAP7_75t_L       g17358(.A(\a[59] ), .B(new_n17614), .Y(new_n17615));
  INVx1_ASAP7_75t_L         g17359(.A(new_n17446), .Y(new_n17616));
  NOR2xp33_ASAP7_75t_L      g17360(.A(new_n2180), .B(new_n12671), .Y(new_n17617));
  O2A1O1Ixp33_ASAP7_75t_L   g17361(.A1(new_n12353), .A2(new_n12355), .B(\b[26] ), .C(new_n17617), .Y(new_n17618));
  A2O1A1Ixp33_ASAP7_75t_L   g17362(.A1(new_n12669), .A2(\b[25] ), .B(new_n17436), .C(new_n17618), .Y(new_n17619));
  A2O1A1Ixp33_ASAP7_75t_L   g17363(.A1(\b[26] ), .A2(new_n12669), .B(new_n17617), .C(new_n17439), .Y(new_n17620));
  NAND2xp33_ASAP7_75t_L     g17364(.A(new_n17620), .B(new_n17619), .Y(new_n17621));
  AOI22xp33_ASAP7_75t_L     g17365(.A1(new_n11647), .A2(\b[28] ), .B1(\b[29] ), .B2(new_n11656), .Y(new_n17622));
  OAI221xp5_ASAP7_75t_L     g17366(.A1(new_n13003), .A2(new_n2650), .B1(new_n12022), .B2(new_n2881), .C(new_n17622), .Y(new_n17623));
  XNOR2x2_ASAP7_75t_L       g17367(.A(\a[62] ), .B(new_n17623), .Y(new_n17624));
  NOR2xp33_ASAP7_75t_L      g17368(.A(new_n17621), .B(new_n17624), .Y(new_n17625));
  AND2x2_ASAP7_75t_L        g17369(.A(new_n17621), .B(new_n17624), .Y(new_n17626));
  NOR2xp33_ASAP7_75t_L      g17370(.A(new_n17625), .B(new_n17626), .Y(new_n17627));
  A2O1A1Ixp33_ASAP7_75t_L   g17371(.A1(new_n17616), .A2(new_n17438), .B(new_n17441), .C(new_n17627), .Y(new_n17628));
  OAI211xp5_ASAP7_75t_L     g17372(.A1(new_n17625), .A2(new_n17626), .B(new_n17448), .C(new_n17442), .Y(new_n17629));
  NAND2xp33_ASAP7_75t_L     g17373(.A(new_n17629), .B(new_n17628), .Y(new_n17630));
  OR2x4_ASAP7_75t_L         g17374(.A(new_n17615), .B(new_n17630), .Y(new_n17631));
  NAND2xp33_ASAP7_75t_L     g17375(.A(new_n17615), .B(new_n17630), .Y(new_n17632));
  AND2x2_ASAP7_75t_L        g17376(.A(new_n17632), .B(new_n17631), .Y(new_n17633));
  INVx1_ASAP7_75t_L         g17377(.A(new_n17633), .Y(new_n17634));
  A2O1A1Ixp33_ASAP7_75t_L   g17378(.A1(new_n17448), .A2(new_n17449), .B(new_n17453), .C(new_n17459), .Y(new_n17635));
  NOR2xp33_ASAP7_75t_L      g17379(.A(new_n17635), .B(new_n17634), .Y(new_n17636));
  O2A1O1Ixp33_ASAP7_75t_L   g17380(.A1(new_n17453), .A2(new_n17450), .B(new_n17459), .C(new_n17633), .Y(new_n17637));
  NOR2xp33_ASAP7_75t_L      g17381(.A(new_n17637), .B(new_n17636), .Y(new_n17638));
  NAND2xp33_ASAP7_75t_L     g17382(.A(new_n17612), .B(new_n17638), .Y(new_n17639));
  INVx1_ASAP7_75t_L         g17383(.A(new_n17639), .Y(new_n17640));
  NOR2xp33_ASAP7_75t_L      g17384(.A(new_n17612), .B(new_n17638), .Y(new_n17641));
  NOR2xp33_ASAP7_75t_L      g17385(.A(new_n17641), .B(new_n17640), .Y(new_n17642));
  NAND3xp33_ASAP7_75t_L     g17386(.A(new_n17471), .B(new_n17464), .C(new_n17642), .Y(new_n17643));
  O2A1O1Ixp33_ASAP7_75t_L   g17387(.A1(new_n17466), .A2(new_n17472), .B(new_n17464), .C(new_n17642), .Y(new_n17644));
  INVx1_ASAP7_75t_L         g17388(.A(new_n17644), .Y(new_n17645));
  AOI22xp33_ASAP7_75t_L     g17389(.A1(new_n8645), .A2(\b[38] ), .B1(new_n8642), .B2(new_n4923), .Y(new_n17646));
  OAI221xp5_ASAP7_75t_L     g17390(.A1(new_n9322), .A2(new_n4701), .B1(new_n4465), .B2(new_n8965), .C(new_n17646), .Y(new_n17647));
  XNOR2x2_ASAP7_75t_L       g17391(.A(\a[53] ), .B(new_n17647), .Y(new_n17648));
  NAND3xp33_ASAP7_75t_L     g17392(.A(new_n17645), .B(new_n17643), .C(new_n17648), .Y(new_n17649));
  AO21x2_ASAP7_75t_L        g17393(.A1(new_n17643), .A2(new_n17645), .B(new_n17648), .Y(new_n17650));
  AND2x2_ASAP7_75t_L        g17394(.A(new_n17649), .B(new_n17650), .Y(new_n17651));
  O2A1O1Ixp33_ASAP7_75t_L   g17395(.A1(new_n17483), .A2(new_n17480), .B(new_n17478), .C(new_n17651), .Y(new_n17652));
  O2A1O1Ixp33_ASAP7_75t_L   g17396(.A1(new_n17334), .A2(new_n17340), .B(new_n17477), .C(new_n17485), .Y(new_n17653));
  AND2x2_ASAP7_75t_L        g17397(.A(new_n17651), .B(new_n17653), .Y(new_n17654));
  NOR2xp33_ASAP7_75t_L      g17398(.A(new_n17652), .B(new_n17654), .Y(new_n17655));
  XOR2x2_ASAP7_75t_L        g17399(.A(new_n17608), .B(new_n17655), .Y(new_n17656));
  O2A1O1Ixp33_ASAP7_75t_L   g17400(.A1(new_n17432), .A2(new_n17489), .B(new_n17487), .C(new_n17656), .Y(new_n17657));
  INVx1_ASAP7_75t_L         g17401(.A(new_n17657), .Y(new_n17658));
  INVx1_ASAP7_75t_L         g17402(.A(new_n17491), .Y(new_n17659));
  A2O1A1O1Ixp25_ASAP7_75t_L g17403(.A1(new_n17346), .A2(new_n17342), .B(new_n17350), .C(new_n17486), .D(new_n17659), .Y(new_n17660));
  NAND2xp33_ASAP7_75t_L     g17404(.A(new_n17656), .B(new_n17660), .Y(new_n17661));
  NAND3xp33_ASAP7_75t_L     g17405(.A(new_n17661), .B(new_n17658), .C(new_n17605), .Y(new_n17662));
  INVx1_ASAP7_75t_L         g17406(.A(new_n17662), .Y(new_n17663));
  AOI21xp33_ASAP7_75t_L     g17407(.A1(new_n17661), .A2(new_n17658), .B(new_n17605), .Y(new_n17664));
  NOR2xp33_ASAP7_75t_L      g17408(.A(new_n17664), .B(new_n17663), .Y(new_n17665));
  NAND3xp33_ASAP7_75t_L     g17409(.A(new_n17665), .B(new_n17502), .C(new_n17498), .Y(new_n17666));
  O2A1O1Ixp33_ASAP7_75t_L   g17410(.A1(new_n17496), .A2(new_n17493), .B(new_n17502), .C(new_n17665), .Y(new_n17667));
  INVx1_ASAP7_75t_L         g17411(.A(new_n17667), .Y(new_n17668));
  AOI22xp33_ASAP7_75t_L     g17412(.A1(new_n6002), .A2(\b[47] ), .B1(new_n5999), .B2(new_n7323), .Y(new_n17669));
  OAI221xp5_ASAP7_75t_L     g17413(.A1(new_n6544), .A2(new_n7033), .B1(new_n6756), .B2(new_n6309), .C(new_n17669), .Y(new_n17670));
  XNOR2x2_ASAP7_75t_L       g17414(.A(\a[44] ), .B(new_n17670), .Y(new_n17671));
  NAND3xp33_ASAP7_75t_L     g17415(.A(new_n17668), .B(new_n17666), .C(new_n17671), .Y(new_n17672));
  INVx1_ASAP7_75t_L         g17416(.A(new_n17672), .Y(new_n17673));
  AOI21xp33_ASAP7_75t_L     g17417(.A1(new_n17668), .A2(new_n17666), .B(new_n17671), .Y(new_n17674));
  NOR2xp33_ASAP7_75t_L      g17418(.A(new_n17674), .B(new_n17673), .Y(new_n17675));
  A2O1A1Ixp33_ASAP7_75t_L   g17419(.A1(new_n17508), .A2(new_n17511), .B(new_n17506), .C(new_n17675), .Y(new_n17676));
  NAND2xp33_ASAP7_75t_L     g17420(.A(new_n17507), .B(new_n17512), .Y(new_n17677));
  NOR2xp33_ASAP7_75t_L      g17421(.A(new_n17677), .B(new_n17675), .Y(new_n17678));
  INVx1_ASAP7_75t_L         g17422(.A(new_n17678), .Y(new_n17679));
  NAND2xp33_ASAP7_75t_L     g17423(.A(new_n17676), .B(new_n17679), .Y(new_n17680));
  AOI22xp33_ASAP7_75t_L     g17424(.A1(new_n5249), .A2(\b[50] ), .B1(new_n5247), .B2(new_n8235), .Y(new_n17681));
  OAI221xp5_ASAP7_75t_L     g17425(.A1(new_n5241), .A2(new_n7907), .B1(new_n7333), .B2(new_n5521), .C(new_n17681), .Y(new_n17682));
  XNOR2x2_ASAP7_75t_L       g17426(.A(\a[41] ), .B(new_n17682), .Y(new_n17683));
  NAND2xp33_ASAP7_75t_L     g17427(.A(new_n17683), .B(new_n17680), .Y(new_n17684));
  NOR2xp33_ASAP7_75t_L      g17428(.A(new_n17683), .B(new_n17680), .Y(new_n17685));
  INVx1_ASAP7_75t_L         g17429(.A(new_n17685), .Y(new_n17686));
  NAND2xp33_ASAP7_75t_L     g17430(.A(new_n17684), .B(new_n17686), .Y(new_n17687));
  NAND2xp33_ASAP7_75t_L     g17431(.A(new_n17514), .B(new_n17523), .Y(new_n17688));
  XOR2x2_ASAP7_75t_L        g17432(.A(new_n17688), .B(new_n17687), .Y(new_n17689));
  AND2x2_ASAP7_75t_L        g17433(.A(new_n17601), .B(new_n17689), .Y(new_n17690));
  NOR2xp33_ASAP7_75t_L      g17434(.A(new_n17601), .B(new_n17689), .Y(new_n17691));
  NOR2xp33_ASAP7_75t_L      g17435(.A(new_n17691), .B(new_n17690), .Y(new_n17692));
  INVx1_ASAP7_75t_L         g17436(.A(new_n17692), .Y(new_n17693));
  NOR3xp33_ASAP7_75t_L      g17437(.A(new_n17693), .B(new_n17535), .C(new_n17527), .Y(new_n17694));
  O2A1O1Ixp33_ASAP7_75t_L   g17438(.A1(new_n17530), .A2(new_n17534), .B(new_n17528), .C(new_n17692), .Y(new_n17695));
  NOR2xp33_ASAP7_75t_L      g17439(.A(new_n17695), .B(new_n17694), .Y(new_n17696));
  NOR2xp33_ASAP7_75t_L      g17440(.A(new_n17597), .B(new_n17696), .Y(new_n17697));
  AND2x2_ASAP7_75t_L        g17441(.A(new_n17597), .B(new_n17696), .Y(new_n17698));
  OR2x4_ASAP7_75t_L         g17442(.A(new_n17697), .B(new_n17698), .Y(new_n17699));
  OR3x1_ASAP7_75t_L         g17443(.A(new_n17699), .B(new_n17593), .C(new_n17594), .Y(new_n17700));
  OAI21xp33_ASAP7_75t_L     g17444(.A1(new_n17593), .A2(new_n17594), .B(new_n17699), .Y(new_n17701));
  NAND2xp33_ASAP7_75t_L     g17445(.A(new_n17701), .B(new_n17700), .Y(new_n17702));
  NOR2xp33_ASAP7_75t_L      g17446(.A(new_n17586), .B(new_n17702), .Y(new_n17703));
  NAND2xp33_ASAP7_75t_L     g17447(.A(new_n17586), .B(new_n17702), .Y(new_n17704));
  INVx1_ASAP7_75t_L         g17448(.A(new_n17704), .Y(new_n17705));
  NOR2xp33_ASAP7_75t_L      g17449(.A(new_n17703), .B(new_n17705), .Y(new_n17706));
  INVx1_ASAP7_75t_L         g17450(.A(new_n17417), .Y(new_n17707));
  MAJIxp5_ASAP7_75t_L       g17451(.A(new_n17556), .B(new_n17416), .C(new_n17707), .Y(new_n17708));
  O2A1O1Ixp33_ASAP7_75t_L   g17452(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n2233), .Y(new_n17709));
  O2A1O1Ixp33_ASAP7_75t_L   g17453(.A1(new_n2386), .A2(new_n17709), .B(\b[63] ), .C(new_n2223), .Y(new_n17710));
  A2O1A1O1Ixp25_ASAP7_75t_L g17454(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n2226), .D(new_n2386), .Y(new_n17711));
  NOR3xp33_ASAP7_75t_L      g17455(.A(new_n17711), .B(new_n12599), .C(\a[26] ), .Y(new_n17712));
  NOR2xp33_ASAP7_75t_L      g17456(.A(new_n17710), .B(new_n17712), .Y(new_n17713));
  INVx1_ASAP7_75t_L         g17457(.A(new_n17713), .Y(new_n17714));
  NAND2xp33_ASAP7_75t_L     g17458(.A(new_n17714), .B(new_n17708), .Y(new_n17715));
  INVx1_ASAP7_75t_L         g17459(.A(new_n17715), .Y(new_n17716));
  NOR2xp33_ASAP7_75t_L      g17460(.A(new_n17714), .B(new_n17708), .Y(new_n17717));
  NOR2xp33_ASAP7_75t_L      g17461(.A(new_n17717), .B(new_n17716), .Y(new_n17718));
  NAND2xp33_ASAP7_75t_L     g17462(.A(new_n17718), .B(new_n17706), .Y(new_n17719));
  OAI22xp33_ASAP7_75t_L     g17463(.A1(new_n17705), .A2(new_n17703), .B1(new_n17717), .B2(new_n17716), .Y(new_n17720));
  NAND2xp33_ASAP7_75t_L     g17464(.A(new_n17720), .B(new_n17719), .Y(new_n17721));
  INVx1_ASAP7_75t_L         g17465(.A(new_n17721), .Y(new_n17722));
  NAND2xp33_ASAP7_75t_L     g17466(.A(new_n17578), .B(new_n17722), .Y(new_n17723));
  INVx1_ASAP7_75t_L         g17467(.A(new_n17723), .Y(new_n17724));
  NOR2xp33_ASAP7_75t_L      g17468(.A(new_n17578), .B(new_n17722), .Y(new_n17725));
  NOR2xp33_ASAP7_75t_L      g17469(.A(new_n17725), .B(new_n17724), .Y(new_n17726));
  A2O1A1Ixp33_ASAP7_75t_L   g17470(.A1(new_n17573), .A2(new_n17574), .B(new_n17568), .C(new_n17726), .Y(new_n17727));
  INVx1_ASAP7_75t_L         g17471(.A(new_n17727), .Y(new_n17728));
  A2O1A1Ixp33_ASAP7_75t_L   g17472(.A1(new_n17406), .A2(new_n17402), .B(new_n17571), .C(new_n17569), .Y(new_n17729));
  NOR2xp33_ASAP7_75t_L      g17473(.A(new_n17726), .B(new_n17729), .Y(new_n17730));
  NOR2xp33_ASAP7_75t_L      g17474(.A(new_n17728), .B(new_n17730), .Y(\f[89] ));
  NAND2xp33_ASAP7_75t_L     g17475(.A(new_n17715), .B(new_n17719), .Y(new_n17732));
  NAND2xp33_ASAP7_75t_L     g17476(.A(\b[63] ), .B(new_n2702), .Y(new_n17733));
  A2O1A1Ixp33_ASAP7_75t_L   g17477(.A1(new_n12607), .A2(new_n12603), .B(new_n2707), .C(new_n17733), .Y(new_n17734));
  AOI221xp5_ASAP7_75t_L     g17478(.A1(\b[61] ), .A2(new_n2931), .B1(\b[62] ), .B2(new_n2706), .C(new_n17734), .Y(new_n17735));
  XNOR2x2_ASAP7_75t_L       g17479(.A(new_n2697), .B(new_n17735), .Y(new_n17736));
  A2O1A1Ixp33_ASAP7_75t_L   g17480(.A1(new_n17702), .A2(new_n17586), .B(new_n17585), .C(new_n17736), .Y(new_n17737));
  INVx1_ASAP7_75t_L         g17481(.A(new_n17585), .Y(new_n17738));
  A2O1A1Ixp33_ASAP7_75t_L   g17482(.A1(new_n17700), .A2(new_n17701), .B(new_n17584), .C(new_n17738), .Y(new_n17739));
  INVx1_ASAP7_75t_L         g17483(.A(new_n17739), .Y(new_n17740));
  INVx1_ASAP7_75t_L         g17484(.A(new_n17736), .Y(new_n17741));
  NAND2xp33_ASAP7_75t_L     g17485(.A(new_n17741), .B(new_n17740), .Y(new_n17742));
  NAND2xp33_ASAP7_75t_L     g17486(.A(new_n17742), .B(new_n17737), .Y(new_n17743));
  INVx1_ASAP7_75t_L         g17487(.A(new_n17690), .Y(new_n17744));
  AOI22xp33_ASAP7_75t_L     g17488(.A1(new_n4544), .A2(\b[54] ), .B1(new_n4542), .B2(new_n9208), .Y(new_n17745));
  OAI221xp5_ASAP7_75t_L     g17489(.A1(new_n4536), .A2(new_n8882), .B1(new_n8569), .B2(new_n4781), .C(new_n17745), .Y(new_n17746));
  XNOR2x2_ASAP7_75t_L       g17490(.A(\a[38] ), .B(new_n17746), .Y(new_n17747));
  INVx1_ASAP7_75t_L         g17491(.A(new_n17747), .Y(new_n17748));
  INVx1_ASAP7_75t_L         g17492(.A(new_n17677), .Y(new_n17749));
  O2A1O1Ixp33_ASAP7_75t_L   g17493(.A1(new_n17673), .A2(new_n17674), .B(new_n17749), .C(new_n17685), .Y(new_n17750));
  INVx1_ASAP7_75t_L         g17494(.A(new_n17750), .Y(new_n17751));
  AOI22xp33_ASAP7_75t_L     g17495(.A1(new_n6822), .A2(\b[45] ), .B1(new_n6819), .B2(new_n6764), .Y(new_n17752));
  OAI221xp5_ASAP7_75t_L     g17496(.A1(new_n7392), .A2(new_n6220), .B1(new_n6195), .B2(new_n7115), .C(new_n17752), .Y(new_n17753));
  XNOR2x2_ASAP7_75t_L       g17497(.A(new_n6816), .B(new_n17753), .Y(new_n17754));
  AOI22xp33_ASAP7_75t_L     g17498(.A1(new_n10594), .A2(\b[33] ), .B1(new_n10591), .B2(new_n3813), .Y(new_n17755));
  OAI221xp5_ASAP7_75t_L     g17499(.A1(new_n11335), .A2(new_n3443), .B1(new_n3419), .B2(new_n11330), .C(new_n17755), .Y(new_n17756));
  XNOR2x2_ASAP7_75t_L       g17500(.A(\a[59] ), .B(new_n17756), .Y(new_n17757));
  AND3x1_ASAP7_75t_L        g17501(.A(new_n17631), .B(new_n17757), .C(new_n17628), .Y(new_n17758));
  O2A1O1Ixp33_ASAP7_75t_L   g17502(.A1(new_n17615), .A2(new_n17630), .B(new_n17628), .C(new_n17757), .Y(new_n17759));
  NOR2xp33_ASAP7_75t_L      g17503(.A(new_n17759), .B(new_n17758), .Y(new_n17760));
  NOR2xp33_ASAP7_75t_L      g17504(.A(new_n2477), .B(new_n12671), .Y(new_n17761));
  A2O1A1Ixp33_ASAP7_75t_L   g17505(.A1(new_n12669), .A2(\b[27] ), .B(new_n17761), .C(new_n2223), .Y(new_n17762));
  INVx1_ASAP7_75t_L         g17506(.A(new_n17762), .Y(new_n17763));
  O2A1O1Ixp33_ASAP7_75t_L   g17507(.A1(new_n12353), .A2(new_n12355), .B(\b[27] ), .C(new_n17761), .Y(new_n17764));
  NAND2xp33_ASAP7_75t_L     g17508(.A(\a[26] ), .B(new_n17764), .Y(new_n17765));
  INVx1_ASAP7_75t_L         g17509(.A(new_n17765), .Y(new_n17766));
  NOR2xp33_ASAP7_75t_L      g17510(.A(new_n17763), .B(new_n17766), .Y(new_n17767));
  A2O1A1Ixp33_ASAP7_75t_L   g17511(.A1(new_n12669), .A2(\b[26] ), .B(new_n17617), .C(new_n17767), .Y(new_n17768));
  OAI21xp33_ASAP7_75t_L     g17512(.A1(new_n17763), .A2(new_n17766), .B(new_n17618), .Y(new_n17769));
  NAND2xp33_ASAP7_75t_L     g17513(.A(new_n17769), .B(new_n17768), .Y(new_n17770));
  O2A1O1Ixp33_ASAP7_75t_L   g17514(.A1(new_n17621), .A2(new_n17624), .B(new_n17619), .C(new_n17770), .Y(new_n17771));
  A2O1A1O1Ixp25_ASAP7_75t_L g17515(.A1(new_n12669), .A2(\b[25] ), .B(new_n17436), .C(new_n17618), .D(new_n17625), .Y(new_n17772));
  NAND2xp33_ASAP7_75t_L     g17516(.A(new_n17770), .B(new_n17772), .Y(new_n17773));
  INVx1_ASAP7_75t_L         g17517(.A(new_n17773), .Y(new_n17774));
  NOR2xp33_ASAP7_75t_L      g17518(.A(new_n17771), .B(new_n17774), .Y(new_n17775));
  INVx1_ASAP7_75t_L         g17519(.A(new_n17775), .Y(new_n17776));
  AOI22xp33_ASAP7_75t_L     g17520(.A1(new_n11656), .A2(\b[30] ), .B1(new_n11654), .B2(new_n3219), .Y(new_n17777));
  OAI221xp5_ASAP7_75t_L     g17521(.A1(new_n12364), .A2(new_n2871), .B1(new_n2852), .B2(new_n13003), .C(new_n17777), .Y(new_n17778));
  XNOR2x2_ASAP7_75t_L       g17522(.A(\a[62] ), .B(new_n17778), .Y(new_n17779));
  INVx1_ASAP7_75t_L         g17523(.A(new_n17779), .Y(new_n17780));
  NOR2xp33_ASAP7_75t_L      g17524(.A(new_n17780), .B(new_n17776), .Y(new_n17781));
  INVx1_ASAP7_75t_L         g17525(.A(new_n17781), .Y(new_n17782));
  NAND2xp33_ASAP7_75t_L     g17526(.A(new_n17780), .B(new_n17776), .Y(new_n17783));
  AND2x2_ASAP7_75t_L        g17527(.A(new_n17783), .B(new_n17782), .Y(new_n17784));
  XNOR2x2_ASAP7_75t_L       g17528(.A(new_n17760), .B(new_n17784), .Y(new_n17785));
  AOI22xp33_ASAP7_75t_L     g17529(.A1(new_n9623), .A2(\b[36] ), .B1(new_n9620), .B2(new_n4473), .Y(new_n17786));
  OAI221xp5_ASAP7_75t_L     g17530(.A1(new_n10280), .A2(new_n4053), .B1(new_n3827), .B2(new_n12010), .C(new_n17786), .Y(new_n17787));
  XNOR2x2_ASAP7_75t_L       g17531(.A(\a[56] ), .B(new_n17787), .Y(new_n17788));
  INVx1_ASAP7_75t_L         g17532(.A(new_n17788), .Y(new_n17789));
  XNOR2x2_ASAP7_75t_L       g17533(.A(new_n17789), .B(new_n17785), .Y(new_n17790));
  INVx1_ASAP7_75t_L         g17534(.A(new_n17790), .Y(new_n17791));
  NOR3xp33_ASAP7_75t_L      g17535(.A(new_n17791), .B(new_n17640), .C(new_n17636), .Y(new_n17792));
  O2A1O1Ixp33_ASAP7_75t_L   g17536(.A1(new_n17634), .A2(new_n17635), .B(new_n17639), .C(new_n17790), .Y(new_n17793));
  NOR2xp33_ASAP7_75t_L      g17537(.A(new_n17793), .B(new_n17792), .Y(new_n17794));
  AOI22xp33_ASAP7_75t_L     g17538(.A1(new_n8645), .A2(\b[39] ), .B1(new_n8642), .B2(new_n5174), .Y(new_n17795));
  OAI221xp5_ASAP7_75t_L     g17539(.A1(new_n9322), .A2(new_n4915), .B1(new_n4701), .B2(new_n8965), .C(new_n17795), .Y(new_n17796));
  XNOR2x2_ASAP7_75t_L       g17540(.A(\a[53] ), .B(new_n17796), .Y(new_n17797));
  INVx1_ASAP7_75t_L         g17541(.A(new_n17797), .Y(new_n17798));
  XNOR2x2_ASAP7_75t_L       g17542(.A(new_n17798), .B(new_n17794), .Y(new_n17799));
  A2O1A1Ixp33_ASAP7_75t_L   g17543(.A1(new_n17648), .A2(new_n17643), .B(new_n17644), .C(new_n17799), .Y(new_n17800));
  A2O1A1Ixp33_ASAP7_75t_L   g17544(.A1(new_n17471), .A2(new_n17464), .B(new_n17642), .C(new_n17649), .Y(new_n17801));
  NOR2xp33_ASAP7_75t_L      g17545(.A(new_n17801), .B(new_n17799), .Y(new_n17802));
  INVx1_ASAP7_75t_L         g17546(.A(new_n17802), .Y(new_n17803));
  NAND2xp33_ASAP7_75t_L     g17547(.A(new_n17800), .B(new_n17803), .Y(new_n17804));
  AOI22xp33_ASAP7_75t_L     g17548(.A1(new_n7659), .A2(\b[42] ), .B1(new_n7656), .B2(new_n5688), .Y(new_n17805));
  OAI221xp5_ASAP7_75t_L     g17549(.A1(new_n8326), .A2(new_n5666), .B1(new_n5186), .B2(new_n7994), .C(new_n17805), .Y(new_n17806));
  XNOR2x2_ASAP7_75t_L       g17550(.A(\a[50] ), .B(new_n17806), .Y(new_n17807));
  XNOR2x2_ASAP7_75t_L       g17551(.A(new_n17807), .B(new_n17804), .Y(new_n17808));
  AOI21xp33_ASAP7_75t_L     g17552(.A1(new_n17655), .A2(new_n17608), .B(new_n17654), .Y(new_n17809));
  XNOR2x2_ASAP7_75t_L       g17553(.A(new_n17808), .B(new_n17809), .Y(new_n17810));
  XOR2x2_ASAP7_75t_L        g17554(.A(new_n17754), .B(new_n17810), .Y(new_n17811));
  INVx1_ASAP7_75t_L         g17555(.A(new_n17811), .Y(new_n17812));
  NAND3xp33_ASAP7_75t_L     g17556(.A(new_n17812), .B(new_n17662), .C(new_n17658), .Y(new_n17813));
  O2A1O1Ixp33_ASAP7_75t_L   g17557(.A1(new_n17660), .A2(new_n17656), .B(new_n17662), .C(new_n17812), .Y(new_n17814));
  INVx1_ASAP7_75t_L         g17558(.A(new_n17814), .Y(new_n17815));
  NAND2xp33_ASAP7_75t_L     g17559(.A(new_n17813), .B(new_n17815), .Y(new_n17816));
  AOI22xp33_ASAP7_75t_L     g17560(.A1(new_n6002), .A2(\b[48] ), .B1(new_n5999), .B2(new_n7341), .Y(new_n17817));
  OAI221xp5_ASAP7_75t_L     g17561(.A1(new_n6544), .A2(new_n7316), .B1(new_n7033), .B2(new_n6309), .C(new_n17817), .Y(new_n17818));
  XNOR2x2_ASAP7_75t_L       g17562(.A(\a[44] ), .B(new_n17818), .Y(new_n17819));
  XNOR2x2_ASAP7_75t_L       g17563(.A(new_n17819), .B(new_n17816), .Y(new_n17820));
  A2O1A1Ixp33_ASAP7_75t_L   g17564(.A1(new_n17671), .A2(new_n17666), .B(new_n17667), .C(new_n17820), .Y(new_n17821));
  OR3x1_ASAP7_75t_L         g17565(.A(new_n17673), .B(new_n17667), .C(new_n17820), .Y(new_n17822));
  NAND2xp33_ASAP7_75t_L     g17566(.A(new_n17821), .B(new_n17822), .Y(new_n17823));
  AOI22xp33_ASAP7_75t_L     g17567(.A1(new_n5249), .A2(\b[51] ), .B1(new_n5247), .B2(new_n8257), .Y(new_n17824));
  OAI221xp5_ASAP7_75t_L     g17568(.A1(new_n5241), .A2(new_n8228), .B1(new_n7907), .B2(new_n5521), .C(new_n17824), .Y(new_n17825));
  XNOR2x2_ASAP7_75t_L       g17569(.A(\a[41] ), .B(new_n17825), .Y(new_n17826));
  NOR2xp33_ASAP7_75t_L      g17570(.A(new_n17826), .B(new_n17823), .Y(new_n17827));
  INVx1_ASAP7_75t_L         g17571(.A(new_n17827), .Y(new_n17828));
  NAND2xp33_ASAP7_75t_L     g17572(.A(new_n17826), .B(new_n17823), .Y(new_n17829));
  AOI21xp33_ASAP7_75t_L     g17573(.A1(new_n17829), .A2(new_n17828), .B(new_n17751), .Y(new_n17830));
  NAND2xp33_ASAP7_75t_L     g17574(.A(new_n17829), .B(new_n17828), .Y(new_n17831));
  O2A1O1Ixp33_ASAP7_75t_L   g17575(.A1(new_n17680), .A2(new_n17683), .B(new_n17679), .C(new_n17831), .Y(new_n17832));
  NOR2xp33_ASAP7_75t_L      g17576(.A(new_n17832), .B(new_n17830), .Y(new_n17833));
  XNOR2x2_ASAP7_75t_L       g17577(.A(new_n17748), .B(new_n17833), .Y(new_n17834));
  O2A1O1Ixp33_ASAP7_75t_L   g17578(.A1(new_n17687), .A2(new_n17688), .B(new_n17744), .C(new_n17834), .Y(new_n17835));
  OA211x2_ASAP7_75t_L       g17579(.A1(new_n17688), .A2(new_n17687), .B(new_n17834), .C(new_n17744), .Y(new_n17836));
  NOR2xp33_ASAP7_75t_L      g17580(.A(new_n17835), .B(new_n17836), .Y(new_n17837));
  AOI22xp33_ASAP7_75t_L     g17581(.A1(new_n3884), .A2(\b[57] ), .B1(new_n3881), .B2(new_n10495), .Y(new_n17838));
  OAI221xp5_ASAP7_75t_L     g17582(.A1(new_n4312), .A2(new_n10178), .B1(new_n9534), .B2(new_n4986), .C(new_n17838), .Y(new_n17839));
  XNOR2x2_ASAP7_75t_L       g17583(.A(\a[35] ), .B(new_n17839), .Y(new_n17840));
  INVx1_ASAP7_75t_L         g17584(.A(new_n17840), .Y(new_n17841));
  XNOR2x2_ASAP7_75t_L       g17585(.A(new_n17841), .B(new_n17837), .Y(new_n17842));
  A2O1A1Ixp33_ASAP7_75t_L   g17586(.A1(new_n17696), .A2(new_n17597), .B(new_n17695), .C(new_n17842), .Y(new_n17843));
  OR3x1_ASAP7_75t_L         g17587(.A(new_n17842), .B(new_n17695), .C(new_n17698), .Y(new_n17844));
  NAND2xp33_ASAP7_75t_L     g17588(.A(new_n17843), .B(new_n17844), .Y(new_n17845));
  AOI22xp33_ASAP7_75t_L     g17589(.A1(new_n3256), .A2(\b[60] ), .B1(new_n3254), .B2(new_n11234), .Y(new_n17846));
  OAI221xp5_ASAP7_75t_L     g17590(.A1(new_n3248), .A2(new_n10881), .B1(new_n10848), .B2(new_n3492), .C(new_n17846), .Y(new_n17847));
  XNOR2x2_ASAP7_75t_L       g17591(.A(\a[32] ), .B(new_n17847), .Y(new_n17848));
  OAI21xp33_ASAP7_75t_L     g17592(.A1(new_n17590), .A2(new_n17592), .B(new_n17700), .Y(new_n17849));
  NAND2xp33_ASAP7_75t_L     g17593(.A(new_n17848), .B(new_n17849), .Y(new_n17850));
  INVx1_ASAP7_75t_L         g17594(.A(new_n17850), .Y(new_n17851));
  NOR2xp33_ASAP7_75t_L      g17595(.A(new_n17848), .B(new_n17849), .Y(new_n17852));
  NOR2xp33_ASAP7_75t_L      g17596(.A(new_n17852), .B(new_n17851), .Y(new_n17853));
  NOR2xp33_ASAP7_75t_L      g17597(.A(new_n17845), .B(new_n17853), .Y(new_n17854));
  NAND2xp33_ASAP7_75t_L     g17598(.A(new_n17845), .B(new_n17853), .Y(new_n17855));
  INVx1_ASAP7_75t_L         g17599(.A(new_n17855), .Y(new_n17856));
  NOR2xp33_ASAP7_75t_L      g17600(.A(new_n17854), .B(new_n17856), .Y(new_n17857));
  XNOR2x2_ASAP7_75t_L       g17601(.A(new_n17743), .B(new_n17857), .Y(new_n17858));
  NOR2xp33_ASAP7_75t_L      g17602(.A(new_n17732), .B(new_n17858), .Y(new_n17859));
  A2O1A1Ixp33_ASAP7_75t_L   g17603(.A1(new_n17718), .A2(new_n17706), .B(new_n17716), .C(new_n17858), .Y(new_n17860));
  INVx1_ASAP7_75t_L         g17604(.A(new_n17860), .Y(new_n17861));
  NOR2xp33_ASAP7_75t_L      g17605(.A(new_n17859), .B(new_n17861), .Y(new_n17862));
  A2O1A1Ixp33_ASAP7_75t_L   g17606(.A1(new_n17722), .A2(new_n17578), .B(new_n17728), .C(new_n17862), .Y(new_n17863));
  INVx1_ASAP7_75t_L         g17607(.A(new_n17863), .Y(new_n17864));
  NOR3xp33_ASAP7_75t_L      g17608(.A(new_n17862), .B(new_n17728), .C(new_n17724), .Y(new_n17865));
  NOR2xp33_ASAP7_75t_L      g17609(.A(new_n17865), .B(new_n17864), .Y(\f[90] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17610(.A1(new_n17574), .A2(new_n17573), .B(new_n17568), .C(new_n17726), .D(new_n17724), .Y(new_n17867));
  A2O1A1O1Ixp25_ASAP7_75t_L g17611(.A1(new_n17701), .A2(new_n17700), .B(new_n17584), .C(new_n17738), .D(new_n17736), .Y(new_n17868));
  O2A1O1Ixp33_ASAP7_75t_L   g17612(.A1(new_n17854), .A2(new_n17856), .B(new_n17743), .C(new_n17868), .Y(new_n17869));
  A2O1A1Ixp33_ASAP7_75t_L   g17613(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n2700), .Y(new_n17870));
  AOI22xp33_ASAP7_75t_L     g17614(.A1(new_n2706), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2931), .Y(new_n17871));
  NAND3xp33_ASAP7_75t_L     g17615(.A(new_n17870), .B(\a[29] ), .C(new_n17871), .Y(new_n17872));
  INVx1_ASAP7_75t_L         g17616(.A(new_n17872), .Y(new_n17873));
  A2O1A1O1Ixp25_ASAP7_75t_L g17617(.A1(new_n13507), .A2(new_n13506), .B(new_n2707), .C(new_n17871), .D(\a[29] ), .Y(new_n17874));
  NOR2xp33_ASAP7_75t_L      g17618(.A(new_n17874), .B(new_n17873), .Y(new_n17875));
  A2O1A1Ixp33_ASAP7_75t_L   g17619(.A1(new_n17843), .A2(new_n17844), .B(new_n17852), .C(new_n17850), .Y(new_n17876));
  NOR2xp33_ASAP7_75t_L      g17620(.A(new_n17875), .B(new_n17876), .Y(new_n17877));
  INVx1_ASAP7_75t_L         g17621(.A(new_n17877), .Y(new_n17878));
  A2O1A1Ixp33_ASAP7_75t_L   g17622(.A1(new_n17853), .A2(new_n17845), .B(new_n17851), .C(new_n17875), .Y(new_n17879));
  AND2x2_ASAP7_75t_L        g17623(.A(new_n17878), .B(new_n17879), .Y(new_n17880));
  AOI22xp33_ASAP7_75t_L     g17624(.A1(new_n3256), .A2(\b[61] ), .B1(new_n3254), .B2(new_n11919), .Y(new_n17881));
  OAI221xp5_ASAP7_75t_L     g17625(.A1(new_n3248), .A2(new_n11226), .B1(new_n10881), .B2(new_n3492), .C(new_n17881), .Y(new_n17882));
  XNOR2x2_ASAP7_75t_L       g17626(.A(\a[32] ), .B(new_n17882), .Y(new_n17883));
  O2A1O1Ixp33_ASAP7_75t_L   g17627(.A1(new_n17527), .A2(new_n17535), .B(new_n17693), .C(new_n17698), .Y(new_n17884));
  INVx1_ASAP7_75t_L         g17628(.A(new_n17884), .Y(new_n17885));
  NOR2xp33_ASAP7_75t_L      g17629(.A(new_n17842), .B(new_n17885), .Y(new_n17886));
  AOI21xp33_ASAP7_75t_L     g17630(.A1(new_n17841), .A2(new_n17837), .B(new_n17886), .Y(new_n17887));
  NAND2xp33_ASAP7_75t_L     g17631(.A(new_n17883), .B(new_n17887), .Y(new_n17888));
  INVx1_ASAP7_75t_L         g17632(.A(new_n17883), .Y(new_n17889));
  A2O1A1Ixp33_ASAP7_75t_L   g17633(.A1(new_n17841), .A2(new_n17837), .B(new_n17886), .C(new_n17889), .Y(new_n17890));
  NAND2xp33_ASAP7_75t_L     g17634(.A(new_n17754), .B(new_n17810), .Y(new_n17891));
  AOI22xp33_ASAP7_75t_L     g17635(.A1(new_n8645), .A2(\b[40] ), .B1(new_n8642), .B2(new_n5194), .Y(new_n17892));
  OAI221xp5_ASAP7_75t_L     g17636(.A1(new_n9322), .A2(new_n5166), .B1(new_n4915), .B2(new_n8965), .C(new_n17892), .Y(new_n17893));
  XNOR2x2_ASAP7_75t_L       g17637(.A(\a[53] ), .B(new_n17893), .Y(new_n17894));
  AOI22xp33_ASAP7_75t_L     g17638(.A1(new_n9623), .A2(\b[37] ), .B1(new_n9620), .B2(new_n4709), .Y(new_n17895));
  OAI221xp5_ASAP7_75t_L     g17639(.A1(new_n10280), .A2(new_n4465), .B1(new_n4053), .B2(new_n12010), .C(new_n17895), .Y(new_n17896));
  XNOR2x2_ASAP7_75t_L       g17640(.A(\a[56] ), .B(new_n17896), .Y(new_n17897));
  INVx1_ASAP7_75t_L         g17641(.A(new_n17759), .Y(new_n17898));
  NOR2xp33_ASAP7_75t_L      g17642(.A(new_n2650), .B(new_n12671), .Y(new_n17899));
  A2O1A1O1Ixp25_ASAP7_75t_L g17643(.A1(new_n12669), .A2(\b[26] ), .B(new_n17617), .C(new_n17765), .D(new_n17763), .Y(new_n17900));
  A2O1A1Ixp33_ASAP7_75t_L   g17644(.A1(new_n12669), .A2(\b[28] ), .B(new_n17899), .C(new_n17900), .Y(new_n17901));
  O2A1O1Ixp33_ASAP7_75t_L   g17645(.A1(new_n12353), .A2(new_n12355), .B(\b[28] ), .C(new_n17899), .Y(new_n17902));
  INVx1_ASAP7_75t_L         g17646(.A(new_n17902), .Y(new_n17903));
  O2A1O1Ixp33_ASAP7_75t_L   g17647(.A1(new_n17618), .A2(new_n17766), .B(new_n17762), .C(new_n17903), .Y(new_n17904));
  INVx1_ASAP7_75t_L         g17648(.A(new_n17904), .Y(new_n17905));
  NAND2xp33_ASAP7_75t_L     g17649(.A(new_n17901), .B(new_n17905), .Y(new_n17906));
  NAND2xp33_ASAP7_75t_L     g17650(.A(\b[31] ), .B(new_n11656), .Y(new_n17907));
  OAI221xp5_ASAP7_75t_L     g17651(.A1(new_n3212), .A2(new_n12364), .B1(new_n12022), .B2(new_n4030), .C(new_n17907), .Y(new_n17908));
  AOI21xp33_ASAP7_75t_L     g17652(.A1(new_n12021), .A2(\b[29] ), .B(new_n17908), .Y(new_n17909));
  NAND2xp33_ASAP7_75t_L     g17653(.A(\a[62] ), .B(new_n17909), .Y(new_n17910));
  A2O1A1Ixp33_ASAP7_75t_L   g17654(.A1(\b[29] ), .A2(new_n12021), .B(new_n17908), .C(new_n11651), .Y(new_n17911));
  AND2x2_ASAP7_75t_L        g17655(.A(new_n17911), .B(new_n17910), .Y(new_n17912));
  NAND2xp33_ASAP7_75t_L     g17656(.A(new_n17906), .B(new_n17912), .Y(new_n17913));
  NOR2xp33_ASAP7_75t_L      g17657(.A(new_n17906), .B(new_n17912), .Y(new_n17914));
  INVx1_ASAP7_75t_L         g17658(.A(new_n17914), .Y(new_n17915));
  AND2x2_ASAP7_75t_L        g17659(.A(new_n17913), .B(new_n17915), .Y(new_n17916));
  NOR2xp33_ASAP7_75t_L      g17660(.A(new_n17774), .B(new_n17781), .Y(new_n17917));
  NAND2xp33_ASAP7_75t_L     g17661(.A(new_n17916), .B(new_n17917), .Y(new_n17918));
  O2A1O1Ixp33_ASAP7_75t_L   g17662(.A1(new_n17771), .A2(new_n17780), .B(new_n17773), .C(new_n17916), .Y(new_n17919));
  INVx1_ASAP7_75t_L         g17663(.A(new_n17919), .Y(new_n17920));
  AOI22xp33_ASAP7_75t_L     g17664(.A1(new_n10594), .A2(\b[34] ), .B1(new_n10591), .B2(new_n3833), .Y(new_n17921));
  OAI221xp5_ASAP7_75t_L     g17665(.A1(new_n11335), .A2(new_n3807), .B1(new_n3443), .B2(new_n11330), .C(new_n17921), .Y(new_n17922));
  XNOR2x2_ASAP7_75t_L       g17666(.A(\a[59] ), .B(new_n17922), .Y(new_n17923));
  NAND3xp33_ASAP7_75t_L     g17667(.A(new_n17918), .B(new_n17920), .C(new_n17923), .Y(new_n17924));
  AO21x2_ASAP7_75t_L        g17668(.A1(new_n17920), .A2(new_n17918), .B(new_n17923), .Y(new_n17925));
  AND2x2_ASAP7_75t_L        g17669(.A(new_n17924), .B(new_n17925), .Y(new_n17926));
  O2A1O1Ixp33_ASAP7_75t_L   g17670(.A1(new_n17758), .A2(new_n17784), .B(new_n17898), .C(new_n17926), .Y(new_n17927));
  INVx1_ASAP7_75t_L         g17671(.A(new_n17926), .Y(new_n17928));
  A2O1A1Ixp33_ASAP7_75t_L   g17672(.A1(new_n17782), .A2(new_n17783), .B(new_n17758), .C(new_n17898), .Y(new_n17929));
  NOR2xp33_ASAP7_75t_L      g17673(.A(new_n17929), .B(new_n17928), .Y(new_n17930));
  NOR2xp33_ASAP7_75t_L      g17674(.A(new_n17927), .B(new_n17930), .Y(new_n17931));
  NAND2xp33_ASAP7_75t_L     g17675(.A(new_n17897), .B(new_n17931), .Y(new_n17932));
  INVx1_ASAP7_75t_L         g17676(.A(new_n17897), .Y(new_n17933));
  OAI21xp33_ASAP7_75t_L     g17677(.A1(new_n17927), .A2(new_n17930), .B(new_n17933), .Y(new_n17934));
  AND2x2_ASAP7_75t_L        g17678(.A(new_n17934), .B(new_n17932), .Y(new_n17935));
  A2O1A1Ixp33_ASAP7_75t_L   g17679(.A1(new_n17789), .A2(new_n17785), .B(new_n17793), .C(new_n17935), .Y(new_n17936));
  AOI21xp33_ASAP7_75t_L     g17680(.A1(new_n17789), .A2(new_n17785), .B(new_n17793), .Y(new_n17937));
  INVx1_ASAP7_75t_L         g17681(.A(new_n17935), .Y(new_n17938));
  NAND2xp33_ASAP7_75t_L     g17682(.A(new_n17937), .B(new_n17938), .Y(new_n17939));
  AND2x2_ASAP7_75t_L        g17683(.A(new_n17936), .B(new_n17939), .Y(new_n17940));
  XOR2x2_ASAP7_75t_L        g17684(.A(new_n17894), .B(new_n17940), .Y(new_n17941));
  A2O1A1Ixp33_ASAP7_75t_L   g17685(.A1(new_n17798), .A2(new_n17794), .B(new_n17802), .C(new_n17941), .Y(new_n17942));
  AOI211xp5_ASAP7_75t_L     g17686(.A1(new_n17794), .A2(new_n17798), .B(new_n17802), .C(new_n17941), .Y(new_n17943));
  INVx1_ASAP7_75t_L         g17687(.A(new_n17943), .Y(new_n17944));
  NAND2xp33_ASAP7_75t_L     g17688(.A(new_n17942), .B(new_n17944), .Y(new_n17945));
  NAND2xp33_ASAP7_75t_L     g17689(.A(\b[43] ), .B(new_n7659), .Y(new_n17946));
  OAI221xp5_ASAP7_75t_L     g17690(.A1(new_n5680), .A2(new_n8326), .B1(new_n7996), .B2(new_n9799), .C(new_n17946), .Y(new_n17947));
  AOI21xp33_ASAP7_75t_L     g17691(.A1(new_n7993), .A2(\b[41] ), .B(new_n17947), .Y(new_n17948));
  NAND2xp33_ASAP7_75t_L     g17692(.A(\a[50] ), .B(new_n17948), .Y(new_n17949));
  A2O1A1Ixp33_ASAP7_75t_L   g17693(.A1(\b[41] ), .A2(new_n7993), .B(new_n17947), .C(new_n7653), .Y(new_n17950));
  NAND2xp33_ASAP7_75t_L     g17694(.A(new_n17950), .B(new_n17949), .Y(new_n17951));
  NOR2xp33_ASAP7_75t_L      g17695(.A(new_n17951), .B(new_n17945), .Y(new_n17952));
  AOI22xp33_ASAP7_75t_L     g17696(.A1(new_n17949), .A2(new_n17950), .B1(new_n17942), .B2(new_n17944), .Y(new_n17953));
  NOR2xp33_ASAP7_75t_L      g17697(.A(new_n17953), .B(new_n17952), .Y(new_n17954));
  INVx1_ASAP7_75t_L         g17698(.A(new_n17804), .Y(new_n17955));
  INVx1_ASAP7_75t_L         g17699(.A(new_n17807), .Y(new_n17956));
  AOI211xp5_ASAP7_75t_L     g17700(.A1(new_n17655), .A2(new_n17608), .B(new_n17654), .C(new_n17808), .Y(new_n17957));
  AOI21xp33_ASAP7_75t_L     g17701(.A1(new_n17956), .A2(new_n17955), .B(new_n17957), .Y(new_n17958));
  NAND2xp33_ASAP7_75t_L     g17702(.A(new_n17958), .B(new_n17954), .Y(new_n17959));
  INVx1_ASAP7_75t_L         g17703(.A(new_n17954), .Y(new_n17960));
  A2O1A1Ixp33_ASAP7_75t_L   g17704(.A1(new_n17956), .A2(new_n17955), .B(new_n17957), .C(new_n17960), .Y(new_n17961));
  AOI22xp33_ASAP7_75t_L     g17705(.A1(new_n6822), .A2(\b[46] ), .B1(new_n6819), .B2(new_n7041), .Y(new_n17962));
  OAI221xp5_ASAP7_75t_L     g17706(.A1(new_n7392), .A2(new_n6756), .B1(new_n6220), .B2(new_n7115), .C(new_n17962), .Y(new_n17963));
  XNOR2x2_ASAP7_75t_L       g17707(.A(\a[47] ), .B(new_n17963), .Y(new_n17964));
  NAND3xp33_ASAP7_75t_L     g17708(.A(new_n17961), .B(new_n17959), .C(new_n17964), .Y(new_n17965));
  AO21x2_ASAP7_75t_L        g17709(.A1(new_n17959), .A2(new_n17961), .B(new_n17964), .Y(new_n17966));
  NAND4xp25_ASAP7_75t_L     g17710(.A(new_n17815), .B(new_n17965), .C(new_n17966), .D(new_n17891), .Y(new_n17967));
  NAND2xp33_ASAP7_75t_L     g17711(.A(new_n17965), .B(new_n17966), .Y(new_n17968));
  A2O1A1Ixp33_ASAP7_75t_L   g17712(.A1(new_n17810), .A2(new_n17754), .B(new_n17814), .C(new_n17968), .Y(new_n17969));
  NAND2xp33_ASAP7_75t_L     g17713(.A(new_n5999), .B(new_n7914), .Y(new_n17970));
  OAI221xp5_ASAP7_75t_L     g17714(.A1(new_n6312), .A2(new_n7907), .B1(new_n7333), .B2(new_n6544), .C(new_n17970), .Y(new_n17971));
  AOI21xp33_ASAP7_75t_L     g17715(.A1(new_n6308), .A2(\b[47] ), .B(new_n17971), .Y(new_n17972));
  NAND2xp33_ASAP7_75t_L     g17716(.A(\a[44] ), .B(new_n17972), .Y(new_n17973));
  A2O1A1Ixp33_ASAP7_75t_L   g17717(.A1(\b[47] ), .A2(new_n6308), .B(new_n17971), .C(new_n5996), .Y(new_n17974));
  AND2x2_ASAP7_75t_L        g17718(.A(new_n17974), .B(new_n17973), .Y(new_n17975));
  NAND3xp33_ASAP7_75t_L     g17719(.A(new_n17969), .B(new_n17967), .C(new_n17975), .Y(new_n17976));
  AO21x2_ASAP7_75t_L        g17720(.A1(new_n17967), .A2(new_n17969), .B(new_n17975), .Y(new_n17977));
  NAND2xp33_ASAP7_75t_L     g17721(.A(new_n17976), .B(new_n17977), .Y(new_n17978));
  OAI21xp33_ASAP7_75t_L     g17722(.A1(new_n17816), .A2(new_n17819), .B(new_n17822), .Y(new_n17979));
  XNOR2x2_ASAP7_75t_L       g17723(.A(new_n17978), .B(new_n17979), .Y(new_n17980));
  AOI22xp33_ASAP7_75t_L     g17724(.A1(new_n5249), .A2(\b[52] ), .B1(new_n5247), .B2(new_n8577), .Y(new_n17981));
  OAI221xp5_ASAP7_75t_L     g17725(.A1(new_n5241), .A2(new_n8249), .B1(new_n8228), .B2(new_n5521), .C(new_n17981), .Y(new_n17982));
  XNOR2x2_ASAP7_75t_L       g17726(.A(\a[41] ), .B(new_n17982), .Y(new_n17983));
  INVx1_ASAP7_75t_L         g17727(.A(new_n17983), .Y(new_n17984));
  NOR2xp33_ASAP7_75t_L      g17728(.A(new_n17984), .B(new_n17980), .Y(new_n17985));
  AND2x2_ASAP7_75t_L        g17729(.A(new_n17984), .B(new_n17980), .Y(new_n17986));
  NOR2xp33_ASAP7_75t_L      g17730(.A(new_n17985), .B(new_n17986), .Y(new_n17987));
  A2O1A1Ixp33_ASAP7_75t_L   g17731(.A1(new_n17829), .A2(new_n17751), .B(new_n17827), .C(new_n17987), .Y(new_n17988));
  INVx1_ASAP7_75t_L         g17732(.A(new_n17987), .Y(new_n17989));
  O2A1O1Ixp33_ASAP7_75t_L   g17733(.A1(new_n17678), .A2(new_n17685), .B(new_n17829), .C(new_n17827), .Y(new_n17990));
  NAND2xp33_ASAP7_75t_L     g17734(.A(new_n17990), .B(new_n17989), .Y(new_n17991));
  AND2x2_ASAP7_75t_L        g17735(.A(new_n17988), .B(new_n17991), .Y(new_n17992));
  NAND2xp33_ASAP7_75t_L     g17736(.A(new_n4542), .B(new_n9542), .Y(new_n17993));
  OAI221xp5_ASAP7_75t_L     g17737(.A1(new_n4550), .A2(new_n9534), .B1(new_n9199), .B2(new_n4536), .C(new_n17993), .Y(new_n17994));
  AOI21xp33_ASAP7_75t_L     g17738(.A1(new_n4780), .A2(\b[53] ), .B(new_n17994), .Y(new_n17995));
  NAND2xp33_ASAP7_75t_L     g17739(.A(\a[38] ), .B(new_n17995), .Y(new_n17996));
  A2O1A1Ixp33_ASAP7_75t_L   g17740(.A1(\b[53] ), .A2(new_n4780), .B(new_n17994), .C(new_n4539), .Y(new_n17997));
  AND2x2_ASAP7_75t_L        g17741(.A(new_n17997), .B(new_n17996), .Y(new_n17998));
  INVx1_ASAP7_75t_L         g17742(.A(new_n17998), .Y(new_n17999));
  XNOR2x2_ASAP7_75t_L       g17743(.A(new_n17999), .B(new_n17992), .Y(new_n18000));
  A2O1A1Ixp33_ASAP7_75t_L   g17744(.A1(new_n17833), .A2(new_n17748), .B(new_n17835), .C(new_n18000), .Y(new_n18001));
  AOI21xp33_ASAP7_75t_L     g17745(.A1(new_n17833), .A2(new_n17748), .B(new_n17835), .Y(new_n18002));
  INVx1_ASAP7_75t_L         g17746(.A(new_n18000), .Y(new_n18003));
  NAND2xp33_ASAP7_75t_L     g17747(.A(new_n18003), .B(new_n18002), .Y(new_n18004));
  AOI22xp33_ASAP7_75t_L     g17748(.A1(new_n3884), .A2(\b[58] ), .B1(new_n3881), .B2(new_n10857), .Y(new_n18005));
  OAI221xp5_ASAP7_75t_L     g17749(.A1(new_n4312), .A2(new_n10488), .B1(new_n10178), .B2(new_n4986), .C(new_n18005), .Y(new_n18006));
  XNOR2x2_ASAP7_75t_L       g17750(.A(\a[35] ), .B(new_n18006), .Y(new_n18007));
  NAND3xp33_ASAP7_75t_L     g17751(.A(new_n18004), .B(new_n18001), .C(new_n18007), .Y(new_n18008));
  AO21x2_ASAP7_75t_L        g17752(.A1(new_n18001), .A2(new_n18004), .B(new_n18007), .Y(new_n18009));
  NAND2xp33_ASAP7_75t_L     g17753(.A(new_n18008), .B(new_n18009), .Y(new_n18010));
  NAND3xp33_ASAP7_75t_L     g17754(.A(new_n17888), .B(new_n17890), .C(new_n18010), .Y(new_n18011));
  AO21x2_ASAP7_75t_L        g17755(.A1(new_n17890), .A2(new_n17888), .B(new_n18010), .Y(new_n18012));
  AND3x1_ASAP7_75t_L        g17756(.A(new_n17880), .B(new_n18012), .C(new_n18011), .Y(new_n18013));
  AOI21xp33_ASAP7_75t_L     g17757(.A1(new_n18012), .A2(new_n18011), .B(new_n17880), .Y(new_n18014));
  NOR2xp33_ASAP7_75t_L      g17758(.A(new_n18014), .B(new_n18013), .Y(new_n18015));
  XNOR2x2_ASAP7_75t_L       g17759(.A(new_n17869), .B(new_n18015), .Y(new_n18016));
  INVx1_ASAP7_75t_L         g17760(.A(new_n18016), .Y(new_n18017));
  O2A1O1Ixp33_ASAP7_75t_L   g17761(.A1(new_n17859), .A2(new_n17867), .B(new_n17860), .C(new_n18017), .Y(new_n18018));
  A2O1A1Ixp33_ASAP7_75t_L   g17762(.A1(new_n17727), .A2(new_n17723), .B(new_n17859), .C(new_n17860), .Y(new_n18019));
  NOR2xp33_ASAP7_75t_L      g17763(.A(new_n18016), .B(new_n18019), .Y(new_n18020));
  NOR2xp33_ASAP7_75t_L      g17764(.A(new_n18020), .B(new_n18018), .Y(\f[91] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17765(.A1(new_n17702), .A2(new_n17586), .B(new_n17585), .C(new_n17741), .Y(new_n18022));
  INVx1_ASAP7_75t_L         g17766(.A(new_n18015), .Y(new_n18023));
  A2O1A1O1Ixp25_ASAP7_75t_L g17767(.A1(new_n17742), .A2(new_n17737), .B(new_n17857), .C(new_n18022), .D(new_n18023), .Y(new_n18024));
  INVx1_ASAP7_75t_L         g17768(.A(new_n18024), .Y(new_n18025));
  A2O1A1Ixp33_ASAP7_75t_L   g17769(.A1(new_n17863), .A2(new_n17860), .B(new_n18017), .C(new_n18025), .Y(new_n18026));
  INVx1_ASAP7_75t_L         g17770(.A(new_n18004), .Y(new_n18027));
  AOI22xp33_ASAP7_75t_L     g17771(.A1(new_n3256), .A2(\b[62] ), .B1(new_n3254), .B2(new_n12280), .Y(new_n18028));
  OAI221xp5_ASAP7_75t_L     g17772(.A1(new_n3248), .A2(new_n11911), .B1(new_n11226), .B2(new_n3492), .C(new_n18028), .Y(new_n18029));
  XNOR2x2_ASAP7_75t_L       g17773(.A(\a[32] ), .B(new_n18029), .Y(new_n18030));
  A2O1A1Ixp33_ASAP7_75t_L   g17774(.A1(new_n18007), .A2(new_n18001), .B(new_n18027), .C(new_n18030), .Y(new_n18031));
  INVx1_ASAP7_75t_L         g17775(.A(new_n18030), .Y(new_n18032));
  NAND3xp33_ASAP7_75t_L     g17776(.A(new_n18008), .B(new_n18004), .C(new_n18032), .Y(new_n18033));
  NAND2xp33_ASAP7_75t_L     g17777(.A(new_n18031), .B(new_n18033), .Y(new_n18034));
  INVx1_ASAP7_75t_L         g17778(.A(new_n17992), .Y(new_n18035));
  O2A1O1Ixp33_ASAP7_75t_L   g17779(.A1(new_n17750), .A2(new_n17831), .B(new_n17828), .C(new_n17987), .Y(new_n18036));
  AOI22xp33_ASAP7_75t_L     g17780(.A1(new_n4544), .A2(\b[56] ), .B1(new_n4542), .B2(new_n10185), .Y(new_n18037));
  OAI221xp5_ASAP7_75t_L     g17781(.A1(new_n4536), .A2(new_n9534), .B1(new_n9199), .B2(new_n4781), .C(new_n18037), .Y(new_n18038));
  XNOR2x2_ASAP7_75t_L       g17782(.A(\a[38] ), .B(new_n18038), .Y(new_n18039));
  INVx1_ASAP7_75t_L         g17783(.A(new_n18039), .Y(new_n18040));
  AOI22xp33_ASAP7_75t_L     g17784(.A1(new_n5249), .A2(\b[53] ), .B1(new_n5247), .B2(new_n8889), .Y(new_n18041));
  OAI221xp5_ASAP7_75t_L     g17785(.A1(new_n5241), .A2(new_n8569), .B1(new_n8249), .B2(new_n5521), .C(new_n18041), .Y(new_n18042));
  XNOR2x2_ASAP7_75t_L       g17786(.A(\a[41] ), .B(new_n18042), .Y(new_n18043));
  INVx1_ASAP7_75t_L         g17787(.A(new_n18043), .Y(new_n18044));
  AOI22xp33_ASAP7_75t_L     g17788(.A1(new_n7659), .A2(\b[44] ), .B1(new_n7656), .B2(new_n7055), .Y(new_n18045));
  OAI221xp5_ASAP7_75t_L     g17789(.A1(new_n8326), .A2(new_n6195), .B1(new_n5680), .B2(new_n7994), .C(new_n18045), .Y(new_n18046));
  XNOR2x2_ASAP7_75t_L       g17790(.A(\a[50] ), .B(new_n18046), .Y(new_n18047));
  INVx1_ASAP7_75t_L         g17791(.A(new_n18047), .Y(new_n18048));
  A2O1A1Ixp33_ASAP7_75t_L   g17792(.A1(new_n17789), .A2(new_n17785), .B(new_n17793), .C(new_n17938), .Y(new_n18049));
  AOI22xp33_ASAP7_75t_L     g17793(.A1(new_n8645), .A2(\b[41] ), .B1(new_n8642), .B2(new_n5669), .Y(new_n18050));
  OAI221xp5_ASAP7_75t_L     g17794(.A1(new_n9322), .A2(new_n5186), .B1(new_n5166), .B2(new_n8965), .C(new_n18050), .Y(new_n18051));
  XNOR2x2_ASAP7_75t_L       g17795(.A(\a[53] ), .B(new_n18051), .Y(new_n18052));
  AOI22xp33_ASAP7_75t_L     g17796(.A1(new_n10594), .A2(\b[35] ), .B1(new_n10591), .B2(new_n5649), .Y(new_n18053));
  OAI221xp5_ASAP7_75t_L     g17797(.A1(new_n11335), .A2(new_n3827), .B1(new_n3807), .B2(new_n11330), .C(new_n18053), .Y(new_n18054));
  XNOR2x2_ASAP7_75t_L       g17798(.A(\a[59] ), .B(new_n18054), .Y(new_n18055));
  INVx1_ASAP7_75t_L         g17799(.A(new_n18055), .Y(new_n18056));
  AOI22xp33_ASAP7_75t_L     g17800(.A1(new_n11656), .A2(\b[32] ), .B1(new_n11654), .B2(new_n3450), .Y(new_n18057));
  OAI221xp5_ASAP7_75t_L     g17801(.A1(new_n12364), .A2(new_n3419), .B1(new_n3212), .B2(new_n13003), .C(new_n18057), .Y(new_n18058));
  XNOR2x2_ASAP7_75t_L       g17802(.A(\a[62] ), .B(new_n18058), .Y(new_n18059));
  INVx1_ASAP7_75t_L         g17803(.A(new_n18059), .Y(new_n18060));
  A2O1A1Ixp33_ASAP7_75t_L   g17804(.A1(new_n17910), .A2(new_n17911), .B(new_n17906), .C(new_n17905), .Y(new_n18061));
  NOR2xp33_ASAP7_75t_L      g17805(.A(new_n2852), .B(new_n12671), .Y(new_n18062));
  A2O1A1Ixp33_ASAP7_75t_L   g17806(.A1(\b[29] ), .A2(new_n12669), .B(new_n18062), .C(new_n17902), .Y(new_n18063));
  O2A1O1Ixp33_ASAP7_75t_L   g17807(.A1(new_n12353), .A2(new_n12355), .B(\b[29] ), .C(new_n18062), .Y(new_n18064));
  A2O1A1Ixp33_ASAP7_75t_L   g17808(.A1(new_n12669), .A2(\b[28] ), .B(new_n17899), .C(new_n18064), .Y(new_n18065));
  AND2x2_ASAP7_75t_L        g17809(.A(new_n18063), .B(new_n18065), .Y(new_n18066));
  XOR2x2_ASAP7_75t_L        g17810(.A(new_n18066), .B(new_n18061), .Y(new_n18067));
  NAND2xp33_ASAP7_75t_L     g17811(.A(new_n18060), .B(new_n18067), .Y(new_n18068));
  INVx1_ASAP7_75t_L         g17812(.A(new_n18067), .Y(new_n18069));
  NAND2xp33_ASAP7_75t_L     g17813(.A(new_n18059), .B(new_n18069), .Y(new_n18070));
  NAND3xp33_ASAP7_75t_L     g17814(.A(new_n18056), .B(new_n18068), .C(new_n18070), .Y(new_n18071));
  INVx1_ASAP7_75t_L         g17815(.A(new_n18071), .Y(new_n18072));
  AOI21xp33_ASAP7_75t_L     g17816(.A1(new_n18070), .A2(new_n18068), .B(new_n18056), .Y(new_n18073));
  NOR2xp33_ASAP7_75t_L      g17817(.A(new_n18073), .B(new_n18072), .Y(new_n18074));
  NAND3xp33_ASAP7_75t_L     g17818(.A(new_n18074), .B(new_n17924), .C(new_n17920), .Y(new_n18075));
  O2A1O1Ixp33_ASAP7_75t_L   g17819(.A1(new_n17916), .A2(new_n17917), .B(new_n17924), .C(new_n18074), .Y(new_n18076));
  INVx1_ASAP7_75t_L         g17820(.A(new_n18076), .Y(new_n18077));
  AOI22xp33_ASAP7_75t_L     g17821(.A1(new_n9623), .A2(\b[38] ), .B1(new_n9620), .B2(new_n4923), .Y(new_n18078));
  OAI221xp5_ASAP7_75t_L     g17822(.A1(new_n10280), .A2(new_n4701), .B1(new_n4465), .B2(new_n12010), .C(new_n18078), .Y(new_n18079));
  XNOR2x2_ASAP7_75t_L       g17823(.A(\a[56] ), .B(new_n18079), .Y(new_n18080));
  NAND3xp33_ASAP7_75t_L     g17824(.A(new_n18077), .B(new_n18075), .C(new_n18080), .Y(new_n18081));
  INVx1_ASAP7_75t_L         g17825(.A(new_n18081), .Y(new_n18082));
  AOI21xp33_ASAP7_75t_L     g17826(.A1(new_n18077), .A2(new_n18075), .B(new_n18080), .Y(new_n18083));
  NOR2xp33_ASAP7_75t_L      g17827(.A(new_n18083), .B(new_n18082), .Y(new_n18084));
  INVx1_ASAP7_75t_L         g17828(.A(new_n18084), .Y(new_n18085));
  OAI211xp5_ASAP7_75t_L     g17829(.A1(new_n17928), .A2(new_n17929), .B(new_n18085), .C(new_n17932), .Y(new_n18086));
  O2A1O1Ixp33_ASAP7_75t_L   g17830(.A1(new_n17928), .A2(new_n17929), .B(new_n17932), .C(new_n18085), .Y(new_n18087));
  INVx1_ASAP7_75t_L         g17831(.A(new_n18087), .Y(new_n18088));
  AND2x2_ASAP7_75t_L        g17832(.A(new_n18086), .B(new_n18088), .Y(new_n18089));
  NAND2xp33_ASAP7_75t_L     g17833(.A(new_n18052), .B(new_n18089), .Y(new_n18090));
  AO21x2_ASAP7_75t_L        g17834(.A1(new_n18086), .A2(new_n18088), .B(new_n18052), .Y(new_n18091));
  AND2x2_ASAP7_75t_L        g17835(.A(new_n18091), .B(new_n18090), .Y(new_n18092));
  O2A1O1Ixp33_ASAP7_75t_L   g17836(.A1(new_n17894), .A2(new_n17940), .B(new_n18049), .C(new_n18092), .Y(new_n18093));
  INVx1_ASAP7_75t_L         g17837(.A(new_n18093), .Y(new_n18094));
  A2O1A1Ixp33_ASAP7_75t_L   g17838(.A1(new_n17939), .A2(new_n17936), .B(new_n17894), .C(new_n18049), .Y(new_n18095));
  INVx1_ASAP7_75t_L         g17839(.A(new_n18095), .Y(new_n18096));
  NAND2xp33_ASAP7_75t_L     g17840(.A(new_n18096), .B(new_n18092), .Y(new_n18097));
  NAND3xp33_ASAP7_75t_L     g17841(.A(new_n18094), .B(new_n18048), .C(new_n18097), .Y(new_n18098));
  INVx1_ASAP7_75t_L         g17842(.A(new_n18098), .Y(new_n18099));
  AOI21xp33_ASAP7_75t_L     g17843(.A1(new_n18094), .A2(new_n18097), .B(new_n18048), .Y(new_n18100));
  NOR4xp25_ASAP7_75t_L      g17844(.A(new_n18099), .B(new_n17943), .C(new_n18100), .D(new_n17952), .Y(new_n18101));
  NOR2xp33_ASAP7_75t_L      g17845(.A(new_n18100), .B(new_n18099), .Y(new_n18102));
  O2A1O1Ixp33_ASAP7_75t_L   g17846(.A1(new_n17945), .A2(new_n17951), .B(new_n17944), .C(new_n18102), .Y(new_n18103));
  NOR2xp33_ASAP7_75t_L      g17847(.A(new_n18101), .B(new_n18103), .Y(new_n18104));
  AOI22xp33_ASAP7_75t_L     g17848(.A1(new_n6822), .A2(\b[47] ), .B1(new_n6819), .B2(new_n7323), .Y(new_n18105));
  OAI221xp5_ASAP7_75t_L     g17849(.A1(new_n7392), .A2(new_n7033), .B1(new_n6756), .B2(new_n7115), .C(new_n18105), .Y(new_n18106));
  XNOR2x2_ASAP7_75t_L       g17850(.A(\a[47] ), .B(new_n18106), .Y(new_n18107));
  AND2x2_ASAP7_75t_L        g17851(.A(new_n18107), .B(new_n18104), .Y(new_n18108));
  NOR2xp33_ASAP7_75t_L      g17852(.A(new_n18107), .B(new_n18104), .Y(new_n18109));
  NAND2xp33_ASAP7_75t_L     g17853(.A(new_n17959), .B(new_n17965), .Y(new_n18110));
  INVx1_ASAP7_75t_L         g17854(.A(new_n18110), .Y(new_n18111));
  NOR3xp33_ASAP7_75t_L      g17855(.A(new_n18111), .B(new_n18109), .C(new_n18108), .Y(new_n18112));
  NOR2xp33_ASAP7_75t_L      g17856(.A(new_n18109), .B(new_n18108), .Y(new_n18113));
  NOR2xp33_ASAP7_75t_L      g17857(.A(new_n18110), .B(new_n18113), .Y(new_n18114));
  NOR2xp33_ASAP7_75t_L      g17858(.A(new_n18112), .B(new_n18114), .Y(new_n18115));
  INVx1_ASAP7_75t_L         g17859(.A(new_n18115), .Y(new_n18116));
  AOI22xp33_ASAP7_75t_L     g17860(.A1(new_n6002), .A2(\b[50] ), .B1(new_n5999), .B2(new_n8235), .Y(new_n18117));
  OAI221xp5_ASAP7_75t_L     g17861(.A1(new_n6544), .A2(new_n7907), .B1(new_n7333), .B2(new_n6309), .C(new_n18117), .Y(new_n18118));
  XNOR2x2_ASAP7_75t_L       g17862(.A(\a[44] ), .B(new_n18118), .Y(new_n18119));
  NAND2xp33_ASAP7_75t_L     g17863(.A(new_n18119), .B(new_n18116), .Y(new_n18120));
  NOR2xp33_ASAP7_75t_L      g17864(.A(new_n18119), .B(new_n18116), .Y(new_n18121));
  INVx1_ASAP7_75t_L         g17865(.A(new_n18121), .Y(new_n18122));
  AND2x2_ASAP7_75t_L        g17866(.A(new_n18120), .B(new_n18122), .Y(new_n18123));
  INVx1_ASAP7_75t_L         g17867(.A(new_n18123), .Y(new_n18124));
  NAND2xp33_ASAP7_75t_L     g17868(.A(new_n17967), .B(new_n17976), .Y(new_n18125));
  NOR2xp33_ASAP7_75t_L      g17869(.A(new_n18125), .B(new_n18124), .Y(new_n18126));
  A2O1A1Ixp33_ASAP7_75t_L   g17870(.A1(new_n17662), .A2(new_n17658), .B(new_n17812), .C(new_n17891), .Y(new_n18127));
  O2A1O1Ixp33_ASAP7_75t_L   g17871(.A1(new_n17968), .A2(new_n18127), .B(new_n17976), .C(new_n18123), .Y(new_n18128));
  NOR2xp33_ASAP7_75t_L      g17872(.A(new_n18128), .B(new_n18126), .Y(new_n18129));
  NAND2xp33_ASAP7_75t_L     g17873(.A(new_n18044), .B(new_n18129), .Y(new_n18130));
  INVx1_ASAP7_75t_L         g17874(.A(new_n18130), .Y(new_n18131));
  NOR2xp33_ASAP7_75t_L      g17875(.A(new_n18044), .B(new_n18129), .Y(new_n18132));
  NOR2xp33_ASAP7_75t_L      g17876(.A(new_n18132), .B(new_n18131), .Y(new_n18133));
  NOR2xp33_ASAP7_75t_L      g17877(.A(new_n17978), .B(new_n17979), .Y(new_n18134));
  NOR2xp33_ASAP7_75t_L      g17878(.A(new_n18134), .B(new_n17985), .Y(new_n18135));
  XNOR2x2_ASAP7_75t_L       g17879(.A(new_n18135), .B(new_n18133), .Y(new_n18136));
  XNOR2x2_ASAP7_75t_L       g17880(.A(new_n18040), .B(new_n18136), .Y(new_n18137));
  A2O1A1Ixp33_ASAP7_75t_L   g17881(.A1(new_n17999), .A2(new_n18035), .B(new_n18036), .C(new_n18137), .Y(new_n18138));
  INVx1_ASAP7_75t_L         g17882(.A(new_n18036), .Y(new_n18139));
  A2O1A1Ixp33_ASAP7_75t_L   g17883(.A1(new_n17991), .A2(new_n17988), .B(new_n17998), .C(new_n18139), .Y(new_n18140));
  NOR2xp33_ASAP7_75t_L      g17884(.A(new_n18140), .B(new_n18137), .Y(new_n18141));
  INVx1_ASAP7_75t_L         g17885(.A(new_n18141), .Y(new_n18142));
  AOI22xp33_ASAP7_75t_L     g17886(.A1(new_n3884), .A2(\b[59] ), .B1(new_n3881), .B2(new_n10887), .Y(new_n18143));
  OAI221xp5_ASAP7_75t_L     g17887(.A1(new_n4312), .A2(new_n10848), .B1(new_n10488), .B2(new_n4986), .C(new_n18143), .Y(new_n18144));
  XNOR2x2_ASAP7_75t_L       g17888(.A(\a[35] ), .B(new_n18144), .Y(new_n18145));
  NAND3xp33_ASAP7_75t_L     g17889(.A(new_n18142), .B(new_n18138), .C(new_n18145), .Y(new_n18146));
  AO21x2_ASAP7_75t_L        g17890(.A1(new_n18138), .A2(new_n18142), .B(new_n18145), .Y(new_n18147));
  AND2x2_ASAP7_75t_L        g17891(.A(new_n18146), .B(new_n18147), .Y(new_n18148));
  NAND2xp33_ASAP7_75t_L     g17892(.A(new_n18034), .B(new_n18148), .Y(new_n18149));
  AO21x2_ASAP7_75t_L        g17893(.A1(new_n18147), .A2(new_n18146), .B(new_n18034), .Y(new_n18150));
  AND2x2_ASAP7_75t_L        g17894(.A(new_n18149), .B(new_n18150), .Y(new_n18151));
  A2O1A1Ixp33_ASAP7_75t_L   g17895(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n2700), .Y(new_n18152));
  A2O1A1Ixp33_ASAP7_75t_L   g17896(.A1(new_n18152), .A2(new_n2932), .B(new_n12599), .C(\a[29] ), .Y(new_n18153));
  O2A1O1Ixp33_ASAP7_75t_L   g17897(.A1(new_n2707), .A2(new_n13934), .B(new_n2932), .C(new_n12599), .Y(new_n18154));
  NAND2xp33_ASAP7_75t_L     g17898(.A(new_n2697), .B(new_n18154), .Y(new_n18155));
  AND2x2_ASAP7_75t_L        g17899(.A(new_n18155), .B(new_n18153), .Y(new_n18156));
  O2A1O1Ixp33_ASAP7_75t_L   g17900(.A1(new_n17883), .A2(new_n17887), .B(new_n18011), .C(new_n18156), .Y(new_n18157));
  INVx1_ASAP7_75t_L         g17901(.A(new_n18157), .Y(new_n18158));
  NAND3xp33_ASAP7_75t_L     g17902(.A(new_n18011), .B(new_n17890), .C(new_n18156), .Y(new_n18159));
  NAND3xp33_ASAP7_75t_L     g17903(.A(new_n18158), .B(new_n18151), .C(new_n18159), .Y(new_n18160));
  AO21x2_ASAP7_75t_L        g17904(.A1(new_n18159), .A2(new_n18158), .B(new_n18151), .Y(new_n18161));
  AND2x2_ASAP7_75t_L        g17905(.A(new_n18160), .B(new_n18161), .Y(new_n18162));
  OAI21xp33_ASAP7_75t_L     g17906(.A1(new_n17877), .A2(new_n18013), .B(new_n18162), .Y(new_n18163));
  INVx1_ASAP7_75t_L         g17907(.A(new_n18163), .Y(new_n18164));
  NOR3xp33_ASAP7_75t_L      g17908(.A(new_n18013), .B(new_n18162), .C(new_n17877), .Y(new_n18165));
  NOR2xp33_ASAP7_75t_L      g17909(.A(new_n18165), .B(new_n18164), .Y(new_n18166));
  XOR2x2_ASAP7_75t_L        g17910(.A(new_n18166), .B(new_n18026), .Y(\f[92] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17911(.A1(new_n18016), .A2(new_n18019), .B(new_n18024), .C(new_n18166), .D(new_n18164), .Y(new_n18168));
  AOI22xp33_ASAP7_75t_L     g17912(.A1(new_n5249), .A2(\b[54] ), .B1(new_n5247), .B2(new_n9208), .Y(new_n18169));
  OAI221xp5_ASAP7_75t_L     g17913(.A1(new_n5241), .A2(new_n8882), .B1(new_n8569), .B2(new_n5521), .C(new_n18169), .Y(new_n18170));
  XNOR2x2_ASAP7_75t_L       g17914(.A(\a[41] ), .B(new_n18170), .Y(new_n18171));
  INVx1_ASAP7_75t_L         g17915(.A(new_n18171), .Y(new_n18172));
  O2A1O1Ixp33_ASAP7_75t_L   g17916(.A1(new_n18108), .A2(new_n18109), .B(new_n18111), .C(new_n18121), .Y(new_n18173));
  AOI22xp33_ASAP7_75t_L     g17917(.A1(new_n7659), .A2(\b[45] ), .B1(new_n7656), .B2(new_n6764), .Y(new_n18174));
  OAI221xp5_ASAP7_75t_L     g17918(.A1(new_n8326), .A2(new_n6220), .B1(new_n6195), .B2(new_n7994), .C(new_n18174), .Y(new_n18175));
  XNOR2x2_ASAP7_75t_L       g17919(.A(new_n7653), .B(new_n18175), .Y(new_n18176));
  INVx1_ASAP7_75t_L         g17920(.A(new_n18090), .Y(new_n18177));
  AOI22xp33_ASAP7_75t_L     g17921(.A1(new_n10594), .A2(\b[36] ), .B1(new_n10591), .B2(new_n4473), .Y(new_n18178));
  OAI221xp5_ASAP7_75t_L     g17922(.A1(new_n11335), .A2(new_n4053), .B1(new_n3827), .B2(new_n11330), .C(new_n18178), .Y(new_n18179));
  XNOR2x2_ASAP7_75t_L       g17923(.A(\a[59] ), .B(new_n18179), .Y(new_n18180));
  INVx1_ASAP7_75t_L         g17924(.A(new_n18180), .Y(new_n18181));
  AOI22xp33_ASAP7_75t_L     g17925(.A1(new_n11656), .A2(\b[33] ), .B1(new_n11654), .B2(new_n3813), .Y(new_n18182));
  OAI221xp5_ASAP7_75t_L     g17926(.A1(new_n12364), .A2(new_n3443), .B1(new_n3419), .B2(new_n13003), .C(new_n18182), .Y(new_n18183));
  XNOR2x2_ASAP7_75t_L       g17927(.A(\a[62] ), .B(new_n18183), .Y(new_n18184));
  NOR2xp33_ASAP7_75t_L      g17928(.A(new_n2871), .B(new_n12671), .Y(new_n18185));
  A2O1A1Ixp33_ASAP7_75t_L   g17929(.A1(new_n12669), .A2(\b[30] ), .B(new_n18185), .C(new_n2697), .Y(new_n18186));
  INVx1_ASAP7_75t_L         g17930(.A(new_n18186), .Y(new_n18187));
  O2A1O1Ixp33_ASAP7_75t_L   g17931(.A1(new_n12353), .A2(new_n12355), .B(\b[30] ), .C(new_n18185), .Y(new_n18188));
  NAND2xp33_ASAP7_75t_L     g17932(.A(\a[29] ), .B(new_n18188), .Y(new_n18189));
  INVx1_ASAP7_75t_L         g17933(.A(new_n18189), .Y(new_n18190));
  NOR2xp33_ASAP7_75t_L      g17934(.A(new_n18187), .B(new_n18190), .Y(new_n18191));
  XNOR2x2_ASAP7_75t_L       g17935(.A(new_n18064), .B(new_n18191), .Y(new_n18192));
  A2O1A1O1Ixp25_ASAP7_75t_L g17936(.A1(new_n12669), .A2(\b[28] ), .B(new_n17899), .C(new_n18064), .D(new_n18061), .Y(new_n18193));
  A2O1A1O1Ixp25_ASAP7_75t_L g17937(.A1(new_n12669), .A2(\b[29] ), .B(new_n18062), .C(new_n17902), .D(new_n18193), .Y(new_n18194));
  NAND2xp33_ASAP7_75t_L     g17938(.A(new_n18192), .B(new_n18194), .Y(new_n18195));
  INVx1_ASAP7_75t_L         g17939(.A(new_n18195), .Y(new_n18196));
  INVx1_ASAP7_75t_L         g17940(.A(new_n18065), .Y(new_n18197));
  O2A1O1Ixp33_ASAP7_75t_L   g17941(.A1(new_n18197), .A2(new_n18061), .B(new_n18063), .C(new_n18192), .Y(new_n18198));
  NOR2xp33_ASAP7_75t_L      g17942(.A(new_n18198), .B(new_n18196), .Y(new_n18199));
  INVx1_ASAP7_75t_L         g17943(.A(new_n18199), .Y(new_n18200));
  NOR2xp33_ASAP7_75t_L      g17944(.A(new_n18184), .B(new_n18200), .Y(new_n18201));
  INVx1_ASAP7_75t_L         g17945(.A(new_n18201), .Y(new_n18202));
  NAND2xp33_ASAP7_75t_L     g17946(.A(new_n18184), .B(new_n18200), .Y(new_n18203));
  NAND3xp33_ASAP7_75t_L     g17947(.A(new_n18202), .B(new_n18181), .C(new_n18203), .Y(new_n18204));
  INVx1_ASAP7_75t_L         g17948(.A(new_n18204), .Y(new_n18205));
  AOI21xp33_ASAP7_75t_L     g17949(.A1(new_n18202), .A2(new_n18203), .B(new_n18181), .Y(new_n18206));
  NOR2xp33_ASAP7_75t_L      g17950(.A(new_n18206), .B(new_n18205), .Y(new_n18207));
  INVx1_ASAP7_75t_L         g17951(.A(new_n18207), .Y(new_n18208));
  O2A1O1Ixp33_ASAP7_75t_L   g17952(.A1(new_n18059), .A2(new_n18069), .B(new_n18071), .C(new_n18208), .Y(new_n18209));
  NAND2xp33_ASAP7_75t_L     g17953(.A(new_n18068), .B(new_n18071), .Y(new_n18210));
  NOR2xp33_ASAP7_75t_L      g17954(.A(new_n18210), .B(new_n18207), .Y(new_n18211));
  NOR2xp33_ASAP7_75t_L      g17955(.A(new_n18211), .B(new_n18209), .Y(new_n18212));
  AOI22xp33_ASAP7_75t_L     g17956(.A1(new_n9623), .A2(\b[39] ), .B1(new_n9620), .B2(new_n5174), .Y(new_n18213));
  OAI221xp5_ASAP7_75t_L     g17957(.A1(new_n10280), .A2(new_n4915), .B1(new_n4701), .B2(new_n12010), .C(new_n18213), .Y(new_n18214));
  XNOR2x2_ASAP7_75t_L       g17958(.A(\a[56] ), .B(new_n18214), .Y(new_n18215));
  INVx1_ASAP7_75t_L         g17959(.A(new_n18215), .Y(new_n18216));
  XNOR2x2_ASAP7_75t_L       g17960(.A(new_n18216), .B(new_n18212), .Y(new_n18217));
  A2O1A1Ixp33_ASAP7_75t_L   g17961(.A1(new_n18080), .A2(new_n18075), .B(new_n18076), .C(new_n18217), .Y(new_n18218));
  A2O1A1Ixp33_ASAP7_75t_L   g17962(.A1(new_n17924), .A2(new_n17920), .B(new_n18074), .C(new_n18081), .Y(new_n18219));
  NOR2xp33_ASAP7_75t_L      g17963(.A(new_n18219), .B(new_n18217), .Y(new_n18220));
  INVx1_ASAP7_75t_L         g17964(.A(new_n18220), .Y(new_n18221));
  NAND2xp33_ASAP7_75t_L     g17965(.A(new_n18218), .B(new_n18221), .Y(new_n18222));
  AOI22xp33_ASAP7_75t_L     g17966(.A1(new_n8645), .A2(\b[42] ), .B1(new_n8642), .B2(new_n5688), .Y(new_n18223));
  OAI221xp5_ASAP7_75t_L     g17967(.A1(new_n9322), .A2(new_n5666), .B1(new_n5186), .B2(new_n8965), .C(new_n18223), .Y(new_n18224));
  XNOR2x2_ASAP7_75t_L       g17968(.A(\a[53] ), .B(new_n18224), .Y(new_n18225));
  XNOR2x2_ASAP7_75t_L       g17969(.A(new_n18225), .B(new_n18222), .Y(new_n18226));
  NOR3xp33_ASAP7_75t_L      g17970(.A(new_n18226), .B(new_n18177), .C(new_n18087), .Y(new_n18227));
  OA21x2_ASAP7_75t_L        g17971(.A1(new_n18087), .A2(new_n18177), .B(new_n18226), .Y(new_n18228));
  NOR2xp33_ASAP7_75t_L      g17972(.A(new_n18227), .B(new_n18228), .Y(new_n18229));
  XOR2x2_ASAP7_75t_L        g17973(.A(new_n18176), .B(new_n18229), .Y(new_n18230));
  INVx1_ASAP7_75t_L         g17974(.A(new_n18230), .Y(new_n18231));
  NAND3xp33_ASAP7_75t_L     g17975(.A(new_n18231), .B(new_n18098), .C(new_n18094), .Y(new_n18232));
  O2A1O1Ixp33_ASAP7_75t_L   g17976(.A1(new_n18096), .A2(new_n18092), .B(new_n18098), .C(new_n18231), .Y(new_n18233));
  INVx1_ASAP7_75t_L         g17977(.A(new_n18233), .Y(new_n18234));
  NAND2xp33_ASAP7_75t_L     g17978(.A(new_n18232), .B(new_n18234), .Y(new_n18235));
  AOI22xp33_ASAP7_75t_L     g17979(.A1(new_n6822), .A2(\b[48] ), .B1(new_n6819), .B2(new_n7341), .Y(new_n18236));
  OAI221xp5_ASAP7_75t_L     g17980(.A1(new_n7392), .A2(new_n7316), .B1(new_n7033), .B2(new_n7115), .C(new_n18236), .Y(new_n18237));
  XNOR2x2_ASAP7_75t_L       g17981(.A(\a[47] ), .B(new_n18237), .Y(new_n18238));
  XNOR2x2_ASAP7_75t_L       g17982(.A(new_n18238), .B(new_n18235), .Y(new_n18239));
  A2O1A1Ixp33_ASAP7_75t_L   g17983(.A1(new_n18104), .A2(new_n18107), .B(new_n18103), .C(new_n18239), .Y(new_n18240));
  OR3x1_ASAP7_75t_L         g17984(.A(new_n18239), .B(new_n18103), .C(new_n18108), .Y(new_n18241));
  NAND2xp33_ASAP7_75t_L     g17985(.A(new_n18240), .B(new_n18241), .Y(new_n18242));
  AOI22xp33_ASAP7_75t_L     g17986(.A1(new_n6002), .A2(\b[51] ), .B1(new_n5999), .B2(new_n8257), .Y(new_n18243));
  OAI221xp5_ASAP7_75t_L     g17987(.A1(new_n6544), .A2(new_n8228), .B1(new_n7907), .B2(new_n6309), .C(new_n18243), .Y(new_n18244));
  XNOR2x2_ASAP7_75t_L       g17988(.A(\a[44] ), .B(new_n18244), .Y(new_n18245));
  NOR2xp33_ASAP7_75t_L      g17989(.A(new_n18245), .B(new_n18242), .Y(new_n18246));
  INVx1_ASAP7_75t_L         g17990(.A(new_n18246), .Y(new_n18247));
  NAND2xp33_ASAP7_75t_L     g17991(.A(new_n18245), .B(new_n18242), .Y(new_n18248));
  AND2x2_ASAP7_75t_L        g17992(.A(new_n18248), .B(new_n18247), .Y(new_n18249));
  INVx1_ASAP7_75t_L         g17993(.A(new_n18249), .Y(new_n18250));
  NAND2xp33_ASAP7_75t_L     g17994(.A(new_n18173), .B(new_n18250), .Y(new_n18251));
  O2A1O1Ixp33_ASAP7_75t_L   g17995(.A1(new_n18113), .A2(new_n18110), .B(new_n18122), .C(new_n18250), .Y(new_n18252));
  INVx1_ASAP7_75t_L         g17996(.A(new_n18252), .Y(new_n18253));
  AO21x2_ASAP7_75t_L        g17997(.A1(new_n18251), .A2(new_n18253), .B(new_n18172), .Y(new_n18254));
  AND2x2_ASAP7_75t_L        g17998(.A(new_n18251), .B(new_n18253), .Y(new_n18255));
  NAND2xp33_ASAP7_75t_L     g17999(.A(new_n18172), .B(new_n18255), .Y(new_n18256));
  AND2x2_ASAP7_75t_L        g18000(.A(new_n18254), .B(new_n18256), .Y(new_n18257));
  A2O1A1Ixp33_ASAP7_75t_L   g18001(.A1(new_n18129), .A2(new_n18044), .B(new_n18126), .C(new_n18257), .Y(new_n18258));
  OR3x1_ASAP7_75t_L         g18002(.A(new_n18257), .B(new_n18126), .C(new_n18131), .Y(new_n18259));
  NAND2xp33_ASAP7_75t_L     g18003(.A(new_n18258), .B(new_n18259), .Y(new_n18260));
  AOI22xp33_ASAP7_75t_L     g18004(.A1(new_n4544), .A2(\b[57] ), .B1(new_n4542), .B2(new_n10495), .Y(new_n18261));
  OAI221xp5_ASAP7_75t_L     g18005(.A1(new_n4536), .A2(new_n10178), .B1(new_n9534), .B2(new_n4781), .C(new_n18261), .Y(new_n18262));
  XNOR2x2_ASAP7_75t_L       g18006(.A(\a[38] ), .B(new_n18262), .Y(new_n18263));
  XOR2x2_ASAP7_75t_L        g18007(.A(new_n18263), .B(new_n18260), .Y(new_n18264));
  MAJx2_ASAP7_75t_L         g18008(.A(new_n18133), .B(new_n18040), .C(new_n18135), .Y(new_n18265));
  XOR2x2_ASAP7_75t_L        g18009(.A(new_n18265), .B(new_n18264), .Y(new_n18266));
  AOI22xp33_ASAP7_75t_L     g18010(.A1(new_n3884), .A2(\b[60] ), .B1(new_n3881), .B2(new_n11234), .Y(new_n18267));
  OAI221xp5_ASAP7_75t_L     g18011(.A1(new_n4312), .A2(new_n10881), .B1(new_n10848), .B2(new_n4986), .C(new_n18267), .Y(new_n18268));
  XNOR2x2_ASAP7_75t_L       g18012(.A(\a[35] ), .B(new_n18268), .Y(new_n18269));
  INVx1_ASAP7_75t_L         g18013(.A(new_n18269), .Y(new_n18270));
  XNOR2x2_ASAP7_75t_L       g18014(.A(new_n18270), .B(new_n18266), .Y(new_n18271));
  A2O1A1Ixp33_ASAP7_75t_L   g18015(.A1(new_n18145), .A2(new_n18138), .B(new_n18141), .C(new_n18271), .Y(new_n18272));
  NAND2xp33_ASAP7_75t_L     g18016(.A(new_n18142), .B(new_n18146), .Y(new_n18273));
  OR2x4_ASAP7_75t_L         g18017(.A(new_n18273), .B(new_n18271), .Y(new_n18274));
  AND2x2_ASAP7_75t_L        g18018(.A(new_n18272), .B(new_n18274), .Y(new_n18275));
  NAND2xp33_ASAP7_75t_L     g18019(.A(\b[63] ), .B(new_n3256), .Y(new_n18276));
  A2O1A1Ixp33_ASAP7_75t_L   g18020(.A1(new_n12607), .A2(new_n12603), .B(new_n3261), .C(new_n18276), .Y(new_n18277));
  AOI221xp5_ASAP7_75t_L     g18021(.A1(\b[61] ), .A2(new_n3491), .B1(\b[62] ), .B2(new_n3260), .C(new_n18277), .Y(new_n18278));
  XNOR2x2_ASAP7_75t_L       g18022(.A(new_n3251), .B(new_n18278), .Y(new_n18279));
  INVx1_ASAP7_75t_L         g18023(.A(new_n18279), .Y(new_n18280));
  A2O1A1O1Ixp25_ASAP7_75t_L g18024(.A1(new_n18147), .A2(new_n18146), .B(new_n18034), .C(new_n18033), .D(new_n18280), .Y(new_n18281));
  A2O1A1Ixp33_ASAP7_75t_L   g18025(.A1(new_n18146), .A2(new_n18147), .B(new_n18034), .C(new_n18033), .Y(new_n18282));
  NOR2xp33_ASAP7_75t_L      g18026(.A(new_n18279), .B(new_n18282), .Y(new_n18283));
  OR3x1_ASAP7_75t_L         g18027(.A(new_n18275), .B(new_n18281), .C(new_n18283), .Y(new_n18284));
  OAI21xp33_ASAP7_75t_L     g18028(.A1(new_n18281), .A2(new_n18283), .B(new_n18275), .Y(new_n18285));
  AND2x2_ASAP7_75t_L        g18029(.A(new_n18285), .B(new_n18284), .Y(new_n18286));
  A2O1A1Ixp33_ASAP7_75t_L   g18030(.A1(new_n18159), .A2(new_n18151), .B(new_n18157), .C(new_n18286), .Y(new_n18287));
  A2O1A1Ixp33_ASAP7_75t_L   g18031(.A1(new_n18011), .A2(new_n17890), .B(new_n18156), .C(new_n18160), .Y(new_n18288));
  AO21x2_ASAP7_75t_L        g18032(.A1(new_n18285), .A2(new_n18284), .B(new_n18288), .Y(new_n18289));
  NAND2xp33_ASAP7_75t_L     g18033(.A(new_n18289), .B(new_n18287), .Y(new_n18290));
  XOR2x2_ASAP7_75t_L        g18034(.A(new_n18290), .B(new_n18168), .Y(\f[93] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18035(.A1(new_n18019), .A2(new_n18016), .B(new_n18024), .C(new_n18166), .Y(new_n18292));
  NAND2xp33_ASAP7_75t_L     g18036(.A(new_n18270), .B(new_n18266), .Y(new_n18293));
  A2O1A1Ixp33_ASAP7_75t_L   g18037(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n3254), .Y(new_n18294));
  AOI22xp33_ASAP7_75t_L     g18038(.A1(new_n3260), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3491), .Y(new_n18295));
  NAND3xp33_ASAP7_75t_L     g18039(.A(new_n18294), .B(\a[32] ), .C(new_n18295), .Y(new_n18296));
  INVx1_ASAP7_75t_L         g18040(.A(new_n18296), .Y(new_n18297));
  A2O1A1O1Ixp25_ASAP7_75t_L g18041(.A1(new_n13507), .A2(new_n13506), .B(new_n3261), .C(new_n18295), .D(\a[32] ), .Y(new_n18298));
  NOR2xp33_ASAP7_75t_L      g18042(.A(new_n18298), .B(new_n18297), .Y(new_n18299));
  O2A1O1Ixp33_ASAP7_75t_L   g18043(.A1(new_n18273), .A2(new_n18271), .B(new_n18293), .C(new_n18299), .Y(new_n18300));
  INVx1_ASAP7_75t_L         g18044(.A(new_n18300), .Y(new_n18301));
  NAND3xp33_ASAP7_75t_L     g18045(.A(new_n18274), .B(new_n18293), .C(new_n18299), .Y(new_n18302));
  NAND2xp33_ASAP7_75t_L     g18046(.A(new_n18301), .B(new_n18302), .Y(new_n18303));
  INVx1_ASAP7_75t_L         g18047(.A(new_n18258), .Y(new_n18304));
  INVx1_ASAP7_75t_L         g18048(.A(new_n18173), .Y(new_n18305));
  NAND2xp33_ASAP7_75t_L     g18049(.A(new_n18176), .B(new_n18229), .Y(new_n18306));
  AOI22xp33_ASAP7_75t_L     g18050(.A1(new_n9623), .A2(\b[40] ), .B1(new_n9620), .B2(new_n5194), .Y(new_n18307));
  OAI221xp5_ASAP7_75t_L     g18051(.A1(new_n10280), .A2(new_n5166), .B1(new_n4915), .B2(new_n12010), .C(new_n18307), .Y(new_n18308));
  XNOR2x2_ASAP7_75t_L       g18052(.A(\a[56] ), .B(new_n18308), .Y(new_n18309));
  INVx1_ASAP7_75t_L         g18053(.A(new_n18309), .Y(new_n18310));
  AOI22xp33_ASAP7_75t_L     g18054(.A1(new_n10594), .A2(\b[37] ), .B1(new_n10591), .B2(new_n4709), .Y(new_n18311));
  OAI221xp5_ASAP7_75t_L     g18055(.A1(new_n11335), .A2(new_n4465), .B1(new_n4053), .B2(new_n11330), .C(new_n18311), .Y(new_n18312));
  XNOR2x2_ASAP7_75t_L       g18056(.A(\a[59] ), .B(new_n18312), .Y(new_n18313));
  INVx1_ASAP7_75t_L         g18057(.A(new_n18313), .Y(new_n18314));
  NOR2xp33_ASAP7_75t_L      g18058(.A(new_n3212), .B(new_n12671), .Y(new_n18315));
  A2O1A1O1Ixp25_ASAP7_75t_L g18059(.A1(new_n12669), .A2(\b[29] ), .B(new_n18062), .C(new_n18189), .D(new_n18187), .Y(new_n18316));
  A2O1A1Ixp33_ASAP7_75t_L   g18060(.A1(new_n12669), .A2(\b[31] ), .B(new_n18315), .C(new_n18316), .Y(new_n18317));
  O2A1O1Ixp33_ASAP7_75t_L   g18061(.A1(new_n12353), .A2(new_n12355), .B(\b[31] ), .C(new_n18315), .Y(new_n18318));
  INVx1_ASAP7_75t_L         g18062(.A(new_n18318), .Y(new_n18319));
  O2A1O1Ixp33_ASAP7_75t_L   g18063(.A1(new_n18064), .A2(new_n18190), .B(new_n18186), .C(new_n18319), .Y(new_n18320));
  INVx1_ASAP7_75t_L         g18064(.A(new_n18320), .Y(new_n18321));
  NAND2xp33_ASAP7_75t_L     g18065(.A(new_n18317), .B(new_n18321), .Y(new_n18322));
  NAND2xp33_ASAP7_75t_L     g18066(.A(new_n11654), .B(new_n3833), .Y(new_n18323));
  OAI221xp5_ASAP7_75t_L     g18067(.A1(new_n12023), .A2(new_n3827), .B1(new_n3807), .B2(new_n12364), .C(new_n18323), .Y(new_n18324));
  AOI21xp33_ASAP7_75t_L     g18068(.A1(new_n12021), .A2(\b[32] ), .B(new_n18324), .Y(new_n18325));
  NAND2xp33_ASAP7_75t_L     g18069(.A(\a[62] ), .B(new_n18325), .Y(new_n18326));
  A2O1A1Ixp33_ASAP7_75t_L   g18070(.A1(\b[32] ), .A2(new_n12021), .B(new_n18324), .C(new_n11651), .Y(new_n18327));
  AND3x1_ASAP7_75t_L        g18071(.A(new_n18326), .B(new_n18327), .C(new_n18322), .Y(new_n18328));
  AND2x2_ASAP7_75t_L        g18072(.A(new_n18327), .B(new_n18326), .Y(new_n18329));
  NOR2xp33_ASAP7_75t_L      g18073(.A(new_n18322), .B(new_n18329), .Y(new_n18330));
  NOR2xp33_ASAP7_75t_L      g18074(.A(new_n18328), .B(new_n18330), .Y(new_n18331));
  INVx1_ASAP7_75t_L         g18075(.A(new_n18331), .Y(new_n18332));
  O2A1O1Ixp33_ASAP7_75t_L   g18076(.A1(new_n18184), .A2(new_n18198), .B(new_n18195), .C(new_n18332), .Y(new_n18333));
  INVx1_ASAP7_75t_L         g18077(.A(new_n18333), .Y(new_n18334));
  NOR2xp33_ASAP7_75t_L      g18078(.A(new_n18196), .B(new_n18201), .Y(new_n18335));
  NAND2xp33_ASAP7_75t_L     g18079(.A(new_n18332), .B(new_n18335), .Y(new_n18336));
  NAND3xp33_ASAP7_75t_L     g18080(.A(new_n18336), .B(new_n18334), .C(new_n18314), .Y(new_n18337));
  INVx1_ASAP7_75t_L         g18081(.A(new_n18337), .Y(new_n18338));
  AOI21xp33_ASAP7_75t_L     g18082(.A1(new_n18336), .A2(new_n18334), .B(new_n18314), .Y(new_n18339));
  NOR2xp33_ASAP7_75t_L      g18083(.A(new_n18339), .B(new_n18338), .Y(new_n18340));
  INVx1_ASAP7_75t_L         g18084(.A(new_n18340), .Y(new_n18341));
  A2O1A1O1Ixp25_ASAP7_75t_L g18085(.A1(new_n18071), .A2(new_n18068), .B(new_n18206), .C(new_n18204), .D(new_n18341), .Y(new_n18342));
  INVx1_ASAP7_75t_L         g18086(.A(new_n18342), .Y(new_n18343));
  INVx1_ASAP7_75t_L         g18087(.A(new_n18209), .Y(new_n18344));
  NAND3xp33_ASAP7_75t_L     g18088(.A(new_n18344), .B(new_n18204), .C(new_n18341), .Y(new_n18345));
  NAND3xp33_ASAP7_75t_L     g18089(.A(new_n18343), .B(new_n18310), .C(new_n18345), .Y(new_n18346));
  INVx1_ASAP7_75t_L         g18090(.A(new_n18346), .Y(new_n18347));
  AOI21xp33_ASAP7_75t_L     g18091(.A1(new_n18343), .A2(new_n18345), .B(new_n18310), .Y(new_n18348));
  NOR2xp33_ASAP7_75t_L      g18092(.A(new_n18348), .B(new_n18347), .Y(new_n18349));
  A2O1A1Ixp33_ASAP7_75t_L   g18093(.A1(new_n18216), .A2(new_n18212), .B(new_n18220), .C(new_n18349), .Y(new_n18350));
  AOI211xp5_ASAP7_75t_L     g18094(.A1(new_n18212), .A2(new_n18216), .B(new_n18220), .C(new_n18349), .Y(new_n18351));
  INVx1_ASAP7_75t_L         g18095(.A(new_n18351), .Y(new_n18352));
  NAND2xp33_ASAP7_75t_L     g18096(.A(new_n18350), .B(new_n18352), .Y(new_n18353));
  NAND2xp33_ASAP7_75t_L     g18097(.A(\b[43] ), .B(new_n8645), .Y(new_n18354));
  OAI221xp5_ASAP7_75t_L     g18098(.A1(new_n5680), .A2(new_n9322), .B1(new_n8967), .B2(new_n9799), .C(new_n18354), .Y(new_n18355));
  AOI21xp33_ASAP7_75t_L     g18099(.A1(new_n8964), .A2(\b[41] ), .B(new_n18355), .Y(new_n18356));
  NAND2xp33_ASAP7_75t_L     g18100(.A(\a[53] ), .B(new_n18356), .Y(new_n18357));
  A2O1A1Ixp33_ASAP7_75t_L   g18101(.A1(\b[41] ), .A2(new_n8964), .B(new_n18355), .C(new_n8639), .Y(new_n18358));
  NAND2xp33_ASAP7_75t_L     g18102(.A(new_n18358), .B(new_n18357), .Y(new_n18359));
  NOR2xp33_ASAP7_75t_L      g18103(.A(new_n18359), .B(new_n18353), .Y(new_n18360));
  INVx1_ASAP7_75t_L         g18104(.A(new_n18360), .Y(new_n18361));
  NAND2xp33_ASAP7_75t_L     g18105(.A(new_n18359), .B(new_n18353), .Y(new_n18362));
  AND2x2_ASAP7_75t_L        g18106(.A(new_n18362), .B(new_n18361), .Y(new_n18363));
  INVx1_ASAP7_75t_L         g18107(.A(new_n18222), .Y(new_n18364));
  INVx1_ASAP7_75t_L         g18108(.A(new_n18225), .Y(new_n18365));
  AOI21xp33_ASAP7_75t_L     g18109(.A1(new_n18365), .A2(new_n18364), .B(new_n18227), .Y(new_n18366));
  NAND2xp33_ASAP7_75t_L     g18110(.A(new_n18366), .B(new_n18363), .Y(new_n18367));
  INVx1_ASAP7_75t_L         g18111(.A(new_n18363), .Y(new_n18368));
  A2O1A1Ixp33_ASAP7_75t_L   g18112(.A1(new_n18365), .A2(new_n18364), .B(new_n18227), .C(new_n18368), .Y(new_n18369));
  AOI22xp33_ASAP7_75t_L     g18113(.A1(new_n7659), .A2(\b[46] ), .B1(new_n7656), .B2(new_n7041), .Y(new_n18370));
  OAI221xp5_ASAP7_75t_L     g18114(.A1(new_n8326), .A2(new_n6756), .B1(new_n6220), .B2(new_n7994), .C(new_n18370), .Y(new_n18371));
  XNOR2x2_ASAP7_75t_L       g18115(.A(\a[50] ), .B(new_n18371), .Y(new_n18372));
  NAND3xp33_ASAP7_75t_L     g18116(.A(new_n18369), .B(new_n18367), .C(new_n18372), .Y(new_n18373));
  AO21x2_ASAP7_75t_L        g18117(.A1(new_n18367), .A2(new_n18369), .B(new_n18372), .Y(new_n18374));
  NAND4xp25_ASAP7_75t_L     g18118(.A(new_n18234), .B(new_n18373), .C(new_n18374), .D(new_n18306), .Y(new_n18375));
  NAND2xp33_ASAP7_75t_L     g18119(.A(new_n18373), .B(new_n18374), .Y(new_n18376));
  A2O1A1Ixp33_ASAP7_75t_L   g18120(.A1(new_n18229), .A2(new_n18176), .B(new_n18233), .C(new_n18376), .Y(new_n18377));
  NAND2xp33_ASAP7_75t_L     g18121(.A(new_n6819), .B(new_n7914), .Y(new_n18378));
  OAI221xp5_ASAP7_75t_L     g18122(.A1(new_n7118), .A2(new_n7907), .B1(new_n7333), .B2(new_n7392), .C(new_n18378), .Y(new_n18379));
  AOI21xp33_ASAP7_75t_L     g18123(.A1(new_n7124), .A2(\b[47] ), .B(new_n18379), .Y(new_n18380));
  NAND2xp33_ASAP7_75t_L     g18124(.A(\a[47] ), .B(new_n18380), .Y(new_n18381));
  A2O1A1Ixp33_ASAP7_75t_L   g18125(.A1(\b[47] ), .A2(new_n7124), .B(new_n18379), .C(new_n6816), .Y(new_n18382));
  AND2x2_ASAP7_75t_L        g18126(.A(new_n18382), .B(new_n18381), .Y(new_n18383));
  NAND3xp33_ASAP7_75t_L     g18127(.A(new_n18377), .B(new_n18375), .C(new_n18383), .Y(new_n18384));
  AO21x2_ASAP7_75t_L        g18128(.A1(new_n18375), .A2(new_n18377), .B(new_n18383), .Y(new_n18385));
  NAND2xp33_ASAP7_75t_L     g18129(.A(new_n18384), .B(new_n18385), .Y(new_n18386));
  OAI21xp33_ASAP7_75t_L     g18130(.A1(new_n18235), .A2(new_n18238), .B(new_n18241), .Y(new_n18387));
  XNOR2x2_ASAP7_75t_L       g18131(.A(new_n18386), .B(new_n18387), .Y(new_n18388));
  AOI22xp33_ASAP7_75t_L     g18132(.A1(new_n6002), .A2(\b[52] ), .B1(new_n5999), .B2(new_n8577), .Y(new_n18389));
  OAI221xp5_ASAP7_75t_L     g18133(.A1(new_n6544), .A2(new_n8249), .B1(new_n8228), .B2(new_n6309), .C(new_n18389), .Y(new_n18390));
  XNOR2x2_ASAP7_75t_L       g18134(.A(\a[44] ), .B(new_n18390), .Y(new_n18391));
  INVx1_ASAP7_75t_L         g18135(.A(new_n18391), .Y(new_n18392));
  NOR2xp33_ASAP7_75t_L      g18136(.A(new_n18392), .B(new_n18388), .Y(new_n18393));
  AND2x2_ASAP7_75t_L        g18137(.A(new_n18392), .B(new_n18388), .Y(new_n18394));
  NOR2xp33_ASAP7_75t_L      g18138(.A(new_n18393), .B(new_n18394), .Y(new_n18395));
  A2O1A1Ixp33_ASAP7_75t_L   g18139(.A1(new_n18248), .A2(new_n18305), .B(new_n18246), .C(new_n18395), .Y(new_n18396));
  INVx1_ASAP7_75t_L         g18140(.A(new_n18395), .Y(new_n18397));
  O2A1O1Ixp33_ASAP7_75t_L   g18141(.A1(new_n18114), .A2(new_n18121), .B(new_n18248), .C(new_n18246), .Y(new_n18398));
  NAND2xp33_ASAP7_75t_L     g18142(.A(new_n18398), .B(new_n18397), .Y(new_n18399));
  AND2x2_ASAP7_75t_L        g18143(.A(new_n18396), .B(new_n18399), .Y(new_n18400));
  NAND2xp33_ASAP7_75t_L     g18144(.A(new_n5247), .B(new_n9542), .Y(new_n18401));
  OAI221xp5_ASAP7_75t_L     g18145(.A1(new_n5253), .A2(new_n9534), .B1(new_n9199), .B2(new_n5241), .C(new_n18401), .Y(new_n18402));
  AOI21xp33_ASAP7_75t_L     g18146(.A1(new_n5526), .A2(\b[53] ), .B(new_n18402), .Y(new_n18403));
  NAND2xp33_ASAP7_75t_L     g18147(.A(\a[41] ), .B(new_n18403), .Y(new_n18404));
  A2O1A1Ixp33_ASAP7_75t_L   g18148(.A1(\b[53] ), .A2(new_n5526), .B(new_n18402), .C(new_n5244), .Y(new_n18405));
  AND2x2_ASAP7_75t_L        g18149(.A(new_n18405), .B(new_n18404), .Y(new_n18406));
  INVx1_ASAP7_75t_L         g18150(.A(new_n18406), .Y(new_n18407));
  XNOR2x2_ASAP7_75t_L       g18151(.A(new_n18407), .B(new_n18400), .Y(new_n18408));
  A2O1A1Ixp33_ASAP7_75t_L   g18152(.A1(new_n18255), .A2(new_n18172), .B(new_n18304), .C(new_n18408), .Y(new_n18409));
  NAND2xp33_ASAP7_75t_L     g18153(.A(new_n18256), .B(new_n18258), .Y(new_n18410));
  NOR2xp33_ASAP7_75t_L      g18154(.A(new_n18408), .B(new_n18410), .Y(new_n18411));
  INVx1_ASAP7_75t_L         g18155(.A(new_n18411), .Y(new_n18412));
  AND2x2_ASAP7_75t_L        g18156(.A(new_n18409), .B(new_n18412), .Y(new_n18413));
  AOI22xp33_ASAP7_75t_L     g18157(.A1(new_n4544), .A2(\b[58] ), .B1(new_n4542), .B2(new_n10857), .Y(new_n18414));
  OAI221xp5_ASAP7_75t_L     g18158(.A1(new_n4536), .A2(new_n10488), .B1(new_n10178), .B2(new_n4781), .C(new_n18414), .Y(new_n18415));
  XNOR2x2_ASAP7_75t_L       g18159(.A(\a[38] ), .B(new_n18415), .Y(new_n18416));
  NAND2xp33_ASAP7_75t_L     g18160(.A(new_n18416), .B(new_n18413), .Y(new_n18417));
  AO21x2_ASAP7_75t_L        g18161(.A1(new_n18409), .A2(new_n18412), .B(new_n18416), .Y(new_n18418));
  NAND2xp33_ASAP7_75t_L     g18162(.A(new_n18418), .B(new_n18417), .Y(new_n18419));
  NAND2xp33_ASAP7_75t_L     g18163(.A(new_n18265), .B(new_n18264), .Y(new_n18420));
  OAI21xp33_ASAP7_75t_L     g18164(.A1(new_n18260), .A2(new_n18263), .B(new_n18420), .Y(new_n18421));
  NOR2xp33_ASAP7_75t_L      g18165(.A(new_n18421), .B(new_n18419), .Y(new_n18422));
  AND2x2_ASAP7_75t_L        g18166(.A(new_n18421), .B(new_n18419), .Y(new_n18423));
  NAND2xp33_ASAP7_75t_L     g18167(.A(\b[61] ), .B(new_n3884), .Y(new_n18424));
  OAI221xp5_ASAP7_75t_L     g18168(.A1(new_n11226), .A2(new_n4312), .B1(new_n4114), .B2(new_n11920), .C(new_n18424), .Y(new_n18425));
  AOI21xp33_ASAP7_75t_L     g18169(.A1(new_n4111), .A2(\b[59] ), .B(new_n18425), .Y(new_n18426));
  NAND2xp33_ASAP7_75t_L     g18170(.A(\a[35] ), .B(new_n18426), .Y(new_n18427));
  A2O1A1Ixp33_ASAP7_75t_L   g18171(.A1(\b[59] ), .A2(new_n4111), .B(new_n18425), .C(new_n3878), .Y(new_n18428));
  AOI211xp5_ASAP7_75t_L     g18172(.A1(new_n18428), .A2(new_n18427), .B(new_n18422), .C(new_n18423), .Y(new_n18429));
  OA211x2_ASAP7_75t_L       g18173(.A1(new_n18422), .A2(new_n18423), .B(new_n18427), .C(new_n18428), .Y(new_n18430));
  NOR2xp33_ASAP7_75t_L      g18174(.A(new_n18429), .B(new_n18430), .Y(new_n18431));
  INVx1_ASAP7_75t_L         g18175(.A(new_n18431), .Y(new_n18432));
  NOR2xp33_ASAP7_75t_L      g18176(.A(new_n18432), .B(new_n18303), .Y(new_n18433));
  INVx1_ASAP7_75t_L         g18177(.A(new_n18433), .Y(new_n18434));
  NAND2xp33_ASAP7_75t_L     g18178(.A(new_n18432), .B(new_n18303), .Y(new_n18435));
  NAND2xp33_ASAP7_75t_L     g18179(.A(new_n18435), .B(new_n18434), .Y(new_n18436));
  A2O1A1O1Ixp25_ASAP7_75t_L g18180(.A1(new_n18150), .A2(new_n18033), .B(new_n18279), .C(new_n18285), .D(new_n18436), .Y(new_n18437));
  A2O1A1O1Ixp25_ASAP7_75t_L g18181(.A1(new_n18147), .A2(new_n18146), .B(new_n18034), .C(new_n18033), .D(new_n18279), .Y(new_n18438));
  O2A1O1Ixp33_ASAP7_75t_L   g18182(.A1(new_n18281), .A2(new_n18283), .B(new_n18275), .C(new_n18438), .Y(new_n18439));
  AND2x2_ASAP7_75t_L        g18183(.A(new_n18439), .B(new_n18436), .Y(new_n18440));
  NOR2xp33_ASAP7_75t_L      g18184(.A(new_n18437), .B(new_n18440), .Y(new_n18441));
  INVx1_ASAP7_75t_L         g18185(.A(new_n18441), .Y(new_n18442));
  A2O1A1O1Ixp25_ASAP7_75t_L g18186(.A1(new_n18163), .A2(new_n18292), .B(new_n18290), .C(new_n18287), .D(new_n18442), .Y(new_n18443));
  A2O1A1Ixp33_ASAP7_75t_L   g18187(.A1(new_n18292), .A2(new_n18163), .B(new_n18290), .C(new_n18287), .Y(new_n18444));
  NOR2xp33_ASAP7_75t_L      g18188(.A(new_n18441), .B(new_n18444), .Y(new_n18445));
  NOR2xp33_ASAP7_75t_L      g18189(.A(new_n18443), .B(new_n18445), .Y(\f[94] ));
  INVx1_ASAP7_75t_L         g18190(.A(new_n18400), .Y(new_n18447));
  O2A1O1Ixp33_ASAP7_75t_L   g18191(.A1(new_n18173), .A2(new_n18250), .B(new_n18247), .C(new_n18395), .Y(new_n18448));
  AOI22xp33_ASAP7_75t_L     g18192(.A1(new_n5249), .A2(\b[56] ), .B1(new_n5247), .B2(new_n10185), .Y(new_n18449));
  OAI221xp5_ASAP7_75t_L     g18193(.A1(new_n5241), .A2(new_n9534), .B1(new_n9199), .B2(new_n5521), .C(new_n18449), .Y(new_n18450));
  XNOR2x2_ASAP7_75t_L       g18194(.A(\a[41] ), .B(new_n18450), .Y(new_n18451));
  INVx1_ASAP7_75t_L         g18195(.A(new_n18451), .Y(new_n18452));
  AOI22xp33_ASAP7_75t_L     g18196(.A1(new_n6002), .A2(\b[53] ), .B1(new_n5999), .B2(new_n8889), .Y(new_n18453));
  OAI221xp5_ASAP7_75t_L     g18197(.A1(new_n6544), .A2(new_n8569), .B1(new_n8249), .B2(new_n6309), .C(new_n18453), .Y(new_n18454));
  XNOR2x2_ASAP7_75t_L       g18198(.A(\a[44] ), .B(new_n18454), .Y(new_n18455));
  INVx1_ASAP7_75t_L         g18199(.A(new_n18455), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18367), .Y(new_n18457));
  AOI22xp33_ASAP7_75t_L     g18201(.A1(new_n8645), .A2(\b[44] ), .B1(new_n8642), .B2(new_n7055), .Y(new_n18458));
  OAI221xp5_ASAP7_75t_L     g18202(.A1(new_n9322), .A2(new_n6195), .B1(new_n5680), .B2(new_n8965), .C(new_n18458), .Y(new_n18459));
  XNOR2x2_ASAP7_75t_L       g18203(.A(\a[53] ), .B(new_n18459), .Y(new_n18460));
  INVx1_ASAP7_75t_L         g18204(.A(new_n18460), .Y(new_n18461));
  AOI22xp33_ASAP7_75t_L     g18205(.A1(new_n9623), .A2(\b[41] ), .B1(new_n9620), .B2(new_n5669), .Y(new_n18462));
  OAI221xp5_ASAP7_75t_L     g18206(.A1(new_n10280), .A2(new_n5186), .B1(new_n5166), .B2(new_n12010), .C(new_n18462), .Y(new_n18463));
  XNOR2x2_ASAP7_75t_L       g18207(.A(\a[56] ), .B(new_n18463), .Y(new_n18464));
  INVx1_ASAP7_75t_L         g18208(.A(new_n18464), .Y(new_n18465));
  AOI22xp33_ASAP7_75t_L     g18209(.A1(new_n10594), .A2(\b[38] ), .B1(new_n10591), .B2(new_n4923), .Y(new_n18466));
  OAI221xp5_ASAP7_75t_L     g18210(.A1(new_n11335), .A2(new_n4701), .B1(new_n4465), .B2(new_n11330), .C(new_n18466), .Y(new_n18467));
  XNOR2x2_ASAP7_75t_L       g18211(.A(\a[59] ), .B(new_n18467), .Y(new_n18468));
  AOI22xp33_ASAP7_75t_L     g18212(.A1(new_n11656), .A2(\b[35] ), .B1(new_n11654), .B2(new_n5649), .Y(new_n18469));
  OAI221xp5_ASAP7_75t_L     g18213(.A1(new_n12364), .A2(new_n3827), .B1(new_n3807), .B2(new_n13003), .C(new_n18469), .Y(new_n18470));
  XNOR2x2_ASAP7_75t_L       g18214(.A(\a[62] ), .B(new_n18470), .Y(new_n18471));
  A2O1A1Ixp33_ASAP7_75t_L   g18215(.A1(new_n18326), .A2(new_n18327), .B(new_n18322), .C(new_n18321), .Y(new_n18472));
  NOR2xp33_ASAP7_75t_L      g18216(.A(new_n3419), .B(new_n12671), .Y(new_n18473));
  A2O1A1Ixp33_ASAP7_75t_L   g18217(.A1(\b[32] ), .A2(new_n12669), .B(new_n18473), .C(new_n18318), .Y(new_n18474));
  INVx1_ASAP7_75t_L         g18218(.A(new_n18474), .Y(new_n18475));
  O2A1O1Ixp33_ASAP7_75t_L   g18219(.A1(new_n12353), .A2(new_n12355), .B(\b[32] ), .C(new_n18473), .Y(new_n18476));
  A2O1A1Ixp33_ASAP7_75t_L   g18220(.A1(new_n12669), .A2(\b[31] ), .B(new_n18315), .C(new_n18476), .Y(new_n18477));
  INVx1_ASAP7_75t_L         g18221(.A(new_n18477), .Y(new_n18478));
  NOR3xp33_ASAP7_75t_L      g18222(.A(new_n18472), .B(new_n18475), .C(new_n18478), .Y(new_n18479));
  NOR2xp33_ASAP7_75t_L      g18223(.A(new_n18475), .B(new_n18478), .Y(new_n18480));
  A2O1A1O1Ixp25_ASAP7_75t_L g18224(.A1(new_n18327), .A2(new_n18326), .B(new_n18322), .C(new_n18321), .D(new_n18480), .Y(new_n18481));
  NOR2xp33_ASAP7_75t_L      g18225(.A(new_n18481), .B(new_n18479), .Y(new_n18482));
  NOR2xp33_ASAP7_75t_L      g18226(.A(new_n18471), .B(new_n18482), .Y(new_n18483));
  INVx1_ASAP7_75t_L         g18227(.A(new_n18471), .Y(new_n18484));
  NOR3xp33_ASAP7_75t_L      g18228(.A(new_n18484), .B(new_n18479), .C(new_n18481), .Y(new_n18485));
  NOR2xp33_ASAP7_75t_L      g18229(.A(new_n18485), .B(new_n18483), .Y(new_n18486));
  INVx1_ASAP7_75t_L         g18230(.A(new_n18486), .Y(new_n18487));
  NOR2xp33_ASAP7_75t_L      g18231(.A(new_n18468), .B(new_n18487), .Y(new_n18488));
  AND2x2_ASAP7_75t_L        g18232(.A(new_n18468), .B(new_n18487), .Y(new_n18489));
  NOR2xp33_ASAP7_75t_L      g18233(.A(new_n18488), .B(new_n18489), .Y(new_n18490));
  INVx1_ASAP7_75t_L         g18234(.A(new_n18490), .Y(new_n18491));
  O2A1O1Ixp33_ASAP7_75t_L   g18235(.A1(new_n18335), .A2(new_n18332), .B(new_n18337), .C(new_n18491), .Y(new_n18492));
  INVx1_ASAP7_75t_L         g18236(.A(new_n18492), .Y(new_n18493));
  A2O1A1Ixp33_ASAP7_75t_L   g18237(.A1(new_n18202), .A2(new_n18195), .B(new_n18332), .C(new_n18337), .Y(new_n18494));
  INVx1_ASAP7_75t_L         g18238(.A(new_n18494), .Y(new_n18495));
  NAND2xp33_ASAP7_75t_L     g18239(.A(new_n18491), .B(new_n18495), .Y(new_n18496));
  NAND3xp33_ASAP7_75t_L     g18240(.A(new_n18493), .B(new_n18465), .C(new_n18496), .Y(new_n18497));
  INVx1_ASAP7_75t_L         g18241(.A(new_n18497), .Y(new_n18498));
  AOI21xp33_ASAP7_75t_L     g18242(.A1(new_n18493), .A2(new_n18496), .B(new_n18465), .Y(new_n18499));
  NOR2xp33_ASAP7_75t_L      g18243(.A(new_n18499), .B(new_n18498), .Y(new_n18500));
  INVx1_ASAP7_75t_L         g18244(.A(new_n18500), .Y(new_n18501));
  A2O1A1O1Ixp25_ASAP7_75t_L g18245(.A1(new_n18344), .A2(new_n18204), .B(new_n18341), .C(new_n18346), .D(new_n18501), .Y(new_n18502));
  INVx1_ASAP7_75t_L         g18246(.A(new_n18502), .Y(new_n18503));
  NAND3xp33_ASAP7_75t_L     g18247(.A(new_n18501), .B(new_n18346), .C(new_n18343), .Y(new_n18504));
  NAND3xp33_ASAP7_75t_L     g18248(.A(new_n18503), .B(new_n18461), .C(new_n18504), .Y(new_n18505));
  INVx1_ASAP7_75t_L         g18249(.A(new_n18505), .Y(new_n18506));
  AOI21xp33_ASAP7_75t_L     g18250(.A1(new_n18503), .A2(new_n18504), .B(new_n18461), .Y(new_n18507));
  NOR2xp33_ASAP7_75t_L      g18251(.A(new_n18507), .B(new_n18506), .Y(new_n18508));
  NAND3xp33_ASAP7_75t_L     g18252(.A(new_n18361), .B(new_n18352), .C(new_n18508), .Y(new_n18509));
  O2A1O1Ixp33_ASAP7_75t_L   g18253(.A1(new_n18353), .A2(new_n18359), .B(new_n18352), .C(new_n18508), .Y(new_n18510));
  INVx1_ASAP7_75t_L         g18254(.A(new_n18510), .Y(new_n18511));
  AOI22xp33_ASAP7_75t_L     g18255(.A1(new_n7659), .A2(\b[47] ), .B1(new_n7656), .B2(new_n7323), .Y(new_n18512));
  OAI221xp5_ASAP7_75t_L     g18256(.A1(new_n8326), .A2(new_n7033), .B1(new_n6756), .B2(new_n7994), .C(new_n18512), .Y(new_n18513));
  XNOR2x2_ASAP7_75t_L       g18257(.A(\a[50] ), .B(new_n18513), .Y(new_n18514));
  NAND3xp33_ASAP7_75t_L     g18258(.A(new_n18511), .B(new_n18509), .C(new_n18514), .Y(new_n18515));
  AO21x2_ASAP7_75t_L        g18259(.A1(new_n18509), .A2(new_n18511), .B(new_n18514), .Y(new_n18516));
  AND2x2_ASAP7_75t_L        g18260(.A(new_n18515), .B(new_n18516), .Y(new_n18517));
  A2O1A1Ixp33_ASAP7_75t_L   g18261(.A1(new_n18369), .A2(new_n18372), .B(new_n18457), .C(new_n18517), .Y(new_n18518));
  NAND2xp33_ASAP7_75t_L     g18262(.A(new_n18367), .B(new_n18373), .Y(new_n18519));
  NOR2xp33_ASAP7_75t_L      g18263(.A(new_n18517), .B(new_n18519), .Y(new_n18520));
  INVx1_ASAP7_75t_L         g18264(.A(new_n18520), .Y(new_n18521));
  AND2x2_ASAP7_75t_L        g18265(.A(new_n18518), .B(new_n18521), .Y(new_n18522));
  INVx1_ASAP7_75t_L         g18266(.A(new_n18522), .Y(new_n18523));
  AOI22xp33_ASAP7_75t_L     g18267(.A1(new_n6822), .A2(\b[50] ), .B1(new_n6819), .B2(new_n8235), .Y(new_n18524));
  OAI221xp5_ASAP7_75t_L     g18268(.A1(new_n7392), .A2(new_n7907), .B1(new_n7333), .B2(new_n7115), .C(new_n18524), .Y(new_n18525));
  XNOR2x2_ASAP7_75t_L       g18269(.A(\a[47] ), .B(new_n18525), .Y(new_n18526));
  NAND2xp33_ASAP7_75t_L     g18270(.A(new_n18526), .B(new_n18523), .Y(new_n18527));
  NOR2xp33_ASAP7_75t_L      g18271(.A(new_n18526), .B(new_n18523), .Y(new_n18528));
  INVx1_ASAP7_75t_L         g18272(.A(new_n18528), .Y(new_n18529));
  AND2x2_ASAP7_75t_L        g18273(.A(new_n18527), .B(new_n18529), .Y(new_n18530));
  INVx1_ASAP7_75t_L         g18274(.A(new_n18530), .Y(new_n18531));
  NAND2xp33_ASAP7_75t_L     g18275(.A(new_n18375), .B(new_n18384), .Y(new_n18532));
  NOR2xp33_ASAP7_75t_L      g18276(.A(new_n18532), .B(new_n18531), .Y(new_n18533));
  A2O1A1Ixp33_ASAP7_75t_L   g18277(.A1(new_n18094), .A2(new_n18098), .B(new_n18231), .C(new_n18306), .Y(new_n18534));
  O2A1O1Ixp33_ASAP7_75t_L   g18278(.A1(new_n18376), .A2(new_n18534), .B(new_n18384), .C(new_n18530), .Y(new_n18535));
  NOR2xp33_ASAP7_75t_L      g18279(.A(new_n18535), .B(new_n18533), .Y(new_n18536));
  NAND2xp33_ASAP7_75t_L     g18280(.A(new_n18456), .B(new_n18536), .Y(new_n18537));
  INVx1_ASAP7_75t_L         g18281(.A(new_n18537), .Y(new_n18538));
  NOR2xp33_ASAP7_75t_L      g18282(.A(new_n18456), .B(new_n18536), .Y(new_n18539));
  NOR2xp33_ASAP7_75t_L      g18283(.A(new_n18539), .B(new_n18538), .Y(new_n18540));
  NOR2xp33_ASAP7_75t_L      g18284(.A(new_n18386), .B(new_n18387), .Y(new_n18541));
  NOR2xp33_ASAP7_75t_L      g18285(.A(new_n18541), .B(new_n18393), .Y(new_n18542));
  XNOR2x2_ASAP7_75t_L       g18286(.A(new_n18542), .B(new_n18540), .Y(new_n18543));
  XNOR2x2_ASAP7_75t_L       g18287(.A(new_n18452), .B(new_n18543), .Y(new_n18544));
  A2O1A1Ixp33_ASAP7_75t_L   g18288(.A1(new_n18407), .A2(new_n18447), .B(new_n18448), .C(new_n18544), .Y(new_n18545));
  INVx1_ASAP7_75t_L         g18289(.A(new_n18448), .Y(new_n18546));
  A2O1A1Ixp33_ASAP7_75t_L   g18290(.A1(new_n18399), .A2(new_n18396), .B(new_n18406), .C(new_n18546), .Y(new_n18547));
  NOR2xp33_ASAP7_75t_L      g18291(.A(new_n18547), .B(new_n18544), .Y(new_n18548));
  INVx1_ASAP7_75t_L         g18292(.A(new_n18548), .Y(new_n18549));
  AOI22xp33_ASAP7_75t_L     g18293(.A1(new_n4544), .A2(\b[59] ), .B1(new_n4542), .B2(new_n10887), .Y(new_n18550));
  OAI221xp5_ASAP7_75t_L     g18294(.A1(new_n4536), .A2(new_n10848), .B1(new_n10488), .B2(new_n4781), .C(new_n18550), .Y(new_n18551));
  XNOR2x2_ASAP7_75t_L       g18295(.A(\a[38] ), .B(new_n18551), .Y(new_n18552));
  NAND3xp33_ASAP7_75t_L     g18296(.A(new_n18549), .B(new_n18545), .C(new_n18552), .Y(new_n18553));
  AO21x2_ASAP7_75t_L        g18297(.A1(new_n18545), .A2(new_n18549), .B(new_n18552), .Y(new_n18554));
  NAND2xp33_ASAP7_75t_L     g18298(.A(new_n18553), .B(new_n18554), .Y(new_n18555));
  O2A1O1Ixp33_ASAP7_75t_L   g18299(.A1(new_n18410), .A2(new_n18408), .B(new_n18417), .C(new_n18555), .Y(new_n18556));
  INVx1_ASAP7_75t_L         g18300(.A(new_n18556), .Y(new_n18557));
  NAND2xp33_ASAP7_75t_L     g18301(.A(new_n18412), .B(new_n18417), .Y(new_n18558));
  INVx1_ASAP7_75t_L         g18302(.A(new_n18558), .Y(new_n18559));
  NAND2xp33_ASAP7_75t_L     g18303(.A(new_n18555), .B(new_n18559), .Y(new_n18560));
  AOI22xp33_ASAP7_75t_L     g18304(.A1(new_n3884), .A2(\b[62] ), .B1(new_n3881), .B2(new_n12280), .Y(new_n18561));
  OAI221xp5_ASAP7_75t_L     g18305(.A1(new_n4312), .A2(new_n11911), .B1(new_n11226), .B2(new_n4986), .C(new_n18561), .Y(new_n18562));
  XNOR2x2_ASAP7_75t_L       g18306(.A(\a[35] ), .B(new_n18562), .Y(new_n18563));
  AND3x1_ASAP7_75t_L        g18307(.A(new_n18560), .B(new_n18563), .C(new_n18557), .Y(new_n18564));
  AOI21xp33_ASAP7_75t_L     g18308(.A1(new_n18560), .A2(new_n18557), .B(new_n18563), .Y(new_n18565));
  NOR2xp33_ASAP7_75t_L      g18309(.A(new_n18565), .B(new_n18564), .Y(new_n18566));
  INVx1_ASAP7_75t_L         g18310(.A(new_n18423), .Y(new_n18567));
  O2A1O1Ixp33_ASAP7_75t_L   g18311(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n3261), .Y(new_n18568));
  O2A1O1Ixp33_ASAP7_75t_L   g18312(.A1(new_n3491), .A2(new_n18568), .B(\b[63] ), .C(new_n3251), .Y(new_n18569));
  A2O1A1O1Ixp25_ASAP7_75t_L g18313(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n3254), .D(new_n3491), .Y(new_n18570));
  NOR3xp33_ASAP7_75t_L      g18314(.A(new_n18570), .B(new_n12599), .C(\a[32] ), .Y(new_n18571));
  NOR2xp33_ASAP7_75t_L      g18315(.A(new_n18569), .B(new_n18571), .Y(new_n18572));
  A2O1A1O1Ixp25_ASAP7_75t_L g18316(.A1(new_n18427), .A2(new_n18428), .B(new_n18422), .C(new_n18567), .D(new_n18572), .Y(new_n18573));
  INVx1_ASAP7_75t_L         g18317(.A(new_n18573), .Y(new_n18574));
  INVx1_ASAP7_75t_L         g18318(.A(new_n18429), .Y(new_n18575));
  NAND3xp33_ASAP7_75t_L     g18319(.A(new_n18575), .B(new_n18567), .C(new_n18572), .Y(new_n18576));
  NAND2xp33_ASAP7_75t_L     g18320(.A(new_n18574), .B(new_n18576), .Y(new_n18577));
  XNOR2x2_ASAP7_75t_L       g18321(.A(new_n18566), .B(new_n18577), .Y(new_n18578));
  O2A1O1Ixp33_ASAP7_75t_L   g18322(.A1(new_n18303), .A2(new_n18432), .B(new_n18301), .C(new_n18578), .Y(new_n18579));
  A2O1A1Ixp33_ASAP7_75t_L   g18323(.A1(new_n18293), .A2(new_n18274), .B(new_n18299), .C(new_n18434), .Y(new_n18580));
  INVx1_ASAP7_75t_L         g18324(.A(new_n18578), .Y(new_n18581));
  NOR2xp33_ASAP7_75t_L      g18325(.A(new_n18580), .B(new_n18581), .Y(new_n18582));
  NOR2xp33_ASAP7_75t_L      g18326(.A(new_n18579), .B(new_n18582), .Y(new_n18583));
  A2O1A1Ixp33_ASAP7_75t_L   g18327(.A1(new_n18444), .A2(new_n18441), .B(new_n18437), .C(new_n18583), .Y(new_n18584));
  INVx1_ASAP7_75t_L         g18328(.A(new_n18584), .Y(new_n18585));
  NOR3xp33_ASAP7_75t_L      g18329(.A(new_n18443), .B(new_n18583), .C(new_n18437), .Y(new_n18586));
  NOR2xp33_ASAP7_75t_L      g18330(.A(new_n18586), .B(new_n18585), .Y(\f[95] ));
  AOI22xp33_ASAP7_75t_L     g18331(.A1(new_n6002), .A2(\b[54] ), .B1(new_n5999), .B2(new_n9208), .Y(new_n18588));
  OAI221xp5_ASAP7_75t_L     g18332(.A1(new_n6544), .A2(new_n8882), .B1(new_n8569), .B2(new_n6309), .C(new_n18588), .Y(new_n18589));
  XNOR2x2_ASAP7_75t_L       g18333(.A(\a[44] ), .B(new_n18589), .Y(new_n18590));
  INVx1_ASAP7_75t_L         g18334(.A(new_n18483), .Y(new_n18591));
  AOI22xp33_ASAP7_75t_L     g18335(.A1(new_n10594), .A2(\b[39] ), .B1(new_n10591), .B2(new_n5174), .Y(new_n18592));
  OAI221xp5_ASAP7_75t_L     g18336(.A1(new_n11335), .A2(new_n4915), .B1(new_n4701), .B2(new_n11330), .C(new_n18592), .Y(new_n18593));
  XNOR2x2_ASAP7_75t_L       g18337(.A(\a[59] ), .B(new_n18593), .Y(new_n18594));
  INVx1_ASAP7_75t_L         g18338(.A(new_n18594), .Y(new_n18595));
  AOI22xp33_ASAP7_75t_L     g18339(.A1(new_n11656), .A2(\b[36] ), .B1(new_n11654), .B2(new_n4473), .Y(new_n18596));
  OAI221xp5_ASAP7_75t_L     g18340(.A1(new_n12364), .A2(new_n4053), .B1(new_n3827), .B2(new_n13003), .C(new_n18596), .Y(new_n18597));
  XNOR2x2_ASAP7_75t_L       g18341(.A(\a[62] ), .B(new_n18597), .Y(new_n18598));
  INVx1_ASAP7_75t_L         g18342(.A(new_n18472), .Y(new_n18599));
  NOR2xp33_ASAP7_75t_L      g18343(.A(new_n3443), .B(new_n12671), .Y(new_n18600));
  A2O1A1Ixp33_ASAP7_75t_L   g18344(.A1(new_n12669), .A2(\b[33] ), .B(new_n18600), .C(new_n3251), .Y(new_n18601));
  INVx1_ASAP7_75t_L         g18345(.A(new_n18601), .Y(new_n18602));
  O2A1O1Ixp33_ASAP7_75t_L   g18346(.A1(new_n12353), .A2(new_n12355), .B(\b[33] ), .C(new_n18600), .Y(new_n18603));
  NAND2xp33_ASAP7_75t_L     g18347(.A(\a[32] ), .B(new_n18603), .Y(new_n18604));
  INVx1_ASAP7_75t_L         g18348(.A(new_n18604), .Y(new_n18605));
  OAI21xp33_ASAP7_75t_L     g18349(.A1(new_n18602), .A2(new_n18605), .B(new_n18476), .Y(new_n18606));
  NOR2xp33_ASAP7_75t_L      g18350(.A(new_n18602), .B(new_n18605), .Y(new_n18607));
  A2O1A1Ixp33_ASAP7_75t_L   g18351(.A1(new_n12669), .A2(\b[32] ), .B(new_n18473), .C(new_n18607), .Y(new_n18608));
  AND2x2_ASAP7_75t_L        g18352(.A(new_n18606), .B(new_n18608), .Y(new_n18609));
  INVx1_ASAP7_75t_L         g18353(.A(new_n18609), .Y(new_n18610));
  O2A1O1Ixp33_ASAP7_75t_L   g18354(.A1(new_n18475), .A2(new_n18599), .B(new_n18477), .C(new_n18610), .Y(new_n18611));
  INVx1_ASAP7_75t_L         g18355(.A(new_n18611), .Y(new_n18612));
  A2O1A1O1Ixp25_ASAP7_75t_L g18356(.A1(new_n18327), .A2(new_n18326), .B(new_n18322), .C(new_n18321), .D(new_n18475), .Y(new_n18613));
  A2O1A1O1Ixp25_ASAP7_75t_L g18357(.A1(new_n12669), .A2(\b[31] ), .B(new_n18315), .C(new_n18476), .D(new_n18613), .Y(new_n18614));
  NAND2xp33_ASAP7_75t_L     g18358(.A(new_n18610), .B(new_n18614), .Y(new_n18615));
  NAND2xp33_ASAP7_75t_L     g18359(.A(new_n18615), .B(new_n18612), .Y(new_n18616));
  NOR2xp33_ASAP7_75t_L      g18360(.A(new_n18598), .B(new_n18616), .Y(new_n18617));
  INVx1_ASAP7_75t_L         g18361(.A(new_n18617), .Y(new_n18618));
  NAND2xp33_ASAP7_75t_L     g18362(.A(new_n18598), .B(new_n18616), .Y(new_n18619));
  AND2x2_ASAP7_75t_L        g18363(.A(new_n18619), .B(new_n18618), .Y(new_n18620));
  NAND2xp33_ASAP7_75t_L     g18364(.A(new_n18595), .B(new_n18620), .Y(new_n18621));
  INVx1_ASAP7_75t_L         g18365(.A(new_n18621), .Y(new_n18622));
  NOR2xp33_ASAP7_75t_L      g18366(.A(new_n18595), .B(new_n18620), .Y(new_n18623));
  NOR2xp33_ASAP7_75t_L      g18367(.A(new_n18623), .B(new_n18622), .Y(new_n18624));
  INVx1_ASAP7_75t_L         g18368(.A(new_n18624), .Y(new_n18625));
  O2A1O1Ixp33_ASAP7_75t_L   g18369(.A1(new_n18468), .A2(new_n18487), .B(new_n18591), .C(new_n18625), .Y(new_n18626));
  NOR3xp33_ASAP7_75t_L      g18370(.A(new_n18624), .B(new_n18488), .C(new_n18483), .Y(new_n18627));
  NOR2xp33_ASAP7_75t_L      g18371(.A(new_n18627), .B(new_n18626), .Y(new_n18628));
  AOI22xp33_ASAP7_75t_L     g18372(.A1(new_n9623), .A2(\b[42] ), .B1(new_n9620), .B2(new_n5688), .Y(new_n18629));
  OAI221xp5_ASAP7_75t_L     g18373(.A1(new_n10280), .A2(new_n5666), .B1(new_n5186), .B2(new_n12010), .C(new_n18629), .Y(new_n18630));
  XNOR2x2_ASAP7_75t_L       g18374(.A(\a[56] ), .B(new_n18630), .Y(new_n18631));
  INVx1_ASAP7_75t_L         g18375(.A(new_n18631), .Y(new_n18632));
  XNOR2x2_ASAP7_75t_L       g18376(.A(new_n18632), .B(new_n18628), .Y(new_n18633));
  A2O1A1Ixp33_ASAP7_75t_L   g18377(.A1(new_n18337), .A2(new_n18334), .B(new_n18491), .C(new_n18497), .Y(new_n18634));
  INVx1_ASAP7_75t_L         g18378(.A(new_n18634), .Y(new_n18635));
  AND2x2_ASAP7_75t_L        g18379(.A(new_n18635), .B(new_n18633), .Y(new_n18636));
  O2A1O1Ixp33_ASAP7_75t_L   g18380(.A1(new_n18495), .A2(new_n18491), .B(new_n18497), .C(new_n18633), .Y(new_n18637));
  NOR2xp33_ASAP7_75t_L      g18381(.A(new_n18637), .B(new_n18636), .Y(new_n18638));
  AOI22xp33_ASAP7_75t_L     g18382(.A1(new_n8645), .A2(\b[45] ), .B1(new_n8642), .B2(new_n6764), .Y(new_n18639));
  OAI221xp5_ASAP7_75t_L     g18383(.A1(new_n9322), .A2(new_n6220), .B1(new_n6195), .B2(new_n8965), .C(new_n18639), .Y(new_n18640));
  XNOR2x2_ASAP7_75t_L       g18384(.A(\a[53] ), .B(new_n18640), .Y(new_n18641));
  INVx1_ASAP7_75t_L         g18385(.A(new_n18641), .Y(new_n18642));
  XNOR2x2_ASAP7_75t_L       g18386(.A(new_n18642), .B(new_n18638), .Y(new_n18643));
  A2O1A1Ixp33_ASAP7_75t_L   g18387(.A1(new_n18346), .A2(new_n18343), .B(new_n18501), .C(new_n18505), .Y(new_n18644));
  INVx1_ASAP7_75t_L         g18388(.A(new_n18644), .Y(new_n18645));
  AND2x2_ASAP7_75t_L        g18389(.A(new_n18645), .B(new_n18643), .Y(new_n18646));
  A2O1A1O1Ixp25_ASAP7_75t_L g18390(.A1(new_n18346), .A2(new_n18343), .B(new_n18501), .C(new_n18505), .D(new_n18643), .Y(new_n18647));
  NOR2xp33_ASAP7_75t_L      g18391(.A(new_n18647), .B(new_n18646), .Y(new_n18648));
  AOI22xp33_ASAP7_75t_L     g18392(.A1(new_n7659), .A2(\b[48] ), .B1(new_n7656), .B2(new_n7341), .Y(new_n18649));
  OAI221xp5_ASAP7_75t_L     g18393(.A1(new_n8326), .A2(new_n7316), .B1(new_n7033), .B2(new_n7994), .C(new_n18649), .Y(new_n18650));
  XNOR2x2_ASAP7_75t_L       g18394(.A(\a[50] ), .B(new_n18650), .Y(new_n18651));
  INVx1_ASAP7_75t_L         g18395(.A(new_n18651), .Y(new_n18652));
  XNOR2x2_ASAP7_75t_L       g18396(.A(new_n18652), .B(new_n18648), .Y(new_n18653));
  A2O1A1Ixp33_ASAP7_75t_L   g18397(.A1(new_n18361), .A2(new_n18352), .B(new_n18508), .C(new_n18515), .Y(new_n18654));
  AND2x2_ASAP7_75t_L        g18398(.A(new_n18654), .B(new_n18653), .Y(new_n18655));
  NOR2xp33_ASAP7_75t_L      g18399(.A(new_n18654), .B(new_n18653), .Y(new_n18656));
  NOR2xp33_ASAP7_75t_L      g18400(.A(new_n18656), .B(new_n18655), .Y(new_n18657));
  AOI22xp33_ASAP7_75t_L     g18401(.A1(new_n6822), .A2(\b[51] ), .B1(new_n6819), .B2(new_n8257), .Y(new_n18658));
  OAI221xp5_ASAP7_75t_L     g18402(.A1(new_n7392), .A2(new_n8228), .B1(new_n7907), .B2(new_n7115), .C(new_n18658), .Y(new_n18659));
  XNOR2x2_ASAP7_75t_L       g18403(.A(new_n6816), .B(new_n18659), .Y(new_n18660));
  XOR2x2_ASAP7_75t_L        g18404(.A(new_n18660), .B(new_n18657), .Y(new_n18661));
  INVx1_ASAP7_75t_L         g18405(.A(new_n18661), .Y(new_n18662));
  NAND3xp33_ASAP7_75t_L     g18406(.A(new_n18529), .B(new_n18521), .C(new_n18662), .Y(new_n18663));
  O2A1O1Ixp33_ASAP7_75t_L   g18407(.A1(new_n18523), .A2(new_n18526), .B(new_n18521), .C(new_n18662), .Y(new_n18664));
  INVx1_ASAP7_75t_L         g18408(.A(new_n18664), .Y(new_n18665));
  AND2x2_ASAP7_75t_L        g18409(.A(new_n18665), .B(new_n18663), .Y(new_n18666));
  INVx1_ASAP7_75t_L         g18410(.A(new_n18666), .Y(new_n18667));
  NAND2xp33_ASAP7_75t_L     g18411(.A(new_n18590), .B(new_n18667), .Y(new_n18668));
  NOR2xp33_ASAP7_75t_L      g18412(.A(new_n18590), .B(new_n18667), .Y(new_n18669));
  INVx1_ASAP7_75t_L         g18413(.A(new_n18669), .Y(new_n18670));
  AND2x2_ASAP7_75t_L        g18414(.A(new_n18668), .B(new_n18670), .Y(new_n18671));
  A2O1A1Ixp33_ASAP7_75t_L   g18415(.A1(new_n18536), .A2(new_n18456), .B(new_n18533), .C(new_n18671), .Y(new_n18672));
  OR3x1_ASAP7_75t_L         g18416(.A(new_n18671), .B(new_n18533), .C(new_n18538), .Y(new_n18673));
  NAND2xp33_ASAP7_75t_L     g18417(.A(new_n18672), .B(new_n18673), .Y(new_n18674));
  AOI22xp33_ASAP7_75t_L     g18418(.A1(new_n5249), .A2(\b[57] ), .B1(new_n5247), .B2(new_n10495), .Y(new_n18675));
  OAI221xp5_ASAP7_75t_L     g18419(.A1(new_n5241), .A2(new_n10178), .B1(new_n9534), .B2(new_n5521), .C(new_n18675), .Y(new_n18676));
  XNOR2x2_ASAP7_75t_L       g18420(.A(\a[41] ), .B(new_n18676), .Y(new_n18677));
  XNOR2x2_ASAP7_75t_L       g18421(.A(new_n18677), .B(new_n18674), .Y(new_n18678));
  MAJx2_ASAP7_75t_L         g18422(.A(new_n18540), .B(new_n18452), .C(new_n18542), .Y(new_n18679));
  XNOR2x2_ASAP7_75t_L       g18423(.A(new_n18679), .B(new_n18678), .Y(new_n18680));
  AOI22xp33_ASAP7_75t_L     g18424(.A1(new_n4544), .A2(\b[60] ), .B1(new_n4542), .B2(new_n11234), .Y(new_n18681));
  OAI221xp5_ASAP7_75t_L     g18425(.A1(new_n4536), .A2(new_n10881), .B1(new_n10848), .B2(new_n4781), .C(new_n18681), .Y(new_n18682));
  XNOR2x2_ASAP7_75t_L       g18426(.A(\a[38] ), .B(new_n18682), .Y(new_n18683));
  INVx1_ASAP7_75t_L         g18427(.A(new_n18683), .Y(new_n18684));
  XNOR2x2_ASAP7_75t_L       g18428(.A(new_n18684), .B(new_n18680), .Y(new_n18685));
  A2O1A1Ixp33_ASAP7_75t_L   g18429(.A1(new_n18552), .A2(new_n18545), .B(new_n18548), .C(new_n18685), .Y(new_n18686));
  NAND2xp33_ASAP7_75t_L     g18430(.A(new_n18549), .B(new_n18553), .Y(new_n18687));
  OR2x4_ASAP7_75t_L         g18431(.A(new_n18687), .B(new_n18685), .Y(new_n18688));
  AND2x2_ASAP7_75t_L        g18432(.A(new_n18686), .B(new_n18688), .Y(new_n18689));
  NAND2xp33_ASAP7_75t_L     g18433(.A(\b[63] ), .B(new_n3884), .Y(new_n18690));
  A2O1A1Ixp33_ASAP7_75t_L   g18434(.A1(new_n12607), .A2(new_n12603), .B(new_n4114), .C(new_n18690), .Y(new_n18691));
  AOI221xp5_ASAP7_75t_L     g18435(.A1(\b[61] ), .A2(new_n4111), .B1(\b[62] ), .B2(new_n3874), .C(new_n18691), .Y(new_n18692));
  XNOR2x2_ASAP7_75t_L       g18436(.A(new_n3878), .B(new_n18692), .Y(new_n18693));
  INVx1_ASAP7_75t_L         g18437(.A(new_n18693), .Y(new_n18694));
  INVx1_ASAP7_75t_L         g18438(.A(new_n18555), .Y(new_n18695));
  A2O1A1O1Ixp25_ASAP7_75t_L g18439(.A1(new_n18413), .A2(new_n18416), .B(new_n18411), .C(new_n18695), .D(new_n18564), .Y(new_n18696));
  NAND2xp33_ASAP7_75t_L     g18440(.A(new_n18694), .B(new_n18696), .Y(new_n18697));
  A2O1A1Ixp33_ASAP7_75t_L   g18441(.A1(new_n18560), .A2(new_n18563), .B(new_n18556), .C(new_n18693), .Y(new_n18698));
  AND2x2_ASAP7_75t_L        g18442(.A(new_n18698), .B(new_n18697), .Y(new_n18699));
  NOR2xp33_ASAP7_75t_L      g18443(.A(new_n18689), .B(new_n18699), .Y(new_n18700));
  NAND2xp33_ASAP7_75t_L     g18444(.A(new_n18689), .B(new_n18699), .Y(new_n18701));
  INVx1_ASAP7_75t_L         g18445(.A(new_n18701), .Y(new_n18702));
  NOR2xp33_ASAP7_75t_L      g18446(.A(new_n18700), .B(new_n18702), .Y(new_n18703));
  A2O1A1Ixp33_ASAP7_75t_L   g18447(.A1(new_n18567), .A2(new_n18575), .B(new_n18572), .C(new_n18566), .Y(new_n18704));
  AND2x2_ASAP7_75t_L        g18448(.A(new_n18576), .B(new_n18704), .Y(new_n18705));
  NAND2xp33_ASAP7_75t_L     g18449(.A(new_n18705), .B(new_n18703), .Y(new_n18706));
  INVx1_ASAP7_75t_L         g18450(.A(new_n18576), .Y(new_n18707));
  INVx1_ASAP7_75t_L         g18451(.A(new_n18703), .Y(new_n18708));
  A2O1A1Ixp33_ASAP7_75t_L   g18452(.A1(new_n18574), .A2(new_n18566), .B(new_n18707), .C(new_n18708), .Y(new_n18709));
  NAND2xp33_ASAP7_75t_L     g18453(.A(new_n18709), .B(new_n18706), .Y(new_n18710));
  A2O1A1O1Ixp25_ASAP7_75t_L g18454(.A1(new_n18434), .A2(new_n18301), .B(new_n18578), .C(new_n18584), .D(new_n18710), .Y(new_n18711));
  A2O1A1Ixp33_ASAP7_75t_L   g18455(.A1(new_n18434), .A2(new_n18301), .B(new_n18578), .C(new_n18584), .Y(new_n18712));
  AOI21xp33_ASAP7_75t_L     g18456(.A1(new_n18709), .A2(new_n18706), .B(new_n18712), .Y(new_n18713));
  NOR2xp33_ASAP7_75t_L      g18457(.A(new_n18711), .B(new_n18713), .Y(\f[96] ));
  INVx1_ASAP7_75t_L         g18458(.A(new_n18696), .Y(new_n18715));
  NAND2xp33_ASAP7_75t_L     g18459(.A(new_n18684), .B(new_n18680), .Y(new_n18716));
  A2O1A1Ixp33_ASAP7_75t_L   g18460(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n3881), .Y(new_n18717));
  AOI22xp33_ASAP7_75t_L     g18461(.A1(new_n3874), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4111), .Y(new_n18718));
  NAND3xp33_ASAP7_75t_L     g18462(.A(new_n18717), .B(\a[35] ), .C(new_n18718), .Y(new_n18719));
  INVx1_ASAP7_75t_L         g18463(.A(new_n18719), .Y(new_n18720));
  A2O1A1O1Ixp25_ASAP7_75t_L g18464(.A1(new_n13507), .A2(new_n13506), .B(new_n4114), .C(new_n18718), .D(\a[35] ), .Y(new_n18721));
  NOR2xp33_ASAP7_75t_L      g18465(.A(new_n18721), .B(new_n18720), .Y(new_n18722));
  O2A1O1Ixp33_ASAP7_75t_L   g18466(.A1(new_n18687), .A2(new_n18685), .B(new_n18716), .C(new_n18722), .Y(new_n18723));
  INVx1_ASAP7_75t_L         g18467(.A(new_n18723), .Y(new_n18724));
  NAND3xp33_ASAP7_75t_L     g18468(.A(new_n18688), .B(new_n18716), .C(new_n18722), .Y(new_n18725));
  AND2x2_ASAP7_75t_L        g18469(.A(new_n18724), .B(new_n18725), .Y(new_n18726));
  INVx1_ASAP7_75t_L         g18470(.A(new_n18678), .Y(new_n18727));
  A2O1A1O1Ixp25_ASAP7_75t_L g18471(.A1(new_n18456), .A2(new_n18536), .B(new_n18533), .C(new_n18668), .D(new_n18669), .Y(new_n18728));
  INVx1_ASAP7_75t_L         g18472(.A(new_n18728), .Y(new_n18729));
  AOI22xp33_ASAP7_75t_L     g18473(.A1(new_n10594), .A2(\b[40] ), .B1(new_n10591), .B2(new_n5194), .Y(new_n18730));
  OAI221xp5_ASAP7_75t_L     g18474(.A1(new_n11335), .A2(new_n5166), .B1(new_n4915), .B2(new_n11330), .C(new_n18730), .Y(new_n18731));
  XNOR2x2_ASAP7_75t_L       g18475(.A(\a[59] ), .B(new_n18731), .Y(new_n18732));
  INVx1_ASAP7_75t_L         g18476(.A(new_n18732), .Y(new_n18733));
  NOR2xp33_ASAP7_75t_L      g18477(.A(new_n3807), .B(new_n12671), .Y(new_n18734));
  A2O1A1O1Ixp25_ASAP7_75t_L g18478(.A1(new_n12669), .A2(\b[32] ), .B(new_n18473), .C(new_n18604), .D(new_n18602), .Y(new_n18735));
  A2O1A1Ixp33_ASAP7_75t_L   g18479(.A1(new_n12669), .A2(\b[34] ), .B(new_n18734), .C(new_n18735), .Y(new_n18736));
  O2A1O1Ixp33_ASAP7_75t_L   g18480(.A1(new_n12353), .A2(new_n12355), .B(\b[34] ), .C(new_n18734), .Y(new_n18737));
  INVx1_ASAP7_75t_L         g18481(.A(new_n18737), .Y(new_n18738));
  O2A1O1Ixp33_ASAP7_75t_L   g18482(.A1(new_n18476), .A2(new_n18605), .B(new_n18601), .C(new_n18738), .Y(new_n18739));
  INVx1_ASAP7_75t_L         g18483(.A(new_n18739), .Y(new_n18740));
  NAND2xp33_ASAP7_75t_L     g18484(.A(new_n18736), .B(new_n18740), .Y(new_n18741));
  NAND2xp33_ASAP7_75t_L     g18485(.A(\b[37] ), .B(new_n11656), .Y(new_n18742));
  OAI221xp5_ASAP7_75t_L     g18486(.A1(new_n4465), .A2(new_n12364), .B1(new_n12022), .B2(new_n13559), .C(new_n18742), .Y(new_n18743));
  AOI21xp33_ASAP7_75t_L     g18487(.A1(new_n12021), .A2(\b[35] ), .B(new_n18743), .Y(new_n18744));
  NAND2xp33_ASAP7_75t_L     g18488(.A(\a[62] ), .B(new_n18744), .Y(new_n18745));
  A2O1A1Ixp33_ASAP7_75t_L   g18489(.A1(\b[35] ), .A2(new_n12021), .B(new_n18743), .C(new_n11651), .Y(new_n18746));
  AND3x1_ASAP7_75t_L        g18490(.A(new_n18745), .B(new_n18746), .C(new_n18741), .Y(new_n18747));
  AND2x2_ASAP7_75t_L        g18491(.A(new_n18746), .B(new_n18745), .Y(new_n18748));
  NOR2xp33_ASAP7_75t_L      g18492(.A(new_n18741), .B(new_n18748), .Y(new_n18749));
  NOR2xp33_ASAP7_75t_L      g18493(.A(new_n18747), .B(new_n18749), .Y(new_n18750));
  INVx1_ASAP7_75t_L         g18494(.A(new_n18750), .Y(new_n18751));
  O2A1O1Ixp33_ASAP7_75t_L   g18495(.A1(new_n18598), .A2(new_n18616), .B(new_n18612), .C(new_n18751), .Y(new_n18752));
  INVx1_ASAP7_75t_L         g18496(.A(new_n18752), .Y(new_n18753));
  O2A1O1Ixp33_ASAP7_75t_L   g18497(.A1(new_n18478), .A2(new_n18613), .B(new_n18609), .C(new_n18617), .Y(new_n18754));
  NAND2xp33_ASAP7_75t_L     g18498(.A(new_n18754), .B(new_n18751), .Y(new_n18755));
  NAND3xp33_ASAP7_75t_L     g18499(.A(new_n18753), .B(new_n18733), .C(new_n18755), .Y(new_n18756));
  AO21x2_ASAP7_75t_L        g18500(.A1(new_n18755), .A2(new_n18753), .B(new_n18733), .Y(new_n18757));
  AND2x2_ASAP7_75t_L        g18501(.A(new_n18756), .B(new_n18757), .Y(new_n18758));
  A2O1A1Ixp33_ASAP7_75t_L   g18502(.A1(new_n18620), .A2(new_n18595), .B(new_n18626), .C(new_n18758), .Y(new_n18759));
  INVx1_ASAP7_75t_L         g18503(.A(new_n18488), .Y(new_n18760));
  A2O1A1Ixp33_ASAP7_75t_L   g18504(.A1(new_n18591), .A2(new_n18760), .B(new_n18623), .C(new_n18621), .Y(new_n18761));
  NOR2xp33_ASAP7_75t_L      g18505(.A(new_n18761), .B(new_n18758), .Y(new_n18762));
  INVx1_ASAP7_75t_L         g18506(.A(new_n18762), .Y(new_n18763));
  AOI22xp33_ASAP7_75t_L     g18507(.A1(new_n9623), .A2(\b[43] ), .B1(new_n9620), .B2(new_n6202), .Y(new_n18764));
  OAI221xp5_ASAP7_75t_L     g18508(.A1(new_n10280), .A2(new_n5680), .B1(new_n5666), .B2(new_n12010), .C(new_n18764), .Y(new_n18765));
  XNOR2x2_ASAP7_75t_L       g18509(.A(\a[56] ), .B(new_n18765), .Y(new_n18766));
  NAND3xp33_ASAP7_75t_L     g18510(.A(new_n18759), .B(new_n18763), .C(new_n18766), .Y(new_n18767));
  AO21x2_ASAP7_75t_L        g18511(.A1(new_n18763), .A2(new_n18759), .B(new_n18766), .Y(new_n18768));
  AND2x2_ASAP7_75t_L        g18512(.A(new_n18767), .B(new_n18768), .Y(new_n18769));
  INVx1_ASAP7_75t_L         g18513(.A(new_n18769), .Y(new_n18770));
  NAND2xp33_ASAP7_75t_L     g18514(.A(new_n18632), .B(new_n18628), .Y(new_n18771));
  A2O1A1Ixp33_ASAP7_75t_L   g18515(.A1(new_n18497), .A2(new_n18493), .B(new_n18633), .C(new_n18771), .Y(new_n18772));
  NOR2xp33_ASAP7_75t_L      g18516(.A(new_n18772), .B(new_n18770), .Y(new_n18773));
  INVx1_ASAP7_75t_L         g18517(.A(new_n18773), .Y(new_n18774));
  O2A1O1Ixp33_ASAP7_75t_L   g18518(.A1(new_n18635), .A2(new_n18633), .B(new_n18771), .C(new_n18769), .Y(new_n18775));
  INVx1_ASAP7_75t_L         g18519(.A(new_n18775), .Y(new_n18776));
  AOI22xp33_ASAP7_75t_L     g18520(.A1(new_n8645), .A2(\b[46] ), .B1(new_n8642), .B2(new_n7041), .Y(new_n18777));
  OAI221xp5_ASAP7_75t_L     g18521(.A1(new_n9322), .A2(new_n6756), .B1(new_n6220), .B2(new_n8965), .C(new_n18777), .Y(new_n18778));
  XNOR2x2_ASAP7_75t_L       g18522(.A(\a[53] ), .B(new_n18778), .Y(new_n18779));
  NAND3xp33_ASAP7_75t_L     g18523(.A(new_n18774), .B(new_n18776), .C(new_n18779), .Y(new_n18780));
  AO21x2_ASAP7_75t_L        g18524(.A1(new_n18776), .A2(new_n18774), .B(new_n18779), .Y(new_n18781));
  AND2x2_ASAP7_75t_L        g18525(.A(new_n18780), .B(new_n18781), .Y(new_n18782));
  INVx1_ASAP7_75t_L         g18526(.A(new_n18782), .Y(new_n18783));
  NAND2xp33_ASAP7_75t_L     g18527(.A(new_n18642), .B(new_n18638), .Y(new_n18784));
  A2O1A1Ixp33_ASAP7_75t_L   g18528(.A1(new_n18505), .A2(new_n18503), .B(new_n18643), .C(new_n18784), .Y(new_n18785));
  NOR2xp33_ASAP7_75t_L      g18529(.A(new_n18785), .B(new_n18783), .Y(new_n18786));
  INVx1_ASAP7_75t_L         g18530(.A(new_n18786), .Y(new_n18787));
  O2A1O1Ixp33_ASAP7_75t_L   g18531(.A1(new_n18645), .A2(new_n18643), .B(new_n18784), .C(new_n18782), .Y(new_n18788));
  INVx1_ASAP7_75t_L         g18532(.A(new_n18788), .Y(new_n18789));
  AOI22xp33_ASAP7_75t_L     g18533(.A1(new_n7659), .A2(\b[49] ), .B1(new_n7656), .B2(new_n7914), .Y(new_n18790));
  OAI221xp5_ASAP7_75t_L     g18534(.A1(new_n8326), .A2(new_n7333), .B1(new_n7316), .B2(new_n7994), .C(new_n18790), .Y(new_n18791));
  XNOR2x2_ASAP7_75t_L       g18535(.A(\a[50] ), .B(new_n18791), .Y(new_n18792));
  NAND3xp33_ASAP7_75t_L     g18536(.A(new_n18787), .B(new_n18789), .C(new_n18792), .Y(new_n18793));
  AO21x2_ASAP7_75t_L        g18537(.A1(new_n18789), .A2(new_n18787), .B(new_n18792), .Y(new_n18794));
  AND2x2_ASAP7_75t_L        g18538(.A(new_n18793), .B(new_n18794), .Y(new_n18795));
  AOI21xp33_ASAP7_75t_L     g18539(.A1(new_n18652), .A2(new_n18648), .B(new_n18656), .Y(new_n18796));
  NAND2xp33_ASAP7_75t_L     g18540(.A(new_n18796), .B(new_n18795), .Y(new_n18797));
  INVx1_ASAP7_75t_L         g18541(.A(new_n18795), .Y(new_n18798));
  A2O1A1Ixp33_ASAP7_75t_L   g18542(.A1(new_n18652), .A2(new_n18648), .B(new_n18656), .C(new_n18798), .Y(new_n18799));
  AOI22xp33_ASAP7_75t_L     g18543(.A1(new_n6822), .A2(\b[52] ), .B1(new_n6819), .B2(new_n8577), .Y(new_n18800));
  OAI221xp5_ASAP7_75t_L     g18544(.A1(new_n7392), .A2(new_n8249), .B1(new_n8228), .B2(new_n7115), .C(new_n18800), .Y(new_n18801));
  XNOR2x2_ASAP7_75t_L       g18545(.A(\a[47] ), .B(new_n18801), .Y(new_n18802));
  NAND3xp33_ASAP7_75t_L     g18546(.A(new_n18799), .B(new_n18797), .C(new_n18802), .Y(new_n18803));
  AO21x2_ASAP7_75t_L        g18547(.A1(new_n18797), .A2(new_n18799), .B(new_n18802), .Y(new_n18804));
  AND2x2_ASAP7_75t_L        g18548(.A(new_n18803), .B(new_n18804), .Y(new_n18805));
  A2O1A1Ixp33_ASAP7_75t_L   g18549(.A1(new_n18660), .A2(new_n18657), .B(new_n18664), .C(new_n18805), .Y(new_n18806));
  NAND2xp33_ASAP7_75t_L     g18550(.A(new_n18660), .B(new_n18657), .Y(new_n18807));
  INVx1_ASAP7_75t_L         g18551(.A(new_n18805), .Y(new_n18808));
  NAND3xp33_ASAP7_75t_L     g18552(.A(new_n18808), .B(new_n18665), .C(new_n18807), .Y(new_n18809));
  AND2x2_ASAP7_75t_L        g18553(.A(new_n18806), .B(new_n18809), .Y(new_n18810));
  NAND2xp33_ASAP7_75t_L     g18554(.A(new_n5999), .B(new_n9542), .Y(new_n18811));
  OAI221xp5_ASAP7_75t_L     g18555(.A1(new_n6312), .A2(new_n9534), .B1(new_n9199), .B2(new_n6544), .C(new_n18811), .Y(new_n18812));
  AOI21xp33_ASAP7_75t_L     g18556(.A1(new_n6308), .A2(\b[53] ), .B(new_n18812), .Y(new_n18813));
  NAND2xp33_ASAP7_75t_L     g18557(.A(\a[44] ), .B(new_n18813), .Y(new_n18814));
  A2O1A1Ixp33_ASAP7_75t_L   g18558(.A1(\b[53] ), .A2(new_n6308), .B(new_n18812), .C(new_n5996), .Y(new_n18815));
  AND2x2_ASAP7_75t_L        g18559(.A(new_n18815), .B(new_n18814), .Y(new_n18816));
  INVx1_ASAP7_75t_L         g18560(.A(new_n18816), .Y(new_n18817));
  XNOR2x2_ASAP7_75t_L       g18561(.A(new_n18817), .B(new_n18810), .Y(new_n18818));
  NAND2xp33_ASAP7_75t_L     g18562(.A(new_n18818), .B(new_n18729), .Y(new_n18819));
  NOR2xp33_ASAP7_75t_L      g18563(.A(new_n18818), .B(new_n18729), .Y(new_n18820));
  INVx1_ASAP7_75t_L         g18564(.A(new_n18820), .Y(new_n18821));
  AOI22xp33_ASAP7_75t_L     g18565(.A1(new_n5249), .A2(\b[58] ), .B1(new_n5247), .B2(new_n10857), .Y(new_n18822));
  OAI221xp5_ASAP7_75t_L     g18566(.A1(new_n5241), .A2(new_n10488), .B1(new_n10178), .B2(new_n5521), .C(new_n18822), .Y(new_n18823));
  XNOR2x2_ASAP7_75t_L       g18567(.A(\a[41] ), .B(new_n18823), .Y(new_n18824));
  NAND3xp33_ASAP7_75t_L     g18568(.A(new_n18821), .B(new_n18819), .C(new_n18824), .Y(new_n18825));
  AO21x2_ASAP7_75t_L        g18569(.A1(new_n18819), .A2(new_n18821), .B(new_n18824), .Y(new_n18826));
  NAND2xp33_ASAP7_75t_L     g18570(.A(new_n18825), .B(new_n18826), .Y(new_n18827));
  NOR2xp33_ASAP7_75t_L      g18571(.A(new_n18677), .B(new_n18674), .Y(new_n18828));
  AOI211xp5_ASAP7_75t_L     g18572(.A1(new_n18727), .A2(new_n18679), .B(new_n18827), .C(new_n18828), .Y(new_n18829));
  A2O1A1Ixp33_ASAP7_75t_L   g18573(.A1(new_n18727), .A2(new_n18679), .B(new_n18828), .C(new_n18827), .Y(new_n18830));
  INVx1_ASAP7_75t_L         g18574(.A(new_n18830), .Y(new_n18831));
  NOR2xp33_ASAP7_75t_L      g18575(.A(new_n18829), .B(new_n18831), .Y(new_n18832));
  NAND2xp33_ASAP7_75t_L     g18576(.A(\b[61] ), .B(new_n4544), .Y(new_n18833));
  OAI221xp5_ASAP7_75t_L     g18577(.A1(new_n11226), .A2(new_n4536), .B1(new_n4549), .B2(new_n11920), .C(new_n18833), .Y(new_n18834));
  AOI21xp33_ASAP7_75t_L     g18578(.A1(new_n4780), .A2(\b[59] ), .B(new_n18834), .Y(new_n18835));
  NAND2xp33_ASAP7_75t_L     g18579(.A(\a[38] ), .B(new_n18835), .Y(new_n18836));
  A2O1A1Ixp33_ASAP7_75t_L   g18580(.A1(\b[59] ), .A2(new_n4780), .B(new_n18834), .C(new_n4539), .Y(new_n18837));
  NAND2xp33_ASAP7_75t_L     g18581(.A(new_n18837), .B(new_n18836), .Y(new_n18838));
  NAND2xp33_ASAP7_75t_L     g18582(.A(new_n18838), .B(new_n18832), .Y(new_n18839));
  OAI211xp5_ASAP7_75t_L     g18583(.A1(new_n18829), .A2(new_n18831), .B(new_n18836), .C(new_n18837), .Y(new_n18840));
  AND2x2_ASAP7_75t_L        g18584(.A(new_n18840), .B(new_n18839), .Y(new_n18841));
  NAND2xp33_ASAP7_75t_L     g18585(.A(new_n18841), .B(new_n18726), .Y(new_n18842));
  INVx1_ASAP7_75t_L         g18586(.A(new_n18726), .Y(new_n18843));
  INVx1_ASAP7_75t_L         g18587(.A(new_n18841), .Y(new_n18844));
  NAND2xp33_ASAP7_75t_L     g18588(.A(new_n18844), .B(new_n18843), .Y(new_n18845));
  NAND2xp33_ASAP7_75t_L     g18589(.A(new_n18842), .B(new_n18845), .Y(new_n18846));
  O2A1O1Ixp33_ASAP7_75t_L   g18590(.A1(new_n18693), .A2(new_n18715), .B(new_n18701), .C(new_n18846), .Y(new_n18847));
  AND3x1_ASAP7_75t_L        g18591(.A(new_n18701), .B(new_n18846), .C(new_n18697), .Y(new_n18848));
  NOR2xp33_ASAP7_75t_L      g18592(.A(new_n18847), .B(new_n18848), .Y(new_n18849));
  A2O1A1Ixp33_ASAP7_75t_L   g18593(.A1(new_n18705), .A2(new_n18703), .B(new_n18711), .C(new_n18849), .Y(new_n18850));
  INVx1_ASAP7_75t_L         g18594(.A(new_n18850), .Y(new_n18851));
  INVx1_ASAP7_75t_L         g18595(.A(new_n18579), .Y(new_n18852));
  A2O1A1Ixp33_ASAP7_75t_L   g18596(.A1(new_n18584), .A2(new_n18852), .B(new_n18710), .C(new_n18706), .Y(new_n18853));
  NOR2xp33_ASAP7_75t_L      g18597(.A(new_n18849), .B(new_n18853), .Y(new_n18854));
  NOR2xp33_ASAP7_75t_L      g18598(.A(new_n18854), .B(new_n18851), .Y(\f[97] ));
  INVx1_ASAP7_75t_L         g18599(.A(new_n18810), .Y(new_n18856));
  A2O1A1O1Ixp25_ASAP7_75t_L g18600(.A1(new_n18529), .A2(new_n18521), .B(new_n18662), .C(new_n18807), .D(new_n18805), .Y(new_n18857));
  AOI22xp33_ASAP7_75t_L     g18601(.A1(new_n6002), .A2(\b[56] ), .B1(new_n5999), .B2(new_n10185), .Y(new_n18858));
  OAI221xp5_ASAP7_75t_L     g18602(.A1(new_n6544), .A2(new_n9534), .B1(new_n9199), .B2(new_n6309), .C(new_n18858), .Y(new_n18859));
  XNOR2x2_ASAP7_75t_L       g18603(.A(\a[44] ), .B(new_n18859), .Y(new_n18860));
  INVx1_ASAP7_75t_L         g18604(.A(new_n18860), .Y(new_n18861));
  AOI22xp33_ASAP7_75t_L     g18605(.A1(new_n6822), .A2(\b[53] ), .B1(new_n6819), .B2(new_n8889), .Y(new_n18862));
  OAI221xp5_ASAP7_75t_L     g18606(.A1(new_n7392), .A2(new_n8569), .B1(new_n8249), .B2(new_n7115), .C(new_n18862), .Y(new_n18863));
  XNOR2x2_ASAP7_75t_L       g18607(.A(\a[47] ), .B(new_n18863), .Y(new_n18864));
  INVx1_ASAP7_75t_L         g18608(.A(new_n18864), .Y(new_n18865));
  AOI22xp33_ASAP7_75t_L     g18609(.A1(new_n9623), .A2(\b[44] ), .B1(new_n9620), .B2(new_n7055), .Y(new_n18866));
  OAI221xp5_ASAP7_75t_L     g18610(.A1(new_n10280), .A2(new_n6195), .B1(new_n5680), .B2(new_n12010), .C(new_n18866), .Y(new_n18867));
  XNOR2x2_ASAP7_75t_L       g18611(.A(\a[56] ), .B(new_n18867), .Y(new_n18868));
  INVx1_ASAP7_75t_L         g18612(.A(new_n18868), .Y(new_n18869));
  AOI22xp33_ASAP7_75t_L     g18613(.A1(new_n10594), .A2(\b[41] ), .B1(new_n10591), .B2(new_n5669), .Y(new_n18870));
  OAI221xp5_ASAP7_75t_L     g18614(.A1(new_n11335), .A2(new_n5186), .B1(new_n5166), .B2(new_n11330), .C(new_n18870), .Y(new_n18871));
  XNOR2x2_ASAP7_75t_L       g18615(.A(\a[59] ), .B(new_n18871), .Y(new_n18872));
  AOI22xp33_ASAP7_75t_L     g18616(.A1(new_n11656), .A2(\b[38] ), .B1(new_n11654), .B2(new_n4923), .Y(new_n18873));
  OAI221xp5_ASAP7_75t_L     g18617(.A1(new_n12364), .A2(new_n4701), .B1(new_n4465), .B2(new_n13003), .C(new_n18873), .Y(new_n18874));
  XNOR2x2_ASAP7_75t_L       g18618(.A(\a[62] ), .B(new_n18874), .Y(new_n18875));
  A2O1A1Ixp33_ASAP7_75t_L   g18619(.A1(new_n18745), .A2(new_n18746), .B(new_n18741), .C(new_n18740), .Y(new_n18876));
  NOR2xp33_ASAP7_75t_L      g18620(.A(new_n3827), .B(new_n12671), .Y(new_n18877));
  INVx1_ASAP7_75t_L         g18621(.A(new_n18877), .Y(new_n18878));
  O2A1O1Ixp33_ASAP7_75t_L   g18622(.A1(new_n12356), .A2(new_n4053), .B(new_n18878), .C(new_n18738), .Y(new_n18879));
  O2A1O1Ixp33_ASAP7_75t_L   g18623(.A1(new_n12353), .A2(new_n12355), .B(\b[35] ), .C(new_n18877), .Y(new_n18880));
  A2O1A1Ixp33_ASAP7_75t_L   g18624(.A1(new_n12669), .A2(\b[34] ), .B(new_n18734), .C(new_n18880), .Y(new_n18881));
  INVx1_ASAP7_75t_L         g18625(.A(new_n18881), .Y(new_n18882));
  NOR3xp33_ASAP7_75t_L      g18626(.A(new_n18876), .B(new_n18879), .C(new_n18882), .Y(new_n18883));
  NOR2xp33_ASAP7_75t_L      g18627(.A(new_n18882), .B(new_n18879), .Y(new_n18884));
  A2O1A1O1Ixp25_ASAP7_75t_L g18628(.A1(new_n18746), .A2(new_n18745), .B(new_n18741), .C(new_n18740), .D(new_n18884), .Y(new_n18885));
  NOR2xp33_ASAP7_75t_L      g18629(.A(new_n18885), .B(new_n18883), .Y(new_n18886));
  NOR2xp33_ASAP7_75t_L      g18630(.A(new_n18875), .B(new_n18886), .Y(new_n18887));
  INVx1_ASAP7_75t_L         g18631(.A(new_n18887), .Y(new_n18888));
  NAND2xp33_ASAP7_75t_L     g18632(.A(new_n18875), .B(new_n18886), .Y(new_n18889));
  NAND2xp33_ASAP7_75t_L     g18633(.A(new_n18889), .B(new_n18888), .Y(new_n18890));
  NOR2xp33_ASAP7_75t_L      g18634(.A(new_n18872), .B(new_n18890), .Y(new_n18891));
  INVx1_ASAP7_75t_L         g18635(.A(new_n18872), .Y(new_n18892));
  AOI21xp33_ASAP7_75t_L     g18636(.A1(new_n18888), .A2(new_n18889), .B(new_n18892), .Y(new_n18893));
  NOR2xp33_ASAP7_75t_L      g18637(.A(new_n18893), .B(new_n18891), .Y(new_n18894));
  INVx1_ASAP7_75t_L         g18638(.A(new_n18894), .Y(new_n18895));
  O2A1O1Ixp33_ASAP7_75t_L   g18639(.A1(new_n18754), .A2(new_n18751), .B(new_n18756), .C(new_n18895), .Y(new_n18896));
  INVx1_ASAP7_75t_L         g18640(.A(new_n18896), .Y(new_n18897));
  NAND3xp33_ASAP7_75t_L     g18641(.A(new_n18895), .B(new_n18756), .C(new_n18753), .Y(new_n18898));
  NAND3xp33_ASAP7_75t_L     g18642(.A(new_n18897), .B(new_n18869), .C(new_n18898), .Y(new_n18899));
  INVx1_ASAP7_75t_L         g18643(.A(new_n18899), .Y(new_n18900));
  AOI21xp33_ASAP7_75t_L     g18644(.A1(new_n18897), .A2(new_n18898), .B(new_n18869), .Y(new_n18901));
  NOR2xp33_ASAP7_75t_L      g18645(.A(new_n18901), .B(new_n18900), .Y(new_n18902));
  NAND3xp33_ASAP7_75t_L     g18646(.A(new_n18902), .B(new_n18767), .C(new_n18763), .Y(new_n18903));
  O2A1O1Ixp33_ASAP7_75t_L   g18647(.A1(new_n18761), .A2(new_n18758), .B(new_n18767), .C(new_n18902), .Y(new_n18904));
  INVx1_ASAP7_75t_L         g18648(.A(new_n18904), .Y(new_n18905));
  AOI22xp33_ASAP7_75t_L     g18649(.A1(new_n8645), .A2(\b[47] ), .B1(new_n8642), .B2(new_n7323), .Y(new_n18906));
  OAI221xp5_ASAP7_75t_L     g18650(.A1(new_n9322), .A2(new_n7033), .B1(new_n6756), .B2(new_n8965), .C(new_n18906), .Y(new_n18907));
  XNOR2x2_ASAP7_75t_L       g18651(.A(\a[53] ), .B(new_n18907), .Y(new_n18908));
  NAND3xp33_ASAP7_75t_L     g18652(.A(new_n18905), .B(new_n18903), .C(new_n18908), .Y(new_n18909));
  AO21x2_ASAP7_75t_L        g18653(.A1(new_n18903), .A2(new_n18905), .B(new_n18908), .Y(new_n18910));
  AND2x2_ASAP7_75t_L        g18654(.A(new_n18909), .B(new_n18910), .Y(new_n18911));
  INVx1_ASAP7_75t_L         g18655(.A(new_n18911), .Y(new_n18912));
  O2A1O1Ixp33_ASAP7_75t_L   g18656(.A1(new_n18770), .A2(new_n18772), .B(new_n18780), .C(new_n18912), .Y(new_n18913));
  INVx1_ASAP7_75t_L         g18657(.A(new_n18913), .Y(new_n18914));
  NAND3xp33_ASAP7_75t_L     g18658(.A(new_n18912), .B(new_n18780), .C(new_n18774), .Y(new_n18915));
  NAND2xp33_ASAP7_75t_L     g18659(.A(new_n18915), .B(new_n18914), .Y(new_n18916));
  AOI22xp33_ASAP7_75t_L     g18660(.A1(new_n7659), .A2(\b[50] ), .B1(new_n7656), .B2(new_n8235), .Y(new_n18917));
  OAI221xp5_ASAP7_75t_L     g18661(.A1(new_n8326), .A2(new_n7907), .B1(new_n7333), .B2(new_n7994), .C(new_n18917), .Y(new_n18918));
  XNOR2x2_ASAP7_75t_L       g18662(.A(\a[50] ), .B(new_n18918), .Y(new_n18919));
  NAND2xp33_ASAP7_75t_L     g18663(.A(new_n18919), .B(new_n18916), .Y(new_n18920));
  INVx1_ASAP7_75t_L         g18664(.A(new_n18919), .Y(new_n18921));
  NAND3xp33_ASAP7_75t_L     g18665(.A(new_n18914), .B(new_n18915), .C(new_n18921), .Y(new_n18922));
  AND2x2_ASAP7_75t_L        g18666(.A(new_n18922), .B(new_n18920), .Y(new_n18923));
  INVx1_ASAP7_75t_L         g18667(.A(new_n18923), .Y(new_n18924));
  NAND2xp33_ASAP7_75t_L     g18668(.A(new_n18787), .B(new_n18793), .Y(new_n18925));
  NOR2xp33_ASAP7_75t_L      g18669(.A(new_n18925), .B(new_n18924), .Y(new_n18926));
  O2A1O1Ixp33_ASAP7_75t_L   g18670(.A1(new_n18783), .A2(new_n18785), .B(new_n18793), .C(new_n18923), .Y(new_n18927));
  NOR2xp33_ASAP7_75t_L      g18671(.A(new_n18927), .B(new_n18926), .Y(new_n18928));
  NAND2xp33_ASAP7_75t_L     g18672(.A(new_n18865), .B(new_n18928), .Y(new_n18929));
  INVx1_ASAP7_75t_L         g18673(.A(new_n18929), .Y(new_n18930));
  NOR2xp33_ASAP7_75t_L      g18674(.A(new_n18865), .B(new_n18928), .Y(new_n18931));
  NOR2xp33_ASAP7_75t_L      g18675(.A(new_n18931), .B(new_n18930), .Y(new_n18932));
  INVx1_ASAP7_75t_L         g18676(.A(new_n18932), .Y(new_n18933));
  NAND2xp33_ASAP7_75t_L     g18677(.A(new_n18797), .B(new_n18803), .Y(new_n18934));
  NOR2xp33_ASAP7_75t_L      g18678(.A(new_n18934), .B(new_n18933), .Y(new_n18935));
  INVx1_ASAP7_75t_L         g18679(.A(new_n18935), .Y(new_n18936));
  INVx1_ASAP7_75t_L         g18680(.A(new_n18797), .Y(new_n18937));
  A2O1A1Ixp33_ASAP7_75t_L   g18681(.A1(new_n18799), .A2(new_n18802), .B(new_n18937), .C(new_n18933), .Y(new_n18938));
  NAND3xp33_ASAP7_75t_L     g18682(.A(new_n18936), .B(new_n18861), .C(new_n18938), .Y(new_n18939));
  AO21x2_ASAP7_75t_L        g18683(.A1(new_n18938), .A2(new_n18936), .B(new_n18861), .Y(new_n18940));
  AND2x2_ASAP7_75t_L        g18684(.A(new_n18939), .B(new_n18940), .Y(new_n18941));
  A2O1A1Ixp33_ASAP7_75t_L   g18685(.A1(new_n18817), .A2(new_n18856), .B(new_n18857), .C(new_n18941), .Y(new_n18942));
  INVx1_ASAP7_75t_L         g18686(.A(new_n18857), .Y(new_n18943));
  A2O1A1Ixp33_ASAP7_75t_L   g18687(.A1(new_n18809), .A2(new_n18806), .B(new_n18816), .C(new_n18943), .Y(new_n18944));
  NOR2xp33_ASAP7_75t_L      g18688(.A(new_n18944), .B(new_n18941), .Y(new_n18945));
  INVx1_ASAP7_75t_L         g18689(.A(new_n18945), .Y(new_n18946));
  AOI22xp33_ASAP7_75t_L     g18690(.A1(new_n5249), .A2(\b[59] ), .B1(new_n5247), .B2(new_n10887), .Y(new_n18947));
  OAI221xp5_ASAP7_75t_L     g18691(.A1(new_n5241), .A2(new_n10848), .B1(new_n10488), .B2(new_n5521), .C(new_n18947), .Y(new_n18948));
  XNOR2x2_ASAP7_75t_L       g18692(.A(\a[41] ), .B(new_n18948), .Y(new_n18949));
  NAND3xp33_ASAP7_75t_L     g18693(.A(new_n18946), .B(new_n18942), .C(new_n18949), .Y(new_n18950));
  INVx1_ASAP7_75t_L         g18694(.A(new_n18950), .Y(new_n18951));
  AOI21xp33_ASAP7_75t_L     g18695(.A1(new_n18946), .A2(new_n18942), .B(new_n18949), .Y(new_n18952));
  NOR2xp33_ASAP7_75t_L      g18696(.A(new_n18952), .B(new_n18951), .Y(new_n18953));
  INVx1_ASAP7_75t_L         g18697(.A(new_n18953), .Y(new_n18954));
  O2A1O1Ixp33_ASAP7_75t_L   g18698(.A1(new_n18729), .A2(new_n18818), .B(new_n18825), .C(new_n18954), .Y(new_n18955));
  INVx1_ASAP7_75t_L         g18699(.A(new_n18955), .Y(new_n18956));
  NAND3xp33_ASAP7_75t_L     g18700(.A(new_n18954), .B(new_n18825), .C(new_n18821), .Y(new_n18957));
  AOI22xp33_ASAP7_75t_L     g18701(.A1(new_n4544), .A2(\b[62] ), .B1(new_n4542), .B2(new_n12280), .Y(new_n18958));
  OAI221xp5_ASAP7_75t_L     g18702(.A1(new_n4536), .A2(new_n11911), .B1(new_n11226), .B2(new_n4781), .C(new_n18958), .Y(new_n18959));
  XNOR2x2_ASAP7_75t_L       g18703(.A(\a[38] ), .B(new_n18959), .Y(new_n18960));
  NAND3xp33_ASAP7_75t_L     g18704(.A(new_n18956), .B(new_n18957), .C(new_n18960), .Y(new_n18961));
  INVx1_ASAP7_75t_L         g18705(.A(new_n18961), .Y(new_n18962));
  AOI21xp33_ASAP7_75t_L     g18706(.A1(new_n18956), .A2(new_n18957), .B(new_n18960), .Y(new_n18963));
  NOR2xp33_ASAP7_75t_L      g18707(.A(new_n18963), .B(new_n18962), .Y(new_n18964));
  O2A1O1Ixp33_ASAP7_75t_L   g18708(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n4114), .Y(new_n18965));
  O2A1O1Ixp33_ASAP7_75t_L   g18709(.A1(new_n4111), .A2(new_n18965), .B(\b[63] ), .C(new_n3878), .Y(new_n18966));
  A2O1A1O1Ixp25_ASAP7_75t_L g18710(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n3881), .D(new_n4111), .Y(new_n18967));
  NOR3xp33_ASAP7_75t_L      g18711(.A(new_n18967), .B(new_n12599), .C(\a[35] ), .Y(new_n18968));
  NOR2xp33_ASAP7_75t_L      g18712(.A(new_n18966), .B(new_n18968), .Y(new_n18969));
  A2O1A1O1Ixp25_ASAP7_75t_L g18713(.A1(new_n18836), .A2(new_n18837), .B(new_n18829), .C(new_n18830), .D(new_n18969), .Y(new_n18970));
  INVx1_ASAP7_75t_L         g18714(.A(new_n18970), .Y(new_n18971));
  NAND3xp33_ASAP7_75t_L     g18715(.A(new_n18839), .B(new_n18830), .C(new_n18969), .Y(new_n18972));
  NAND2xp33_ASAP7_75t_L     g18716(.A(new_n18971), .B(new_n18972), .Y(new_n18973));
  XOR2x2_ASAP7_75t_L        g18717(.A(new_n18973), .B(new_n18964), .Y(new_n18974));
  INVx1_ASAP7_75t_L         g18718(.A(new_n18974), .Y(new_n18975));
  O2A1O1Ixp33_ASAP7_75t_L   g18719(.A1(new_n18843), .A2(new_n18844), .B(new_n18724), .C(new_n18975), .Y(new_n18976));
  A2O1A1Ixp33_ASAP7_75t_L   g18720(.A1(new_n18716), .A2(new_n18688), .B(new_n18722), .C(new_n18842), .Y(new_n18977));
  NOR2xp33_ASAP7_75t_L      g18721(.A(new_n18974), .B(new_n18977), .Y(new_n18978));
  NOR2xp33_ASAP7_75t_L      g18722(.A(new_n18976), .B(new_n18978), .Y(new_n18979));
  A2O1A1Ixp33_ASAP7_75t_L   g18723(.A1(new_n18853), .A2(new_n18849), .B(new_n18847), .C(new_n18979), .Y(new_n18980));
  INVx1_ASAP7_75t_L         g18724(.A(new_n18980), .Y(new_n18981));
  A2O1A1Ixp33_ASAP7_75t_L   g18725(.A1(new_n18701), .A2(new_n18697), .B(new_n18846), .C(new_n18850), .Y(new_n18982));
  NOR2xp33_ASAP7_75t_L      g18726(.A(new_n18979), .B(new_n18982), .Y(new_n18983));
  NOR2xp33_ASAP7_75t_L      g18727(.A(new_n18981), .B(new_n18983), .Y(\f[98] ));
  INVx1_ASAP7_75t_L         g18728(.A(new_n18972), .Y(new_n18985));
  AOI22xp33_ASAP7_75t_L     g18729(.A1(new_n6822), .A2(\b[54] ), .B1(new_n6819), .B2(new_n9208), .Y(new_n18986));
  OAI221xp5_ASAP7_75t_L     g18730(.A1(new_n7392), .A2(new_n8882), .B1(new_n8569), .B2(new_n7115), .C(new_n18986), .Y(new_n18987));
  XNOR2x2_ASAP7_75t_L       g18731(.A(\a[47] ), .B(new_n18987), .Y(new_n18988));
  INVx1_ASAP7_75t_L         g18732(.A(new_n18988), .Y(new_n18989));
  AOI22xp33_ASAP7_75t_L     g18733(.A1(new_n9623), .A2(\b[45] ), .B1(new_n9620), .B2(new_n6764), .Y(new_n18990));
  OAI221xp5_ASAP7_75t_L     g18734(.A1(new_n10280), .A2(new_n6220), .B1(new_n6195), .B2(new_n12010), .C(new_n18990), .Y(new_n18991));
  XNOR2x2_ASAP7_75t_L       g18735(.A(\a[56] ), .B(new_n18991), .Y(new_n18992));
  INVx1_ASAP7_75t_L         g18736(.A(new_n18992), .Y(new_n18993));
  INVx1_ASAP7_75t_L         g18737(.A(new_n18876), .Y(new_n18994));
  NOR2xp33_ASAP7_75t_L      g18738(.A(new_n4053), .B(new_n12671), .Y(new_n18995));
  O2A1O1Ixp33_ASAP7_75t_L   g18739(.A1(new_n4053), .A2(new_n12356), .B(new_n18878), .C(new_n3878), .Y(new_n18996));
  AOI211xp5_ASAP7_75t_L     g18740(.A1(new_n12669), .A2(\b[35] ), .B(new_n18877), .C(\a[35] ), .Y(new_n18997));
  NOR2xp33_ASAP7_75t_L      g18741(.A(new_n18997), .B(new_n18996), .Y(new_n18998));
  INVx1_ASAP7_75t_L         g18742(.A(new_n18998), .Y(new_n18999));
  A2O1A1Ixp33_ASAP7_75t_L   g18743(.A1(new_n12669), .A2(\b[36] ), .B(new_n18995), .C(new_n18999), .Y(new_n19000));
  O2A1O1Ixp33_ASAP7_75t_L   g18744(.A1(new_n12353), .A2(new_n12355), .B(\b[36] ), .C(new_n18995), .Y(new_n19001));
  NAND2xp33_ASAP7_75t_L     g18745(.A(new_n19001), .B(new_n18998), .Y(new_n19002));
  AND2x2_ASAP7_75t_L        g18746(.A(new_n19002), .B(new_n19000), .Y(new_n19003));
  INVx1_ASAP7_75t_L         g18747(.A(new_n19003), .Y(new_n19004));
  O2A1O1Ixp33_ASAP7_75t_L   g18748(.A1(new_n18879), .A2(new_n18994), .B(new_n18881), .C(new_n19004), .Y(new_n19005));
  INVx1_ASAP7_75t_L         g18749(.A(new_n19005), .Y(new_n19006));
  A2O1A1O1Ixp25_ASAP7_75t_L g18750(.A1(new_n18746), .A2(new_n18745), .B(new_n18741), .C(new_n18740), .D(new_n18879), .Y(new_n19007));
  A2O1A1O1Ixp25_ASAP7_75t_L g18751(.A1(new_n12669), .A2(\b[34] ), .B(new_n18734), .C(new_n18880), .D(new_n19007), .Y(new_n19008));
  NAND2xp33_ASAP7_75t_L     g18752(.A(new_n19004), .B(new_n19008), .Y(new_n19009));
  NAND2xp33_ASAP7_75t_L     g18753(.A(new_n19009), .B(new_n19006), .Y(new_n19010));
  AOI22xp33_ASAP7_75t_L     g18754(.A1(new_n11656), .A2(\b[39] ), .B1(new_n11654), .B2(new_n5174), .Y(new_n19011));
  OAI221xp5_ASAP7_75t_L     g18755(.A1(new_n12364), .A2(new_n4915), .B1(new_n4701), .B2(new_n13003), .C(new_n19011), .Y(new_n19012));
  XNOR2x2_ASAP7_75t_L       g18756(.A(\a[62] ), .B(new_n19012), .Y(new_n19013));
  AND2x2_ASAP7_75t_L        g18757(.A(new_n19013), .B(new_n19010), .Y(new_n19014));
  NOR2xp33_ASAP7_75t_L      g18758(.A(new_n19013), .B(new_n19010), .Y(new_n19015));
  NOR2xp33_ASAP7_75t_L      g18759(.A(new_n19015), .B(new_n19014), .Y(new_n19016));
  AOI22xp33_ASAP7_75t_L     g18760(.A1(new_n10594), .A2(\b[42] ), .B1(new_n10591), .B2(new_n5688), .Y(new_n19017));
  OAI221xp5_ASAP7_75t_L     g18761(.A1(new_n11335), .A2(new_n5666), .B1(new_n5186), .B2(new_n11330), .C(new_n19017), .Y(new_n19018));
  XNOR2x2_ASAP7_75t_L       g18762(.A(\a[59] ), .B(new_n19018), .Y(new_n19019));
  INVx1_ASAP7_75t_L         g18763(.A(new_n19019), .Y(new_n19020));
  XNOR2x2_ASAP7_75t_L       g18764(.A(new_n19020), .B(new_n19016), .Y(new_n19021));
  O2A1O1Ixp33_ASAP7_75t_L   g18765(.A1(new_n18872), .A2(new_n18890), .B(new_n18888), .C(new_n19021), .Y(new_n19022));
  INVx1_ASAP7_75t_L         g18766(.A(new_n18875), .Y(new_n19023));
  O2A1O1Ixp33_ASAP7_75t_L   g18767(.A1(new_n18883), .A2(new_n18885), .B(new_n19023), .C(new_n18891), .Y(new_n19024));
  AND2x2_ASAP7_75t_L        g18768(.A(new_n19024), .B(new_n19021), .Y(new_n19025));
  NOR2xp33_ASAP7_75t_L      g18769(.A(new_n19022), .B(new_n19025), .Y(new_n19026));
  XNOR2x2_ASAP7_75t_L       g18770(.A(new_n18993), .B(new_n19026), .Y(new_n19027));
  A2O1A1Ixp33_ASAP7_75t_L   g18771(.A1(new_n18756), .A2(new_n18753), .B(new_n18895), .C(new_n18899), .Y(new_n19028));
  INVx1_ASAP7_75t_L         g18772(.A(new_n19028), .Y(new_n19029));
  AND2x2_ASAP7_75t_L        g18773(.A(new_n19029), .B(new_n19027), .Y(new_n19030));
  A2O1A1O1Ixp25_ASAP7_75t_L g18774(.A1(new_n18756), .A2(new_n18753), .B(new_n18895), .C(new_n18899), .D(new_n19027), .Y(new_n19031));
  NOR2xp33_ASAP7_75t_L      g18775(.A(new_n19031), .B(new_n19030), .Y(new_n19032));
  AOI22xp33_ASAP7_75t_L     g18776(.A1(new_n8645), .A2(\b[48] ), .B1(new_n8642), .B2(new_n7341), .Y(new_n19033));
  OAI221xp5_ASAP7_75t_L     g18777(.A1(new_n9322), .A2(new_n7316), .B1(new_n7033), .B2(new_n8965), .C(new_n19033), .Y(new_n19034));
  XNOR2x2_ASAP7_75t_L       g18778(.A(\a[53] ), .B(new_n19034), .Y(new_n19035));
  INVx1_ASAP7_75t_L         g18779(.A(new_n19035), .Y(new_n19036));
  XNOR2x2_ASAP7_75t_L       g18780(.A(new_n19036), .B(new_n19032), .Y(new_n19037));
  A2O1A1Ixp33_ASAP7_75t_L   g18781(.A1(new_n18767), .A2(new_n18763), .B(new_n18902), .C(new_n18909), .Y(new_n19038));
  AND2x2_ASAP7_75t_L        g18782(.A(new_n19038), .B(new_n19037), .Y(new_n19039));
  NOR2xp33_ASAP7_75t_L      g18783(.A(new_n19038), .B(new_n19037), .Y(new_n19040));
  NOR2xp33_ASAP7_75t_L      g18784(.A(new_n19040), .B(new_n19039), .Y(new_n19041));
  AOI22xp33_ASAP7_75t_L     g18785(.A1(new_n7659), .A2(\b[51] ), .B1(new_n7656), .B2(new_n8257), .Y(new_n19042));
  OAI221xp5_ASAP7_75t_L     g18786(.A1(new_n8326), .A2(new_n8228), .B1(new_n7907), .B2(new_n7994), .C(new_n19042), .Y(new_n19043));
  XNOR2x2_ASAP7_75t_L       g18787(.A(new_n7653), .B(new_n19043), .Y(new_n19044));
  XOR2x2_ASAP7_75t_L        g18788(.A(new_n19044), .B(new_n19041), .Y(new_n19045));
  INVx1_ASAP7_75t_L         g18789(.A(new_n19045), .Y(new_n19046));
  O2A1O1Ixp33_ASAP7_75t_L   g18790(.A1(new_n18913), .A2(new_n18919), .B(new_n18915), .C(new_n19046), .Y(new_n19047));
  AND3x1_ASAP7_75t_L        g18791(.A(new_n19046), .B(new_n18922), .C(new_n18915), .Y(new_n19048));
  NOR2xp33_ASAP7_75t_L      g18792(.A(new_n19047), .B(new_n19048), .Y(new_n19049));
  NAND2xp33_ASAP7_75t_L     g18793(.A(new_n18989), .B(new_n19049), .Y(new_n19050));
  OAI21xp33_ASAP7_75t_L     g18794(.A1(new_n19047), .A2(new_n19048), .B(new_n18988), .Y(new_n19051));
  AND2x2_ASAP7_75t_L        g18795(.A(new_n19051), .B(new_n19050), .Y(new_n19052));
  A2O1A1Ixp33_ASAP7_75t_L   g18796(.A1(new_n18928), .A2(new_n18865), .B(new_n18926), .C(new_n19052), .Y(new_n19053));
  OR3x1_ASAP7_75t_L         g18797(.A(new_n18930), .B(new_n18926), .C(new_n19052), .Y(new_n19054));
  NAND2xp33_ASAP7_75t_L     g18798(.A(new_n19053), .B(new_n19054), .Y(new_n19055));
  AOI22xp33_ASAP7_75t_L     g18799(.A1(new_n6002), .A2(\b[57] ), .B1(new_n5999), .B2(new_n10495), .Y(new_n19056));
  OAI221xp5_ASAP7_75t_L     g18800(.A1(new_n6544), .A2(new_n10178), .B1(new_n9534), .B2(new_n6309), .C(new_n19056), .Y(new_n19057));
  XNOR2x2_ASAP7_75t_L       g18801(.A(\a[44] ), .B(new_n19057), .Y(new_n19058));
  XNOR2x2_ASAP7_75t_L       g18802(.A(new_n19058), .B(new_n19055), .Y(new_n19059));
  AND3x1_ASAP7_75t_L        g18803(.A(new_n18939), .B(new_n19059), .C(new_n18936), .Y(new_n19060));
  O2A1O1Ixp33_ASAP7_75t_L   g18804(.A1(new_n18933), .A2(new_n18934), .B(new_n18939), .C(new_n19059), .Y(new_n19061));
  NOR2xp33_ASAP7_75t_L      g18805(.A(new_n19061), .B(new_n19060), .Y(new_n19062));
  AOI22xp33_ASAP7_75t_L     g18806(.A1(new_n5249), .A2(\b[60] ), .B1(new_n5247), .B2(new_n11234), .Y(new_n19063));
  OAI221xp5_ASAP7_75t_L     g18807(.A1(new_n5241), .A2(new_n10881), .B1(new_n10848), .B2(new_n5521), .C(new_n19063), .Y(new_n19064));
  XNOR2x2_ASAP7_75t_L       g18808(.A(\a[41] ), .B(new_n19064), .Y(new_n19065));
  INVx1_ASAP7_75t_L         g18809(.A(new_n19065), .Y(new_n19066));
  XNOR2x2_ASAP7_75t_L       g18810(.A(new_n19066), .B(new_n19062), .Y(new_n19067));
  A2O1A1Ixp33_ASAP7_75t_L   g18811(.A1(new_n18949), .A2(new_n18942), .B(new_n18945), .C(new_n19067), .Y(new_n19068));
  A2O1A1Ixp33_ASAP7_75t_L   g18812(.A1(new_n18939), .A2(new_n18940), .B(new_n18944), .C(new_n18950), .Y(new_n19069));
  NOR2xp33_ASAP7_75t_L      g18813(.A(new_n19067), .B(new_n19069), .Y(new_n19070));
  INVx1_ASAP7_75t_L         g18814(.A(new_n19070), .Y(new_n19071));
  NAND2xp33_ASAP7_75t_L     g18815(.A(new_n19068), .B(new_n19071), .Y(new_n19072));
  NAND2xp33_ASAP7_75t_L     g18816(.A(\b[63] ), .B(new_n4544), .Y(new_n19073));
  A2O1A1Ixp33_ASAP7_75t_L   g18817(.A1(new_n12607), .A2(new_n12603), .B(new_n4549), .C(new_n19073), .Y(new_n19074));
  AOI221xp5_ASAP7_75t_L     g18818(.A1(\b[61] ), .A2(new_n4780), .B1(\b[62] ), .B2(new_n4548), .C(new_n19074), .Y(new_n19075));
  XNOR2x2_ASAP7_75t_L       g18819(.A(new_n4539), .B(new_n19075), .Y(new_n19076));
  XNOR2x2_ASAP7_75t_L       g18820(.A(new_n19076), .B(new_n19072), .Y(new_n19077));
  A2O1A1Ixp33_ASAP7_75t_L   g18821(.A1(new_n18957), .A2(new_n18960), .B(new_n18955), .C(new_n19077), .Y(new_n19078));
  A2O1A1Ixp33_ASAP7_75t_L   g18822(.A1(new_n18825), .A2(new_n18821), .B(new_n18954), .C(new_n18961), .Y(new_n19079));
  NOR2xp33_ASAP7_75t_L      g18823(.A(new_n19077), .B(new_n19079), .Y(new_n19080));
  INVx1_ASAP7_75t_L         g18824(.A(new_n19080), .Y(new_n19081));
  NAND2xp33_ASAP7_75t_L     g18825(.A(new_n19078), .B(new_n19081), .Y(new_n19082));
  AOI211xp5_ASAP7_75t_L     g18826(.A1(new_n18964), .A2(new_n18971), .B(new_n18985), .C(new_n19082), .Y(new_n19083));
  INVx1_ASAP7_75t_L         g18827(.A(new_n19083), .Y(new_n19084));
  A2O1A1Ixp33_ASAP7_75t_L   g18828(.A1(new_n18971), .A2(new_n18964), .B(new_n18985), .C(new_n19082), .Y(new_n19085));
  AND2x2_ASAP7_75t_L        g18829(.A(new_n19085), .B(new_n19084), .Y(new_n19086));
  INVx1_ASAP7_75t_L         g18830(.A(new_n19086), .Y(new_n19087));
  A2O1A1O1Ixp25_ASAP7_75t_L g18831(.A1(new_n18842), .A2(new_n18724), .B(new_n18975), .C(new_n18980), .D(new_n19087), .Y(new_n19088));
  A2O1A1Ixp33_ASAP7_75t_L   g18832(.A1(new_n18842), .A2(new_n18724), .B(new_n18975), .C(new_n18980), .Y(new_n19089));
  NOR2xp33_ASAP7_75t_L      g18833(.A(new_n19086), .B(new_n19089), .Y(new_n19090));
  NOR2xp33_ASAP7_75t_L      g18834(.A(new_n19088), .B(new_n19090), .Y(\f[99] ));
  INVx1_ASAP7_75t_L         g18835(.A(new_n18976), .Y(new_n19092));
  A2O1A1Ixp33_ASAP7_75t_L   g18836(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n4542), .Y(new_n19093));
  AOI22xp33_ASAP7_75t_L     g18837(.A1(new_n4548), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4780), .Y(new_n19094));
  NAND3xp33_ASAP7_75t_L     g18838(.A(new_n19093), .B(\a[38] ), .C(new_n19094), .Y(new_n19095));
  A2O1A1O1Ixp25_ASAP7_75t_L g18839(.A1(new_n13507), .A2(new_n13506), .B(new_n4549), .C(new_n19094), .D(\a[38] ), .Y(new_n19096));
  INVx1_ASAP7_75t_L         g18840(.A(new_n19096), .Y(new_n19097));
  AND2x2_ASAP7_75t_L        g18841(.A(new_n19095), .B(new_n19097), .Y(new_n19098));
  INVx1_ASAP7_75t_L         g18842(.A(new_n19098), .Y(new_n19099));
  A2O1A1Ixp33_ASAP7_75t_L   g18843(.A1(new_n19066), .A2(new_n19062), .B(new_n19070), .C(new_n19099), .Y(new_n19100));
  AOI21xp33_ASAP7_75t_L     g18844(.A1(new_n19066), .A2(new_n19062), .B(new_n19070), .Y(new_n19101));
  NAND2xp33_ASAP7_75t_L     g18845(.A(new_n19098), .B(new_n19101), .Y(new_n19102));
  NAND2xp33_ASAP7_75t_L     g18846(.A(\b[40] ), .B(new_n11656), .Y(new_n19103));
  OAI221xp5_ASAP7_75t_L     g18847(.A1(new_n5166), .A2(new_n12364), .B1(new_n12022), .B2(new_n11823), .C(new_n19103), .Y(new_n19104));
  AOI21xp33_ASAP7_75t_L     g18848(.A1(new_n12021), .A2(\b[38] ), .B(new_n19104), .Y(new_n19105));
  NAND2xp33_ASAP7_75t_L     g18849(.A(\a[62] ), .B(new_n19105), .Y(new_n19106));
  A2O1A1Ixp33_ASAP7_75t_L   g18850(.A1(\b[38] ), .A2(new_n12021), .B(new_n19104), .C(new_n11651), .Y(new_n19107));
  NAND2xp33_ASAP7_75t_L     g18851(.A(new_n19107), .B(new_n19106), .Y(new_n19108));
  NOR2xp33_ASAP7_75t_L      g18852(.A(new_n4465), .B(new_n12671), .Y(new_n19109));
  O2A1O1Ixp33_ASAP7_75t_L   g18853(.A1(new_n12353), .A2(new_n12355), .B(\b[37] ), .C(new_n19109), .Y(new_n19110));
  INVx1_ASAP7_75t_L         g18854(.A(new_n19001), .Y(new_n19111));
  O2A1O1Ixp33_ASAP7_75t_L   g18855(.A1(new_n4053), .A2(new_n12356), .B(new_n18878), .C(\a[35] ), .Y(new_n19112));
  O2A1O1Ixp33_ASAP7_75t_L   g18856(.A1(new_n18997), .A2(new_n18996), .B(new_n19111), .C(new_n19112), .Y(new_n19113));
  NAND2xp33_ASAP7_75t_L     g18857(.A(new_n19110), .B(new_n19113), .Y(new_n19114));
  INVx1_ASAP7_75t_L         g18858(.A(new_n19110), .Y(new_n19115));
  A2O1A1Ixp33_ASAP7_75t_L   g18859(.A1(new_n18999), .A2(new_n19111), .B(new_n19112), .C(new_n19115), .Y(new_n19116));
  AND2x2_ASAP7_75t_L        g18860(.A(new_n19114), .B(new_n19116), .Y(new_n19117));
  XOR2x2_ASAP7_75t_L        g18861(.A(new_n19117), .B(new_n19108), .Y(new_n19118));
  INVx1_ASAP7_75t_L         g18862(.A(new_n19118), .Y(new_n19119));
  O2A1O1Ixp33_ASAP7_75t_L   g18863(.A1(new_n18882), .A2(new_n19007), .B(new_n19003), .C(new_n19015), .Y(new_n19120));
  INVx1_ASAP7_75t_L         g18864(.A(new_n19120), .Y(new_n19121));
  NOR2xp33_ASAP7_75t_L      g18865(.A(new_n19119), .B(new_n19121), .Y(new_n19122));
  O2A1O1Ixp33_ASAP7_75t_L   g18866(.A1(new_n19013), .A2(new_n19010), .B(new_n19006), .C(new_n19118), .Y(new_n19123));
  NOR2xp33_ASAP7_75t_L      g18867(.A(new_n19123), .B(new_n19122), .Y(new_n19124));
  AOI22xp33_ASAP7_75t_L     g18868(.A1(new_n10594), .A2(\b[43] ), .B1(new_n10591), .B2(new_n6202), .Y(new_n19125));
  OAI221xp5_ASAP7_75t_L     g18869(.A1(new_n11335), .A2(new_n5680), .B1(new_n5666), .B2(new_n11330), .C(new_n19125), .Y(new_n19126));
  XNOR2x2_ASAP7_75t_L       g18870(.A(\a[59] ), .B(new_n19126), .Y(new_n19127));
  NAND2xp33_ASAP7_75t_L     g18871(.A(new_n19127), .B(new_n19124), .Y(new_n19128));
  INVx1_ASAP7_75t_L         g18872(.A(new_n19127), .Y(new_n19129));
  OAI21xp33_ASAP7_75t_L     g18873(.A1(new_n19123), .A2(new_n19122), .B(new_n19129), .Y(new_n19130));
  AND2x2_ASAP7_75t_L        g18874(.A(new_n19130), .B(new_n19128), .Y(new_n19131));
  INVx1_ASAP7_75t_L         g18875(.A(new_n19131), .Y(new_n19132));
  INVx1_ASAP7_75t_L         g18876(.A(new_n18891), .Y(new_n19133));
  NAND2xp33_ASAP7_75t_L     g18877(.A(new_n19020), .B(new_n19016), .Y(new_n19134));
  A2O1A1Ixp33_ASAP7_75t_L   g18878(.A1(new_n19133), .A2(new_n18888), .B(new_n19021), .C(new_n19134), .Y(new_n19135));
  NOR2xp33_ASAP7_75t_L      g18879(.A(new_n19135), .B(new_n19132), .Y(new_n19136));
  INVx1_ASAP7_75t_L         g18880(.A(new_n19136), .Y(new_n19137));
  O2A1O1Ixp33_ASAP7_75t_L   g18881(.A1(new_n19024), .A2(new_n19021), .B(new_n19134), .C(new_n19131), .Y(new_n19138));
  INVx1_ASAP7_75t_L         g18882(.A(new_n19138), .Y(new_n19139));
  AOI22xp33_ASAP7_75t_L     g18883(.A1(new_n9623), .A2(\b[46] ), .B1(new_n9620), .B2(new_n7041), .Y(new_n19140));
  OAI221xp5_ASAP7_75t_L     g18884(.A1(new_n10280), .A2(new_n6756), .B1(new_n6220), .B2(new_n12010), .C(new_n19140), .Y(new_n19141));
  XNOR2x2_ASAP7_75t_L       g18885(.A(\a[56] ), .B(new_n19141), .Y(new_n19142));
  NAND3xp33_ASAP7_75t_L     g18886(.A(new_n19137), .B(new_n19139), .C(new_n19142), .Y(new_n19143));
  AO21x2_ASAP7_75t_L        g18887(.A1(new_n19139), .A2(new_n19137), .B(new_n19142), .Y(new_n19144));
  AND2x2_ASAP7_75t_L        g18888(.A(new_n19143), .B(new_n19144), .Y(new_n19145));
  INVx1_ASAP7_75t_L         g18889(.A(new_n19145), .Y(new_n19146));
  NAND2xp33_ASAP7_75t_L     g18890(.A(new_n18993), .B(new_n19026), .Y(new_n19147));
  A2O1A1Ixp33_ASAP7_75t_L   g18891(.A1(new_n18899), .A2(new_n18897), .B(new_n19027), .C(new_n19147), .Y(new_n19148));
  NOR2xp33_ASAP7_75t_L      g18892(.A(new_n19148), .B(new_n19146), .Y(new_n19149));
  INVx1_ASAP7_75t_L         g18893(.A(new_n19149), .Y(new_n19150));
  O2A1O1Ixp33_ASAP7_75t_L   g18894(.A1(new_n19029), .A2(new_n19027), .B(new_n19147), .C(new_n19145), .Y(new_n19151));
  INVx1_ASAP7_75t_L         g18895(.A(new_n19151), .Y(new_n19152));
  AOI22xp33_ASAP7_75t_L     g18896(.A1(new_n8645), .A2(\b[49] ), .B1(new_n8642), .B2(new_n7914), .Y(new_n19153));
  OAI221xp5_ASAP7_75t_L     g18897(.A1(new_n9322), .A2(new_n7333), .B1(new_n7316), .B2(new_n8965), .C(new_n19153), .Y(new_n19154));
  XNOR2x2_ASAP7_75t_L       g18898(.A(\a[53] ), .B(new_n19154), .Y(new_n19155));
  NAND3xp33_ASAP7_75t_L     g18899(.A(new_n19150), .B(new_n19152), .C(new_n19155), .Y(new_n19156));
  AO21x2_ASAP7_75t_L        g18900(.A1(new_n19152), .A2(new_n19150), .B(new_n19155), .Y(new_n19157));
  AND2x2_ASAP7_75t_L        g18901(.A(new_n19156), .B(new_n19157), .Y(new_n19158));
  AOI21xp33_ASAP7_75t_L     g18902(.A1(new_n19036), .A2(new_n19032), .B(new_n19040), .Y(new_n19159));
  NAND2xp33_ASAP7_75t_L     g18903(.A(new_n19159), .B(new_n19158), .Y(new_n19160));
  INVx1_ASAP7_75t_L         g18904(.A(new_n19158), .Y(new_n19161));
  A2O1A1Ixp33_ASAP7_75t_L   g18905(.A1(new_n19036), .A2(new_n19032), .B(new_n19040), .C(new_n19161), .Y(new_n19162));
  AOI22xp33_ASAP7_75t_L     g18906(.A1(new_n7659), .A2(\b[52] ), .B1(new_n7656), .B2(new_n8577), .Y(new_n19163));
  OAI221xp5_ASAP7_75t_L     g18907(.A1(new_n8326), .A2(new_n8249), .B1(new_n8228), .B2(new_n7994), .C(new_n19163), .Y(new_n19164));
  XNOR2x2_ASAP7_75t_L       g18908(.A(\a[50] ), .B(new_n19164), .Y(new_n19165));
  NAND3xp33_ASAP7_75t_L     g18909(.A(new_n19162), .B(new_n19160), .C(new_n19165), .Y(new_n19166));
  AO21x2_ASAP7_75t_L        g18910(.A1(new_n19160), .A2(new_n19162), .B(new_n19165), .Y(new_n19167));
  NAND2xp33_ASAP7_75t_L     g18911(.A(new_n19044), .B(new_n19041), .Y(new_n19168));
  A2O1A1Ixp33_ASAP7_75t_L   g18912(.A1(new_n18915), .A2(new_n18922), .B(new_n19046), .C(new_n19168), .Y(new_n19169));
  AO21x2_ASAP7_75t_L        g18913(.A1(new_n19166), .A2(new_n19167), .B(new_n19169), .Y(new_n19170));
  AND2x2_ASAP7_75t_L        g18914(.A(new_n19166), .B(new_n19167), .Y(new_n19171));
  A2O1A1Ixp33_ASAP7_75t_L   g18915(.A1(new_n19044), .A2(new_n19041), .B(new_n19047), .C(new_n19171), .Y(new_n19172));
  AND2x2_ASAP7_75t_L        g18916(.A(new_n19170), .B(new_n19172), .Y(new_n19173));
  NAND2xp33_ASAP7_75t_L     g18917(.A(new_n6819), .B(new_n9542), .Y(new_n19174));
  OAI221xp5_ASAP7_75t_L     g18918(.A1(new_n7118), .A2(new_n9534), .B1(new_n9199), .B2(new_n7392), .C(new_n19174), .Y(new_n19175));
  AOI21xp33_ASAP7_75t_L     g18919(.A1(new_n7124), .A2(\b[53] ), .B(new_n19175), .Y(new_n19176));
  NAND2xp33_ASAP7_75t_L     g18920(.A(\a[47] ), .B(new_n19176), .Y(new_n19177));
  A2O1A1Ixp33_ASAP7_75t_L   g18921(.A1(\b[53] ), .A2(new_n7124), .B(new_n19175), .C(new_n6816), .Y(new_n19178));
  AND2x2_ASAP7_75t_L        g18922(.A(new_n19178), .B(new_n19177), .Y(new_n19179));
  INVx1_ASAP7_75t_L         g18923(.A(new_n19179), .Y(new_n19180));
  XNOR2x2_ASAP7_75t_L       g18924(.A(new_n19180), .B(new_n19173), .Y(new_n19181));
  INVx1_ASAP7_75t_L         g18925(.A(new_n19181), .Y(new_n19182));
  NAND3xp33_ASAP7_75t_L     g18926(.A(new_n19182), .B(new_n19053), .C(new_n19050), .Y(new_n19183));
  INVx1_ASAP7_75t_L         g18927(.A(new_n19053), .Y(new_n19184));
  A2O1A1Ixp33_ASAP7_75t_L   g18928(.A1(new_n19049), .A2(new_n18989), .B(new_n19184), .C(new_n19181), .Y(new_n19185));
  NAND2xp33_ASAP7_75t_L     g18929(.A(\b[58] ), .B(new_n6002), .Y(new_n19186));
  OAI221xp5_ASAP7_75t_L     g18930(.A1(new_n10488), .A2(new_n6544), .B1(new_n6311), .B2(new_n10856), .C(new_n19186), .Y(new_n19187));
  AOI21xp33_ASAP7_75t_L     g18931(.A1(new_n6308), .A2(\b[56] ), .B(new_n19187), .Y(new_n19188));
  NAND2xp33_ASAP7_75t_L     g18932(.A(\a[44] ), .B(new_n19188), .Y(new_n19189));
  A2O1A1Ixp33_ASAP7_75t_L   g18933(.A1(\b[56] ), .A2(new_n6308), .B(new_n19187), .C(new_n5996), .Y(new_n19190));
  AND2x2_ASAP7_75t_L        g18934(.A(new_n19190), .B(new_n19189), .Y(new_n19191));
  NAND3xp33_ASAP7_75t_L     g18935(.A(new_n19183), .B(new_n19185), .C(new_n19191), .Y(new_n19192));
  AO21x2_ASAP7_75t_L        g18936(.A1(new_n19185), .A2(new_n19183), .B(new_n19191), .Y(new_n19193));
  NAND2xp33_ASAP7_75t_L     g18937(.A(new_n19192), .B(new_n19193), .Y(new_n19194));
  OR2x4_ASAP7_75t_L         g18938(.A(new_n19058), .B(new_n19055), .Y(new_n19195));
  A2O1A1Ixp33_ASAP7_75t_L   g18939(.A1(new_n18939), .A2(new_n18936), .B(new_n19059), .C(new_n19195), .Y(new_n19196));
  NOR2xp33_ASAP7_75t_L      g18940(.A(new_n19196), .B(new_n19194), .Y(new_n19197));
  NAND2xp33_ASAP7_75t_L     g18941(.A(new_n19196), .B(new_n19194), .Y(new_n19198));
  INVx1_ASAP7_75t_L         g18942(.A(new_n19198), .Y(new_n19199));
  NOR2xp33_ASAP7_75t_L      g18943(.A(new_n19197), .B(new_n19199), .Y(new_n19200));
  NAND2xp33_ASAP7_75t_L     g18944(.A(\b[61] ), .B(new_n5249), .Y(new_n19201));
  OAI221xp5_ASAP7_75t_L     g18945(.A1(new_n11226), .A2(new_n5241), .B1(new_n5252), .B2(new_n11920), .C(new_n19201), .Y(new_n19202));
  AOI21xp33_ASAP7_75t_L     g18946(.A1(new_n5526), .A2(\b[59] ), .B(new_n19202), .Y(new_n19203));
  NAND2xp33_ASAP7_75t_L     g18947(.A(\a[41] ), .B(new_n19203), .Y(new_n19204));
  A2O1A1Ixp33_ASAP7_75t_L   g18948(.A1(\b[59] ), .A2(new_n5526), .B(new_n19202), .C(new_n5244), .Y(new_n19205));
  NAND2xp33_ASAP7_75t_L     g18949(.A(new_n19205), .B(new_n19204), .Y(new_n19206));
  NAND2xp33_ASAP7_75t_L     g18950(.A(new_n19206), .B(new_n19200), .Y(new_n19207));
  INVx1_ASAP7_75t_L         g18951(.A(new_n19207), .Y(new_n19208));
  NOR2xp33_ASAP7_75t_L      g18952(.A(new_n19206), .B(new_n19200), .Y(new_n19209));
  NOR2xp33_ASAP7_75t_L      g18953(.A(new_n19209), .B(new_n19208), .Y(new_n19210));
  NAND3xp33_ASAP7_75t_L     g18954(.A(new_n19102), .B(new_n19100), .C(new_n19210), .Y(new_n19211));
  AO21x2_ASAP7_75t_L        g18955(.A1(new_n19100), .A2(new_n19102), .B(new_n19210), .Y(new_n19212));
  AND2x2_ASAP7_75t_L        g18956(.A(new_n19211), .B(new_n19212), .Y(new_n19213));
  INVx1_ASAP7_75t_L         g18957(.A(new_n19213), .Y(new_n19214));
  OA211x2_ASAP7_75t_L       g18958(.A1(new_n19072), .A2(new_n19076), .B(new_n19081), .C(new_n19214), .Y(new_n19215));
  O2A1O1Ixp33_ASAP7_75t_L   g18959(.A1(new_n19072), .A2(new_n19076), .B(new_n19081), .C(new_n19214), .Y(new_n19216));
  NOR2xp33_ASAP7_75t_L      g18960(.A(new_n19216), .B(new_n19215), .Y(new_n19217));
  INVx1_ASAP7_75t_L         g18961(.A(new_n19217), .Y(new_n19218));
  A2O1A1O1Ixp25_ASAP7_75t_L g18962(.A1(new_n19092), .A2(new_n18980), .B(new_n19087), .C(new_n19084), .D(new_n19218), .Y(new_n19219));
  A2O1A1Ixp33_ASAP7_75t_L   g18963(.A1(new_n18980), .A2(new_n19092), .B(new_n19087), .C(new_n19084), .Y(new_n19220));
  NOR2xp33_ASAP7_75t_L      g18964(.A(new_n19217), .B(new_n19220), .Y(new_n19221));
  NOR2xp33_ASAP7_75t_L      g18965(.A(new_n19219), .B(new_n19221), .Y(\f[100] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18966(.A1(new_n19083), .A2(new_n19088), .B(new_n19217), .C(new_n19216), .Y(new_n19223));
  AOI211xp5_ASAP7_75t_L     g18967(.A1(new_n18989), .A2(new_n19049), .B(new_n19184), .C(new_n19181), .Y(new_n19224));
  INVx1_ASAP7_75t_L         g18968(.A(new_n19173), .Y(new_n19225));
  A2O1A1O1Ixp25_ASAP7_75t_L g18969(.A1(new_n18922), .A2(new_n18915), .B(new_n19046), .C(new_n19168), .D(new_n19171), .Y(new_n19226));
  AOI22xp33_ASAP7_75t_L     g18970(.A1(new_n6822), .A2(\b[56] ), .B1(new_n6819), .B2(new_n10185), .Y(new_n19227));
  OAI221xp5_ASAP7_75t_L     g18971(.A1(new_n7392), .A2(new_n9534), .B1(new_n9199), .B2(new_n7115), .C(new_n19227), .Y(new_n19228));
  XNOR2x2_ASAP7_75t_L       g18972(.A(\a[47] ), .B(new_n19228), .Y(new_n19229));
  INVx1_ASAP7_75t_L         g18973(.A(new_n19229), .Y(new_n19230));
  AOI22xp33_ASAP7_75t_L     g18974(.A1(new_n7659), .A2(\b[53] ), .B1(new_n7656), .B2(new_n8889), .Y(new_n19231));
  OAI221xp5_ASAP7_75t_L     g18975(.A1(new_n8326), .A2(new_n8569), .B1(new_n8249), .B2(new_n7994), .C(new_n19231), .Y(new_n19232));
  XNOR2x2_ASAP7_75t_L       g18976(.A(\a[50] ), .B(new_n19232), .Y(new_n19233));
  INVx1_ASAP7_75t_L         g18977(.A(new_n19233), .Y(new_n19234));
  AOI22xp33_ASAP7_75t_L     g18978(.A1(new_n10594), .A2(\b[44] ), .B1(new_n10591), .B2(new_n7055), .Y(new_n19235));
  OAI221xp5_ASAP7_75t_L     g18979(.A1(new_n11335), .A2(new_n6195), .B1(new_n5680), .B2(new_n11330), .C(new_n19235), .Y(new_n19236));
  XNOR2x2_ASAP7_75t_L       g18980(.A(\a[59] ), .B(new_n19236), .Y(new_n19237));
  A2O1A1Ixp33_ASAP7_75t_L   g18981(.A1(new_n18999), .A2(new_n19111), .B(new_n19112), .C(new_n19110), .Y(new_n19238));
  NAND2xp33_ASAP7_75t_L     g18982(.A(\b[37] ), .B(new_n12670), .Y(new_n19239));
  OAI211xp5_ASAP7_75t_L     g18983(.A1(new_n12356), .A2(new_n4915), .B(new_n19110), .C(new_n19239), .Y(new_n19240));
  INVx1_ASAP7_75t_L         g18984(.A(new_n12353), .Y(new_n19241));
  INVx1_ASAP7_75t_L         g18985(.A(new_n12355), .Y(new_n19242));
  A2O1A1Ixp33_ASAP7_75t_L   g18986(.A1(new_n19241), .A2(new_n19242), .B(new_n4915), .C(new_n19239), .Y(new_n19243));
  A2O1A1Ixp33_ASAP7_75t_L   g18987(.A1(new_n12669), .A2(\b[37] ), .B(new_n19109), .C(new_n19243), .Y(new_n19244));
  AND2x2_ASAP7_75t_L        g18988(.A(new_n19244), .B(new_n19240), .Y(new_n19245));
  INVx1_ASAP7_75t_L         g18989(.A(new_n19245), .Y(new_n19246));
  A2O1A1O1Ixp25_ASAP7_75t_L g18990(.A1(new_n19107), .A2(new_n19106), .B(new_n19117), .C(new_n19238), .D(new_n19246), .Y(new_n19247));
  A2O1A1Ixp33_ASAP7_75t_L   g18991(.A1(new_n19106), .A2(new_n19107), .B(new_n19117), .C(new_n19238), .Y(new_n19248));
  NOR2xp33_ASAP7_75t_L      g18992(.A(new_n19245), .B(new_n19248), .Y(new_n19249));
  NOR2xp33_ASAP7_75t_L      g18993(.A(new_n19247), .B(new_n19249), .Y(new_n19250));
  INVx1_ASAP7_75t_L         g18994(.A(new_n19250), .Y(new_n19251));
  AOI22xp33_ASAP7_75t_L     g18995(.A1(new_n11656), .A2(\b[41] ), .B1(new_n11654), .B2(new_n5669), .Y(new_n19252));
  OAI221xp5_ASAP7_75t_L     g18996(.A1(new_n12364), .A2(new_n5186), .B1(new_n5166), .B2(new_n13003), .C(new_n19252), .Y(new_n19253));
  XNOR2x2_ASAP7_75t_L       g18997(.A(\a[62] ), .B(new_n19253), .Y(new_n19254));
  INVx1_ASAP7_75t_L         g18998(.A(new_n19254), .Y(new_n19255));
  NAND2xp33_ASAP7_75t_L     g18999(.A(new_n19255), .B(new_n19251), .Y(new_n19256));
  NAND2xp33_ASAP7_75t_L     g19000(.A(new_n19254), .B(new_n19250), .Y(new_n19257));
  NAND3xp33_ASAP7_75t_L     g19001(.A(new_n19256), .B(new_n19237), .C(new_n19257), .Y(new_n19258));
  AO21x2_ASAP7_75t_L        g19002(.A1(new_n19257), .A2(new_n19256), .B(new_n19237), .Y(new_n19259));
  AND2x2_ASAP7_75t_L        g19003(.A(new_n19258), .B(new_n19259), .Y(new_n19260));
  INVx1_ASAP7_75t_L         g19004(.A(new_n19260), .Y(new_n19261));
  O2A1O1Ixp33_ASAP7_75t_L   g19005(.A1(new_n19119), .A2(new_n19121), .B(new_n19128), .C(new_n19261), .Y(new_n19262));
  INVx1_ASAP7_75t_L         g19006(.A(new_n19262), .Y(new_n19263));
  OAI211xp5_ASAP7_75t_L     g19007(.A1(new_n19119), .A2(new_n19121), .B(new_n19261), .C(new_n19128), .Y(new_n19264));
  AND2x2_ASAP7_75t_L        g19008(.A(new_n19264), .B(new_n19263), .Y(new_n19265));
  AOI22xp33_ASAP7_75t_L     g19009(.A1(new_n9623), .A2(\b[47] ), .B1(new_n9620), .B2(new_n7323), .Y(new_n19266));
  OAI221xp5_ASAP7_75t_L     g19010(.A1(new_n10280), .A2(new_n7033), .B1(new_n6756), .B2(new_n12010), .C(new_n19266), .Y(new_n19267));
  XNOR2x2_ASAP7_75t_L       g19011(.A(\a[56] ), .B(new_n19267), .Y(new_n19268));
  NAND2xp33_ASAP7_75t_L     g19012(.A(new_n19268), .B(new_n19265), .Y(new_n19269));
  AO21x2_ASAP7_75t_L        g19013(.A1(new_n19264), .A2(new_n19263), .B(new_n19268), .Y(new_n19270));
  AND2x2_ASAP7_75t_L        g19014(.A(new_n19270), .B(new_n19269), .Y(new_n19271));
  INVx1_ASAP7_75t_L         g19015(.A(new_n19271), .Y(new_n19272));
  O2A1O1Ixp33_ASAP7_75t_L   g19016(.A1(new_n19132), .A2(new_n19135), .B(new_n19143), .C(new_n19272), .Y(new_n19273));
  INVx1_ASAP7_75t_L         g19017(.A(new_n19273), .Y(new_n19274));
  NAND3xp33_ASAP7_75t_L     g19018(.A(new_n19272), .B(new_n19143), .C(new_n19137), .Y(new_n19275));
  NAND2xp33_ASAP7_75t_L     g19019(.A(new_n19275), .B(new_n19274), .Y(new_n19276));
  AOI22xp33_ASAP7_75t_L     g19020(.A1(new_n8645), .A2(\b[50] ), .B1(new_n8642), .B2(new_n8235), .Y(new_n19277));
  OAI221xp5_ASAP7_75t_L     g19021(.A1(new_n9322), .A2(new_n7907), .B1(new_n7333), .B2(new_n8965), .C(new_n19277), .Y(new_n19278));
  XNOR2x2_ASAP7_75t_L       g19022(.A(\a[53] ), .B(new_n19278), .Y(new_n19279));
  NAND2xp33_ASAP7_75t_L     g19023(.A(new_n19279), .B(new_n19276), .Y(new_n19280));
  INVx1_ASAP7_75t_L         g19024(.A(new_n19279), .Y(new_n19281));
  NAND3xp33_ASAP7_75t_L     g19025(.A(new_n19274), .B(new_n19275), .C(new_n19281), .Y(new_n19282));
  AND2x2_ASAP7_75t_L        g19026(.A(new_n19282), .B(new_n19280), .Y(new_n19283));
  INVx1_ASAP7_75t_L         g19027(.A(new_n19283), .Y(new_n19284));
  NAND2xp33_ASAP7_75t_L     g19028(.A(new_n19150), .B(new_n19156), .Y(new_n19285));
  NOR2xp33_ASAP7_75t_L      g19029(.A(new_n19285), .B(new_n19284), .Y(new_n19286));
  INVx1_ASAP7_75t_L         g19030(.A(new_n19286), .Y(new_n19287));
  O2A1O1Ixp33_ASAP7_75t_L   g19031(.A1(new_n19146), .A2(new_n19148), .B(new_n19156), .C(new_n19283), .Y(new_n19288));
  INVx1_ASAP7_75t_L         g19032(.A(new_n19288), .Y(new_n19289));
  NAND3xp33_ASAP7_75t_L     g19033(.A(new_n19287), .B(new_n19234), .C(new_n19289), .Y(new_n19290));
  OAI21xp33_ASAP7_75t_L     g19034(.A1(new_n19288), .A2(new_n19286), .B(new_n19233), .Y(new_n19291));
  AND2x2_ASAP7_75t_L        g19035(.A(new_n19291), .B(new_n19290), .Y(new_n19292));
  INVx1_ASAP7_75t_L         g19036(.A(new_n19292), .Y(new_n19293));
  NAND2xp33_ASAP7_75t_L     g19037(.A(new_n19160), .B(new_n19166), .Y(new_n19294));
  NOR2xp33_ASAP7_75t_L      g19038(.A(new_n19294), .B(new_n19293), .Y(new_n19295));
  INVx1_ASAP7_75t_L         g19039(.A(new_n19295), .Y(new_n19296));
  INVx1_ASAP7_75t_L         g19040(.A(new_n19160), .Y(new_n19297));
  A2O1A1Ixp33_ASAP7_75t_L   g19041(.A1(new_n19162), .A2(new_n19165), .B(new_n19297), .C(new_n19293), .Y(new_n19298));
  AND2x2_ASAP7_75t_L        g19042(.A(new_n19298), .B(new_n19296), .Y(new_n19299));
  NAND2xp33_ASAP7_75t_L     g19043(.A(new_n19230), .B(new_n19299), .Y(new_n19300));
  AO21x2_ASAP7_75t_L        g19044(.A1(new_n19298), .A2(new_n19296), .B(new_n19230), .Y(new_n19301));
  AND2x2_ASAP7_75t_L        g19045(.A(new_n19301), .B(new_n19300), .Y(new_n19302));
  A2O1A1Ixp33_ASAP7_75t_L   g19046(.A1(new_n19180), .A2(new_n19225), .B(new_n19226), .C(new_n19302), .Y(new_n19303));
  INVx1_ASAP7_75t_L         g19047(.A(new_n19226), .Y(new_n19304));
  A2O1A1Ixp33_ASAP7_75t_L   g19048(.A1(new_n19170), .A2(new_n19172), .B(new_n19179), .C(new_n19304), .Y(new_n19305));
  NOR2xp33_ASAP7_75t_L      g19049(.A(new_n19305), .B(new_n19302), .Y(new_n19306));
  INVx1_ASAP7_75t_L         g19050(.A(new_n19306), .Y(new_n19307));
  AOI22xp33_ASAP7_75t_L     g19051(.A1(new_n6002), .A2(\b[59] ), .B1(new_n5999), .B2(new_n10887), .Y(new_n19308));
  OAI221xp5_ASAP7_75t_L     g19052(.A1(new_n6544), .A2(new_n10848), .B1(new_n10488), .B2(new_n6309), .C(new_n19308), .Y(new_n19309));
  XNOR2x2_ASAP7_75t_L       g19053(.A(\a[44] ), .B(new_n19309), .Y(new_n19310));
  NAND3xp33_ASAP7_75t_L     g19054(.A(new_n19307), .B(new_n19303), .C(new_n19310), .Y(new_n19311));
  AO21x2_ASAP7_75t_L        g19055(.A1(new_n19303), .A2(new_n19307), .B(new_n19310), .Y(new_n19312));
  AND2x2_ASAP7_75t_L        g19056(.A(new_n19311), .B(new_n19312), .Y(new_n19313));
  A2O1A1Ixp33_ASAP7_75t_L   g19057(.A1(new_n19185), .A2(new_n19191), .B(new_n19224), .C(new_n19313), .Y(new_n19314));
  INVx1_ASAP7_75t_L         g19058(.A(new_n19313), .Y(new_n19315));
  NAND3xp33_ASAP7_75t_L     g19059(.A(new_n19315), .B(new_n19192), .C(new_n19183), .Y(new_n19316));
  AOI22xp33_ASAP7_75t_L     g19060(.A1(new_n5249), .A2(\b[62] ), .B1(new_n5247), .B2(new_n12280), .Y(new_n19317));
  OAI221xp5_ASAP7_75t_L     g19061(.A1(new_n5241), .A2(new_n11911), .B1(new_n11226), .B2(new_n5521), .C(new_n19317), .Y(new_n19318));
  XNOR2x2_ASAP7_75t_L       g19062(.A(\a[41] ), .B(new_n19318), .Y(new_n19319));
  NAND3xp33_ASAP7_75t_L     g19063(.A(new_n19316), .B(new_n19314), .C(new_n19319), .Y(new_n19320));
  AO21x2_ASAP7_75t_L        g19064(.A1(new_n19314), .A2(new_n19316), .B(new_n19319), .Y(new_n19321));
  AND2x2_ASAP7_75t_L        g19065(.A(new_n19320), .B(new_n19321), .Y(new_n19322));
  O2A1O1Ixp33_ASAP7_75t_L   g19066(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n4549), .Y(new_n19323));
  O2A1O1Ixp33_ASAP7_75t_L   g19067(.A1(new_n4780), .A2(new_n19323), .B(\b[63] ), .C(new_n4539), .Y(new_n19324));
  A2O1A1O1Ixp25_ASAP7_75t_L g19068(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n4542), .D(new_n4780), .Y(new_n19325));
  NOR3xp33_ASAP7_75t_L      g19069(.A(new_n19325), .B(new_n12599), .C(\a[38] ), .Y(new_n19326));
  NOR2xp33_ASAP7_75t_L      g19070(.A(new_n19324), .B(new_n19326), .Y(new_n19327));
  A2O1A1O1Ixp25_ASAP7_75t_L g19071(.A1(new_n19204), .A2(new_n19205), .B(new_n19197), .C(new_n19198), .D(new_n19327), .Y(new_n19328));
  NAND3xp33_ASAP7_75t_L     g19072(.A(new_n19207), .B(new_n19198), .C(new_n19327), .Y(new_n19329));
  INVx1_ASAP7_75t_L         g19073(.A(new_n19329), .Y(new_n19330));
  NOR2xp33_ASAP7_75t_L      g19074(.A(new_n19328), .B(new_n19330), .Y(new_n19331));
  XNOR2x2_ASAP7_75t_L       g19075(.A(new_n19331), .B(new_n19322), .Y(new_n19332));
  INVx1_ASAP7_75t_L         g19076(.A(new_n19332), .Y(new_n19333));
  O2A1O1Ixp33_ASAP7_75t_L   g19077(.A1(new_n19101), .A2(new_n19098), .B(new_n19211), .C(new_n19333), .Y(new_n19334));
  A2O1A1Ixp33_ASAP7_75t_L   g19078(.A1(new_n19095), .A2(new_n19097), .B(new_n19101), .C(new_n19211), .Y(new_n19335));
  NOR2xp33_ASAP7_75t_L      g19079(.A(new_n19335), .B(new_n19332), .Y(new_n19336));
  NOR2xp33_ASAP7_75t_L      g19080(.A(new_n19336), .B(new_n19334), .Y(new_n19337));
  XNOR2x2_ASAP7_75t_L       g19081(.A(new_n19337), .B(new_n19223), .Y(\f[101] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19082(.A1(new_n19220), .A2(new_n19217), .B(new_n19216), .C(new_n19337), .Y(new_n19339));
  AOI22xp33_ASAP7_75t_L     g19083(.A1(new_n7659), .A2(\b[54] ), .B1(new_n7656), .B2(new_n9208), .Y(new_n19340));
  OAI221xp5_ASAP7_75t_L     g19084(.A1(new_n8326), .A2(new_n8882), .B1(new_n8569), .B2(new_n7994), .C(new_n19340), .Y(new_n19341));
  XNOR2x2_ASAP7_75t_L       g19085(.A(\a[50] ), .B(new_n19341), .Y(new_n19342));
  INVx1_ASAP7_75t_L         g19086(.A(new_n19342), .Y(new_n19343));
  INVx1_ASAP7_75t_L         g19087(.A(new_n19269), .Y(new_n19344));
  AOI22xp33_ASAP7_75t_L     g19088(.A1(new_n9623), .A2(\b[48] ), .B1(new_n9620), .B2(new_n7341), .Y(new_n19345));
  OAI221xp5_ASAP7_75t_L     g19089(.A1(new_n10280), .A2(new_n7316), .B1(new_n7033), .B2(new_n12010), .C(new_n19345), .Y(new_n19346));
  XNOR2x2_ASAP7_75t_L       g19090(.A(new_n9610), .B(new_n19346), .Y(new_n19347));
  O2A1O1Ixp33_ASAP7_75t_L   g19091(.A1(new_n12356), .A2(new_n4915), .B(new_n19239), .C(new_n19115), .Y(new_n19348));
  NOR2xp33_ASAP7_75t_L      g19092(.A(new_n4915), .B(new_n12671), .Y(new_n19349));
  A2O1A1Ixp33_ASAP7_75t_L   g19093(.A1(new_n12669), .A2(\b[37] ), .B(new_n19109), .C(\a[38] ), .Y(new_n19350));
  NOR2xp33_ASAP7_75t_L      g19094(.A(\a[38] ), .B(new_n19115), .Y(new_n19351));
  INVx1_ASAP7_75t_L         g19095(.A(new_n19351), .Y(new_n19352));
  NAND2xp33_ASAP7_75t_L     g19096(.A(new_n19350), .B(new_n19352), .Y(new_n19353));
  A2O1A1Ixp33_ASAP7_75t_L   g19097(.A1(new_n12669), .A2(\b[39] ), .B(new_n19349), .C(new_n19353), .Y(new_n19354));
  INVx1_ASAP7_75t_L         g19098(.A(new_n19354), .Y(new_n19355));
  O2A1O1Ixp33_ASAP7_75t_L   g19099(.A1(new_n12353), .A2(new_n12355), .B(\b[39] ), .C(new_n19349), .Y(new_n19356));
  AND3x1_ASAP7_75t_L        g19100(.A(new_n19352), .B(new_n19350), .C(new_n19356), .Y(new_n19357));
  NOR2xp33_ASAP7_75t_L      g19101(.A(new_n19357), .B(new_n19355), .Y(new_n19358));
  A2O1A1Ixp33_ASAP7_75t_L   g19102(.A1(new_n19248), .A2(new_n19246), .B(new_n19348), .C(new_n19358), .Y(new_n19359));
  A2O1A1O1Ixp25_ASAP7_75t_L g19103(.A1(new_n19107), .A2(new_n19106), .B(new_n19117), .C(new_n19238), .D(new_n19245), .Y(new_n19360));
  OR3x1_ASAP7_75t_L         g19104(.A(new_n19360), .B(new_n19348), .C(new_n19358), .Y(new_n19361));
  NAND2xp33_ASAP7_75t_L     g19105(.A(\b[41] ), .B(new_n11647), .Y(new_n19362));
  OAI221xp5_ASAP7_75t_L     g19106(.A1(new_n12023), .A2(new_n5680), .B1(new_n12022), .B2(new_n5687), .C(new_n19362), .Y(new_n19363));
  AOI21xp33_ASAP7_75t_L     g19107(.A1(new_n12021), .A2(\b[40] ), .B(new_n19363), .Y(new_n19364));
  NAND2xp33_ASAP7_75t_L     g19108(.A(\a[62] ), .B(new_n19364), .Y(new_n19365));
  A2O1A1Ixp33_ASAP7_75t_L   g19109(.A1(\b[40] ), .A2(new_n12021), .B(new_n19363), .C(new_n11651), .Y(new_n19366));
  NAND4xp25_ASAP7_75t_L     g19110(.A(new_n19361), .B(new_n19365), .C(new_n19366), .D(new_n19359), .Y(new_n19367));
  AO22x1_ASAP7_75t_L        g19111(.A1(new_n19366), .A2(new_n19365), .B1(new_n19359), .B2(new_n19361), .Y(new_n19368));
  NAND2xp33_ASAP7_75t_L     g19112(.A(new_n19367), .B(new_n19368), .Y(new_n19369));
  AOI22xp33_ASAP7_75t_L     g19113(.A1(new_n10594), .A2(\b[45] ), .B1(new_n10591), .B2(new_n6764), .Y(new_n19370));
  OAI221xp5_ASAP7_75t_L     g19114(.A1(new_n11335), .A2(new_n6220), .B1(new_n6195), .B2(new_n11330), .C(new_n19370), .Y(new_n19371));
  XNOR2x2_ASAP7_75t_L       g19115(.A(\a[59] ), .B(new_n19371), .Y(new_n19372));
  INVx1_ASAP7_75t_L         g19116(.A(new_n19372), .Y(new_n19373));
  NAND2xp33_ASAP7_75t_L     g19117(.A(new_n19369), .B(new_n19373), .Y(new_n19374));
  NAND3xp33_ASAP7_75t_L     g19118(.A(new_n19372), .B(new_n19368), .C(new_n19367), .Y(new_n19375));
  AND2x2_ASAP7_75t_L        g19119(.A(new_n19375), .B(new_n19374), .Y(new_n19376));
  INVx1_ASAP7_75t_L         g19120(.A(new_n19376), .Y(new_n19377));
  NAND2xp33_ASAP7_75t_L     g19121(.A(new_n19257), .B(new_n19258), .Y(new_n19378));
  NOR2xp33_ASAP7_75t_L      g19122(.A(new_n19378), .B(new_n19377), .Y(new_n19379));
  O2A1O1Ixp33_ASAP7_75t_L   g19123(.A1(new_n19251), .A2(new_n19255), .B(new_n19258), .C(new_n19376), .Y(new_n19380));
  NOR2xp33_ASAP7_75t_L      g19124(.A(new_n19380), .B(new_n19379), .Y(new_n19381));
  XNOR2x2_ASAP7_75t_L       g19125(.A(new_n19347), .B(new_n19381), .Y(new_n19382));
  OA21x2_ASAP7_75t_L        g19126(.A1(new_n19262), .A2(new_n19344), .B(new_n19382), .Y(new_n19383));
  NOR3xp33_ASAP7_75t_L      g19127(.A(new_n19344), .B(new_n19382), .C(new_n19262), .Y(new_n19384));
  NOR2xp33_ASAP7_75t_L      g19128(.A(new_n19384), .B(new_n19383), .Y(new_n19385));
  AOI22xp33_ASAP7_75t_L     g19129(.A1(new_n8645), .A2(\b[51] ), .B1(new_n8642), .B2(new_n8257), .Y(new_n19386));
  OAI221xp5_ASAP7_75t_L     g19130(.A1(new_n9322), .A2(new_n8228), .B1(new_n7907), .B2(new_n8965), .C(new_n19386), .Y(new_n19387));
  XNOR2x2_ASAP7_75t_L       g19131(.A(new_n8639), .B(new_n19387), .Y(new_n19388));
  XOR2x2_ASAP7_75t_L        g19132(.A(new_n19388), .B(new_n19385), .Y(new_n19389));
  INVx1_ASAP7_75t_L         g19133(.A(new_n19389), .Y(new_n19390));
  O2A1O1Ixp33_ASAP7_75t_L   g19134(.A1(new_n19273), .A2(new_n19279), .B(new_n19275), .C(new_n19390), .Y(new_n19391));
  AND3x1_ASAP7_75t_L        g19135(.A(new_n19390), .B(new_n19282), .C(new_n19275), .Y(new_n19392));
  NOR2xp33_ASAP7_75t_L      g19136(.A(new_n19391), .B(new_n19392), .Y(new_n19393));
  NAND2xp33_ASAP7_75t_L     g19137(.A(new_n19343), .B(new_n19393), .Y(new_n19394));
  OAI21xp33_ASAP7_75t_L     g19138(.A1(new_n19391), .A2(new_n19392), .B(new_n19342), .Y(new_n19395));
  AND2x2_ASAP7_75t_L        g19139(.A(new_n19395), .B(new_n19394), .Y(new_n19396));
  INVx1_ASAP7_75t_L         g19140(.A(new_n19396), .Y(new_n19397));
  O2A1O1Ixp33_ASAP7_75t_L   g19141(.A1(new_n19284), .A2(new_n19285), .B(new_n19290), .C(new_n19397), .Y(new_n19398));
  INVx1_ASAP7_75t_L         g19142(.A(new_n19398), .Y(new_n19399));
  NAND3xp33_ASAP7_75t_L     g19143(.A(new_n19397), .B(new_n19290), .C(new_n19287), .Y(new_n19400));
  NAND2xp33_ASAP7_75t_L     g19144(.A(new_n19400), .B(new_n19399), .Y(new_n19401));
  AOI22xp33_ASAP7_75t_L     g19145(.A1(new_n6822), .A2(\b[57] ), .B1(new_n6819), .B2(new_n10495), .Y(new_n19402));
  OAI221xp5_ASAP7_75t_L     g19146(.A1(new_n7392), .A2(new_n10178), .B1(new_n9534), .B2(new_n7115), .C(new_n19402), .Y(new_n19403));
  XNOR2x2_ASAP7_75t_L       g19147(.A(\a[47] ), .B(new_n19403), .Y(new_n19404));
  XNOR2x2_ASAP7_75t_L       g19148(.A(new_n19404), .B(new_n19401), .Y(new_n19405));
  INVx1_ASAP7_75t_L         g19149(.A(new_n19405), .Y(new_n19406));
  NAND2xp33_ASAP7_75t_L     g19150(.A(new_n19296), .B(new_n19300), .Y(new_n19407));
  NOR2xp33_ASAP7_75t_L      g19151(.A(new_n19406), .B(new_n19407), .Y(new_n19408));
  O2A1O1Ixp33_ASAP7_75t_L   g19152(.A1(new_n19293), .A2(new_n19294), .B(new_n19300), .C(new_n19405), .Y(new_n19409));
  NOR2xp33_ASAP7_75t_L      g19153(.A(new_n19409), .B(new_n19408), .Y(new_n19410));
  AOI22xp33_ASAP7_75t_L     g19154(.A1(new_n6002), .A2(\b[60] ), .B1(new_n5999), .B2(new_n11234), .Y(new_n19411));
  OAI221xp5_ASAP7_75t_L     g19155(.A1(new_n6544), .A2(new_n10881), .B1(new_n10848), .B2(new_n6309), .C(new_n19411), .Y(new_n19412));
  XNOR2x2_ASAP7_75t_L       g19156(.A(\a[44] ), .B(new_n19412), .Y(new_n19413));
  INVx1_ASAP7_75t_L         g19157(.A(new_n19413), .Y(new_n19414));
  XNOR2x2_ASAP7_75t_L       g19158(.A(new_n19414), .B(new_n19410), .Y(new_n19415));
  A2O1A1Ixp33_ASAP7_75t_L   g19159(.A1(new_n19310), .A2(new_n19303), .B(new_n19306), .C(new_n19415), .Y(new_n19416));
  A2O1A1Ixp33_ASAP7_75t_L   g19160(.A1(new_n19300), .A2(new_n19301), .B(new_n19305), .C(new_n19311), .Y(new_n19417));
  NOR2xp33_ASAP7_75t_L      g19161(.A(new_n19415), .B(new_n19417), .Y(new_n19418));
  INVx1_ASAP7_75t_L         g19162(.A(new_n19418), .Y(new_n19419));
  NAND2xp33_ASAP7_75t_L     g19163(.A(new_n19416), .B(new_n19419), .Y(new_n19420));
  NAND2xp33_ASAP7_75t_L     g19164(.A(\b[63] ), .B(new_n5249), .Y(new_n19421));
  A2O1A1Ixp33_ASAP7_75t_L   g19165(.A1(new_n12607), .A2(new_n12603), .B(new_n5252), .C(new_n19421), .Y(new_n19422));
  AOI221xp5_ASAP7_75t_L     g19166(.A1(\b[61] ), .A2(new_n5526), .B1(\b[62] ), .B2(new_n5240), .C(new_n19422), .Y(new_n19423));
  XNOR2x2_ASAP7_75t_L       g19167(.A(new_n5244), .B(new_n19423), .Y(new_n19424));
  XNOR2x2_ASAP7_75t_L       g19168(.A(new_n19424), .B(new_n19420), .Y(new_n19425));
  INVx1_ASAP7_75t_L         g19169(.A(new_n19425), .Y(new_n19426));
  A2O1A1O1Ixp25_ASAP7_75t_L g19170(.A1(new_n19192), .A2(new_n19183), .B(new_n19315), .C(new_n19320), .D(new_n19426), .Y(new_n19427));
  A2O1A1Ixp33_ASAP7_75t_L   g19171(.A1(new_n19192), .A2(new_n19183), .B(new_n19315), .C(new_n19320), .Y(new_n19428));
  NOR2xp33_ASAP7_75t_L      g19172(.A(new_n19428), .B(new_n19425), .Y(new_n19429));
  NOR2xp33_ASAP7_75t_L      g19173(.A(new_n19429), .B(new_n19427), .Y(new_n19430));
  A2O1A1Ixp33_ASAP7_75t_L   g19174(.A1(new_n19198), .A2(new_n19207), .B(new_n19327), .C(new_n19322), .Y(new_n19431));
  AND3x1_ASAP7_75t_L        g19175(.A(new_n19430), .B(new_n19431), .C(new_n19329), .Y(new_n19432));
  INVx1_ASAP7_75t_L         g19176(.A(new_n19432), .Y(new_n19433));
  INVx1_ASAP7_75t_L         g19177(.A(new_n19328), .Y(new_n19434));
  INVx1_ASAP7_75t_L         g19178(.A(new_n19430), .Y(new_n19435));
  A2O1A1Ixp33_ASAP7_75t_L   g19179(.A1(new_n19434), .A2(new_n19322), .B(new_n19330), .C(new_n19435), .Y(new_n19436));
  AND2x2_ASAP7_75t_L        g19180(.A(new_n19436), .B(new_n19433), .Y(new_n19437));
  INVx1_ASAP7_75t_L         g19181(.A(new_n19437), .Y(new_n19438));
  A2O1A1O1Ixp25_ASAP7_75t_L g19182(.A1(new_n19211), .A2(new_n19100), .B(new_n19333), .C(new_n19339), .D(new_n19438), .Y(new_n19439));
  A2O1A1Ixp33_ASAP7_75t_L   g19183(.A1(new_n19211), .A2(new_n19100), .B(new_n19333), .C(new_n19339), .Y(new_n19440));
  NOR2xp33_ASAP7_75t_L      g19184(.A(new_n19437), .B(new_n19440), .Y(new_n19441));
  NOR2xp33_ASAP7_75t_L      g19185(.A(new_n19439), .B(new_n19441), .Y(\f[102] ));
  INVx1_ASAP7_75t_L         g19186(.A(new_n19334), .Y(new_n19443));
  NOR2xp33_ASAP7_75t_L      g19187(.A(new_n19424), .B(new_n19420), .Y(new_n19444));
  A2O1A1Ixp33_ASAP7_75t_L   g19188(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n5247), .Y(new_n19445));
  AOI22xp33_ASAP7_75t_L     g19189(.A1(new_n5240), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5526), .Y(new_n19446));
  NAND3xp33_ASAP7_75t_L     g19190(.A(new_n19445), .B(\a[41] ), .C(new_n19446), .Y(new_n19447));
  A2O1A1O1Ixp25_ASAP7_75t_L g19191(.A1(new_n13507), .A2(new_n13506), .B(new_n5252), .C(new_n19446), .D(\a[41] ), .Y(new_n19448));
  INVx1_ASAP7_75t_L         g19192(.A(new_n19448), .Y(new_n19449));
  AND2x2_ASAP7_75t_L        g19193(.A(new_n19447), .B(new_n19449), .Y(new_n19450));
  INVx1_ASAP7_75t_L         g19194(.A(new_n19450), .Y(new_n19451));
  A2O1A1Ixp33_ASAP7_75t_L   g19195(.A1(new_n19414), .A2(new_n19410), .B(new_n19418), .C(new_n19451), .Y(new_n19452));
  AOI21xp33_ASAP7_75t_L     g19196(.A1(new_n19414), .A2(new_n19410), .B(new_n19418), .Y(new_n19453));
  NAND2xp33_ASAP7_75t_L     g19197(.A(new_n19450), .B(new_n19453), .Y(new_n19454));
  A2O1A1Ixp33_ASAP7_75t_L   g19198(.A1(new_n19287), .A2(new_n19290), .B(new_n19397), .C(new_n19394), .Y(new_n19455));
  INVx1_ASAP7_75t_L         g19199(.A(new_n19379), .Y(new_n19456));
  NOR2xp33_ASAP7_75t_L      g19200(.A(new_n5166), .B(new_n12671), .Y(new_n19457));
  O2A1O1Ixp33_ASAP7_75t_L   g19201(.A1(new_n12353), .A2(new_n12355), .B(\b[40] ), .C(new_n19457), .Y(new_n19458));
  INVx1_ASAP7_75t_L         g19202(.A(new_n19458), .Y(new_n19459));
  A2O1A1Ixp33_ASAP7_75t_L   g19203(.A1(new_n12669), .A2(\b[37] ), .B(new_n19109), .C(new_n4539), .Y(new_n19460));
  A2O1A1O1Ixp25_ASAP7_75t_L g19204(.A1(new_n19350), .A2(new_n19352), .B(new_n19356), .C(new_n19460), .D(new_n19459), .Y(new_n19461));
  INVx1_ASAP7_75t_L         g19205(.A(new_n19461), .Y(new_n19462));
  A2O1A1O1Ixp25_ASAP7_75t_L g19206(.A1(new_n12669), .A2(\b[37] ), .B(new_n19109), .C(new_n4539), .D(new_n19355), .Y(new_n19463));
  A2O1A1Ixp33_ASAP7_75t_L   g19207(.A1(new_n12669), .A2(\b[40] ), .B(new_n19457), .C(new_n19463), .Y(new_n19464));
  AOI22xp33_ASAP7_75t_L     g19208(.A1(new_n11647), .A2(\b[42] ), .B1(\b[43] ), .B2(new_n11656), .Y(new_n19465));
  OAI221xp5_ASAP7_75t_L     g19209(.A1(new_n13003), .A2(new_n5666), .B1(new_n12022), .B2(new_n9799), .C(new_n19465), .Y(new_n19466));
  XNOR2x2_ASAP7_75t_L       g19210(.A(new_n11651), .B(new_n19466), .Y(new_n19467));
  NAND3xp33_ASAP7_75t_L     g19211(.A(new_n19467), .B(new_n19464), .C(new_n19462), .Y(new_n19468));
  AO21x2_ASAP7_75t_L        g19212(.A1(new_n19462), .A2(new_n19464), .B(new_n19467), .Y(new_n19469));
  AND2x2_ASAP7_75t_L        g19213(.A(new_n19468), .B(new_n19469), .Y(new_n19470));
  NAND3xp33_ASAP7_75t_L     g19214(.A(new_n19470), .B(new_n19367), .C(new_n19361), .Y(new_n19471));
  AO21x2_ASAP7_75t_L        g19215(.A1(new_n19361), .A2(new_n19367), .B(new_n19470), .Y(new_n19472));
  AOI22xp33_ASAP7_75t_L     g19216(.A1(new_n10594), .A2(\b[46] ), .B1(new_n10591), .B2(new_n7041), .Y(new_n19473));
  OAI221xp5_ASAP7_75t_L     g19217(.A1(new_n11335), .A2(new_n6756), .B1(new_n6220), .B2(new_n11330), .C(new_n19473), .Y(new_n19474));
  XNOR2x2_ASAP7_75t_L       g19218(.A(\a[59] ), .B(new_n19474), .Y(new_n19475));
  NAND3xp33_ASAP7_75t_L     g19219(.A(new_n19472), .B(new_n19471), .C(new_n19475), .Y(new_n19476));
  AO21x2_ASAP7_75t_L        g19220(.A1(new_n19471), .A2(new_n19472), .B(new_n19475), .Y(new_n19477));
  AND2x2_ASAP7_75t_L        g19221(.A(new_n19476), .B(new_n19477), .Y(new_n19478));
  NAND3xp33_ASAP7_75t_L     g19222(.A(new_n19456), .B(new_n19374), .C(new_n19478), .Y(new_n19479));
  INVx1_ASAP7_75t_L         g19223(.A(new_n19478), .Y(new_n19480));
  A2O1A1Ixp33_ASAP7_75t_L   g19224(.A1(new_n19373), .A2(new_n19369), .B(new_n19379), .C(new_n19480), .Y(new_n19481));
  NAND2xp33_ASAP7_75t_L     g19225(.A(new_n9620), .B(new_n7914), .Y(new_n19482));
  OAI221xp5_ASAP7_75t_L     g19226(.A1(new_n9950), .A2(new_n7907), .B1(new_n7333), .B2(new_n10280), .C(new_n19482), .Y(new_n19483));
  AOI21xp33_ASAP7_75t_L     g19227(.A1(new_n9948), .A2(\b[47] ), .B(new_n19483), .Y(new_n19484));
  NAND2xp33_ASAP7_75t_L     g19228(.A(\a[56] ), .B(new_n19484), .Y(new_n19485));
  A2O1A1Ixp33_ASAP7_75t_L   g19229(.A1(\b[47] ), .A2(new_n9948), .B(new_n19483), .C(new_n9610), .Y(new_n19486));
  AND2x2_ASAP7_75t_L        g19230(.A(new_n19486), .B(new_n19485), .Y(new_n19487));
  NAND3xp33_ASAP7_75t_L     g19231(.A(new_n19479), .B(new_n19481), .C(new_n19487), .Y(new_n19488));
  AO21x2_ASAP7_75t_L        g19232(.A1(new_n19481), .A2(new_n19479), .B(new_n19487), .Y(new_n19489));
  AND2x2_ASAP7_75t_L        g19233(.A(new_n19488), .B(new_n19489), .Y(new_n19490));
  AOI21xp33_ASAP7_75t_L     g19234(.A1(new_n19381), .A2(new_n19347), .B(new_n19384), .Y(new_n19491));
  NAND2xp33_ASAP7_75t_L     g19235(.A(new_n19490), .B(new_n19491), .Y(new_n19492));
  INVx1_ASAP7_75t_L         g19236(.A(new_n19490), .Y(new_n19493));
  A2O1A1Ixp33_ASAP7_75t_L   g19237(.A1(new_n19381), .A2(new_n19347), .B(new_n19384), .C(new_n19493), .Y(new_n19494));
  NAND2xp33_ASAP7_75t_L     g19238(.A(new_n19494), .B(new_n19492), .Y(new_n19495));
  AOI22xp33_ASAP7_75t_L     g19239(.A1(new_n8645), .A2(\b[52] ), .B1(new_n8642), .B2(new_n8577), .Y(new_n19496));
  OAI221xp5_ASAP7_75t_L     g19240(.A1(new_n9322), .A2(new_n8249), .B1(new_n8228), .B2(new_n8965), .C(new_n19496), .Y(new_n19497));
  XNOR2x2_ASAP7_75t_L       g19241(.A(\a[53] ), .B(new_n19497), .Y(new_n19498));
  INVx1_ASAP7_75t_L         g19242(.A(new_n19498), .Y(new_n19499));
  NOR2xp33_ASAP7_75t_L      g19243(.A(new_n19499), .B(new_n19495), .Y(new_n19500));
  INVx1_ASAP7_75t_L         g19244(.A(new_n19500), .Y(new_n19501));
  NAND2xp33_ASAP7_75t_L     g19245(.A(new_n19499), .B(new_n19495), .Y(new_n19502));
  NAND2xp33_ASAP7_75t_L     g19246(.A(new_n19388), .B(new_n19385), .Y(new_n19503));
  A2O1A1Ixp33_ASAP7_75t_L   g19247(.A1(new_n19275), .A2(new_n19282), .B(new_n19390), .C(new_n19503), .Y(new_n19504));
  AO21x2_ASAP7_75t_L        g19248(.A1(new_n19501), .A2(new_n19502), .B(new_n19504), .Y(new_n19505));
  AND2x2_ASAP7_75t_L        g19249(.A(new_n19502), .B(new_n19501), .Y(new_n19506));
  A2O1A1Ixp33_ASAP7_75t_L   g19250(.A1(new_n19388), .A2(new_n19385), .B(new_n19391), .C(new_n19506), .Y(new_n19507));
  AND2x2_ASAP7_75t_L        g19251(.A(new_n19505), .B(new_n19507), .Y(new_n19508));
  NAND2xp33_ASAP7_75t_L     g19252(.A(new_n7656), .B(new_n9542), .Y(new_n19509));
  OAI221xp5_ASAP7_75t_L     g19253(.A1(new_n7997), .A2(new_n9534), .B1(new_n9199), .B2(new_n8326), .C(new_n19509), .Y(new_n19510));
  AOI21xp33_ASAP7_75t_L     g19254(.A1(new_n7993), .A2(\b[53] ), .B(new_n19510), .Y(new_n19511));
  NAND2xp33_ASAP7_75t_L     g19255(.A(\a[50] ), .B(new_n19511), .Y(new_n19512));
  A2O1A1Ixp33_ASAP7_75t_L   g19256(.A1(\b[53] ), .A2(new_n7993), .B(new_n19510), .C(new_n7653), .Y(new_n19513));
  AND2x2_ASAP7_75t_L        g19257(.A(new_n19513), .B(new_n19512), .Y(new_n19514));
  INVx1_ASAP7_75t_L         g19258(.A(new_n19514), .Y(new_n19515));
  XNOR2x2_ASAP7_75t_L       g19259(.A(new_n19515), .B(new_n19508), .Y(new_n19516));
  OR2x4_ASAP7_75t_L         g19260(.A(new_n19516), .B(new_n19455), .Y(new_n19517));
  A2O1A1Ixp33_ASAP7_75t_L   g19261(.A1(new_n19393), .A2(new_n19343), .B(new_n19398), .C(new_n19516), .Y(new_n19518));
  NAND2xp33_ASAP7_75t_L     g19262(.A(\b[58] ), .B(new_n6822), .Y(new_n19519));
  OAI221xp5_ASAP7_75t_L     g19263(.A1(new_n10488), .A2(new_n7392), .B1(new_n7117), .B2(new_n10856), .C(new_n19519), .Y(new_n19520));
  AOI21xp33_ASAP7_75t_L     g19264(.A1(new_n7124), .A2(\b[56] ), .B(new_n19520), .Y(new_n19521));
  NAND2xp33_ASAP7_75t_L     g19265(.A(\a[47] ), .B(new_n19521), .Y(new_n19522));
  A2O1A1Ixp33_ASAP7_75t_L   g19266(.A1(\b[56] ), .A2(new_n7124), .B(new_n19520), .C(new_n6816), .Y(new_n19523));
  AND2x2_ASAP7_75t_L        g19267(.A(new_n19523), .B(new_n19522), .Y(new_n19524));
  NAND3xp33_ASAP7_75t_L     g19268(.A(new_n19517), .B(new_n19518), .C(new_n19524), .Y(new_n19525));
  AO21x2_ASAP7_75t_L        g19269(.A1(new_n19518), .A2(new_n19517), .B(new_n19524), .Y(new_n19526));
  NAND2xp33_ASAP7_75t_L     g19270(.A(new_n19525), .B(new_n19526), .Y(new_n19527));
  NOR2xp33_ASAP7_75t_L      g19271(.A(new_n19404), .B(new_n19401), .Y(new_n19528));
  A2O1A1O1Ixp25_ASAP7_75t_L g19272(.A1(new_n19230), .A2(new_n19299), .B(new_n19295), .C(new_n19406), .D(new_n19528), .Y(new_n19529));
  XNOR2x2_ASAP7_75t_L       g19273(.A(new_n19527), .B(new_n19529), .Y(new_n19530));
  NAND2xp33_ASAP7_75t_L     g19274(.A(\b[61] ), .B(new_n6002), .Y(new_n19531));
  OAI221xp5_ASAP7_75t_L     g19275(.A1(new_n11226), .A2(new_n6544), .B1(new_n6311), .B2(new_n11920), .C(new_n19531), .Y(new_n19532));
  AOI21xp33_ASAP7_75t_L     g19276(.A1(new_n6308), .A2(\b[59] ), .B(new_n19532), .Y(new_n19533));
  NAND2xp33_ASAP7_75t_L     g19277(.A(\a[44] ), .B(new_n19533), .Y(new_n19534));
  A2O1A1Ixp33_ASAP7_75t_L   g19278(.A1(\b[59] ), .A2(new_n6308), .B(new_n19532), .C(new_n5996), .Y(new_n19535));
  NAND2xp33_ASAP7_75t_L     g19279(.A(new_n19535), .B(new_n19534), .Y(new_n19536));
  NAND2xp33_ASAP7_75t_L     g19280(.A(new_n19536), .B(new_n19530), .Y(new_n19537));
  INVx1_ASAP7_75t_L         g19281(.A(new_n19537), .Y(new_n19538));
  NOR2xp33_ASAP7_75t_L      g19282(.A(new_n19536), .B(new_n19530), .Y(new_n19539));
  NOR2xp33_ASAP7_75t_L      g19283(.A(new_n19539), .B(new_n19538), .Y(new_n19540));
  NAND3xp33_ASAP7_75t_L     g19284(.A(new_n19454), .B(new_n19452), .C(new_n19540), .Y(new_n19541));
  AO21x2_ASAP7_75t_L        g19285(.A1(new_n19452), .A2(new_n19454), .B(new_n19540), .Y(new_n19542));
  AND2x2_ASAP7_75t_L        g19286(.A(new_n19541), .B(new_n19542), .Y(new_n19543));
  NOR3xp33_ASAP7_75t_L      g19287(.A(new_n19543), .B(new_n19429), .C(new_n19444), .Y(new_n19544));
  OA21x2_ASAP7_75t_L        g19288(.A1(new_n19444), .A2(new_n19429), .B(new_n19543), .Y(new_n19545));
  NOR2xp33_ASAP7_75t_L      g19289(.A(new_n19544), .B(new_n19545), .Y(new_n19546));
  INVx1_ASAP7_75t_L         g19290(.A(new_n19546), .Y(new_n19547));
  A2O1A1O1Ixp25_ASAP7_75t_L g19291(.A1(new_n19443), .A2(new_n19339), .B(new_n19438), .C(new_n19433), .D(new_n19547), .Y(new_n19548));
  A2O1A1Ixp33_ASAP7_75t_L   g19292(.A1(new_n19339), .A2(new_n19443), .B(new_n19438), .C(new_n19433), .Y(new_n19549));
  NOR2xp33_ASAP7_75t_L      g19293(.A(new_n19546), .B(new_n19549), .Y(new_n19550));
  NOR2xp33_ASAP7_75t_L      g19294(.A(new_n19548), .B(new_n19550), .Y(\f[103] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19295(.A1(new_n19432), .A2(new_n19439), .B(new_n19546), .C(new_n19545), .Y(new_n19552));
  INVx1_ASAP7_75t_L         g19296(.A(new_n19508), .Y(new_n19553));
  A2O1A1O1Ixp25_ASAP7_75t_L g19297(.A1(new_n19282), .A2(new_n19275), .B(new_n19390), .C(new_n19503), .D(new_n19506), .Y(new_n19554));
  AOI22xp33_ASAP7_75t_L     g19298(.A1(new_n7659), .A2(\b[56] ), .B1(new_n7656), .B2(new_n10185), .Y(new_n19555));
  OAI221xp5_ASAP7_75t_L     g19299(.A1(new_n8326), .A2(new_n9534), .B1(new_n9199), .B2(new_n7994), .C(new_n19555), .Y(new_n19556));
  XNOR2x2_ASAP7_75t_L       g19300(.A(\a[50] ), .B(new_n19556), .Y(new_n19557));
  INVx1_ASAP7_75t_L         g19301(.A(new_n19557), .Y(new_n19558));
  AOI22xp33_ASAP7_75t_L     g19302(.A1(new_n8645), .A2(\b[53] ), .B1(new_n8642), .B2(new_n8889), .Y(new_n19559));
  OAI221xp5_ASAP7_75t_L     g19303(.A1(new_n9322), .A2(new_n8569), .B1(new_n8249), .B2(new_n8965), .C(new_n19559), .Y(new_n19560));
  XNOR2x2_ASAP7_75t_L       g19304(.A(\a[53] ), .B(new_n19560), .Y(new_n19561));
  AOI22xp33_ASAP7_75t_L     g19305(.A1(new_n10594), .A2(\b[47] ), .B1(new_n10591), .B2(new_n7323), .Y(new_n19562));
  OAI221xp5_ASAP7_75t_L     g19306(.A1(new_n11335), .A2(new_n7033), .B1(new_n6756), .B2(new_n11330), .C(new_n19562), .Y(new_n19563));
  XNOR2x2_ASAP7_75t_L       g19307(.A(\a[59] ), .B(new_n19563), .Y(new_n19564));
  INVx1_ASAP7_75t_L         g19308(.A(new_n19564), .Y(new_n19565));
  NAND2xp33_ASAP7_75t_L     g19309(.A(\b[40] ), .B(new_n12670), .Y(new_n19566));
  OAI211xp5_ASAP7_75t_L     g19310(.A1(new_n12356), .A2(new_n5666), .B(new_n19458), .C(new_n19566), .Y(new_n19567));
  A2O1A1Ixp33_ASAP7_75t_L   g19311(.A1(new_n19241), .A2(new_n19242), .B(new_n5666), .C(new_n19566), .Y(new_n19568));
  A2O1A1Ixp33_ASAP7_75t_L   g19312(.A1(new_n12669), .A2(\b[40] ), .B(new_n19457), .C(new_n19568), .Y(new_n19569));
  AND2x2_ASAP7_75t_L        g19313(.A(new_n19569), .B(new_n19567), .Y(new_n19570));
  A2O1A1Ixp33_ASAP7_75t_L   g19314(.A1(new_n19467), .A2(new_n19464), .B(new_n19461), .C(new_n19570), .Y(new_n19571));
  INVx1_ASAP7_75t_L         g19315(.A(new_n19570), .Y(new_n19572));
  NAND3xp33_ASAP7_75t_L     g19316(.A(new_n19468), .B(new_n19462), .C(new_n19572), .Y(new_n19573));
  AND2x2_ASAP7_75t_L        g19317(.A(new_n19571), .B(new_n19573), .Y(new_n19574));
  AOI22xp33_ASAP7_75t_L     g19318(.A1(new_n11656), .A2(\b[44] ), .B1(new_n11654), .B2(new_n7055), .Y(new_n19575));
  OAI221xp5_ASAP7_75t_L     g19319(.A1(new_n12364), .A2(new_n6195), .B1(new_n5680), .B2(new_n13003), .C(new_n19575), .Y(new_n19576));
  XNOR2x2_ASAP7_75t_L       g19320(.A(\a[62] ), .B(new_n19576), .Y(new_n19577));
  NOR2xp33_ASAP7_75t_L      g19321(.A(new_n19577), .B(new_n19574), .Y(new_n19578));
  INVx1_ASAP7_75t_L         g19322(.A(new_n19578), .Y(new_n19579));
  NAND2xp33_ASAP7_75t_L     g19323(.A(new_n19577), .B(new_n19574), .Y(new_n19580));
  NAND3xp33_ASAP7_75t_L     g19324(.A(new_n19579), .B(new_n19565), .C(new_n19580), .Y(new_n19581));
  AO21x2_ASAP7_75t_L        g19325(.A1(new_n19580), .A2(new_n19579), .B(new_n19565), .Y(new_n19582));
  AND2x2_ASAP7_75t_L        g19326(.A(new_n19581), .B(new_n19582), .Y(new_n19583));
  A2O1A1O1Ixp25_ASAP7_75t_L g19327(.A1(new_n19367), .A2(new_n19361), .B(new_n19470), .C(new_n19476), .D(new_n19583), .Y(new_n19584));
  AND3x1_ASAP7_75t_L        g19328(.A(new_n19583), .B(new_n19476), .C(new_n19472), .Y(new_n19585));
  NOR2xp33_ASAP7_75t_L      g19329(.A(new_n19584), .B(new_n19585), .Y(new_n19586));
  INVx1_ASAP7_75t_L         g19330(.A(new_n19586), .Y(new_n19587));
  AOI22xp33_ASAP7_75t_L     g19331(.A1(new_n9623), .A2(\b[50] ), .B1(new_n9620), .B2(new_n8235), .Y(new_n19588));
  OAI221xp5_ASAP7_75t_L     g19332(.A1(new_n10280), .A2(new_n7907), .B1(new_n7333), .B2(new_n12010), .C(new_n19588), .Y(new_n19589));
  XNOR2x2_ASAP7_75t_L       g19333(.A(\a[56] ), .B(new_n19589), .Y(new_n19590));
  AND2x2_ASAP7_75t_L        g19334(.A(new_n19590), .B(new_n19587), .Y(new_n19591));
  NOR2xp33_ASAP7_75t_L      g19335(.A(new_n19590), .B(new_n19587), .Y(new_n19592));
  NOR2xp33_ASAP7_75t_L      g19336(.A(new_n19592), .B(new_n19591), .Y(new_n19593));
  AND3x1_ASAP7_75t_L        g19337(.A(new_n19593), .B(new_n19488), .C(new_n19479), .Y(new_n19594));
  A2O1A1Ixp33_ASAP7_75t_L   g19338(.A1(new_n19368), .A2(new_n19367), .B(new_n19372), .C(new_n19456), .Y(new_n19595));
  O2A1O1Ixp33_ASAP7_75t_L   g19339(.A1(new_n19480), .A2(new_n19595), .B(new_n19488), .C(new_n19593), .Y(new_n19596));
  NOR3xp33_ASAP7_75t_L      g19340(.A(new_n19594), .B(new_n19596), .C(new_n19561), .Y(new_n19597));
  OA21x2_ASAP7_75t_L        g19341(.A1(new_n19596), .A2(new_n19594), .B(new_n19561), .Y(new_n19598));
  NOR2xp33_ASAP7_75t_L      g19342(.A(new_n19597), .B(new_n19598), .Y(new_n19599));
  INVx1_ASAP7_75t_L         g19343(.A(new_n19599), .Y(new_n19600));
  NAND2xp33_ASAP7_75t_L     g19344(.A(new_n19492), .B(new_n19501), .Y(new_n19601));
  NOR2xp33_ASAP7_75t_L      g19345(.A(new_n19601), .B(new_n19600), .Y(new_n19602));
  O2A1O1Ixp33_ASAP7_75t_L   g19346(.A1(new_n19495), .A2(new_n19499), .B(new_n19492), .C(new_n19599), .Y(new_n19603));
  NOR2xp33_ASAP7_75t_L      g19347(.A(new_n19603), .B(new_n19602), .Y(new_n19604));
  NAND2xp33_ASAP7_75t_L     g19348(.A(new_n19558), .B(new_n19604), .Y(new_n19605));
  INVx1_ASAP7_75t_L         g19349(.A(new_n19605), .Y(new_n19606));
  NOR2xp33_ASAP7_75t_L      g19350(.A(new_n19558), .B(new_n19604), .Y(new_n19607));
  NOR2xp33_ASAP7_75t_L      g19351(.A(new_n19607), .B(new_n19606), .Y(new_n19608));
  A2O1A1Ixp33_ASAP7_75t_L   g19352(.A1(new_n19515), .A2(new_n19553), .B(new_n19554), .C(new_n19608), .Y(new_n19609));
  INVx1_ASAP7_75t_L         g19353(.A(new_n19554), .Y(new_n19610));
  A2O1A1Ixp33_ASAP7_75t_L   g19354(.A1(new_n19505), .A2(new_n19507), .B(new_n19514), .C(new_n19610), .Y(new_n19611));
  NOR2xp33_ASAP7_75t_L      g19355(.A(new_n19611), .B(new_n19608), .Y(new_n19612));
  INVx1_ASAP7_75t_L         g19356(.A(new_n19612), .Y(new_n19613));
  AOI22xp33_ASAP7_75t_L     g19357(.A1(new_n6822), .A2(\b[59] ), .B1(new_n6819), .B2(new_n10887), .Y(new_n19614));
  OAI221xp5_ASAP7_75t_L     g19358(.A1(new_n7392), .A2(new_n10848), .B1(new_n10488), .B2(new_n7115), .C(new_n19614), .Y(new_n19615));
  XNOR2x2_ASAP7_75t_L       g19359(.A(\a[47] ), .B(new_n19615), .Y(new_n19616));
  NAND3xp33_ASAP7_75t_L     g19360(.A(new_n19613), .B(new_n19609), .C(new_n19616), .Y(new_n19617));
  AO21x2_ASAP7_75t_L        g19361(.A1(new_n19609), .A2(new_n19613), .B(new_n19616), .Y(new_n19618));
  AND2x2_ASAP7_75t_L        g19362(.A(new_n19617), .B(new_n19618), .Y(new_n19619));
  INVx1_ASAP7_75t_L         g19363(.A(new_n19619), .Y(new_n19620));
  O2A1O1Ixp33_ASAP7_75t_L   g19364(.A1(new_n19455), .A2(new_n19516), .B(new_n19525), .C(new_n19620), .Y(new_n19621));
  AND3x1_ASAP7_75t_L        g19365(.A(new_n19620), .B(new_n19525), .C(new_n19517), .Y(new_n19622));
  NOR2xp33_ASAP7_75t_L      g19366(.A(new_n19621), .B(new_n19622), .Y(new_n19623));
  AOI22xp33_ASAP7_75t_L     g19367(.A1(new_n6002), .A2(\b[62] ), .B1(new_n5999), .B2(new_n12280), .Y(new_n19624));
  OAI221xp5_ASAP7_75t_L     g19368(.A1(new_n6544), .A2(new_n11911), .B1(new_n11226), .B2(new_n6309), .C(new_n19624), .Y(new_n19625));
  XNOR2x2_ASAP7_75t_L       g19369(.A(\a[44] ), .B(new_n19625), .Y(new_n19626));
  XOR2x2_ASAP7_75t_L        g19370(.A(new_n19626), .B(new_n19623), .Y(new_n19627));
  INVx1_ASAP7_75t_L         g19371(.A(new_n19627), .Y(new_n19628));
  O2A1O1Ixp33_ASAP7_75t_L   g19372(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n5252), .Y(new_n19629));
  O2A1O1Ixp33_ASAP7_75t_L   g19373(.A1(new_n5526), .A2(new_n19629), .B(\b[63] ), .C(new_n5244), .Y(new_n19630));
  A2O1A1O1Ixp25_ASAP7_75t_L g19374(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n5247), .D(new_n5526), .Y(new_n19631));
  NOR3xp33_ASAP7_75t_L      g19375(.A(new_n19631), .B(new_n12599), .C(\a[41] ), .Y(new_n19632));
  NOR2xp33_ASAP7_75t_L      g19376(.A(new_n19630), .B(new_n19632), .Y(new_n19633));
  A2O1A1O1Ixp25_ASAP7_75t_L g19377(.A1(new_n19526), .A2(new_n19525), .B(new_n19529), .C(new_n19537), .D(new_n19633), .Y(new_n19634));
  INVx1_ASAP7_75t_L         g19378(.A(new_n19634), .Y(new_n19635));
  O2A1O1Ixp33_ASAP7_75t_L   g19379(.A1(new_n19409), .A2(new_n19528), .B(new_n19527), .C(new_n19538), .Y(new_n19636));
  NAND2xp33_ASAP7_75t_L     g19380(.A(new_n19633), .B(new_n19636), .Y(new_n19637));
  NAND2xp33_ASAP7_75t_L     g19381(.A(new_n19635), .B(new_n19637), .Y(new_n19638));
  XNOR2x2_ASAP7_75t_L       g19382(.A(new_n19628), .B(new_n19638), .Y(new_n19639));
  INVx1_ASAP7_75t_L         g19383(.A(new_n19639), .Y(new_n19640));
  O2A1O1Ixp33_ASAP7_75t_L   g19384(.A1(new_n19453), .A2(new_n19450), .B(new_n19541), .C(new_n19640), .Y(new_n19641));
  A2O1A1Ixp33_ASAP7_75t_L   g19385(.A1(new_n19447), .A2(new_n19449), .B(new_n19453), .C(new_n19541), .Y(new_n19642));
  NOR2xp33_ASAP7_75t_L      g19386(.A(new_n19639), .B(new_n19642), .Y(new_n19643));
  NOR2xp33_ASAP7_75t_L      g19387(.A(new_n19643), .B(new_n19641), .Y(new_n19644));
  XNOR2x2_ASAP7_75t_L       g19388(.A(new_n19644), .B(new_n19552), .Y(\f[104] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19389(.A1(new_n19549), .A2(new_n19546), .B(new_n19545), .C(new_n19644), .Y(new_n19646));
  NAND2xp33_ASAP7_75t_L     g19390(.A(new_n19626), .B(new_n19623), .Y(new_n19647));
  AOI22xp33_ASAP7_75t_L     g19391(.A1(new_n7659), .A2(\b[57] ), .B1(new_n7656), .B2(new_n10495), .Y(new_n19648));
  OAI221xp5_ASAP7_75t_L     g19392(.A1(new_n8326), .A2(new_n10178), .B1(new_n9534), .B2(new_n7994), .C(new_n19648), .Y(new_n19649));
  XNOR2x2_ASAP7_75t_L       g19393(.A(new_n7653), .B(new_n19649), .Y(new_n19650));
  NOR2xp33_ASAP7_75t_L      g19394(.A(new_n19585), .B(new_n19592), .Y(new_n19651));
  AOI22xp33_ASAP7_75t_L     g19395(.A1(new_n9623), .A2(\b[51] ), .B1(new_n9620), .B2(new_n8257), .Y(new_n19652));
  OAI221xp5_ASAP7_75t_L     g19396(.A1(new_n10280), .A2(new_n8228), .B1(new_n7907), .B2(new_n12010), .C(new_n19652), .Y(new_n19653));
  XNOR2x2_ASAP7_75t_L       g19397(.A(\a[56] ), .B(new_n19653), .Y(new_n19654));
  A2O1A1Ixp33_ASAP7_75t_L   g19398(.A1(new_n12669), .A2(\b[40] ), .B(new_n19457), .C(\a[41] ), .Y(new_n19655));
  NOR2xp33_ASAP7_75t_L      g19399(.A(\a[41] ), .B(new_n19459), .Y(new_n19656));
  INVx1_ASAP7_75t_L         g19400(.A(new_n19656), .Y(new_n19657));
  AND2x2_ASAP7_75t_L        g19401(.A(new_n19655), .B(new_n19657), .Y(new_n19658));
  NOR2xp33_ASAP7_75t_L      g19402(.A(new_n5666), .B(new_n12671), .Y(new_n19659));
  O2A1O1Ixp33_ASAP7_75t_L   g19403(.A1(new_n12353), .A2(new_n12355), .B(\b[42] ), .C(new_n19659), .Y(new_n19660));
  NAND2xp33_ASAP7_75t_L     g19404(.A(new_n19660), .B(new_n19658), .Y(new_n19661));
  INVx1_ASAP7_75t_L         g19405(.A(new_n19658), .Y(new_n19662));
  A2O1A1Ixp33_ASAP7_75t_L   g19406(.A1(\b[42] ), .A2(new_n12669), .B(new_n19659), .C(new_n19662), .Y(new_n19663));
  AND2x2_ASAP7_75t_L        g19407(.A(new_n19661), .B(new_n19663), .Y(new_n19664));
  INVx1_ASAP7_75t_L         g19408(.A(new_n19664), .Y(new_n19665));
  AOI22xp33_ASAP7_75t_L     g19409(.A1(new_n11656), .A2(\b[45] ), .B1(new_n11654), .B2(new_n6764), .Y(new_n19666));
  OAI221xp5_ASAP7_75t_L     g19410(.A1(new_n12364), .A2(new_n6220), .B1(new_n6195), .B2(new_n13003), .C(new_n19666), .Y(new_n19667));
  XNOR2x2_ASAP7_75t_L       g19411(.A(\a[62] ), .B(new_n19667), .Y(new_n19668));
  XNOR2x2_ASAP7_75t_L       g19412(.A(new_n19665), .B(new_n19668), .Y(new_n19669));
  O2A1O1Ixp33_ASAP7_75t_L   g19413(.A1(new_n12356), .A2(new_n5666), .B(new_n19566), .C(new_n19459), .Y(new_n19670));
  A2O1A1O1Ixp25_ASAP7_75t_L g19414(.A1(new_n19464), .A2(new_n19467), .B(new_n19461), .C(new_n19572), .D(new_n19670), .Y(new_n19671));
  NAND2xp33_ASAP7_75t_L     g19415(.A(new_n19671), .B(new_n19669), .Y(new_n19672));
  A2O1A1Ixp33_ASAP7_75t_L   g19416(.A1(new_n19460), .A2(new_n19354), .B(new_n19459), .C(new_n19468), .Y(new_n19673));
  INVx1_ASAP7_75t_L         g19417(.A(new_n19669), .Y(new_n19674));
  A2O1A1Ixp33_ASAP7_75t_L   g19418(.A1(new_n19673), .A2(new_n19572), .B(new_n19670), .C(new_n19674), .Y(new_n19675));
  AND2x2_ASAP7_75t_L        g19419(.A(new_n19672), .B(new_n19675), .Y(new_n19676));
  AOI22xp33_ASAP7_75t_L     g19420(.A1(new_n10594), .A2(\b[48] ), .B1(new_n10591), .B2(new_n7341), .Y(new_n19677));
  OAI221xp5_ASAP7_75t_L     g19421(.A1(new_n11335), .A2(new_n7316), .B1(new_n7033), .B2(new_n11330), .C(new_n19677), .Y(new_n19678));
  XNOR2x2_ASAP7_75t_L       g19422(.A(\a[59] ), .B(new_n19678), .Y(new_n19679));
  INVx1_ASAP7_75t_L         g19423(.A(new_n19679), .Y(new_n19680));
  XNOR2x2_ASAP7_75t_L       g19424(.A(new_n19680), .B(new_n19676), .Y(new_n19681));
  O2A1O1Ixp33_ASAP7_75t_L   g19425(.A1(new_n19574), .A2(new_n19577), .B(new_n19581), .C(new_n19681), .Y(new_n19682));
  INVx1_ASAP7_75t_L         g19426(.A(new_n19682), .Y(new_n19683));
  A2O1A1Ixp33_ASAP7_75t_L   g19427(.A1(new_n19573), .A2(new_n19571), .B(new_n19577), .C(new_n19581), .Y(new_n19684));
  INVx1_ASAP7_75t_L         g19428(.A(new_n19684), .Y(new_n19685));
  NAND2xp33_ASAP7_75t_L     g19429(.A(new_n19685), .B(new_n19681), .Y(new_n19686));
  AND2x2_ASAP7_75t_L        g19430(.A(new_n19686), .B(new_n19683), .Y(new_n19687));
  XOR2x2_ASAP7_75t_L        g19431(.A(new_n19654), .B(new_n19687), .Y(new_n19688));
  XNOR2x2_ASAP7_75t_L       g19432(.A(new_n19651), .B(new_n19688), .Y(new_n19689));
  AOI22xp33_ASAP7_75t_L     g19433(.A1(new_n8645), .A2(\b[54] ), .B1(new_n8642), .B2(new_n9208), .Y(new_n19690));
  OAI221xp5_ASAP7_75t_L     g19434(.A1(new_n9322), .A2(new_n8882), .B1(new_n8569), .B2(new_n8965), .C(new_n19690), .Y(new_n19691));
  XNOR2x2_ASAP7_75t_L       g19435(.A(\a[53] ), .B(new_n19691), .Y(new_n19692));
  AND2x2_ASAP7_75t_L        g19436(.A(new_n19692), .B(new_n19689), .Y(new_n19693));
  NOR2xp33_ASAP7_75t_L      g19437(.A(new_n19692), .B(new_n19689), .Y(new_n19694));
  NOR2xp33_ASAP7_75t_L      g19438(.A(new_n19694), .B(new_n19693), .Y(new_n19695));
  OA21x2_ASAP7_75t_L        g19439(.A1(new_n19594), .A2(new_n19597), .B(new_n19695), .Y(new_n19696));
  NOR3xp33_ASAP7_75t_L      g19440(.A(new_n19695), .B(new_n19597), .C(new_n19594), .Y(new_n19697));
  NOR2xp33_ASAP7_75t_L      g19441(.A(new_n19697), .B(new_n19696), .Y(new_n19698));
  XOR2x2_ASAP7_75t_L        g19442(.A(new_n19650), .B(new_n19698), .Y(new_n19699));
  A2O1A1Ixp33_ASAP7_75t_L   g19443(.A1(new_n19604), .A2(new_n19558), .B(new_n19602), .C(new_n19699), .Y(new_n19700));
  OR3x1_ASAP7_75t_L         g19444(.A(new_n19699), .B(new_n19602), .C(new_n19606), .Y(new_n19701));
  NAND2xp33_ASAP7_75t_L     g19445(.A(new_n19700), .B(new_n19701), .Y(new_n19702));
  AOI22xp33_ASAP7_75t_L     g19446(.A1(new_n6822), .A2(\b[60] ), .B1(new_n6819), .B2(new_n11234), .Y(new_n19703));
  OAI221xp5_ASAP7_75t_L     g19447(.A1(new_n7392), .A2(new_n10881), .B1(new_n10848), .B2(new_n7115), .C(new_n19703), .Y(new_n19704));
  XNOR2x2_ASAP7_75t_L       g19448(.A(\a[47] ), .B(new_n19704), .Y(new_n19705));
  XNOR2x2_ASAP7_75t_L       g19449(.A(new_n19705), .B(new_n19702), .Y(new_n19706));
  A2O1A1Ixp33_ASAP7_75t_L   g19450(.A1(new_n19616), .A2(new_n19609), .B(new_n19612), .C(new_n19706), .Y(new_n19707));
  INVx1_ASAP7_75t_L         g19451(.A(new_n19706), .Y(new_n19708));
  NAND3xp33_ASAP7_75t_L     g19452(.A(new_n19708), .B(new_n19617), .C(new_n19613), .Y(new_n19709));
  NAND2xp33_ASAP7_75t_L     g19453(.A(new_n19707), .B(new_n19709), .Y(new_n19710));
  NAND2xp33_ASAP7_75t_L     g19454(.A(\b[63] ), .B(new_n6002), .Y(new_n19711));
  A2O1A1Ixp33_ASAP7_75t_L   g19455(.A1(new_n12607), .A2(new_n12603), .B(new_n6311), .C(new_n19711), .Y(new_n19712));
  AOI221xp5_ASAP7_75t_L     g19456(.A1(\b[61] ), .A2(new_n6308), .B1(\b[62] ), .B2(new_n5992), .C(new_n19712), .Y(new_n19713));
  XNOR2x2_ASAP7_75t_L       g19457(.A(new_n5996), .B(new_n19713), .Y(new_n19714));
  XNOR2x2_ASAP7_75t_L       g19458(.A(new_n19714), .B(new_n19710), .Y(new_n19715));
  INVx1_ASAP7_75t_L         g19459(.A(new_n19715), .Y(new_n19716));
  A2O1A1O1Ixp25_ASAP7_75t_L g19460(.A1(new_n19525), .A2(new_n19517), .B(new_n19620), .C(new_n19647), .D(new_n19716), .Y(new_n19717));
  A2O1A1Ixp33_ASAP7_75t_L   g19461(.A1(new_n19525), .A2(new_n19517), .B(new_n19620), .C(new_n19647), .Y(new_n19718));
  NOR2xp33_ASAP7_75t_L      g19462(.A(new_n19718), .B(new_n19715), .Y(new_n19719));
  NOR2xp33_ASAP7_75t_L      g19463(.A(new_n19719), .B(new_n19717), .Y(new_n19720));
  INVx1_ASAP7_75t_L         g19464(.A(new_n19720), .Y(new_n19721));
  A2O1A1Ixp33_ASAP7_75t_L   g19465(.A1(new_n19407), .A2(new_n19406), .B(new_n19528), .C(new_n19527), .Y(new_n19722));
  A2O1A1Ixp33_ASAP7_75t_L   g19466(.A1(new_n19722), .A2(new_n19537), .B(new_n19633), .C(new_n19627), .Y(new_n19723));
  NAND2xp33_ASAP7_75t_L     g19467(.A(new_n19723), .B(new_n19637), .Y(new_n19724));
  NOR2xp33_ASAP7_75t_L      g19468(.A(new_n19724), .B(new_n19721), .Y(new_n19725));
  O2A1O1Ixp33_ASAP7_75t_L   g19469(.A1(new_n19628), .A2(new_n19634), .B(new_n19637), .C(new_n19720), .Y(new_n19726));
  NOR2xp33_ASAP7_75t_L      g19470(.A(new_n19726), .B(new_n19725), .Y(new_n19727));
  INVx1_ASAP7_75t_L         g19471(.A(new_n19727), .Y(new_n19728));
  A2O1A1O1Ixp25_ASAP7_75t_L g19472(.A1(new_n19541), .A2(new_n19452), .B(new_n19640), .C(new_n19646), .D(new_n19728), .Y(new_n19729));
  A2O1A1Ixp33_ASAP7_75t_L   g19473(.A1(new_n19541), .A2(new_n19452), .B(new_n19640), .C(new_n19646), .Y(new_n19730));
  NOR2xp33_ASAP7_75t_L      g19474(.A(new_n19727), .B(new_n19730), .Y(new_n19731));
  NOR2xp33_ASAP7_75t_L      g19475(.A(new_n19729), .B(new_n19731), .Y(\f[105] ));
  INVx1_ASAP7_75t_L         g19476(.A(new_n19641), .Y(new_n19733));
  INVx1_ASAP7_75t_L         g19477(.A(new_n19725), .Y(new_n19734));
  OAI21xp33_ASAP7_75t_L     g19478(.A1(new_n19702), .A2(new_n19705), .B(new_n19709), .Y(new_n19735));
  OAI22xp33_ASAP7_75t_L     g19479(.A1(new_n6309), .A2(new_n12273), .B1(new_n12599), .B2(new_n6544), .Y(new_n19736));
  A2O1A1O1Ixp25_ASAP7_75t_L g19480(.A1(new_n12600), .A2(new_n12597), .B(new_n12628), .C(new_n5999), .D(new_n19736), .Y(new_n19737));
  NAND2xp33_ASAP7_75t_L     g19481(.A(\a[44] ), .B(new_n19737), .Y(new_n19738));
  A2O1A1Ixp33_ASAP7_75t_L   g19482(.A1(new_n12276), .A2(new_n12605), .B(new_n12627), .C(new_n13507), .Y(new_n19739));
  A2O1A1Ixp33_ASAP7_75t_L   g19483(.A1(new_n19739), .A2(new_n5999), .B(new_n19736), .C(new_n5996), .Y(new_n19740));
  NAND2xp33_ASAP7_75t_L     g19484(.A(new_n19738), .B(new_n19740), .Y(new_n19741));
  XNOR2x2_ASAP7_75t_L       g19485(.A(new_n19741), .B(new_n19735), .Y(new_n19742));
  NAND2xp33_ASAP7_75t_L     g19486(.A(\b[61] ), .B(new_n6822), .Y(new_n19743));
  OAI221xp5_ASAP7_75t_L     g19487(.A1(new_n11226), .A2(new_n7392), .B1(new_n7117), .B2(new_n11920), .C(new_n19743), .Y(new_n19744));
  AOI21xp33_ASAP7_75t_L     g19488(.A1(new_n7124), .A2(\b[59] ), .B(new_n19744), .Y(new_n19745));
  NAND2xp33_ASAP7_75t_L     g19489(.A(\a[47] ), .B(new_n19745), .Y(new_n19746));
  A2O1A1Ixp33_ASAP7_75t_L   g19490(.A1(\b[59] ), .A2(new_n7124), .B(new_n19744), .C(new_n6816), .Y(new_n19747));
  NAND2xp33_ASAP7_75t_L     g19491(.A(new_n19747), .B(new_n19746), .Y(new_n19748));
  INVx1_ASAP7_75t_L         g19492(.A(new_n19700), .Y(new_n19749));
  O2A1O1Ixp33_ASAP7_75t_L   g19493(.A1(new_n19597), .A2(new_n19594), .B(new_n19695), .C(new_n19694), .Y(new_n19750));
  NOR2xp33_ASAP7_75t_L      g19494(.A(new_n5680), .B(new_n12671), .Y(new_n19751));
  O2A1O1Ixp33_ASAP7_75t_L   g19495(.A1(new_n12353), .A2(new_n12355), .B(\b[43] ), .C(new_n19751), .Y(new_n19752));
  INVx1_ASAP7_75t_L         g19496(.A(new_n19663), .Y(new_n19753));
  A2O1A1O1Ixp25_ASAP7_75t_L g19497(.A1(new_n12669), .A2(\b[40] ), .B(new_n19457), .C(new_n5244), .D(new_n19753), .Y(new_n19754));
  NAND2xp33_ASAP7_75t_L     g19498(.A(new_n19752), .B(new_n19754), .Y(new_n19755));
  INVx1_ASAP7_75t_L         g19499(.A(new_n19752), .Y(new_n19756));
  A2O1A1Ixp33_ASAP7_75t_L   g19500(.A1(new_n19459), .A2(new_n5244), .B(new_n19753), .C(new_n19756), .Y(new_n19757));
  AND2x2_ASAP7_75t_L        g19501(.A(new_n19757), .B(new_n19755), .Y(new_n19758));
  AOI22xp33_ASAP7_75t_L     g19502(.A1(new_n11647), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n11656), .Y(new_n19759));
  OAI221xp5_ASAP7_75t_L     g19503(.A1(new_n13003), .A2(new_n6220), .B1(new_n12022), .B2(new_n7887), .C(new_n19759), .Y(new_n19760));
  XNOR2x2_ASAP7_75t_L       g19504(.A(\a[62] ), .B(new_n19760), .Y(new_n19761));
  NOR2xp33_ASAP7_75t_L      g19505(.A(new_n19758), .B(new_n19761), .Y(new_n19762));
  INVx1_ASAP7_75t_L         g19506(.A(new_n19762), .Y(new_n19763));
  NAND2xp33_ASAP7_75t_L     g19507(.A(new_n19758), .B(new_n19761), .Y(new_n19764));
  AND2x2_ASAP7_75t_L        g19508(.A(new_n19764), .B(new_n19763), .Y(new_n19765));
  INVx1_ASAP7_75t_L         g19509(.A(new_n19765), .Y(new_n19766));
  O2A1O1Ixp33_ASAP7_75t_L   g19510(.A1(new_n19665), .A2(new_n19668), .B(new_n19675), .C(new_n19766), .Y(new_n19767));
  OA211x2_ASAP7_75t_L       g19511(.A1(new_n19668), .A2(new_n19665), .B(new_n19766), .C(new_n19675), .Y(new_n19768));
  NOR2xp33_ASAP7_75t_L      g19512(.A(new_n19767), .B(new_n19768), .Y(new_n19769));
  AOI22xp33_ASAP7_75t_L     g19513(.A1(new_n10594), .A2(\b[49] ), .B1(new_n10591), .B2(new_n7914), .Y(new_n19770));
  OAI221xp5_ASAP7_75t_L     g19514(.A1(new_n11335), .A2(new_n7333), .B1(new_n7316), .B2(new_n11330), .C(new_n19770), .Y(new_n19771));
  XNOR2x2_ASAP7_75t_L       g19515(.A(\a[59] ), .B(new_n19771), .Y(new_n19772));
  AND2x2_ASAP7_75t_L        g19516(.A(new_n19772), .B(new_n19769), .Y(new_n19773));
  NOR2xp33_ASAP7_75t_L      g19517(.A(new_n19772), .B(new_n19769), .Y(new_n19774));
  NOR2xp33_ASAP7_75t_L      g19518(.A(new_n19774), .B(new_n19773), .Y(new_n19775));
  INVx1_ASAP7_75t_L         g19519(.A(new_n19775), .Y(new_n19776));
  NAND2xp33_ASAP7_75t_L     g19520(.A(new_n19680), .B(new_n19676), .Y(new_n19777));
  A2O1A1Ixp33_ASAP7_75t_L   g19521(.A1(new_n19581), .A2(new_n19579), .B(new_n19681), .C(new_n19777), .Y(new_n19778));
  NOR2xp33_ASAP7_75t_L      g19522(.A(new_n19778), .B(new_n19776), .Y(new_n19779));
  INVx1_ASAP7_75t_L         g19523(.A(new_n19779), .Y(new_n19780));
  O2A1O1Ixp33_ASAP7_75t_L   g19524(.A1(new_n19685), .A2(new_n19681), .B(new_n19777), .C(new_n19775), .Y(new_n19781));
  INVx1_ASAP7_75t_L         g19525(.A(new_n19781), .Y(new_n19782));
  AOI22xp33_ASAP7_75t_L     g19526(.A1(new_n9623), .A2(\b[52] ), .B1(new_n9620), .B2(new_n8577), .Y(new_n19783));
  OAI221xp5_ASAP7_75t_L     g19527(.A1(new_n10280), .A2(new_n8249), .B1(new_n8228), .B2(new_n12010), .C(new_n19783), .Y(new_n19784));
  XNOR2x2_ASAP7_75t_L       g19528(.A(\a[56] ), .B(new_n19784), .Y(new_n19785));
  NAND3xp33_ASAP7_75t_L     g19529(.A(new_n19780), .B(new_n19782), .C(new_n19785), .Y(new_n19786));
  INVx1_ASAP7_75t_L         g19530(.A(new_n19786), .Y(new_n19787));
  AOI21xp33_ASAP7_75t_L     g19531(.A1(new_n19780), .A2(new_n19782), .B(new_n19785), .Y(new_n19788));
  NOR2xp33_ASAP7_75t_L      g19532(.A(new_n19788), .B(new_n19787), .Y(new_n19789));
  INVx1_ASAP7_75t_L         g19533(.A(new_n19789), .Y(new_n19790));
  INVx1_ASAP7_75t_L         g19534(.A(new_n19687), .Y(new_n19791));
  MAJIxp5_ASAP7_75t_L       g19535(.A(new_n19791), .B(new_n19651), .C(new_n19654), .Y(new_n19792));
  NOR2xp33_ASAP7_75t_L      g19536(.A(new_n19792), .B(new_n19790), .Y(new_n19793));
  AND2x2_ASAP7_75t_L        g19537(.A(new_n19792), .B(new_n19790), .Y(new_n19794));
  NOR2xp33_ASAP7_75t_L      g19538(.A(new_n19793), .B(new_n19794), .Y(new_n19795));
  AOI22xp33_ASAP7_75t_L     g19539(.A1(new_n8645), .A2(\b[55] ), .B1(new_n8642), .B2(new_n9542), .Y(new_n19796));
  OAI221xp5_ASAP7_75t_L     g19540(.A1(new_n9322), .A2(new_n9199), .B1(new_n8882), .B2(new_n8965), .C(new_n19796), .Y(new_n19797));
  XNOR2x2_ASAP7_75t_L       g19541(.A(\a[53] ), .B(new_n19797), .Y(new_n19798));
  AND2x2_ASAP7_75t_L        g19542(.A(new_n19798), .B(new_n19795), .Y(new_n19799));
  NOR2xp33_ASAP7_75t_L      g19543(.A(new_n19798), .B(new_n19795), .Y(new_n19800));
  NOR2xp33_ASAP7_75t_L      g19544(.A(new_n19800), .B(new_n19799), .Y(new_n19801));
  XNOR2x2_ASAP7_75t_L       g19545(.A(new_n19750), .B(new_n19801), .Y(new_n19802));
  AOI22xp33_ASAP7_75t_L     g19546(.A1(new_n7659), .A2(\b[58] ), .B1(new_n7656), .B2(new_n10857), .Y(new_n19803));
  OAI221xp5_ASAP7_75t_L     g19547(.A1(new_n8326), .A2(new_n10488), .B1(new_n10178), .B2(new_n7994), .C(new_n19803), .Y(new_n19804));
  XNOR2x2_ASAP7_75t_L       g19548(.A(\a[50] ), .B(new_n19804), .Y(new_n19805));
  XOR2x2_ASAP7_75t_L        g19549(.A(new_n19805), .B(new_n19802), .Y(new_n19806));
  A2O1A1Ixp33_ASAP7_75t_L   g19550(.A1(new_n19698), .A2(new_n19650), .B(new_n19749), .C(new_n19806), .Y(new_n19807));
  AO21x2_ASAP7_75t_L        g19551(.A1(new_n19650), .A2(new_n19698), .B(new_n19749), .Y(new_n19808));
  NOR2xp33_ASAP7_75t_L      g19552(.A(new_n19806), .B(new_n19808), .Y(new_n19809));
  INVx1_ASAP7_75t_L         g19553(.A(new_n19809), .Y(new_n19810));
  NAND2xp33_ASAP7_75t_L     g19554(.A(new_n19807), .B(new_n19810), .Y(new_n19811));
  XOR2x2_ASAP7_75t_L        g19555(.A(new_n19748), .B(new_n19811), .Y(new_n19812));
  INVx1_ASAP7_75t_L         g19556(.A(new_n19812), .Y(new_n19813));
  NOR2xp33_ASAP7_75t_L      g19557(.A(new_n19813), .B(new_n19742), .Y(new_n19814));
  AND2x2_ASAP7_75t_L        g19558(.A(new_n19813), .B(new_n19742), .Y(new_n19815));
  NOR2xp33_ASAP7_75t_L      g19559(.A(new_n19714), .B(new_n19710), .Y(new_n19816));
  NOR4xp25_ASAP7_75t_L      g19560(.A(new_n19815), .B(new_n19719), .C(new_n19816), .D(new_n19814), .Y(new_n19817));
  NOR2xp33_ASAP7_75t_L      g19561(.A(new_n19814), .B(new_n19815), .Y(new_n19818));
  NOR2xp33_ASAP7_75t_L      g19562(.A(new_n19816), .B(new_n19719), .Y(new_n19819));
  NOR2xp33_ASAP7_75t_L      g19563(.A(new_n19819), .B(new_n19818), .Y(new_n19820));
  NOR2xp33_ASAP7_75t_L      g19564(.A(new_n19817), .B(new_n19820), .Y(new_n19821));
  INVx1_ASAP7_75t_L         g19565(.A(new_n19821), .Y(new_n19822));
  A2O1A1O1Ixp25_ASAP7_75t_L g19566(.A1(new_n19733), .A2(new_n19646), .B(new_n19726), .C(new_n19734), .D(new_n19822), .Y(new_n19823));
  A2O1A1Ixp33_ASAP7_75t_L   g19567(.A1(new_n19646), .A2(new_n19733), .B(new_n19728), .C(new_n19734), .Y(new_n19824));
  NOR2xp33_ASAP7_75t_L      g19568(.A(new_n19821), .B(new_n19824), .Y(new_n19825));
  NOR2xp33_ASAP7_75t_L      g19569(.A(new_n19823), .B(new_n19825), .Y(\f[106] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19570(.A1(new_n19725), .A2(new_n19729), .B(new_n19821), .C(new_n19820), .Y(new_n19827));
  NOR2xp33_ASAP7_75t_L      g19571(.A(new_n19741), .B(new_n19735), .Y(new_n19828));
  NOR2xp33_ASAP7_75t_L      g19572(.A(new_n19828), .B(new_n19814), .Y(new_n19829));
  AOI22xp33_ASAP7_75t_L     g19573(.A1(new_n6822), .A2(\b[62] ), .B1(new_n6819), .B2(new_n12280), .Y(new_n19830));
  OAI221xp5_ASAP7_75t_L     g19574(.A1(new_n7392), .A2(new_n11911), .B1(new_n11226), .B2(new_n7115), .C(new_n19830), .Y(new_n19831));
  XNOR2x2_ASAP7_75t_L       g19575(.A(\a[47] ), .B(new_n19831), .Y(new_n19832));
  AOI22xp33_ASAP7_75t_L     g19576(.A1(new_n8645), .A2(\b[56] ), .B1(new_n8642), .B2(new_n10185), .Y(new_n19833));
  OAI221xp5_ASAP7_75t_L     g19577(.A1(new_n9322), .A2(new_n9534), .B1(new_n9199), .B2(new_n8965), .C(new_n19833), .Y(new_n19834));
  XNOR2x2_ASAP7_75t_L       g19578(.A(\a[53] ), .B(new_n19834), .Y(new_n19835));
  INVx1_ASAP7_75t_L         g19579(.A(new_n19835), .Y(new_n19836));
  AOI22xp33_ASAP7_75t_L     g19580(.A1(new_n9623), .A2(\b[53] ), .B1(new_n9620), .B2(new_n8889), .Y(new_n19837));
  OAI221xp5_ASAP7_75t_L     g19581(.A1(new_n10280), .A2(new_n8569), .B1(new_n8249), .B2(new_n12010), .C(new_n19837), .Y(new_n19838));
  XNOR2x2_ASAP7_75t_L       g19582(.A(\a[56] ), .B(new_n19838), .Y(new_n19839));
  INVx1_ASAP7_75t_L         g19583(.A(new_n19839), .Y(new_n19840));
  AOI22xp33_ASAP7_75t_L     g19584(.A1(new_n10594), .A2(\b[50] ), .B1(new_n10591), .B2(new_n8235), .Y(new_n19841));
  OAI221xp5_ASAP7_75t_L     g19585(.A1(new_n11335), .A2(new_n7907), .B1(new_n7333), .B2(new_n11330), .C(new_n19841), .Y(new_n19842));
  XNOR2x2_ASAP7_75t_L       g19586(.A(\a[59] ), .B(new_n19842), .Y(new_n19843));
  NAND2xp33_ASAP7_75t_L     g19587(.A(\b[43] ), .B(new_n12670), .Y(new_n19844));
  A2O1A1Ixp33_ASAP7_75t_L   g19588(.A1(new_n19241), .A2(new_n19242), .B(new_n6220), .C(new_n19844), .Y(new_n19845));
  XNOR2x2_ASAP7_75t_L       g19589(.A(new_n19845), .B(new_n19752), .Y(new_n19846));
  NAND2xp33_ASAP7_75t_L     g19590(.A(\b[46] ), .B(new_n11647), .Y(new_n19847));
  OAI221xp5_ASAP7_75t_L     g19591(.A1(new_n12023), .A2(new_n7316), .B1(new_n12022), .B2(new_n7322), .C(new_n19847), .Y(new_n19848));
  AOI21xp33_ASAP7_75t_L     g19592(.A1(new_n12021), .A2(\b[45] ), .B(new_n19848), .Y(new_n19849));
  NAND2xp33_ASAP7_75t_L     g19593(.A(\a[62] ), .B(new_n19849), .Y(new_n19850));
  A2O1A1Ixp33_ASAP7_75t_L   g19594(.A1(\b[45] ), .A2(new_n12021), .B(new_n19848), .C(new_n11651), .Y(new_n19851));
  AOI21xp33_ASAP7_75t_L     g19595(.A1(new_n19850), .A2(new_n19851), .B(new_n19846), .Y(new_n19852));
  AND3x1_ASAP7_75t_L        g19596(.A(new_n19850), .B(new_n19851), .C(new_n19846), .Y(new_n19853));
  NOR2xp33_ASAP7_75t_L      g19597(.A(new_n19852), .B(new_n19853), .Y(new_n19854));
  INVx1_ASAP7_75t_L         g19598(.A(new_n19854), .Y(new_n19855));
  O2A1O1Ixp33_ASAP7_75t_L   g19599(.A1(new_n19756), .A2(new_n19754), .B(new_n19763), .C(new_n19855), .Y(new_n19856));
  INVx1_ASAP7_75t_L         g19600(.A(new_n19856), .Y(new_n19857));
  A2O1A1O1Ixp25_ASAP7_75t_L g19601(.A1(new_n19459), .A2(new_n5244), .B(new_n19753), .C(new_n19752), .D(new_n19762), .Y(new_n19858));
  NAND2xp33_ASAP7_75t_L     g19602(.A(new_n19858), .B(new_n19855), .Y(new_n19859));
  NAND2xp33_ASAP7_75t_L     g19603(.A(new_n19859), .B(new_n19857), .Y(new_n19860));
  NOR2xp33_ASAP7_75t_L      g19604(.A(new_n19843), .B(new_n19860), .Y(new_n19861));
  INVx1_ASAP7_75t_L         g19605(.A(new_n19861), .Y(new_n19862));
  NAND2xp33_ASAP7_75t_L     g19606(.A(new_n19843), .B(new_n19860), .Y(new_n19863));
  AND2x2_ASAP7_75t_L        g19607(.A(new_n19863), .B(new_n19862), .Y(new_n19864));
  INVx1_ASAP7_75t_L         g19608(.A(new_n19864), .Y(new_n19865));
  OR3x1_ASAP7_75t_L         g19609(.A(new_n19865), .B(new_n19768), .C(new_n19773), .Y(new_n19866));
  A2O1A1Ixp33_ASAP7_75t_L   g19610(.A1(new_n19769), .A2(new_n19772), .B(new_n19768), .C(new_n19865), .Y(new_n19867));
  NAND3xp33_ASAP7_75t_L     g19611(.A(new_n19866), .B(new_n19840), .C(new_n19867), .Y(new_n19868));
  AO21x2_ASAP7_75t_L        g19612(.A1(new_n19867), .A2(new_n19866), .B(new_n19840), .Y(new_n19869));
  AND2x2_ASAP7_75t_L        g19613(.A(new_n19868), .B(new_n19869), .Y(new_n19870));
  INVx1_ASAP7_75t_L         g19614(.A(new_n19870), .Y(new_n19871));
  NOR3xp33_ASAP7_75t_L      g19615(.A(new_n19871), .B(new_n19787), .C(new_n19779), .Y(new_n19872));
  O2A1O1Ixp33_ASAP7_75t_L   g19616(.A1(new_n19776), .A2(new_n19778), .B(new_n19786), .C(new_n19870), .Y(new_n19873));
  NOR2xp33_ASAP7_75t_L      g19617(.A(new_n19873), .B(new_n19872), .Y(new_n19874));
  NAND2xp33_ASAP7_75t_L     g19618(.A(new_n19836), .B(new_n19874), .Y(new_n19875));
  OAI21xp33_ASAP7_75t_L     g19619(.A1(new_n19873), .A2(new_n19872), .B(new_n19835), .Y(new_n19876));
  AND2x2_ASAP7_75t_L        g19620(.A(new_n19876), .B(new_n19875), .Y(new_n19877));
  NOR2xp33_ASAP7_75t_L      g19621(.A(new_n19793), .B(new_n19799), .Y(new_n19878));
  NAND2xp33_ASAP7_75t_L     g19622(.A(new_n19877), .B(new_n19878), .Y(new_n19879));
  INVx1_ASAP7_75t_L         g19623(.A(new_n19877), .Y(new_n19880));
  A2O1A1Ixp33_ASAP7_75t_L   g19624(.A1(new_n19795), .A2(new_n19798), .B(new_n19793), .C(new_n19880), .Y(new_n19881));
  AOI22xp33_ASAP7_75t_L     g19625(.A1(new_n7659), .A2(\b[59] ), .B1(new_n7656), .B2(new_n10887), .Y(new_n19882));
  OAI221xp5_ASAP7_75t_L     g19626(.A1(new_n8326), .A2(new_n10848), .B1(new_n10488), .B2(new_n7994), .C(new_n19882), .Y(new_n19883));
  XNOR2x2_ASAP7_75t_L       g19627(.A(\a[50] ), .B(new_n19883), .Y(new_n19884));
  AND3x1_ASAP7_75t_L        g19628(.A(new_n19879), .B(new_n19881), .C(new_n19884), .Y(new_n19885));
  AOI21xp33_ASAP7_75t_L     g19629(.A1(new_n19879), .A2(new_n19881), .B(new_n19884), .Y(new_n19886));
  NOR2xp33_ASAP7_75t_L      g19630(.A(new_n19886), .B(new_n19885), .Y(new_n19887));
  OAI22xp33_ASAP7_75t_L     g19631(.A1(new_n19799), .A2(new_n19800), .B1(new_n19694), .B2(new_n19696), .Y(new_n19888));
  O2A1O1Ixp33_ASAP7_75t_L   g19632(.A1(new_n19805), .A2(new_n19802), .B(new_n19888), .C(new_n19887), .Y(new_n19889));
  OA211x2_ASAP7_75t_L       g19633(.A1(new_n19802), .A2(new_n19805), .B(new_n19887), .C(new_n19888), .Y(new_n19890));
  NOR2xp33_ASAP7_75t_L      g19634(.A(new_n19889), .B(new_n19890), .Y(new_n19891));
  AND2x2_ASAP7_75t_L        g19635(.A(new_n19832), .B(new_n19891), .Y(new_n19892));
  NOR2xp33_ASAP7_75t_L      g19636(.A(new_n19832), .B(new_n19891), .Y(new_n19893));
  NOR2xp33_ASAP7_75t_L      g19637(.A(new_n19893), .B(new_n19892), .Y(new_n19894));
  A2O1A1Ixp33_ASAP7_75t_L   g19638(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n5999), .Y(new_n19895));
  A2O1A1Ixp33_ASAP7_75t_L   g19639(.A1(new_n19895), .A2(new_n6309), .B(new_n12599), .C(\a[44] ), .Y(new_n19896));
  O2A1O1Ixp33_ASAP7_75t_L   g19640(.A1(new_n6311), .A2(new_n13934), .B(new_n6309), .C(new_n12599), .Y(new_n19897));
  NAND2xp33_ASAP7_75t_L     g19641(.A(new_n5996), .B(new_n19897), .Y(new_n19898));
  NAND2xp33_ASAP7_75t_L     g19642(.A(new_n19898), .B(new_n19896), .Y(new_n19899));
  AOI31xp33_ASAP7_75t_L     g19643(.A1(new_n19807), .A2(new_n19746), .A3(new_n19747), .B(new_n19809), .Y(new_n19900));
  NAND2xp33_ASAP7_75t_L     g19644(.A(new_n19899), .B(new_n19900), .Y(new_n19901));
  INVx1_ASAP7_75t_L         g19645(.A(new_n19901), .Y(new_n19902));
  O2A1O1Ixp33_ASAP7_75t_L   g19646(.A1(new_n19748), .A2(new_n19811), .B(new_n19810), .C(new_n19899), .Y(new_n19903));
  NOR2xp33_ASAP7_75t_L      g19647(.A(new_n19902), .B(new_n19903), .Y(new_n19904));
  XNOR2x2_ASAP7_75t_L       g19648(.A(new_n19894), .B(new_n19904), .Y(new_n19905));
  XOR2x2_ASAP7_75t_L        g19649(.A(new_n19905), .B(new_n19829), .Y(new_n19906));
  XNOR2x2_ASAP7_75t_L       g19650(.A(new_n19906), .B(new_n19827), .Y(\f[107] ));
  AND2x2_ASAP7_75t_L        g19651(.A(new_n19905), .B(new_n19829), .Y(new_n19908));
  A2O1A1O1Ixp25_ASAP7_75t_L g19652(.A1(new_n19821), .A2(new_n19824), .B(new_n19820), .C(new_n19906), .D(new_n19908), .Y(new_n19909));
  AOI22xp33_ASAP7_75t_L     g19653(.A1(new_n7659), .A2(\b[60] ), .B1(new_n7656), .B2(new_n11234), .Y(new_n19910));
  OAI221xp5_ASAP7_75t_L     g19654(.A1(new_n8326), .A2(new_n10881), .B1(new_n10848), .B2(new_n7994), .C(new_n19910), .Y(new_n19911));
  XNOR2x2_ASAP7_75t_L       g19655(.A(\a[50] ), .B(new_n19911), .Y(new_n19912));
  INVx1_ASAP7_75t_L         g19656(.A(new_n19873), .Y(new_n19913));
  AOI22xp33_ASAP7_75t_L     g19657(.A1(new_n8645), .A2(\b[57] ), .B1(new_n8642), .B2(new_n10495), .Y(new_n19914));
  OAI221xp5_ASAP7_75t_L     g19658(.A1(new_n9322), .A2(new_n10178), .B1(new_n9534), .B2(new_n8965), .C(new_n19914), .Y(new_n19915));
  XNOR2x2_ASAP7_75t_L       g19659(.A(\a[53] ), .B(new_n19915), .Y(new_n19916));
  NOR3xp33_ASAP7_75t_L      g19660(.A(new_n19865), .B(new_n19773), .C(new_n19768), .Y(new_n19917));
  AOI22xp33_ASAP7_75t_L     g19661(.A1(new_n9623), .A2(\b[54] ), .B1(new_n9620), .B2(new_n9208), .Y(new_n19918));
  OAI221xp5_ASAP7_75t_L     g19662(.A1(new_n10280), .A2(new_n8882), .B1(new_n8569), .B2(new_n12010), .C(new_n19918), .Y(new_n19919));
  XNOR2x2_ASAP7_75t_L       g19663(.A(\a[56] ), .B(new_n19919), .Y(new_n19920));
  INVx1_ASAP7_75t_L         g19664(.A(new_n19920), .Y(new_n19921));
  AOI22xp33_ASAP7_75t_L     g19665(.A1(new_n10594), .A2(\b[51] ), .B1(new_n10591), .B2(new_n8257), .Y(new_n19922));
  OAI221xp5_ASAP7_75t_L     g19666(.A1(new_n11335), .A2(new_n8228), .B1(new_n7907), .B2(new_n11330), .C(new_n19922), .Y(new_n19923));
  XNOR2x2_ASAP7_75t_L       g19667(.A(\a[59] ), .B(new_n19923), .Y(new_n19924));
  INVx1_ASAP7_75t_L         g19668(.A(new_n19924), .Y(new_n19925));
  AOI22xp33_ASAP7_75t_L     g19669(.A1(new_n11656), .A2(\b[48] ), .B1(new_n11654), .B2(new_n7341), .Y(new_n19926));
  OAI221xp5_ASAP7_75t_L     g19670(.A1(new_n12364), .A2(new_n7316), .B1(new_n7033), .B2(new_n13003), .C(new_n19926), .Y(new_n19927));
  XNOR2x2_ASAP7_75t_L       g19671(.A(\a[62] ), .B(new_n19927), .Y(new_n19928));
  INVx1_ASAP7_75t_L         g19672(.A(new_n19928), .Y(new_n19929));
  NOR2xp33_ASAP7_75t_L      g19673(.A(new_n6220), .B(new_n12671), .Y(new_n19930));
  A2O1A1Ixp33_ASAP7_75t_L   g19674(.A1(new_n12669), .A2(\b[45] ), .B(new_n19930), .C(new_n5996), .Y(new_n19931));
  O2A1O1Ixp33_ASAP7_75t_L   g19675(.A1(new_n12353), .A2(new_n12355), .B(\b[45] ), .C(new_n19930), .Y(new_n19932));
  NAND2xp33_ASAP7_75t_L     g19676(.A(\a[44] ), .B(new_n19932), .Y(new_n19933));
  NAND2xp33_ASAP7_75t_L     g19677(.A(new_n19931), .B(new_n19933), .Y(new_n19934));
  XNOR2x2_ASAP7_75t_L       g19678(.A(new_n19756), .B(new_n19934), .Y(new_n19935));
  A2O1A1Ixp33_ASAP7_75t_L   g19679(.A1(new_n19845), .A2(new_n19752), .B(new_n19852), .C(new_n19935), .Y(new_n19936));
  O2A1O1Ixp33_ASAP7_75t_L   g19680(.A1(new_n12356), .A2(new_n6220), .B(new_n19844), .C(new_n19756), .Y(new_n19937));
  OR3x1_ASAP7_75t_L         g19681(.A(new_n19852), .B(new_n19937), .C(new_n19935), .Y(new_n19938));
  NAND3xp33_ASAP7_75t_L     g19682(.A(new_n19929), .B(new_n19936), .C(new_n19938), .Y(new_n19939));
  AO21x2_ASAP7_75t_L        g19683(.A1(new_n19936), .A2(new_n19938), .B(new_n19929), .Y(new_n19940));
  AND2x2_ASAP7_75t_L        g19684(.A(new_n19939), .B(new_n19940), .Y(new_n19941));
  NOR2xp33_ASAP7_75t_L      g19685(.A(new_n19941), .B(new_n19925), .Y(new_n19942));
  NAND2xp33_ASAP7_75t_L     g19686(.A(new_n19941), .B(new_n19925), .Y(new_n19943));
  INVx1_ASAP7_75t_L         g19687(.A(new_n19943), .Y(new_n19944));
  NOR2xp33_ASAP7_75t_L      g19688(.A(new_n19942), .B(new_n19944), .Y(new_n19945));
  INVx1_ASAP7_75t_L         g19689(.A(new_n19945), .Y(new_n19946));
  O2A1O1Ixp33_ASAP7_75t_L   g19690(.A1(new_n19858), .A2(new_n19855), .B(new_n19862), .C(new_n19946), .Y(new_n19947));
  INVx1_ASAP7_75t_L         g19691(.A(new_n19947), .Y(new_n19948));
  A2O1A1Ixp33_ASAP7_75t_L   g19692(.A1(new_n12669), .A2(\b[40] ), .B(new_n19457), .C(new_n5244), .Y(new_n19949));
  A2O1A1O1Ixp25_ASAP7_75t_L g19693(.A1(new_n19655), .A2(new_n19657), .B(new_n19660), .C(new_n19949), .D(new_n19756), .Y(new_n19950));
  O2A1O1Ixp33_ASAP7_75t_L   g19694(.A1(new_n19762), .A2(new_n19950), .B(new_n19854), .C(new_n19861), .Y(new_n19951));
  NAND2xp33_ASAP7_75t_L     g19695(.A(new_n19951), .B(new_n19946), .Y(new_n19952));
  AO21x2_ASAP7_75t_L        g19696(.A1(new_n19952), .A2(new_n19948), .B(new_n19921), .Y(new_n19953));
  NAND3xp33_ASAP7_75t_L     g19697(.A(new_n19948), .B(new_n19921), .C(new_n19952), .Y(new_n19954));
  AND2x2_ASAP7_75t_L        g19698(.A(new_n19954), .B(new_n19953), .Y(new_n19955));
  A2O1A1Ixp33_ASAP7_75t_L   g19699(.A1(new_n19867), .A2(new_n19840), .B(new_n19917), .C(new_n19955), .Y(new_n19956));
  INVx1_ASAP7_75t_L         g19700(.A(new_n19955), .Y(new_n19957));
  NAND3xp33_ASAP7_75t_L     g19701(.A(new_n19957), .B(new_n19868), .C(new_n19866), .Y(new_n19958));
  AND2x2_ASAP7_75t_L        g19702(.A(new_n19956), .B(new_n19958), .Y(new_n19959));
  INVx1_ASAP7_75t_L         g19703(.A(new_n19959), .Y(new_n19960));
  NAND2xp33_ASAP7_75t_L     g19704(.A(new_n19916), .B(new_n19960), .Y(new_n19961));
  INVx1_ASAP7_75t_L         g19705(.A(new_n19916), .Y(new_n19962));
  NAND2xp33_ASAP7_75t_L     g19706(.A(new_n19962), .B(new_n19959), .Y(new_n19963));
  AND2x2_ASAP7_75t_L        g19707(.A(new_n19963), .B(new_n19961), .Y(new_n19964));
  A2O1A1Ixp33_ASAP7_75t_L   g19708(.A1(new_n19913), .A2(new_n19836), .B(new_n19872), .C(new_n19964), .Y(new_n19965));
  INVx1_ASAP7_75t_L         g19709(.A(new_n19965), .Y(new_n19966));
  AOI211xp5_ASAP7_75t_L     g19710(.A1(new_n19913), .A2(new_n19836), .B(new_n19872), .C(new_n19964), .Y(new_n19967));
  OAI21xp33_ASAP7_75t_L     g19711(.A1(new_n19967), .A2(new_n19966), .B(new_n19912), .Y(new_n19968));
  OR3x1_ASAP7_75t_L         g19712(.A(new_n19966), .B(new_n19912), .C(new_n19967), .Y(new_n19969));
  AND2x2_ASAP7_75t_L        g19713(.A(new_n19968), .B(new_n19969), .Y(new_n19970));
  O2A1O1Ixp33_ASAP7_75t_L   g19714(.A1(new_n19793), .A2(new_n19799), .B(new_n19880), .C(new_n19885), .Y(new_n19971));
  NAND2xp33_ASAP7_75t_L     g19715(.A(new_n19971), .B(new_n19970), .Y(new_n19972));
  INVx1_ASAP7_75t_L         g19716(.A(new_n19881), .Y(new_n19973));
  INVx1_ASAP7_75t_L         g19717(.A(new_n19970), .Y(new_n19974));
  A2O1A1Ixp33_ASAP7_75t_L   g19718(.A1(new_n19884), .A2(new_n19879), .B(new_n19973), .C(new_n19974), .Y(new_n19975));
  AND2x2_ASAP7_75t_L        g19719(.A(new_n19972), .B(new_n19975), .Y(new_n19976));
  NAND2xp33_ASAP7_75t_L     g19720(.A(\b[63] ), .B(new_n6822), .Y(new_n19977));
  A2O1A1Ixp33_ASAP7_75t_L   g19721(.A1(new_n12607), .A2(new_n12603), .B(new_n7117), .C(new_n19977), .Y(new_n19978));
  AOI221xp5_ASAP7_75t_L     g19722(.A1(\b[61] ), .A2(new_n7124), .B1(\b[62] ), .B2(new_n6812), .C(new_n19978), .Y(new_n19979));
  XNOR2x2_ASAP7_75t_L       g19723(.A(new_n6816), .B(new_n19979), .Y(new_n19980));
  INVx1_ASAP7_75t_L         g19724(.A(new_n19980), .Y(new_n19981));
  XNOR2x2_ASAP7_75t_L       g19725(.A(new_n19981), .B(new_n19976), .Y(new_n19982));
  A2O1A1Ixp33_ASAP7_75t_L   g19726(.A1(new_n19891), .A2(new_n19832), .B(new_n19890), .C(new_n19982), .Y(new_n19983));
  OR3x1_ASAP7_75t_L         g19727(.A(new_n19982), .B(new_n19890), .C(new_n19892), .Y(new_n19984));
  AND2x2_ASAP7_75t_L        g19728(.A(new_n19983), .B(new_n19984), .Y(new_n19985));
  INVx1_ASAP7_75t_L         g19729(.A(new_n19985), .Y(new_n19986));
  O2A1O1Ixp33_ASAP7_75t_L   g19730(.A1(new_n19894), .A2(new_n19903), .B(new_n19901), .C(new_n19986), .Y(new_n19987));
  INVx1_ASAP7_75t_L         g19731(.A(new_n19987), .Y(new_n19988));
  OAI211xp5_ASAP7_75t_L     g19732(.A1(new_n19894), .A2(new_n19903), .B(new_n19986), .C(new_n19901), .Y(new_n19989));
  NAND2xp33_ASAP7_75t_L     g19733(.A(new_n19989), .B(new_n19988), .Y(new_n19990));
  XOR2x2_ASAP7_75t_L        g19734(.A(new_n19990), .B(new_n19909), .Y(\f[108] ));
  INVx1_ASAP7_75t_L         g19735(.A(new_n19909), .Y(new_n19992));
  A2O1A1Ixp33_ASAP7_75t_L   g19736(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n6819), .Y(new_n19993));
  AOI22xp33_ASAP7_75t_L     g19737(.A1(new_n6812), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n7124), .Y(new_n19994));
  NAND3xp33_ASAP7_75t_L     g19738(.A(new_n19993), .B(\a[47] ), .C(new_n19994), .Y(new_n19995));
  A2O1A1O1Ixp25_ASAP7_75t_L g19739(.A1(new_n13507), .A2(new_n13506), .B(new_n7117), .C(new_n19994), .D(\a[47] ), .Y(new_n19996));
  INVx1_ASAP7_75t_L         g19740(.A(new_n19996), .Y(new_n19997));
  AOI22xp33_ASAP7_75t_L     g19741(.A1(new_n19995), .A2(new_n19997), .B1(new_n19969), .B2(new_n19972), .Y(new_n19998));
  NAND2xp33_ASAP7_75t_L     g19742(.A(new_n19969), .B(new_n19972), .Y(new_n19999));
  NAND2xp33_ASAP7_75t_L     g19743(.A(new_n19995), .B(new_n19997), .Y(new_n20000));
  NOR2xp33_ASAP7_75t_L      g19744(.A(new_n20000), .B(new_n19999), .Y(new_n20001));
  NOR2xp33_ASAP7_75t_L      g19745(.A(new_n19998), .B(new_n20001), .Y(new_n20002));
  INVx1_ASAP7_75t_L         g19746(.A(new_n20002), .Y(new_n20003));
  NAND2xp33_ASAP7_75t_L     g19747(.A(\b[61] ), .B(new_n7659), .Y(new_n20004));
  OAI221xp5_ASAP7_75t_L     g19748(.A1(new_n11226), .A2(new_n8326), .B1(new_n7996), .B2(new_n11920), .C(new_n20004), .Y(new_n20005));
  AOI21xp33_ASAP7_75t_L     g19749(.A1(new_n7993), .A2(\b[59] ), .B(new_n20005), .Y(new_n20006));
  NAND2xp33_ASAP7_75t_L     g19750(.A(\a[50] ), .B(new_n20006), .Y(new_n20007));
  A2O1A1Ixp33_ASAP7_75t_L   g19751(.A1(\b[59] ), .A2(new_n7993), .B(new_n20005), .C(new_n7653), .Y(new_n20008));
  AOI22xp33_ASAP7_75t_L     g19752(.A1(new_n8645), .A2(\b[58] ), .B1(new_n8642), .B2(new_n10857), .Y(new_n20009));
  OAI221xp5_ASAP7_75t_L     g19753(.A1(new_n9322), .A2(new_n10488), .B1(new_n10178), .B2(new_n8965), .C(new_n20009), .Y(new_n20010));
  XNOR2x2_ASAP7_75t_L       g19754(.A(\a[53] ), .B(new_n20010), .Y(new_n20011));
  INVx1_ASAP7_75t_L         g19755(.A(new_n20011), .Y(new_n20012));
  AOI22xp33_ASAP7_75t_L     g19756(.A1(new_n10594), .A2(\b[52] ), .B1(new_n10591), .B2(new_n8577), .Y(new_n20013));
  OAI221xp5_ASAP7_75t_L     g19757(.A1(new_n11335), .A2(new_n8249), .B1(new_n8228), .B2(new_n11330), .C(new_n20013), .Y(new_n20014));
  XNOR2x2_ASAP7_75t_L       g19758(.A(\a[59] ), .B(new_n20014), .Y(new_n20015));
  NAND2xp33_ASAP7_75t_L     g19759(.A(new_n19936), .B(new_n19939), .Y(new_n20016));
  NOR2xp33_ASAP7_75t_L      g19760(.A(new_n6756), .B(new_n12671), .Y(new_n20017));
  INVx1_ASAP7_75t_L         g19761(.A(new_n19931), .Y(new_n20018));
  A2O1A1O1Ixp25_ASAP7_75t_L g19762(.A1(new_n12669), .A2(\b[43] ), .B(new_n19751), .C(new_n19933), .D(new_n20018), .Y(new_n20019));
  A2O1A1Ixp33_ASAP7_75t_L   g19763(.A1(new_n12669), .A2(\b[46] ), .B(new_n20017), .C(new_n20019), .Y(new_n20020));
  O2A1O1Ixp33_ASAP7_75t_L   g19764(.A1(new_n12353), .A2(new_n12355), .B(\b[46] ), .C(new_n20017), .Y(new_n20021));
  INVx1_ASAP7_75t_L         g19765(.A(new_n20021), .Y(new_n20022));
  A2O1A1Ixp33_ASAP7_75t_L   g19766(.A1(new_n12669), .A2(\b[43] ), .B(new_n19751), .C(new_n19933), .Y(new_n20023));
  O2A1O1Ixp33_ASAP7_75t_L   g19767(.A1(new_n19932), .A2(\a[44] ), .B(new_n20023), .C(new_n20022), .Y(new_n20024));
  INVx1_ASAP7_75t_L         g19768(.A(new_n20024), .Y(new_n20025));
  NAND2xp33_ASAP7_75t_L     g19769(.A(new_n20020), .B(new_n20025), .Y(new_n20026));
  NAND2xp33_ASAP7_75t_L     g19770(.A(new_n11654), .B(new_n7914), .Y(new_n20027));
  OAI221xp5_ASAP7_75t_L     g19771(.A1(new_n12023), .A2(new_n7907), .B1(new_n7333), .B2(new_n12364), .C(new_n20027), .Y(new_n20028));
  AOI21xp33_ASAP7_75t_L     g19772(.A1(new_n12021), .A2(\b[47] ), .B(new_n20028), .Y(new_n20029));
  NAND2xp33_ASAP7_75t_L     g19773(.A(\a[62] ), .B(new_n20029), .Y(new_n20030));
  A2O1A1Ixp33_ASAP7_75t_L   g19774(.A1(\b[47] ), .A2(new_n12021), .B(new_n20028), .C(new_n11651), .Y(new_n20031));
  AND2x2_ASAP7_75t_L        g19775(.A(new_n20031), .B(new_n20030), .Y(new_n20032));
  NAND2xp33_ASAP7_75t_L     g19776(.A(new_n20026), .B(new_n20032), .Y(new_n20033));
  NOR2xp33_ASAP7_75t_L      g19777(.A(new_n20026), .B(new_n20032), .Y(new_n20034));
  INVx1_ASAP7_75t_L         g19778(.A(new_n20034), .Y(new_n20035));
  AND2x2_ASAP7_75t_L        g19779(.A(new_n20033), .B(new_n20035), .Y(new_n20036));
  XOR2x2_ASAP7_75t_L        g19780(.A(new_n20016), .B(new_n20036), .Y(new_n20037));
  XNOR2x2_ASAP7_75t_L       g19781(.A(new_n20015), .B(new_n20037), .Y(new_n20038));
  A2O1A1Ixp33_ASAP7_75t_L   g19782(.A1(new_n19941), .A2(new_n19925), .B(new_n19947), .C(new_n20038), .Y(new_n20039));
  A2O1A1Ixp33_ASAP7_75t_L   g19783(.A1(new_n19862), .A2(new_n19857), .B(new_n19942), .C(new_n19943), .Y(new_n20040));
  NOR2xp33_ASAP7_75t_L      g19784(.A(new_n20040), .B(new_n20038), .Y(new_n20041));
  INVx1_ASAP7_75t_L         g19785(.A(new_n20041), .Y(new_n20042));
  AOI22xp33_ASAP7_75t_L     g19786(.A1(new_n9623), .A2(\b[55] ), .B1(new_n9620), .B2(new_n9542), .Y(new_n20043));
  OAI221xp5_ASAP7_75t_L     g19787(.A1(new_n10280), .A2(new_n9199), .B1(new_n8882), .B2(new_n12010), .C(new_n20043), .Y(new_n20044));
  XNOR2x2_ASAP7_75t_L       g19788(.A(\a[56] ), .B(new_n20044), .Y(new_n20045));
  NAND3xp33_ASAP7_75t_L     g19789(.A(new_n20042), .B(new_n20039), .C(new_n20045), .Y(new_n20046));
  INVx1_ASAP7_75t_L         g19790(.A(new_n20046), .Y(new_n20047));
  AOI21xp33_ASAP7_75t_L     g19791(.A1(new_n20042), .A2(new_n20039), .B(new_n20045), .Y(new_n20048));
  NOR2xp33_ASAP7_75t_L      g19792(.A(new_n20048), .B(new_n20047), .Y(new_n20049));
  A2O1A1O1Ixp25_ASAP7_75t_L g19793(.A1(new_n19868), .A2(new_n19866), .B(new_n19957), .C(new_n19954), .D(new_n20049), .Y(new_n20050));
  INVx1_ASAP7_75t_L         g19794(.A(new_n20050), .Y(new_n20051));
  NAND3xp33_ASAP7_75t_L     g19795(.A(new_n20049), .B(new_n19956), .C(new_n19954), .Y(new_n20052));
  AO21x2_ASAP7_75t_L        g19796(.A1(new_n20052), .A2(new_n20051), .B(new_n20012), .Y(new_n20053));
  NAND3xp33_ASAP7_75t_L     g19797(.A(new_n20051), .B(new_n20012), .C(new_n20052), .Y(new_n20054));
  AND2x2_ASAP7_75t_L        g19798(.A(new_n20054), .B(new_n20053), .Y(new_n20055));
  INVx1_ASAP7_75t_L         g19799(.A(new_n20055), .Y(new_n20056));
  O2A1O1Ixp33_ASAP7_75t_L   g19800(.A1(new_n19916), .A2(new_n19960), .B(new_n19965), .C(new_n20056), .Y(new_n20057));
  INVx1_ASAP7_75t_L         g19801(.A(new_n19963), .Y(new_n20058));
  A2O1A1O1Ixp25_ASAP7_75t_L g19802(.A1(new_n19836), .A2(new_n19874), .B(new_n19872), .C(new_n19961), .D(new_n20058), .Y(new_n20059));
  NAND2xp33_ASAP7_75t_L     g19803(.A(new_n20059), .B(new_n20056), .Y(new_n20060));
  INVx1_ASAP7_75t_L         g19804(.A(new_n20060), .Y(new_n20061));
  NOR2xp33_ASAP7_75t_L      g19805(.A(new_n20057), .B(new_n20061), .Y(new_n20062));
  AOI21xp33_ASAP7_75t_L     g19806(.A1(new_n20008), .A2(new_n20007), .B(new_n20062), .Y(new_n20063));
  NAND2xp33_ASAP7_75t_L     g19807(.A(new_n20008), .B(new_n20007), .Y(new_n20064));
  INVx1_ASAP7_75t_L         g19808(.A(new_n20062), .Y(new_n20065));
  NOR2xp33_ASAP7_75t_L      g19809(.A(new_n20064), .B(new_n20065), .Y(new_n20066));
  NOR2xp33_ASAP7_75t_L      g19810(.A(new_n20063), .B(new_n20066), .Y(new_n20067));
  INVx1_ASAP7_75t_L         g19811(.A(new_n20067), .Y(new_n20068));
  NOR2xp33_ASAP7_75t_L      g19812(.A(new_n20068), .B(new_n20003), .Y(new_n20069));
  INVx1_ASAP7_75t_L         g19813(.A(new_n20069), .Y(new_n20070));
  NAND2xp33_ASAP7_75t_L     g19814(.A(new_n20068), .B(new_n20003), .Y(new_n20071));
  AND2x2_ASAP7_75t_L        g19815(.A(new_n20071), .B(new_n20070), .Y(new_n20072));
  INVx1_ASAP7_75t_L         g19816(.A(new_n19976), .Y(new_n20073));
  OA21x2_ASAP7_75t_L        g19817(.A1(new_n20073), .A2(new_n19980), .B(new_n19984), .Y(new_n20074));
  AND2x2_ASAP7_75t_L        g19818(.A(new_n20072), .B(new_n20074), .Y(new_n20075));
  O2A1O1Ixp33_ASAP7_75t_L   g19819(.A1(new_n20073), .A2(new_n19980), .B(new_n19984), .C(new_n20072), .Y(new_n20076));
  NOR2xp33_ASAP7_75t_L      g19820(.A(new_n20076), .B(new_n20075), .Y(new_n20077));
  A2O1A1Ixp33_ASAP7_75t_L   g19821(.A1(new_n19992), .A2(new_n19989), .B(new_n19987), .C(new_n20077), .Y(new_n20078));
  INVx1_ASAP7_75t_L         g19822(.A(new_n20078), .Y(new_n20079));
  NAND2xp33_ASAP7_75t_L     g19823(.A(new_n19905), .B(new_n19829), .Y(new_n20080));
  A2O1A1Ixp33_ASAP7_75t_L   g19824(.A1(new_n19824), .A2(new_n19821), .B(new_n19820), .C(new_n19906), .Y(new_n20081));
  A2O1A1Ixp33_ASAP7_75t_L   g19825(.A1(new_n20081), .A2(new_n20080), .B(new_n19990), .C(new_n19988), .Y(new_n20082));
  NOR2xp33_ASAP7_75t_L      g19826(.A(new_n20077), .B(new_n20082), .Y(new_n20083));
  NOR2xp33_ASAP7_75t_L      g19827(.A(new_n20083), .B(new_n20079), .Y(\f[109] ));
  AOI22xp33_ASAP7_75t_L     g19828(.A1(new_n7659), .A2(\b[62] ), .B1(new_n7656), .B2(new_n12280), .Y(new_n20085));
  OAI221xp5_ASAP7_75t_L     g19829(.A1(new_n8326), .A2(new_n11911), .B1(new_n11226), .B2(new_n7994), .C(new_n20085), .Y(new_n20086));
  XNOR2x2_ASAP7_75t_L       g19830(.A(\a[50] ), .B(new_n20086), .Y(new_n20087));
  AOI22xp33_ASAP7_75t_L     g19831(.A1(new_n9623), .A2(\b[56] ), .B1(new_n9620), .B2(new_n10185), .Y(new_n20088));
  OAI221xp5_ASAP7_75t_L     g19832(.A1(new_n10280), .A2(new_n9534), .B1(new_n9199), .B2(new_n12010), .C(new_n20088), .Y(new_n20089));
  XNOR2x2_ASAP7_75t_L       g19833(.A(\a[56] ), .B(new_n20089), .Y(new_n20090));
  INVx1_ASAP7_75t_L         g19834(.A(new_n20036), .Y(new_n20091));
  INVx1_ASAP7_75t_L         g19835(.A(new_n20015), .Y(new_n20092));
  NAND2xp33_ASAP7_75t_L     g19836(.A(new_n20092), .B(new_n20037), .Y(new_n20093));
  AOI22xp33_ASAP7_75t_L     g19837(.A1(new_n10594), .A2(\b[53] ), .B1(new_n10591), .B2(new_n8889), .Y(new_n20094));
  OAI221xp5_ASAP7_75t_L     g19838(.A1(new_n11335), .A2(new_n8569), .B1(new_n8249), .B2(new_n11330), .C(new_n20094), .Y(new_n20095));
  XNOR2x2_ASAP7_75t_L       g19839(.A(\a[59] ), .B(new_n20095), .Y(new_n20096));
  INVx1_ASAP7_75t_L         g19840(.A(new_n20096), .Y(new_n20097));
  AOI22xp33_ASAP7_75t_L     g19841(.A1(new_n11656), .A2(\b[50] ), .B1(new_n11654), .B2(new_n8235), .Y(new_n20098));
  OAI221xp5_ASAP7_75t_L     g19842(.A1(new_n12364), .A2(new_n7907), .B1(new_n7333), .B2(new_n13003), .C(new_n20098), .Y(new_n20099));
  XNOR2x2_ASAP7_75t_L       g19843(.A(\a[62] ), .B(new_n20099), .Y(new_n20100));
  A2O1A1O1Ixp25_ASAP7_75t_L g19844(.A1(new_n19756), .A2(new_n19933), .B(new_n20018), .C(new_n20021), .D(new_n20034), .Y(new_n20101));
  NOR2xp33_ASAP7_75t_L      g19845(.A(new_n7033), .B(new_n12671), .Y(new_n20102));
  A2O1A1Ixp33_ASAP7_75t_L   g19846(.A1(\b[47] ), .A2(new_n12669), .B(new_n20102), .C(new_n20021), .Y(new_n20103));
  O2A1O1Ixp33_ASAP7_75t_L   g19847(.A1(new_n12353), .A2(new_n12355), .B(\b[47] ), .C(new_n20102), .Y(new_n20104));
  A2O1A1Ixp33_ASAP7_75t_L   g19848(.A1(new_n12669), .A2(\b[46] ), .B(new_n20017), .C(new_n20104), .Y(new_n20105));
  NAND2xp33_ASAP7_75t_L     g19849(.A(new_n20105), .B(new_n20103), .Y(new_n20106));
  XOR2x2_ASAP7_75t_L        g19850(.A(new_n20106), .B(new_n20101), .Y(new_n20107));
  INVx1_ASAP7_75t_L         g19851(.A(new_n20107), .Y(new_n20108));
  NOR2xp33_ASAP7_75t_L      g19852(.A(new_n20100), .B(new_n20108), .Y(new_n20109));
  INVx1_ASAP7_75t_L         g19853(.A(new_n20109), .Y(new_n20110));
  NAND2xp33_ASAP7_75t_L     g19854(.A(new_n20100), .B(new_n20108), .Y(new_n20111));
  NAND3xp33_ASAP7_75t_L     g19855(.A(new_n20110), .B(new_n20097), .C(new_n20111), .Y(new_n20112));
  AO21x2_ASAP7_75t_L        g19856(.A1(new_n20111), .A2(new_n20110), .B(new_n20097), .Y(new_n20113));
  AND2x2_ASAP7_75t_L        g19857(.A(new_n20112), .B(new_n20113), .Y(new_n20114));
  INVx1_ASAP7_75t_L         g19858(.A(new_n20114), .Y(new_n20115));
  A2O1A1O1Ixp25_ASAP7_75t_L g19859(.A1(new_n19939), .A2(new_n19936), .B(new_n20091), .C(new_n20093), .D(new_n20115), .Y(new_n20116));
  A2O1A1Ixp33_ASAP7_75t_L   g19860(.A1(new_n19939), .A2(new_n19936), .B(new_n20091), .C(new_n20093), .Y(new_n20117));
  NOR2xp33_ASAP7_75t_L      g19861(.A(new_n20117), .B(new_n20114), .Y(new_n20118));
  OR3x1_ASAP7_75t_L         g19862(.A(new_n20116), .B(new_n20090), .C(new_n20118), .Y(new_n20119));
  OAI21xp33_ASAP7_75t_L     g19863(.A1(new_n20118), .A2(new_n20116), .B(new_n20090), .Y(new_n20120));
  AND2x2_ASAP7_75t_L        g19864(.A(new_n20120), .B(new_n20119), .Y(new_n20121));
  NAND2xp33_ASAP7_75t_L     g19865(.A(new_n20042), .B(new_n20046), .Y(new_n20122));
  INVx1_ASAP7_75t_L         g19866(.A(new_n20122), .Y(new_n20123));
  NAND2xp33_ASAP7_75t_L     g19867(.A(new_n20123), .B(new_n20121), .Y(new_n20124));
  O2A1O1Ixp33_ASAP7_75t_L   g19868(.A1(new_n20040), .A2(new_n20038), .B(new_n20046), .C(new_n20121), .Y(new_n20125));
  INVx1_ASAP7_75t_L         g19869(.A(new_n20125), .Y(new_n20126));
  AOI22xp33_ASAP7_75t_L     g19870(.A1(new_n8645), .A2(\b[59] ), .B1(new_n8642), .B2(new_n10887), .Y(new_n20127));
  OAI221xp5_ASAP7_75t_L     g19871(.A1(new_n9322), .A2(new_n10848), .B1(new_n10488), .B2(new_n8965), .C(new_n20127), .Y(new_n20128));
  XNOR2x2_ASAP7_75t_L       g19872(.A(\a[53] ), .B(new_n20128), .Y(new_n20129));
  NAND3xp33_ASAP7_75t_L     g19873(.A(new_n20126), .B(new_n20124), .C(new_n20129), .Y(new_n20130));
  AO21x2_ASAP7_75t_L        g19874(.A1(new_n20124), .A2(new_n20126), .B(new_n20129), .Y(new_n20131));
  AND2x2_ASAP7_75t_L        g19875(.A(new_n20130), .B(new_n20131), .Y(new_n20132));
  INVx1_ASAP7_75t_L         g19876(.A(new_n20132), .Y(new_n20133));
  A2O1A1Ixp33_ASAP7_75t_L   g19877(.A1(new_n20052), .A2(new_n20012), .B(new_n20050), .C(new_n20133), .Y(new_n20134));
  NAND3xp33_ASAP7_75t_L     g19878(.A(new_n20132), .B(new_n20054), .C(new_n20051), .Y(new_n20135));
  NAND3xp33_ASAP7_75t_L     g19879(.A(new_n20134), .B(new_n20087), .C(new_n20135), .Y(new_n20136));
  AO21x2_ASAP7_75t_L        g19880(.A1(new_n20135), .A2(new_n20134), .B(new_n20087), .Y(new_n20137));
  NAND2xp33_ASAP7_75t_L     g19881(.A(new_n20136), .B(new_n20137), .Y(new_n20138));
  INVx1_ASAP7_75t_L         g19882(.A(new_n20066), .Y(new_n20139));
  A2O1A1Ixp33_ASAP7_75t_L   g19883(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n6819), .Y(new_n20140));
  A2O1A1Ixp33_ASAP7_75t_L   g19884(.A1(new_n20140), .A2(new_n7115), .B(new_n12599), .C(\a[47] ), .Y(new_n20141));
  O2A1O1Ixp33_ASAP7_75t_L   g19885(.A1(new_n7117), .A2(new_n13934), .B(new_n7115), .C(new_n12599), .Y(new_n20142));
  NAND2xp33_ASAP7_75t_L     g19886(.A(new_n6816), .B(new_n20142), .Y(new_n20143));
  AND2x2_ASAP7_75t_L        g19887(.A(new_n20143), .B(new_n20141), .Y(new_n20144));
  INVx1_ASAP7_75t_L         g19888(.A(new_n20144), .Y(new_n20145));
  NAND3xp33_ASAP7_75t_L     g19889(.A(new_n20139), .B(new_n20060), .C(new_n20145), .Y(new_n20146));
  A2O1A1Ixp33_ASAP7_75t_L   g19890(.A1(new_n20056), .A2(new_n20059), .B(new_n20066), .C(new_n20144), .Y(new_n20147));
  NAND2xp33_ASAP7_75t_L     g19891(.A(new_n20147), .B(new_n20146), .Y(new_n20148));
  NAND2xp33_ASAP7_75t_L     g19892(.A(new_n20138), .B(new_n20148), .Y(new_n20149));
  NAND4xp25_ASAP7_75t_L     g19893(.A(new_n20146), .B(new_n20136), .C(new_n20137), .D(new_n20147), .Y(new_n20150));
  AND2x2_ASAP7_75t_L        g19894(.A(new_n20150), .B(new_n20149), .Y(new_n20151));
  INVx1_ASAP7_75t_L         g19895(.A(new_n20151), .Y(new_n20152));
  O2A1O1Ixp33_ASAP7_75t_L   g19896(.A1(new_n19999), .A2(new_n20000), .B(new_n20070), .C(new_n20152), .Y(new_n20153));
  NOR2xp33_ASAP7_75t_L      g19897(.A(new_n20001), .B(new_n20069), .Y(new_n20154));
  NAND2xp33_ASAP7_75t_L     g19898(.A(new_n20152), .B(new_n20154), .Y(new_n20155));
  INVx1_ASAP7_75t_L         g19899(.A(new_n20155), .Y(new_n20156));
  NOR2xp33_ASAP7_75t_L      g19900(.A(new_n20153), .B(new_n20156), .Y(new_n20157));
  A2O1A1Ixp33_ASAP7_75t_L   g19901(.A1(new_n20082), .A2(new_n20077), .B(new_n20076), .C(new_n20157), .Y(new_n20158));
  INVx1_ASAP7_75t_L         g19902(.A(new_n20158), .Y(new_n20159));
  NOR3xp33_ASAP7_75t_L      g19903(.A(new_n20079), .B(new_n20157), .C(new_n20076), .Y(new_n20160));
  NOR2xp33_ASAP7_75t_L      g19904(.A(new_n20159), .B(new_n20160), .Y(\f[110] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g19905(.A1(new_n19989), .A2(new_n19992), .B(new_n19987), .C(new_n20077), .D(new_n20076), .Y(new_n20162));
  A2O1A1Ixp33_ASAP7_75t_L   g19906(.A1(new_n19956), .A2(new_n19954), .B(new_n20049), .C(new_n20054), .Y(new_n20163));
  AOI22xp33_ASAP7_75t_L     g19907(.A1(new_n8645), .A2(\b[60] ), .B1(new_n8642), .B2(new_n11234), .Y(new_n20164));
  OAI221xp5_ASAP7_75t_L     g19908(.A1(new_n9322), .A2(new_n10881), .B1(new_n10848), .B2(new_n8965), .C(new_n20164), .Y(new_n20165));
  XNOR2x2_ASAP7_75t_L       g19909(.A(\a[53] ), .B(new_n20165), .Y(new_n20166));
  NAND2xp33_ASAP7_75t_L     g19910(.A(new_n20016), .B(new_n20036), .Y(new_n20167));
  AOI22xp33_ASAP7_75t_L     g19911(.A1(new_n9623), .A2(\b[57] ), .B1(new_n9620), .B2(new_n10495), .Y(new_n20168));
  OAI221xp5_ASAP7_75t_L     g19912(.A1(new_n10280), .A2(new_n10178), .B1(new_n9534), .B2(new_n12010), .C(new_n20168), .Y(new_n20169));
  XNOR2x2_ASAP7_75t_L       g19913(.A(new_n9610), .B(new_n20169), .Y(new_n20170));
  AOI22xp33_ASAP7_75t_L     g19914(.A1(new_n11656), .A2(\b[51] ), .B1(new_n11654), .B2(new_n8257), .Y(new_n20171));
  OAI221xp5_ASAP7_75t_L     g19915(.A1(new_n12364), .A2(new_n8228), .B1(new_n7907), .B2(new_n13003), .C(new_n20171), .Y(new_n20172));
  XNOR2x2_ASAP7_75t_L       g19916(.A(\a[62] ), .B(new_n20172), .Y(new_n20173));
  NOR2xp33_ASAP7_75t_L      g19917(.A(new_n7316), .B(new_n12671), .Y(new_n20174));
  INVx1_ASAP7_75t_L         g19918(.A(new_n20174), .Y(new_n20175));
  A2O1A1Ixp33_ASAP7_75t_L   g19919(.A1(new_n12669), .A2(\b[47] ), .B(new_n20102), .C(\a[47] ), .Y(new_n20176));
  INVx1_ASAP7_75t_L         g19920(.A(new_n20104), .Y(new_n20177));
  NOR2xp33_ASAP7_75t_L      g19921(.A(\a[47] ), .B(new_n20177), .Y(new_n20178));
  INVx1_ASAP7_75t_L         g19922(.A(new_n20178), .Y(new_n20179));
  AND2x2_ASAP7_75t_L        g19923(.A(new_n20176), .B(new_n20179), .Y(new_n20180));
  O2A1O1Ixp33_ASAP7_75t_L   g19924(.A1(new_n7333), .A2(new_n12356), .B(new_n20175), .C(new_n20180), .Y(new_n20181));
  O2A1O1Ixp33_ASAP7_75t_L   g19925(.A1(new_n12353), .A2(new_n12355), .B(\b[48] ), .C(new_n20174), .Y(new_n20182));
  AND3x1_ASAP7_75t_L        g19926(.A(new_n20179), .B(new_n20176), .C(new_n20182), .Y(new_n20183));
  NOR2xp33_ASAP7_75t_L      g19927(.A(new_n20183), .B(new_n20181), .Y(new_n20184));
  XNOR2x2_ASAP7_75t_L       g19928(.A(new_n20184), .B(new_n20173), .Y(new_n20185));
  INVx1_ASAP7_75t_L         g19929(.A(new_n20101), .Y(new_n20186));
  A2O1A1O1Ixp25_ASAP7_75t_L g19930(.A1(new_n12669), .A2(\b[46] ), .B(new_n20017), .C(new_n20104), .D(new_n20186), .Y(new_n20187));
  A2O1A1O1Ixp25_ASAP7_75t_L g19931(.A1(new_n12669), .A2(\b[47] ), .B(new_n20102), .C(new_n20021), .D(new_n20187), .Y(new_n20188));
  XNOR2x2_ASAP7_75t_L       g19932(.A(new_n20185), .B(new_n20188), .Y(new_n20189));
  AOI22xp33_ASAP7_75t_L     g19933(.A1(new_n10594), .A2(\b[54] ), .B1(new_n10591), .B2(new_n9208), .Y(new_n20190));
  OAI221xp5_ASAP7_75t_L     g19934(.A1(new_n11335), .A2(new_n8882), .B1(new_n8569), .B2(new_n11330), .C(new_n20190), .Y(new_n20191));
  XNOR2x2_ASAP7_75t_L       g19935(.A(\a[59] ), .B(new_n20191), .Y(new_n20192));
  XNOR2x2_ASAP7_75t_L       g19936(.A(new_n20192), .B(new_n20189), .Y(new_n20193));
  O2A1O1Ixp33_ASAP7_75t_L   g19937(.A1(new_n20100), .A2(new_n20108), .B(new_n20112), .C(new_n20193), .Y(new_n20194));
  AND3x1_ASAP7_75t_L        g19938(.A(new_n20193), .B(new_n20112), .C(new_n20110), .Y(new_n20195));
  NOR2xp33_ASAP7_75t_L      g19939(.A(new_n20194), .B(new_n20195), .Y(new_n20196));
  XOR2x2_ASAP7_75t_L        g19940(.A(new_n20170), .B(new_n20196), .Y(new_n20197));
  INVx1_ASAP7_75t_L         g19941(.A(new_n20197), .Y(new_n20198));
  A2O1A1O1Ixp25_ASAP7_75t_L g19942(.A1(new_n20093), .A2(new_n20167), .B(new_n20115), .C(new_n20119), .D(new_n20198), .Y(new_n20199));
  A2O1A1Ixp33_ASAP7_75t_L   g19943(.A1(new_n20093), .A2(new_n20167), .B(new_n20115), .C(new_n20119), .Y(new_n20200));
  NOR2xp33_ASAP7_75t_L      g19944(.A(new_n20197), .B(new_n20200), .Y(new_n20201));
  OAI21xp33_ASAP7_75t_L     g19945(.A1(new_n20201), .A2(new_n20199), .B(new_n20166), .Y(new_n20202));
  INVx1_ASAP7_75t_L         g19946(.A(new_n20166), .Y(new_n20203));
  NOR2xp33_ASAP7_75t_L      g19947(.A(new_n20201), .B(new_n20199), .Y(new_n20204));
  NAND2xp33_ASAP7_75t_L     g19948(.A(new_n20203), .B(new_n20204), .Y(new_n20205));
  AND2x2_ASAP7_75t_L        g19949(.A(new_n20202), .B(new_n20205), .Y(new_n20206));
  AND3x1_ASAP7_75t_L        g19950(.A(new_n20206), .B(new_n20130), .C(new_n20126), .Y(new_n20207));
  O2A1O1Ixp33_ASAP7_75t_L   g19951(.A1(new_n20121), .A2(new_n20123), .B(new_n20130), .C(new_n20206), .Y(new_n20208));
  NOR2xp33_ASAP7_75t_L      g19952(.A(new_n20208), .B(new_n20207), .Y(new_n20209));
  NAND2xp33_ASAP7_75t_L     g19953(.A(\b[63] ), .B(new_n7659), .Y(new_n20210));
  A2O1A1Ixp33_ASAP7_75t_L   g19954(.A1(new_n12607), .A2(new_n12603), .B(new_n7996), .C(new_n20210), .Y(new_n20211));
  AOI221xp5_ASAP7_75t_L     g19955(.A1(\b[61] ), .A2(new_n7993), .B1(\b[62] ), .B2(new_n7649), .C(new_n20211), .Y(new_n20212));
  XNOR2x2_ASAP7_75t_L       g19956(.A(new_n7653), .B(new_n20212), .Y(new_n20213));
  INVx1_ASAP7_75t_L         g19957(.A(new_n20213), .Y(new_n20214));
  XNOR2x2_ASAP7_75t_L       g19958(.A(new_n20214), .B(new_n20209), .Y(new_n20215));
  INVx1_ASAP7_75t_L         g19959(.A(new_n20215), .Y(new_n20216));
  O2A1O1Ixp33_ASAP7_75t_L   g19960(.A1(new_n20133), .A2(new_n20163), .B(new_n20136), .C(new_n20216), .Y(new_n20217));
  AND3x1_ASAP7_75t_L        g19961(.A(new_n20216), .B(new_n20136), .C(new_n20135), .Y(new_n20218));
  NOR2xp33_ASAP7_75t_L      g19962(.A(new_n20217), .B(new_n20218), .Y(new_n20219));
  O2A1O1Ixp33_ASAP7_75t_L   g19963(.A1(new_n20138), .A2(new_n20148), .B(new_n20147), .C(new_n20219), .Y(new_n20220));
  INVx1_ASAP7_75t_L         g19964(.A(new_n20219), .Y(new_n20221));
  A2O1A1Ixp33_ASAP7_75t_L   g19965(.A1(new_n20139), .A2(new_n20060), .B(new_n20145), .C(new_n20150), .Y(new_n20222));
  NOR2xp33_ASAP7_75t_L      g19966(.A(new_n20222), .B(new_n20221), .Y(new_n20223));
  NOR2xp33_ASAP7_75t_L      g19967(.A(new_n20220), .B(new_n20223), .Y(new_n20224));
  INVx1_ASAP7_75t_L         g19968(.A(new_n20224), .Y(new_n20225));
  O2A1O1Ixp33_ASAP7_75t_L   g19969(.A1(new_n20153), .A2(new_n20162), .B(new_n20155), .C(new_n20225), .Y(new_n20226));
  NOR3xp33_ASAP7_75t_L      g19970(.A(new_n20159), .B(new_n20224), .C(new_n20156), .Y(new_n20227));
  NOR2xp33_ASAP7_75t_L      g19971(.A(new_n20226), .B(new_n20227), .Y(\f[111] ));
  INVx1_ASAP7_75t_L         g19972(.A(new_n20223), .Y(new_n20229));
  AOI21xp33_ASAP7_75t_L     g19973(.A1(new_n20214), .A2(new_n20209), .B(new_n20218), .Y(new_n20230));
  NAND2xp33_ASAP7_75t_L     g19974(.A(\b[61] ), .B(new_n8645), .Y(new_n20231));
  OAI221xp5_ASAP7_75t_L     g19975(.A1(new_n11226), .A2(new_n9322), .B1(new_n8967), .B2(new_n11920), .C(new_n20231), .Y(new_n20232));
  AOI21xp33_ASAP7_75t_L     g19976(.A1(new_n8964), .A2(\b[59] ), .B(new_n20232), .Y(new_n20233));
  NAND2xp33_ASAP7_75t_L     g19977(.A(\a[53] ), .B(new_n20233), .Y(new_n20234));
  A2O1A1Ixp33_ASAP7_75t_L   g19978(.A1(\b[59] ), .A2(new_n8964), .B(new_n20232), .C(new_n8639), .Y(new_n20235));
  AND2x2_ASAP7_75t_L        g19979(.A(new_n20235), .B(new_n20234), .Y(new_n20236));
  AOI22xp33_ASAP7_75t_L     g19980(.A1(new_n9623), .A2(\b[58] ), .B1(new_n9620), .B2(new_n10857), .Y(new_n20237));
  OAI221xp5_ASAP7_75t_L     g19981(.A1(new_n10280), .A2(new_n10488), .B1(new_n10178), .B2(new_n12010), .C(new_n20237), .Y(new_n20238));
  XNOR2x2_ASAP7_75t_L       g19982(.A(\a[56] ), .B(new_n20238), .Y(new_n20239));
  NOR2xp33_ASAP7_75t_L      g19983(.A(new_n20192), .B(new_n20189), .Y(new_n20240));
  AOI22xp33_ASAP7_75t_L     g19984(.A1(new_n10594), .A2(\b[55] ), .B1(new_n10591), .B2(new_n9542), .Y(new_n20241));
  OAI221xp5_ASAP7_75t_L     g19985(.A1(new_n11335), .A2(new_n9199), .B1(new_n8882), .B2(new_n11330), .C(new_n20241), .Y(new_n20242));
  XNOR2x2_ASAP7_75t_L       g19986(.A(\a[59] ), .B(new_n20242), .Y(new_n20243));
  INVx1_ASAP7_75t_L         g19987(.A(new_n20173), .Y(new_n20244));
  MAJIxp5_ASAP7_75t_L       g19988(.A(new_n20188), .B(new_n20244), .C(new_n20184), .Y(new_n20245));
  NOR2xp33_ASAP7_75t_L      g19989(.A(new_n7333), .B(new_n12671), .Y(new_n20246));
  O2A1O1Ixp33_ASAP7_75t_L   g19990(.A1(new_n12353), .A2(new_n12355), .B(\b[49] ), .C(new_n20246), .Y(new_n20247));
  INVx1_ASAP7_75t_L         g19991(.A(new_n20247), .Y(new_n20248));
  A2O1A1Ixp33_ASAP7_75t_L   g19992(.A1(new_n12669), .A2(\b[47] ), .B(new_n20102), .C(new_n6816), .Y(new_n20249));
  A2O1A1O1Ixp25_ASAP7_75t_L g19993(.A1(new_n20176), .A2(new_n20179), .B(new_n20182), .C(new_n20249), .D(new_n20248), .Y(new_n20250));
  INVx1_ASAP7_75t_L         g19994(.A(new_n20246), .Y(new_n20251));
  A2O1A1Ixp33_ASAP7_75t_L   g19995(.A1(new_n20179), .A2(new_n20176), .B(new_n20182), .C(new_n20249), .Y(new_n20252));
  O2A1O1Ixp33_ASAP7_75t_L   g19996(.A1(new_n7907), .A2(new_n12356), .B(new_n20251), .C(new_n20252), .Y(new_n20253));
  NOR2xp33_ASAP7_75t_L      g19997(.A(new_n20250), .B(new_n20253), .Y(new_n20254));
  INVx1_ASAP7_75t_L         g19998(.A(new_n20254), .Y(new_n20255));
  AOI22xp33_ASAP7_75t_L     g19999(.A1(new_n11647), .A2(\b[51] ), .B1(\b[52] ), .B2(new_n11656), .Y(new_n20256));
  OAI221xp5_ASAP7_75t_L     g20000(.A1(new_n13003), .A2(new_n8228), .B1(new_n12022), .B2(new_n10519), .C(new_n20256), .Y(new_n20257));
  XNOR2x2_ASAP7_75t_L       g20001(.A(\a[62] ), .B(new_n20257), .Y(new_n20258));
  NOR2xp33_ASAP7_75t_L      g20002(.A(new_n20255), .B(new_n20258), .Y(new_n20259));
  INVx1_ASAP7_75t_L         g20003(.A(new_n20259), .Y(new_n20260));
  NAND2xp33_ASAP7_75t_L     g20004(.A(new_n20255), .B(new_n20258), .Y(new_n20261));
  NAND2xp33_ASAP7_75t_L     g20005(.A(new_n20261), .B(new_n20260), .Y(new_n20262));
  XOR2x2_ASAP7_75t_L        g20006(.A(new_n20262), .B(new_n20245), .Y(new_n20263));
  XNOR2x2_ASAP7_75t_L       g20007(.A(new_n20243), .B(new_n20263), .Y(new_n20264));
  OA21x2_ASAP7_75t_L        g20008(.A1(new_n20240), .A2(new_n20194), .B(new_n20264), .Y(new_n20265));
  NOR3xp33_ASAP7_75t_L      g20009(.A(new_n20264), .B(new_n20194), .C(new_n20240), .Y(new_n20266));
  NOR3xp33_ASAP7_75t_L      g20010(.A(new_n20265), .B(new_n20266), .C(new_n20239), .Y(new_n20267));
  INVx1_ASAP7_75t_L         g20011(.A(new_n20239), .Y(new_n20268));
  NOR2xp33_ASAP7_75t_L      g20012(.A(new_n20266), .B(new_n20265), .Y(new_n20269));
  NOR2xp33_ASAP7_75t_L      g20013(.A(new_n20268), .B(new_n20269), .Y(new_n20270));
  NOR2xp33_ASAP7_75t_L      g20014(.A(new_n20267), .B(new_n20270), .Y(new_n20271));
  A2O1A1Ixp33_ASAP7_75t_L   g20015(.A1(new_n20196), .A2(new_n20170), .B(new_n20199), .C(new_n20271), .Y(new_n20272));
  INVx1_ASAP7_75t_L         g20016(.A(new_n20272), .Y(new_n20273));
  AOI211xp5_ASAP7_75t_L     g20017(.A1(new_n20196), .A2(new_n20170), .B(new_n20271), .C(new_n20199), .Y(new_n20274));
  NOR2xp33_ASAP7_75t_L      g20018(.A(new_n20274), .B(new_n20273), .Y(new_n20275));
  XNOR2x2_ASAP7_75t_L       g20019(.A(new_n20236), .B(new_n20275), .Y(new_n20276));
  A2O1A1Ixp33_ASAP7_75t_L   g20020(.A1(new_n20204), .A2(new_n20203), .B(new_n20207), .C(new_n20276), .Y(new_n20277));
  INVx1_ASAP7_75t_L         g20021(.A(new_n20277), .Y(new_n20278));
  AOI211xp5_ASAP7_75t_L     g20022(.A1(new_n20203), .A2(new_n20204), .B(new_n20207), .C(new_n20276), .Y(new_n20279));
  NOR2xp33_ASAP7_75t_L      g20023(.A(new_n20279), .B(new_n20278), .Y(new_n20280));
  A2O1A1Ixp33_ASAP7_75t_L   g20024(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n7656), .Y(new_n20281));
  OAI221xp5_ASAP7_75t_L     g20025(.A1(new_n8326), .A2(new_n12599), .B1(new_n12273), .B2(new_n7994), .C(new_n20281), .Y(new_n20282));
  XNOR2x2_ASAP7_75t_L       g20026(.A(\a[50] ), .B(new_n20282), .Y(new_n20283));
  XNOR2x2_ASAP7_75t_L       g20027(.A(new_n20283), .B(new_n20280), .Y(new_n20284));
  INVx1_ASAP7_75t_L         g20028(.A(new_n20284), .Y(new_n20285));
  NAND2xp33_ASAP7_75t_L     g20029(.A(new_n20285), .B(new_n20230), .Y(new_n20286));
  A2O1A1Ixp33_ASAP7_75t_L   g20030(.A1(new_n20214), .A2(new_n20209), .B(new_n20218), .C(new_n20284), .Y(new_n20287));
  AND2x2_ASAP7_75t_L        g20031(.A(new_n20287), .B(new_n20286), .Y(new_n20288));
  INVx1_ASAP7_75t_L         g20032(.A(new_n20288), .Y(new_n20289));
  A2O1A1O1Ixp25_ASAP7_75t_L g20033(.A1(new_n20155), .A2(new_n20158), .B(new_n20220), .C(new_n20229), .D(new_n20289), .Y(new_n20290));
  A2O1A1Ixp33_ASAP7_75t_L   g20034(.A1(new_n20158), .A2(new_n20155), .B(new_n20225), .C(new_n20229), .Y(new_n20291));
  NOR2xp33_ASAP7_75t_L      g20035(.A(new_n20288), .B(new_n20291), .Y(new_n20292));
  NOR2xp33_ASAP7_75t_L      g20036(.A(new_n20290), .B(new_n20292), .Y(\f[112] ));
  INVx1_ASAP7_75t_L         g20037(.A(new_n20287), .Y(new_n20294));
  MAJIxp5_ASAP7_75t_L       g20038(.A(new_n20245), .B(new_n20243), .C(new_n20262), .Y(new_n20295));
  INVx1_ASAP7_75t_L         g20039(.A(new_n20250), .Y(new_n20296));
  NAND2xp33_ASAP7_75t_L     g20040(.A(\b[53] ), .B(new_n11656), .Y(new_n20297));
  OAI221xp5_ASAP7_75t_L     g20041(.A1(new_n8569), .A2(new_n12364), .B1(new_n12022), .B2(new_n8888), .C(new_n20297), .Y(new_n20298));
  AOI21xp33_ASAP7_75t_L     g20042(.A1(new_n12021), .A2(\b[51] ), .B(new_n20298), .Y(new_n20299));
  NAND2xp33_ASAP7_75t_L     g20043(.A(\a[62] ), .B(new_n20299), .Y(new_n20300));
  A2O1A1Ixp33_ASAP7_75t_L   g20044(.A1(\b[51] ), .A2(new_n12021), .B(new_n20298), .C(new_n11651), .Y(new_n20301));
  NAND2xp33_ASAP7_75t_L     g20045(.A(new_n20301), .B(new_n20300), .Y(new_n20302));
  NOR2xp33_ASAP7_75t_L      g20046(.A(new_n7907), .B(new_n12671), .Y(new_n20303));
  O2A1O1Ixp33_ASAP7_75t_L   g20047(.A1(new_n12353), .A2(new_n12355), .B(\b[50] ), .C(new_n20303), .Y(new_n20304));
  AND2x2_ASAP7_75t_L        g20048(.A(new_n20247), .B(new_n20304), .Y(new_n20305));
  O2A1O1Ixp33_ASAP7_75t_L   g20049(.A1(new_n7907), .A2(new_n12356), .B(new_n20251), .C(new_n20304), .Y(new_n20306));
  NOR2xp33_ASAP7_75t_L      g20050(.A(new_n20306), .B(new_n20305), .Y(new_n20307));
  XOR2x2_ASAP7_75t_L        g20051(.A(new_n20307), .B(new_n20302), .Y(new_n20308));
  NAND3xp33_ASAP7_75t_L     g20052(.A(new_n20260), .B(new_n20296), .C(new_n20308), .Y(new_n20309));
  O2A1O1Ixp33_ASAP7_75t_L   g20053(.A1(new_n20255), .A2(new_n20258), .B(new_n20296), .C(new_n20308), .Y(new_n20310));
  INVx1_ASAP7_75t_L         g20054(.A(new_n20310), .Y(new_n20311));
  AOI22xp33_ASAP7_75t_L     g20055(.A1(new_n10594), .A2(\b[56] ), .B1(new_n10591), .B2(new_n10185), .Y(new_n20312));
  OAI221xp5_ASAP7_75t_L     g20056(.A1(new_n11335), .A2(new_n9534), .B1(new_n9199), .B2(new_n11330), .C(new_n20312), .Y(new_n20313));
  XNOR2x2_ASAP7_75t_L       g20057(.A(\a[59] ), .B(new_n20313), .Y(new_n20314));
  INVx1_ASAP7_75t_L         g20058(.A(new_n20314), .Y(new_n20315));
  AO21x2_ASAP7_75t_L        g20059(.A1(new_n20309), .A2(new_n20311), .B(new_n20315), .Y(new_n20316));
  NAND3xp33_ASAP7_75t_L     g20060(.A(new_n20315), .B(new_n20311), .C(new_n20309), .Y(new_n20317));
  AND3x1_ASAP7_75t_L        g20061(.A(new_n20295), .B(new_n20317), .C(new_n20316), .Y(new_n20318));
  AOI21xp33_ASAP7_75t_L     g20062(.A1(new_n20317), .A2(new_n20316), .B(new_n20295), .Y(new_n20319));
  NOR2xp33_ASAP7_75t_L      g20063(.A(new_n20319), .B(new_n20318), .Y(new_n20320));
  AOI22xp33_ASAP7_75t_L     g20064(.A1(new_n9623), .A2(\b[59] ), .B1(new_n9620), .B2(new_n10887), .Y(new_n20321));
  OAI221xp5_ASAP7_75t_L     g20065(.A1(new_n10280), .A2(new_n10848), .B1(new_n10488), .B2(new_n12010), .C(new_n20321), .Y(new_n20322));
  XNOR2x2_ASAP7_75t_L       g20066(.A(\a[56] ), .B(new_n20322), .Y(new_n20323));
  AND2x2_ASAP7_75t_L        g20067(.A(new_n20323), .B(new_n20320), .Y(new_n20324));
  NOR2xp33_ASAP7_75t_L      g20068(.A(new_n20323), .B(new_n20320), .Y(new_n20325));
  NOR2xp33_ASAP7_75t_L      g20069(.A(new_n20325), .B(new_n20324), .Y(new_n20326));
  O2A1O1Ixp33_ASAP7_75t_L   g20070(.A1(new_n20240), .A2(new_n20194), .B(new_n20264), .C(new_n20267), .Y(new_n20327));
  NAND2xp33_ASAP7_75t_L     g20071(.A(new_n20326), .B(new_n20327), .Y(new_n20328));
  INVx1_ASAP7_75t_L         g20072(.A(new_n20326), .Y(new_n20329));
  A2O1A1Ixp33_ASAP7_75t_L   g20073(.A1(new_n20269), .A2(new_n20268), .B(new_n20265), .C(new_n20329), .Y(new_n20330));
  AOI22xp33_ASAP7_75t_L     g20074(.A1(new_n8645), .A2(\b[62] ), .B1(new_n8642), .B2(new_n12280), .Y(new_n20331));
  OAI221xp5_ASAP7_75t_L     g20075(.A1(new_n9322), .A2(new_n11911), .B1(new_n11226), .B2(new_n8965), .C(new_n20331), .Y(new_n20332));
  XNOR2x2_ASAP7_75t_L       g20076(.A(\a[53] ), .B(new_n20332), .Y(new_n20333));
  NAND3xp33_ASAP7_75t_L     g20077(.A(new_n20328), .B(new_n20330), .C(new_n20333), .Y(new_n20334));
  AO21x2_ASAP7_75t_L        g20078(.A1(new_n20330), .A2(new_n20328), .B(new_n20333), .Y(new_n20335));
  NAND2xp33_ASAP7_75t_L     g20079(.A(new_n20334), .B(new_n20335), .Y(new_n20336));
  INVx1_ASAP7_75t_L         g20080(.A(new_n20236), .Y(new_n20337));
  A2O1A1Ixp33_ASAP7_75t_L   g20081(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n7656), .Y(new_n20338));
  A2O1A1Ixp33_ASAP7_75t_L   g20082(.A1(new_n20338), .A2(new_n7994), .B(new_n12599), .C(\a[50] ), .Y(new_n20339));
  O2A1O1Ixp33_ASAP7_75t_L   g20083(.A1(new_n7996), .A2(new_n13934), .B(new_n7994), .C(new_n12599), .Y(new_n20340));
  NAND2xp33_ASAP7_75t_L     g20084(.A(new_n7653), .B(new_n20340), .Y(new_n20341));
  NAND2xp33_ASAP7_75t_L     g20085(.A(new_n20341), .B(new_n20339), .Y(new_n20342));
  A2O1A1Ixp33_ASAP7_75t_L   g20086(.A1(new_n20275), .A2(new_n20337), .B(new_n20273), .C(new_n20342), .Y(new_n20343));
  A2O1A1Ixp33_ASAP7_75t_L   g20087(.A1(new_n20234), .A2(new_n20235), .B(new_n20274), .C(new_n20272), .Y(new_n20344));
  NOR2xp33_ASAP7_75t_L      g20088(.A(new_n20342), .B(new_n20344), .Y(new_n20345));
  INVx1_ASAP7_75t_L         g20089(.A(new_n20345), .Y(new_n20346));
  NAND2xp33_ASAP7_75t_L     g20090(.A(new_n20346), .B(new_n20343), .Y(new_n20347));
  NAND2xp33_ASAP7_75t_L     g20091(.A(new_n20336), .B(new_n20347), .Y(new_n20348));
  NOR2xp33_ASAP7_75t_L      g20092(.A(new_n20336), .B(new_n20347), .Y(new_n20349));
  INVx1_ASAP7_75t_L         g20093(.A(new_n20349), .Y(new_n20350));
  NAND2xp33_ASAP7_75t_L     g20094(.A(new_n20348), .B(new_n20350), .Y(new_n20351));
  AOI21xp33_ASAP7_75t_L     g20095(.A1(new_n20277), .A2(new_n20283), .B(new_n20279), .Y(new_n20352));
  NOR2xp33_ASAP7_75t_L      g20096(.A(new_n20352), .B(new_n20351), .Y(new_n20353));
  NAND2xp33_ASAP7_75t_L     g20097(.A(new_n20352), .B(new_n20351), .Y(new_n20354));
  INVx1_ASAP7_75t_L         g20098(.A(new_n20354), .Y(new_n20355));
  NOR2xp33_ASAP7_75t_L      g20099(.A(new_n20353), .B(new_n20355), .Y(new_n20356));
  A2O1A1Ixp33_ASAP7_75t_L   g20100(.A1(new_n20291), .A2(new_n20288), .B(new_n20294), .C(new_n20356), .Y(new_n20357));
  INVx1_ASAP7_75t_L         g20101(.A(new_n20357), .Y(new_n20358));
  NOR3xp33_ASAP7_75t_L      g20102(.A(new_n20290), .B(new_n20356), .C(new_n20294), .Y(new_n20359));
  NOR2xp33_ASAP7_75t_L      g20103(.A(new_n20359), .B(new_n20358), .Y(\f[113] ));
  AOI22xp33_ASAP7_75t_L     g20104(.A1(new_n9623), .A2(\b[60] ), .B1(new_n9620), .B2(new_n11234), .Y(new_n20361));
  OAI221xp5_ASAP7_75t_L     g20105(.A1(new_n10280), .A2(new_n10881), .B1(new_n10848), .B2(new_n12010), .C(new_n20361), .Y(new_n20362));
  XNOR2x2_ASAP7_75t_L       g20106(.A(new_n9610), .B(new_n20362), .Y(new_n20363));
  AOI22xp33_ASAP7_75t_L     g20107(.A1(new_n10594), .A2(\b[57] ), .B1(new_n10591), .B2(new_n10495), .Y(new_n20364));
  OAI221xp5_ASAP7_75t_L     g20108(.A1(new_n11335), .A2(new_n10178), .B1(new_n9534), .B2(new_n11330), .C(new_n20364), .Y(new_n20365));
  XNOR2x2_ASAP7_75t_L       g20109(.A(\a[59] ), .B(new_n20365), .Y(new_n20366));
  AOI22xp33_ASAP7_75t_L     g20110(.A1(new_n11656), .A2(\b[54] ), .B1(new_n11654), .B2(new_n9208), .Y(new_n20367));
  OAI221xp5_ASAP7_75t_L     g20111(.A1(new_n12364), .A2(new_n8882), .B1(new_n8569), .B2(new_n13003), .C(new_n20367), .Y(new_n20368));
  XNOR2x2_ASAP7_75t_L       g20112(.A(\a[62] ), .B(new_n20368), .Y(new_n20369));
  A2O1A1Ixp33_ASAP7_75t_L   g20113(.A1(\b[50] ), .A2(new_n12669), .B(new_n20303), .C(new_n20247), .Y(new_n20370));
  NOR2xp33_ASAP7_75t_L      g20114(.A(new_n8228), .B(new_n12671), .Y(new_n20371));
  A2O1A1Ixp33_ASAP7_75t_L   g20115(.A1(new_n12669), .A2(\b[51] ), .B(new_n20371), .C(new_n7653), .Y(new_n20372));
  INVx1_ASAP7_75t_L         g20116(.A(new_n20372), .Y(new_n20373));
  O2A1O1Ixp33_ASAP7_75t_L   g20117(.A1(new_n12353), .A2(new_n12355), .B(\b[51] ), .C(new_n20371), .Y(new_n20374));
  NAND2xp33_ASAP7_75t_L     g20118(.A(\a[50] ), .B(new_n20374), .Y(new_n20375));
  INVx1_ASAP7_75t_L         g20119(.A(new_n20375), .Y(new_n20376));
  NOR2xp33_ASAP7_75t_L      g20120(.A(new_n20373), .B(new_n20376), .Y(new_n20377));
  INVx1_ASAP7_75t_L         g20121(.A(new_n20377), .Y(new_n20378));
  O2A1O1Ixp33_ASAP7_75t_L   g20122(.A1(new_n7907), .A2(new_n12356), .B(new_n20251), .C(new_n20378), .Y(new_n20379));
  INVx1_ASAP7_75t_L         g20123(.A(new_n20379), .Y(new_n20380));
  NAND2xp33_ASAP7_75t_L     g20124(.A(new_n20247), .B(new_n20378), .Y(new_n20381));
  AND2x2_ASAP7_75t_L        g20125(.A(new_n20381), .B(new_n20380), .Y(new_n20382));
  A2O1A1O1Ixp25_ASAP7_75t_L g20126(.A1(new_n20301), .A2(new_n20300), .B(new_n20307), .C(new_n20370), .D(new_n20382), .Y(new_n20383));
  A2O1A1Ixp33_ASAP7_75t_L   g20127(.A1(new_n20300), .A2(new_n20301), .B(new_n20307), .C(new_n20370), .Y(new_n20384));
  INVx1_ASAP7_75t_L         g20128(.A(new_n20382), .Y(new_n20385));
  NOR2xp33_ASAP7_75t_L      g20129(.A(new_n20385), .B(new_n20384), .Y(new_n20386));
  NOR2xp33_ASAP7_75t_L      g20130(.A(new_n20383), .B(new_n20386), .Y(new_n20387));
  NOR2xp33_ASAP7_75t_L      g20131(.A(new_n20369), .B(new_n20387), .Y(new_n20388));
  INVx1_ASAP7_75t_L         g20132(.A(new_n20369), .Y(new_n20389));
  NOR3xp33_ASAP7_75t_L      g20133(.A(new_n20389), .B(new_n20383), .C(new_n20386), .Y(new_n20390));
  NOR2xp33_ASAP7_75t_L      g20134(.A(new_n20388), .B(new_n20390), .Y(new_n20391));
  XOR2x2_ASAP7_75t_L        g20135(.A(new_n20366), .B(new_n20391), .Y(new_n20392));
  A2O1A1O1Ixp25_ASAP7_75t_L g20136(.A1(new_n20260), .A2(new_n20296), .B(new_n20308), .C(new_n20317), .D(new_n20392), .Y(new_n20393));
  AND3x1_ASAP7_75t_L        g20137(.A(new_n20392), .B(new_n20317), .C(new_n20311), .Y(new_n20394));
  NOR2xp33_ASAP7_75t_L      g20138(.A(new_n20393), .B(new_n20394), .Y(new_n20395));
  XOR2x2_ASAP7_75t_L        g20139(.A(new_n20363), .B(new_n20395), .Y(new_n20396));
  INVx1_ASAP7_75t_L         g20140(.A(new_n20396), .Y(new_n20397));
  OR3x1_ASAP7_75t_L         g20141(.A(new_n20397), .B(new_n20319), .C(new_n20324), .Y(new_n20398));
  A2O1A1Ixp33_ASAP7_75t_L   g20142(.A1(new_n20320), .A2(new_n20323), .B(new_n20319), .C(new_n20397), .Y(new_n20399));
  NAND2xp33_ASAP7_75t_L     g20143(.A(new_n20399), .B(new_n20398), .Y(new_n20400));
  NAND2xp33_ASAP7_75t_L     g20144(.A(\b[63] ), .B(new_n8645), .Y(new_n20401));
  A2O1A1Ixp33_ASAP7_75t_L   g20145(.A1(new_n12607), .A2(new_n12603), .B(new_n8967), .C(new_n20401), .Y(new_n20402));
  AOI221xp5_ASAP7_75t_L     g20146(.A1(\b[61] ), .A2(new_n8964), .B1(\b[62] ), .B2(new_n8635), .C(new_n20402), .Y(new_n20403));
  XNOR2x2_ASAP7_75t_L       g20147(.A(new_n8639), .B(new_n20403), .Y(new_n20404));
  XNOR2x2_ASAP7_75t_L       g20148(.A(new_n20404), .B(new_n20400), .Y(new_n20405));
  NAND2xp33_ASAP7_75t_L     g20149(.A(new_n20328), .B(new_n20334), .Y(new_n20406));
  XOR2x2_ASAP7_75t_L        g20150(.A(new_n20406), .B(new_n20405), .Y(new_n20407));
  O2A1O1Ixp33_ASAP7_75t_L   g20151(.A1(new_n20336), .A2(new_n20347), .B(new_n20346), .C(new_n20407), .Y(new_n20408));
  INVx1_ASAP7_75t_L         g20152(.A(new_n20407), .Y(new_n20409));
  NOR2xp33_ASAP7_75t_L      g20153(.A(new_n20345), .B(new_n20349), .Y(new_n20410));
  INVx1_ASAP7_75t_L         g20154(.A(new_n20410), .Y(new_n20411));
  NOR2xp33_ASAP7_75t_L      g20155(.A(new_n20409), .B(new_n20411), .Y(new_n20412));
  NOR2xp33_ASAP7_75t_L      g20156(.A(new_n20408), .B(new_n20412), .Y(new_n20413));
  A2O1A1Ixp33_ASAP7_75t_L   g20157(.A1(new_n20352), .A2(new_n20351), .B(new_n20358), .C(new_n20413), .Y(new_n20414));
  INVx1_ASAP7_75t_L         g20158(.A(new_n20414), .Y(new_n20415));
  NOR3xp33_ASAP7_75t_L      g20159(.A(new_n20358), .B(new_n20413), .C(new_n20355), .Y(new_n20416));
  NOR2xp33_ASAP7_75t_L      g20160(.A(new_n20416), .B(new_n20415), .Y(\f[114] ));
  INVx1_ASAP7_75t_L         g20161(.A(new_n20412), .Y(new_n20418));
  MAJIxp5_ASAP7_75t_L       g20162(.A(new_n20406), .B(new_n20400), .C(new_n20404), .Y(new_n20419));
  NAND2xp33_ASAP7_75t_L     g20163(.A(new_n20363), .B(new_n20395), .Y(new_n20420));
  NAND2xp33_ASAP7_75t_L     g20164(.A(new_n20420), .B(new_n20398), .Y(new_n20421));
  NAND2xp33_ASAP7_75t_L     g20165(.A(\b[61] ), .B(new_n9623), .Y(new_n20422));
  OAI221xp5_ASAP7_75t_L     g20166(.A1(new_n11226), .A2(new_n10280), .B1(new_n9949), .B2(new_n11920), .C(new_n20422), .Y(new_n20423));
  AOI21xp33_ASAP7_75t_L     g20167(.A1(new_n9948), .A2(\b[59] ), .B(new_n20423), .Y(new_n20424));
  NAND2xp33_ASAP7_75t_L     g20168(.A(\a[56] ), .B(new_n20424), .Y(new_n20425));
  A2O1A1Ixp33_ASAP7_75t_L   g20169(.A1(\b[59] ), .A2(new_n9948), .B(new_n20423), .C(new_n9610), .Y(new_n20426));
  AND2x2_ASAP7_75t_L        g20170(.A(new_n20426), .B(new_n20425), .Y(new_n20427));
  OR3x1_ASAP7_75t_L         g20171(.A(new_n20366), .B(new_n20388), .C(new_n20390), .Y(new_n20428));
  AOI22xp33_ASAP7_75t_L     g20172(.A1(new_n10594), .A2(\b[58] ), .B1(new_n10591), .B2(new_n10857), .Y(new_n20429));
  OAI221xp5_ASAP7_75t_L     g20173(.A1(new_n11335), .A2(new_n10488), .B1(new_n10178), .B2(new_n11330), .C(new_n20429), .Y(new_n20430));
  XNOR2x2_ASAP7_75t_L       g20174(.A(\a[59] ), .B(new_n20430), .Y(new_n20431));
  NOR2xp33_ASAP7_75t_L      g20175(.A(new_n8249), .B(new_n12671), .Y(new_n20432));
  A2O1A1O1Ixp25_ASAP7_75t_L g20176(.A1(new_n12669), .A2(\b[49] ), .B(new_n20246), .C(new_n20375), .D(new_n20373), .Y(new_n20433));
  A2O1A1Ixp33_ASAP7_75t_L   g20177(.A1(new_n12669), .A2(\b[52] ), .B(new_n20432), .C(new_n20433), .Y(new_n20434));
  O2A1O1Ixp33_ASAP7_75t_L   g20178(.A1(new_n12353), .A2(new_n12355), .B(\b[52] ), .C(new_n20432), .Y(new_n20435));
  INVx1_ASAP7_75t_L         g20179(.A(new_n20435), .Y(new_n20436));
  O2A1O1Ixp33_ASAP7_75t_L   g20180(.A1(new_n20247), .A2(new_n20376), .B(new_n20372), .C(new_n20436), .Y(new_n20437));
  INVx1_ASAP7_75t_L         g20181(.A(new_n20437), .Y(new_n20438));
  NAND2xp33_ASAP7_75t_L     g20182(.A(new_n20434), .B(new_n20438), .Y(new_n20439));
  NAND2xp33_ASAP7_75t_L     g20183(.A(new_n11654), .B(new_n9542), .Y(new_n20440));
  OAI221xp5_ASAP7_75t_L     g20184(.A1(new_n12023), .A2(new_n9534), .B1(new_n9199), .B2(new_n12364), .C(new_n20440), .Y(new_n20441));
  AOI21xp33_ASAP7_75t_L     g20185(.A1(new_n12021), .A2(\b[53] ), .B(new_n20441), .Y(new_n20442));
  NAND2xp33_ASAP7_75t_L     g20186(.A(\a[62] ), .B(new_n20442), .Y(new_n20443));
  A2O1A1Ixp33_ASAP7_75t_L   g20187(.A1(\b[53] ), .A2(new_n12021), .B(new_n20441), .C(new_n11651), .Y(new_n20444));
  AND2x2_ASAP7_75t_L        g20188(.A(new_n20444), .B(new_n20443), .Y(new_n20445));
  NAND2xp33_ASAP7_75t_L     g20189(.A(new_n20439), .B(new_n20445), .Y(new_n20446));
  NOR2xp33_ASAP7_75t_L      g20190(.A(new_n20439), .B(new_n20445), .Y(new_n20447));
  INVx1_ASAP7_75t_L         g20191(.A(new_n20447), .Y(new_n20448));
  AND2x2_ASAP7_75t_L        g20192(.A(new_n20446), .B(new_n20448), .Y(new_n20449));
  A2O1A1Ixp33_ASAP7_75t_L   g20193(.A1(new_n20382), .A2(new_n20384), .B(new_n20388), .C(new_n20449), .Y(new_n20450));
  INVx1_ASAP7_75t_L         g20194(.A(new_n20450), .Y(new_n20451));
  A2O1A1O1Ixp25_ASAP7_75t_L g20195(.A1(new_n20301), .A2(new_n20300), .B(new_n20307), .C(new_n20370), .D(new_n20385), .Y(new_n20452));
  O2A1O1Ixp33_ASAP7_75t_L   g20196(.A1(new_n20383), .A2(new_n20386), .B(new_n20389), .C(new_n20452), .Y(new_n20453));
  INVx1_ASAP7_75t_L         g20197(.A(new_n20453), .Y(new_n20454));
  NOR2xp33_ASAP7_75t_L      g20198(.A(new_n20454), .B(new_n20449), .Y(new_n20455));
  NOR2xp33_ASAP7_75t_L      g20199(.A(new_n20455), .B(new_n20451), .Y(new_n20456));
  INVx1_ASAP7_75t_L         g20200(.A(new_n20456), .Y(new_n20457));
  NOR2xp33_ASAP7_75t_L      g20201(.A(new_n20431), .B(new_n20457), .Y(new_n20458));
  INVx1_ASAP7_75t_L         g20202(.A(new_n20458), .Y(new_n20459));
  NAND2xp33_ASAP7_75t_L     g20203(.A(new_n20431), .B(new_n20457), .Y(new_n20460));
  AND2x2_ASAP7_75t_L        g20204(.A(new_n20460), .B(new_n20459), .Y(new_n20461));
  INVx1_ASAP7_75t_L         g20205(.A(new_n20461), .Y(new_n20462));
  A2O1A1O1Ixp25_ASAP7_75t_L g20206(.A1(new_n20317), .A2(new_n20311), .B(new_n20392), .C(new_n20428), .D(new_n20462), .Y(new_n20463));
  A2O1A1Ixp33_ASAP7_75t_L   g20207(.A1(new_n20317), .A2(new_n20311), .B(new_n20392), .C(new_n20428), .Y(new_n20464));
  NOR2xp33_ASAP7_75t_L      g20208(.A(new_n20464), .B(new_n20461), .Y(new_n20465));
  NOR2xp33_ASAP7_75t_L      g20209(.A(new_n20465), .B(new_n20463), .Y(new_n20466));
  XNOR2x2_ASAP7_75t_L       g20210(.A(new_n20427), .B(new_n20466), .Y(new_n20467));
  NAND2xp33_ASAP7_75t_L     g20211(.A(new_n20421), .B(new_n20467), .Y(new_n20468));
  INVx1_ASAP7_75t_L         g20212(.A(new_n20468), .Y(new_n20469));
  NOR2xp33_ASAP7_75t_L      g20213(.A(new_n20421), .B(new_n20467), .Y(new_n20470));
  NOR2xp33_ASAP7_75t_L      g20214(.A(new_n20470), .B(new_n20469), .Y(new_n20471));
  A2O1A1Ixp33_ASAP7_75t_L   g20215(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n8642), .Y(new_n20472));
  OAI221xp5_ASAP7_75t_L     g20216(.A1(new_n9322), .A2(new_n12599), .B1(new_n12273), .B2(new_n8965), .C(new_n20472), .Y(new_n20473));
  XNOR2x2_ASAP7_75t_L       g20217(.A(\a[53] ), .B(new_n20473), .Y(new_n20474));
  XNOR2x2_ASAP7_75t_L       g20218(.A(new_n20474), .B(new_n20471), .Y(new_n20475));
  NOR2xp33_ASAP7_75t_L      g20219(.A(new_n20419), .B(new_n20475), .Y(new_n20476));
  NAND2xp33_ASAP7_75t_L     g20220(.A(new_n20419), .B(new_n20475), .Y(new_n20477));
  INVx1_ASAP7_75t_L         g20221(.A(new_n20477), .Y(new_n20478));
  NOR2xp33_ASAP7_75t_L      g20222(.A(new_n20476), .B(new_n20478), .Y(new_n20479));
  INVx1_ASAP7_75t_L         g20223(.A(new_n20479), .Y(new_n20480));
  A2O1A1O1Ixp25_ASAP7_75t_L g20224(.A1(new_n20354), .A2(new_n20357), .B(new_n20408), .C(new_n20418), .D(new_n20480), .Y(new_n20481));
  A2O1A1Ixp33_ASAP7_75t_L   g20225(.A1(new_n20357), .A2(new_n20354), .B(new_n20408), .C(new_n20418), .Y(new_n20482));
  NOR2xp33_ASAP7_75t_L      g20226(.A(new_n20479), .B(new_n20482), .Y(new_n20483));
  NOR2xp33_ASAP7_75t_L      g20227(.A(new_n20481), .B(new_n20483), .Y(\f[115] ));
  O2A1O1Ixp33_ASAP7_75t_L   g20228(.A1(new_n20388), .A2(new_n20452), .B(new_n20449), .C(new_n20458), .Y(new_n20485));
  INVx1_ASAP7_75t_L         g20229(.A(new_n20485), .Y(new_n20486));
  AOI22xp33_ASAP7_75t_L     g20230(.A1(new_n10594), .A2(\b[59] ), .B1(new_n10591), .B2(new_n10887), .Y(new_n20487));
  OAI221xp5_ASAP7_75t_L     g20231(.A1(new_n11335), .A2(new_n10848), .B1(new_n10488), .B2(new_n11330), .C(new_n20487), .Y(new_n20488));
  XNOR2x2_ASAP7_75t_L       g20232(.A(\a[59] ), .B(new_n20488), .Y(new_n20489));
  INVx1_ASAP7_75t_L         g20233(.A(new_n20489), .Y(new_n20490));
  AOI22xp33_ASAP7_75t_L     g20234(.A1(new_n11656), .A2(\b[56] ), .B1(new_n11654), .B2(new_n10185), .Y(new_n20491));
  OAI221xp5_ASAP7_75t_L     g20235(.A1(new_n12364), .A2(new_n9534), .B1(new_n9199), .B2(new_n13003), .C(new_n20491), .Y(new_n20492));
  XNOR2x2_ASAP7_75t_L       g20236(.A(\a[62] ), .B(new_n20492), .Y(new_n20493));
  O2A1O1Ixp33_ASAP7_75t_L   g20237(.A1(new_n20373), .A2(new_n20379), .B(new_n20435), .C(new_n20447), .Y(new_n20494));
  NOR2xp33_ASAP7_75t_L      g20238(.A(new_n8569), .B(new_n12671), .Y(new_n20495));
  A2O1A1Ixp33_ASAP7_75t_L   g20239(.A1(\b[53] ), .A2(new_n12669), .B(new_n20495), .C(new_n20435), .Y(new_n20496));
  O2A1O1Ixp33_ASAP7_75t_L   g20240(.A1(new_n12353), .A2(new_n12355), .B(\b[53] ), .C(new_n20495), .Y(new_n20497));
  A2O1A1Ixp33_ASAP7_75t_L   g20241(.A1(new_n12669), .A2(\b[52] ), .B(new_n20432), .C(new_n20497), .Y(new_n20498));
  NAND2xp33_ASAP7_75t_L     g20242(.A(new_n20498), .B(new_n20496), .Y(new_n20499));
  XOR2x2_ASAP7_75t_L        g20243(.A(new_n20499), .B(new_n20494), .Y(new_n20500));
  INVx1_ASAP7_75t_L         g20244(.A(new_n20500), .Y(new_n20501));
  NOR2xp33_ASAP7_75t_L      g20245(.A(new_n20493), .B(new_n20501), .Y(new_n20502));
  INVx1_ASAP7_75t_L         g20246(.A(new_n20502), .Y(new_n20503));
  NAND2xp33_ASAP7_75t_L     g20247(.A(new_n20493), .B(new_n20501), .Y(new_n20504));
  NAND3xp33_ASAP7_75t_L     g20248(.A(new_n20503), .B(new_n20490), .C(new_n20504), .Y(new_n20505));
  AO21x2_ASAP7_75t_L        g20249(.A1(new_n20504), .A2(new_n20503), .B(new_n20490), .Y(new_n20506));
  AO21x2_ASAP7_75t_L        g20250(.A1(new_n20506), .A2(new_n20505), .B(new_n20486), .Y(new_n20507));
  AND2x2_ASAP7_75t_L        g20251(.A(new_n20505), .B(new_n20506), .Y(new_n20508));
  A2O1A1Ixp33_ASAP7_75t_L   g20252(.A1(new_n20449), .A2(new_n20454), .B(new_n20458), .C(new_n20508), .Y(new_n20509));
  AOI22xp33_ASAP7_75t_L     g20253(.A1(new_n9623), .A2(\b[62] ), .B1(new_n9620), .B2(new_n12280), .Y(new_n20510));
  OAI221xp5_ASAP7_75t_L     g20254(.A1(new_n10280), .A2(new_n11911), .B1(new_n11226), .B2(new_n12010), .C(new_n20510), .Y(new_n20511));
  XNOR2x2_ASAP7_75t_L       g20255(.A(\a[56] ), .B(new_n20511), .Y(new_n20512));
  NAND3xp33_ASAP7_75t_L     g20256(.A(new_n20507), .B(new_n20509), .C(new_n20512), .Y(new_n20513));
  AO21x2_ASAP7_75t_L        g20257(.A1(new_n20509), .A2(new_n20507), .B(new_n20512), .Y(new_n20514));
  NAND2xp33_ASAP7_75t_L     g20258(.A(new_n20513), .B(new_n20514), .Y(new_n20515));
  INVx1_ASAP7_75t_L         g20259(.A(new_n20427), .Y(new_n20516));
  A2O1A1Ixp33_ASAP7_75t_L   g20260(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n8642), .Y(new_n20517));
  A2O1A1Ixp33_ASAP7_75t_L   g20261(.A1(new_n20517), .A2(new_n8965), .B(new_n12599), .C(\a[53] ), .Y(new_n20518));
  O2A1O1Ixp33_ASAP7_75t_L   g20262(.A1(new_n8967), .A2(new_n13934), .B(new_n8965), .C(new_n12599), .Y(new_n20519));
  NAND2xp33_ASAP7_75t_L     g20263(.A(new_n8639), .B(new_n20519), .Y(new_n20520));
  NAND2xp33_ASAP7_75t_L     g20264(.A(new_n20520), .B(new_n20518), .Y(new_n20521));
  A2O1A1Ixp33_ASAP7_75t_L   g20265(.A1(new_n20466), .A2(new_n20516), .B(new_n20463), .C(new_n20521), .Y(new_n20522));
  INVx1_ASAP7_75t_L         g20266(.A(new_n20463), .Y(new_n20523));
  A2O1A1Ixp33_ASAP7_75t_L   g20267(.A1(new_n20425), .A2(new_n20426), .B(new_n20465), .C(new_n20523), .Y(new_n20524));
  NOR2xp33_ASAP7_75t_L      g20268(.A(new_n20521), .B(new_n20524), .Y(new_n20525));
  INVx1_ASAP7_75t_L         g20269(.A(new_n20525), .Y(new_n20526));
  NAND2xp33_ASAP7_75t_L     g20270(.A(new_n20522), .B(new_n20526), .Y(new_n20527));
  NAND2xp33_ASAP7_75t_L     g20271(.A(new_n20515), .B(new_n20527), .Y(new_n20528));
  NOR2xp33_ASAP7_75t_L      g20272(.A(new_n20515), .B(new_n20527), .Y(new_n20529));
  INVx1_ASAP7_75t_L         g20273(.A(new_n20529), .Y(new_n20530));
  AND2x2_ASAP7_75t_L        g20274(.A(new_n20528), .B(new_n20530), .Y(new_n20531));
  A2O1A1Ixp33_ASAP7_75t_L   g20275(.A1(new_n20474), .A2(new_n20468), .B(new_n20470), .C(new_n20531), .Y(new_n20532));
  AO221x2_ASAP7_75t_L       g20276(.A1(new_n20468), .A2(new_n20474), .B1(new_n20530), .B2(new_n20528), .C(new_n20470), .Y(new_n20533));
  NAND2xp33_ASAP7_75t_L     g20277(.A(new_n20533), .B(new_n20532), .Y(new_n20534));
  INVx1_ASAP7_75t_L         g20278(.A(new_n20534), .Y(new_n20535));
  A2O1A1Ixp33_ASAP7_75t_L   g20279(.A1(new_n20482), .A2(new_n20479), .B(new_n20478), .C(new_n20535), .Y(new_n20536));
  INVx1_ASAP7_75t_L         g20280(.A(new_n20536), .Y(new_n20537));
  A2O1A1Ixp33_ASAP7_75t_L   g20281(.A1(new_n20414), .A2(new_n20418), .B(new_n20480), .C(new_n20477), .Y(new_n20538));
  NOR2xp33_ASAP7_75t_L      g20282(.A(new_n20535), .B(new_n20538), .Y(new_n20539));
  NOR2xp33_ASAP7_75t_L      g20283(.A(new_n20537), .B(new_n20539), .Y(\f[116] ));
  INVx1_ASAP7_75t_L         g20284(.A(new_n20481), .Y(new_n20541));
  NAND2xp33_ASAP7_75t_L     g20285(.A(\b[63] ), .B(new_n9623), .Y(new_n20542));
  A2O1A1Ixp33_ASAP7_75t_L   g20286(.A1(new_n12607), .A2(new_n12603), .B(new_n9949), .C(new_n20542), .Y(new_n20543));
  AOI221xp5_ASAP7_75t_L     g20287(.A1(\b[61] ), .A2(new_n9948), .B1(\b[62] ), .B2(new_n9614), .C(new_n20543), .Y(new_n20544));
  XNOR2x2_ASAP7_75t_L       g20288(.A(new_n9610), .B(new_n20544), .Y(new_n20545));
  A2O1A1Ixp33_ASAP7_75t_L   g20289(.A1(new_n20505), .A2(new_n20506), .B(new_n20486), .C(new_n20513), .Y(new_n20546));
  NOR2xp33_ASAP7_75t_L      g20290(.A(new_n20545), .B(new_n20546), .Y(new_n20547));
  INVx1_ASAP7_75t_L         g20291(.A(new_n20545), .Y(new_n20548));
  O2A1O1Ixp33_ASAP7_75t_L   g20292(.A1(new_n20486), .A2(new_n20508), .B(new_n20513), .C(new_n20548), .Y(new_n20549));
  NOR2xp33_ASAP7_75t_L      g20293(.A(new_n20549), .B(new_n20547), .Y(new_n20550));
  AOI22xp33_ASAP7_75t_L     g20294(.A1(new_n10594), .A2(\b[60] ), .B1(new_n10591), .B2(new_n11234), .Y(new_n20551));
  OAI221xp5_ASAP7_75t_L     g20295(.A1(new_n11335), .A2(new_n10881), .B1(new_n10848), .B2(new_n11330), .C(new_n20551), .Y(new_n20552));
  XNOR2x2_ASAP7_75t_L       g20296(.A(\a[59] ), .B(new_n20552), .Y(new_n20553));
  INVx1_ASAP7_75t_L         g20297(.A(new_n20553), .Y(new_n20554));
  A2O1A1Ixp33_ASAP7_75t_L   g20298(.A1(new_n12669), .A2(\b[53] ), .B(new_n20495), .C(\a[53] ), .Y(new_n20555));
  INVx1_ASAP7_75t_L         g20299(.A(new_n20497), .Y(new_n20556));
  NOR2xp33_ASAP7_75t_L      g20300(.A(\a[53] ), .B(new_n20556), .Y(new_n20557));
  INVx1_ASAP7_75t_L         g20301(.A(new_n20557), .Y(new_n20558));
  AND2x2_ASAP7_75t_L        g20302(.A(new_n20555), .B(new_n20558), .Y(new_n20559));
  INVx1_ASAP7_75t_L         g20303(.A(new_n20559), .Y(new_n20560));
  NOR2xp33_ASAP7_75t_L      g20304(.A(new_n8882), .B(new_n12671), .Y(new_n20561));
  INVx1_ASAP7_75t_L         g20305(.A(new_n20561), .Y(new_n20562));
  A2O1A1Ixp33_ASAP7_75t_L   g20306(.A1(new_n19241), .A2(new_n19242), .B(new_n9199), .C(new_n20562), .Y(new_n20563));
  NOR2xp33_ASAP7_75t_L      g20307(.A(new_n20563), .B(new_n20560), .Y(new_n20564));
  O2A1O1Ixp33_ASAP7_75t_L   g20308(.A1(new_n12356), .A2(new_n9199), .B(new_n20562), .C(new_n20559), .Y(new_n20565));
  NOR2xp33_ASAP7_75t_L      g20309(.A(new_n20565), .B(new_n20564), .Y(new_n20566));
  INVx1_ASAP7_75t_L         g20310(.A(new_n20566), .Y(new_n20567));
  AOI22xp33_ASAP7_75t_L     g20311(.A1(new_n11656), .A2(\b[57] ), .B1(new_n11654), .B2(new_n10495), .Y(new_n20568));
  OAI221xp5_ASAP7_75t_L     g20312(.A1(new_n12364), .A2(new_n10178), .B1(new_n9534), .B2(new_n13003), .C(new_n20568), .Y(new_n20569));
  XNOR2x2_ASAP7_75t_L       g20313(.A(\a[62] ), .B(new_n20569), .Y(new_n20570));
  XNOR2x2_ASAP7_75t_L       g20314(.A(new_n20567), .B(new_n20570), .Y(new_n20571));
  INVx1_ASAP7_75t_L         g20315(.A(new_n20571), .Y(new_n20572));
  INVx1_ASAP7_75t_L         g20316(.A(new_n20494), .Y(new_n20573));
  A2O1A1O1Ixp25_ASAP7_75t_L g20317(.A1(new_n12669), .A2(\b[52] ), .B(new_n20432), .C(new_n20497), .D(new_n20573), .Y(new_n20574));
  A2O1A1O1Ixp25_ASAP7_75t_L g20318(.A1(new_n12669), .A2(\b[53] ), .B(new_n20495), .C(new_n20435), .D(new_n20574), .Y(new_n20575));
  NAND2xp33_ASAP7_75t_L     g20319(.A(new_n20572), .B(new_n20575), .Y(new_n20576));
  A2O1A1Ixp33_ASAP7_75t_L   g20320(.A1(new_n20435), .A2(new_n20556), .B(new_n20574), .C(new_n20571), .Y(new_n20577));
  AND2x2_ASAP7_75t_L        g20321(.A(new_n20577), .B(new_n20576), .Y(new_n20578));
  XNOR2x2_ASAP7_75t_L       g20322(.A(new_n20554), .B(new_n20578), .Y(new_n20579));
  O2A1O1Ixp33_ASAP7_75t_L   g20323(.A1(new_n20493), .A2(new_n20501), .B(new_n20505), .C(new_n20579), .Y(new_n20580));
  AND3x1_ASAP7_75t_L        g20324(.A(new_n20579), .B(new_n20505), .C(new_n20503), .Y(new_n20581));
  NOR2xp33_ASAP7_75t_L      g20325(.A(new_n20580), .B(new_n20581), .Y(new_n20582));
  NAND2xp33_ASAP7_75t_L     g20326(.A(new_n20582), .B(new_n20550), .Y(new_n20583));
  INVx1_ASAP7_75t_L         g20327(.A(new_n20583), .Y(new_n20584));
  NOR2xp33_ASAP7_75t_L      g20328(.A(new_n20582), .B(new_n20550), .Y(new_n20585));
  NOR2xp33_ASAP7_75t_L      g20329(.A(new_n20585), .B(new_n20584), .Y(new_n20586));
  INVx1_ASAP7_75t_L         g20330(.A(new_n20586), .Y(new_n20587));
  NOR2xp33_ASAP7_75t_L      g20331(.A(new_n20525), .B(new_n20529), .Y(new_n20588));
  INVx1_ASAP7_75t_L         g20332(.A(new_n20588), .Y(new_n20589));
  NOR2xp33_ASAP7_75t_L      g20333(.A(new_n20587), .B(new_n20589), .Y(new_n20590));
  O2A1O1Ixp33_ASAP7_75t_L   g20334(.A1(new_n20515), .A2(new_n20527), .B(new_n20526), .C(new_n20586), .Y(new_n20591));
  NOR2xp33_ASAP7_75t_L      g20335(.A(new_n20591), .B(new_n20590), .Y(new_n20592));
  INVx1_ASAP7_75t_L         g20336(.A(new_n20592), .Y(new_n20593));
  A2O1A1O1Ixp25_ASAP7_75t_L g20337(.A1(new_n20477), .A2(new_n20541), .B(new_n20534), .C(new_n20533), .D(new_n20593), .Y(new_n20594));
  A2O1A1Ixp33_ASAP7_75t_L   g20338(.A1(new_n20541), .A2(new_n20477), .B(new_n20534), .C(new_n20533), .Y(new_n20595));
  NOR2xp33_ASAP7_75t_L      g20339(.A(new_n20592), .B(new_n20595), .Y(new_n20596));
  NOR2xp33_ASAP7_75t_L      g20340(.A(new_n20594), .B(new_n20596), .Y(\f[117] ));
  INVx1_ASAP7_75t_L         g20341(.A(new_n20590), .Y(new_n20598));
  AOI22xp33_ASAP7_75t_L     g20342(.A1(new_n10594), .A2(\b[61] ), .B1(new_n10591), .B2(new_n11919), .Y(new_n20599));
  OAI221xp5_ASAP7_75t_L     g20343(.A1(new_n11335), .A2(new_n11226), .B1(new_n10881), .B2(new_n11330), .C(new_n20599), .Y(new_n20600));
  XNOR2x2_ASAP7_75t_L       g20344(.A(\a[59] ), .B(new_n20600), .Y(new_n20601));
  NOR2xp33_ASAP7_75t_L      g20345(.A(new_n20567), .B(new_n20570), .Y(new_n20602));
  NOR2xp33_ASAP7_75t_L      g20346(.A(new_n9199), .B(new_n12671), .Y(new_n20603));
  O2A1O1Ixp33_ASAP7_75t_L   g20347(.A1(new_n12353), .A2(new_n12355), .B(\b[55] ), .C(new_n20603), .Y(new_n20604));
  A2O1A1Ixp33_ASAP7_75t_L   g20348(.A1(new_n20556), .A2(new_n8639), .B(new_n20565), .C(new_n20604), .Y(new_n20605));
  A2O1A1O1Ixp25_ASAP7_75t_L g20349(.A1(new_n12669), .A2(\b[53] ), .B(new_n20495), .C(new_n8639), .D(new_n20565), .Y(new_n20606));
  A2O1A1Ixp33_ASAP7_75t_L   g20350(.A1(new_n12669), .A2(\b[55] ), .B(new_n20603), .C(new_n20606), .Y(new_n20607));
  NAND2xp33_ASAP7_75t_L     g20351(.A(new_n20605), .B(new_n20607), .Y(new_n20608));
  AOI22xp33_ASAP7_75t_L     g20352(.A1(new_n11647), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n11656), .Y(new_n20609));
  OAI221xp5_ASAP7_75t_L     g20353(.A1(new_n13003), .A2(new_n10178), .B1(new_n12022), .B2(new_n10856), .C(new_n20609), .Y(new_n20610));
  XNOR2x2_ASAP7_75t_L       g20354(.A(\a[62] ), .B(new_n20610), .Y(new_n20611));
  NOR2xp33_ASAP7_75t_L      g20355(.A(new_n20608), .B(new_n20611), .Y(new_n20612));
  AND2x2_ASAP7_75t_L        g20356(.A(new_n20608), .B(new_n20611), .Y(new_n20613));
  NOR2xp33_ASAP7_75t_L      g20357(.A(new_n20612), .B(new_n20613), .Y(new_n20614));
  A2O1A1Ixp33_ASAP7_75t_L   g20358(.A1(new_n20575), .A2(new_n20572), .B(new_n20602), .C(new_n20614), .Y(new_n20615));
  OAI221xp5_ASAP7_75t_L     g20359(.A1(new_n20570), .A2(new_n20567), .B1(new_n20612), .B2(new_n20613), .C(new_n20576), .Y(new_n20616));
  NAND2xp33_ASAP7_75t_L     g20360(.A(new_n20615), .B(new_n20616), .Y(new_n20617));
  OR2x4_ASAP7_75t_L         g20361(.A(new_n20601), .B(new_n20617), .Y(new_n20618));
  NAND2xp33_ASAP7_75t_L     g20362(.A(new_n20601), .B(new_n20617), .Y(new_n20619));
  AND2x2_ASAP7_75t_L        g20363(.A(new_n20619), .B(new_n20618), .Y(new_n20620));
  A2O1A1Ixp33_ASAP7_75t_L   g20364(.A1(new_n20578), .A2(new_n20554), .B(new_n20580), .C(new_n20620), .Y(new_n20621));
  INVx1_ASAP7_75t_L         g20365(.A(new_n20621), .Y(new_n20622));
  AOI211xp5_ASAP7_75t_L     g20366(.A1(new_n20554), .A2(new_n20578), .B(new_n20580), .C(new_n20620), .Y(new_n20623));
  NOR2xp33_ASAP7_75t_L      g20367(.A(new_n20623), .B(new_n20622), .Y(new_n20624));
  A2O1A1Ixp33_ASAP7_75t_L   g20368(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n9620), .Y(new_n20625));
  OAI221xp5_ASAP7_75t_L     g20369(.A1(new_n10280), .A2(new_n12599), .B1(new_n12273), .B2(new_n12010), .C(new_n20625), .Y(new_n20626));
  XNOR2x2_ASAP7_75t_L       g20370(.A(\a[56] ), .B(new_n20626), .Y(new_n20627));
  XNOR2x2_ASAP7_75t_L       g20371(.A(new_n20627), .B(new_n20624), .Y(new_n20628));
  INVx1_ASAP7_75t_L         g20372(.A(new_n20628), .Y(new_n20629));
  O2A1O1Ixp33_ASAP7_75t_L   g20373(.A1(new_n20545), .A2(new_n20546), .B(new_n20583), .C(new_n20629), .Y(new_n20630));
  INVx1_ASAP7_75t_L         g20374(.A(new_n20630), .Y(new_n20631));
  OAI211xp5_ASAP7_75t_L     g20375(.A1(new_n20545), .A2(new_n20546), .B(new_n20629), .C(new_n20583), .Y(new_n20632));
  AND2x2_ASAP7_75t_L        g20376(.A(new_n20632), .B(new_n20631), .Y(new_n20633));
  INVx1_ASAP7_75t_L         g20377(.A(new_n20633), .Y(new_n20634));
  A2O1A1O1Ixp25_ASAP7_75t_L g20378(.A1(new_n20533), .A2(new_n20536), .B(new_n20591), .C(new_n20598), .D(new_n20634), .Y(new_n20635));
  A2O1A1Ixp33_ASAP7_75t_L   g20379(.A1(new_n20536), .A2(new_n20533), .B(new_n20593), .C(new_n20598), .Y(new_n20636));
  NOR2xp33_ASAP7_75t_L      g20380(.A(new_n20633), .B(new_n20636), .Y(new_n20637));
  NOR2xp33_ASAP7_75t_L      g20381(.A(new_n20635), .B(new_n20637), .Y(\f[118] ));
  NAND2xp33_ASAP7_75t_L     g20382(.A(\b[59] ), .B(new_n11656), .Y(new_n20639));
  OAI221xp5_ASAP7_75t_L     g20383(.A1(new_n10848), .A2(new_n12364), .B1(new_n12022), .B2(new_n10888), .C(new_n20639), .Y(new_n20640));
  AOI21xp33_ASAP7_75t_L     g20384(.A1(new_n12021), .A2(\b[57] ), .B(new_n20640), .Y(new_n20641));
  NAND2xp33_ASAP7_75t_L     g20385(.A(\a[62] ), .B(new_n20641), .Y(new_n20642));
  A2O1A1Ixp33_ASAP7_75t_L   g20386(.A1(\b[57] ), .A2(new_n12021), .B(new_n20640), .C(new_n11651), .Y(new_n20643));
  NAND2xp33_ASAP7_75t_L     g20387(.A(new_n20643), .B(new_n20642), .Y(new_n20644));
  NOR2xp33_ASAP7_75t_L      g20388(.A(new_n9534), .B(new_n12671), .Y(new_n20645));
  O2A1O1Ixp33_ASAP7_75t_L   g20389(.A1(new_n12353), .A2(new_n12355), .B(\b[56] ), .C(new_n20645), .Y(new_n20646));
  NAND2xp33_ASAP7_75t_L     g20390(.A(new_n20646), .B(new_n20604), .Y(new_n20647));
  INVx1_ASAP7_75t_L         g20391(.A(new_n20604), .Y(new_n20648));
  A2O1A1Ixp33_ASAP7_75t_L   g20392(.A1(\b[56] ), .A2(new_n12669), .B(new_n20645), .C(new_n20648), .Y(new_n20649));
  AND2x2_ASAP7_75t_L        g20393(.A(new_n20647), .B(new_n20649), .Y(new_n20650));
  INVx1_ASAP7_75t_L         g20394(.A(new_n20650), .Y(new_n20651));
  XNOR2x2_ASAP7_75t_L       g20395(.A(new_n20651), .B(new_n20644), .Y(new_n20652));
  A2O1A1O1Ixp25_ASAP7_75t_L g20396(.A1(new_n20556), .A2(new_n8639), .B(new_n20565), .C(new_n20604), .D(new_n20612), .Y(new_n20653));
  NAND2xp33_ASAP7_75t_L     g20397(.A(new_n20653), .B(new_n20652), .Y(new_n20654));
  INVx1_ASAP7_75t_L         g20398(.A(new_n20606), .Y(new_n20655));
  INVx1_ASAP7_75t_L         g20399(.A(new_n20652), .Y(new_n20656));
  A2O1A1Ixp33_ASAP7_75t_L   g20400(.A1(new_n20655), .A2(new_n20604), .B(new_n20612), .C(new_n20656), .Y(new_n20657));
  AOI22xp33_ASAP7_75t_L     g20401(.A1(new_n10594), .A2(\b[62] ), .B1(new_n10591), .B2(new_n12280), .Y(new_n20658));
  OAI221xp5_ASAP7_75t_L     g20402(.A1(new_n11335), .A2(new_n11911), .B1(new_n11226), .B2(new_n11330), .C(new_n20658), .Y(new_n20659));
  XNOR2x2_ASAP7_75t_L       g20403(.A(\a[59] ), .B(new_n20659), .Y(new_n20660));
  NAND3xp33_ASAP7_75t_L     g20404(.A(new_n20657), .B(new_n20654), .C(new_n20660), .Y(new_n20661));
  AO21x2_ASAP7_75t_L        g20405(.A1(new_n20654), .A2(new_n20657), .B(new_n20660), .Y(new_n20662));
  NAND2xp33_ASAP7_75t_L     g20406(.A(new_n20661), .B(new_n20662), .Y(new_n20663));
  NAND2xp33_ASAP7_75t_L     g20407(.A(new_n20615), .B(new_n20618), .Y(new_n20664));
  A2O1A1Ixp33_ASAP7_75t_L   g20408(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n9620), .Y(new_n20665));
  A2O1A1Ixp33_ASAP7_75t_L   g20409(.A1(new_n20665), .A2(new_n12010), .B(new_n12599), .C(\a[56] ), .Y(new_n20666));
  O2A1O1Ixp33_ASAP7_75t_L   g20410(.A1(new_n9949), .A2(new_n13934), .B(new_n12010), .C(new_n12599), .Y(new_n20667));
  NAND2xp33_ASAP7_75t_L     g20411(.A(new_n9610), .B(new_n20667), .Y(new_n20668));
  NAND2xp33_ASAP7_75t_L     g20412(.A(new_n20668), .B(new_n20666), .Y(new_n20669));
  NAND2xp33_ASAP7_75t_L     g20413(.A(new_n20669), .B(new_n20664), .Y(new_n20670));
  NOR2xp33_ASAP7_75t_L      g20414(.A(new_n20669), .B(new_n20664), .Y(new_n20671));
  INVx1_ASAP7_75t_L         g20415(.A(new_n20671), .Y(new_n20672));
  NAND2xp33_ASAP7_75t_L     g20416(.A(new_n20670), .B(new_n20672), .Y(new_n20673));
  NAND2xp33_ASAP7_75t_L     g20417(.A(new_n20663), .B(new_n20673), .Y(new_n20674));
  NOR2xp33_ASAP7_75t_L      g20418(.A(new_n20663), .B(new_n20673), .Y(new_n20675));
  INVx1_ASAP7_75t_L         g20419(.A(new_n20675), .Y(new_n20676));
  NAND2xp33_ASAP7_75t_L     g20420(.A(new_n20674), .B(new_n20676), .Y(new_n20677));
  AOI21xp33_ASAP7_75t_L     g20421(.A1(new_n20621), .A2(new_n20627), .B(new_n20623), .Y(new_n20678));
  NOR2xp33_ASAP7_75t_L      g20422(.A(new_n20678), .B(new_n20677), .Y(new_n20679));
  NAND2xp33_ASAP7_75t_L     g20423(.A(new_n20678), .B(new_n20677), .Y(new_n20680));
  INVx1_ASAP7_75t_L         g20424(.A(new_n20680), .Y(new_n20681));
  NOR2xp33_ASAP7_75t_L      g20425(.A(new_n20679), .B(new_n20681), .Y(new_n20682));
  A2O1A1Ixp33_ASAP7_75t_L   g20426(.A1(new_n20636), .A2(new_n20633), .B(new_n20630), .C(new_n20682), .Y(new_n20683));
  INVx1_ASAP7_75t_L         g20427(.A(new_n20683), .Y(new_n20684));
  NOR3xp33_ASAP7_75t_L      g20428(.A(new_n20635), .B(new_n20682), .C(new_n20630), .Y(new_n20685));
  NOR2xp33_ASAP7_75t_L      g20429(.A(new_n20685), .B(new_n20684), .Y(\f[119] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20430(.A1(new_n20595), .A2(new_n20592), .B(new_n20590), .C(new_n20633), .Y(new_n20687));
  A2O1A1Ixp33_ASAP7_75t_L   g20431(.A1(\b[56] ), .A2(new_n12669), .B(new_n20645), .C(new_n20604), .Y(new_n20688));
  A2O1A1Ixp33_ASAP7_75t_L   g20432(.A1(new_n20642), .A2(new_n20643), .B(new_n20650), .C(new_n20688), .Y(new_n20689));
  NOR2xp33_ASAP7_75t_L      g20433(.A(new_n10178), .B(new_n12671), .Y(new_n20690));
  O2A1O1Ixp33_ASAP7_75t_L   g20434(.A1(new_n12353), .A2(new_n12355), .B(\b[57] ), .C(new_n20690), .Y(new_n20691));
  INVx1_ASAP7_75t_L         g20435(.A(new_n20691), .Y(new_n20692));
  NOR2xp33_ASAP7_75t_L      g20436(.A(\a[56] ), .B(new_n20692), .Y(new_n20693));
  INVx1_ASAP7_75t_L         g20437(.A(new_n20693), .Y(new_n20694));
  A2O1A1Ixp33_ASAP7_75t_L   g20438(.A1(new_n12669), .A2(\b[57] ), .B(new_n20690), .C(\a[56] ), .Y(new_n20695));
  NAND2xp33_ASAP7_75t_L     g20439(.A(new_n20695), .B(new_n20694), .Y(new_n20696));
  A2O1A1Ixp33_ASAP7_75t_L   g20440(.A1(new_n12669), .A2(\b[55] ), .B(new_n20603), .C(new_n20696), .Y(new_n20697));
  NAND3xp33_ASAP7_75t_L     g20441(.A(new_n20694), .B(new_n20604), .C(new_n20695), .Y(new_n20698));
  AND2x2_ASAP7_75t_L        g20442(.A(new_n20698), .B(new_n20697), .Y(new_n20699));
  NOR2xp33_ASAP7_75t_L      g20443(.A(new_n20699), .B(new_n20689), .Y(new_n20700));
  INVx1_ASAP7_75t_L         g20444(.A(new_n20699), .Y(new_n20701));
  A2O1A1O1Ixp25_ASAP7_75t_L g20445(.A1(new_n20643), .A2(new_n20642), .B(new_n20650), .C(new_n20688), .D(new_n20701), .Y(new_n20702));
  NOR2xp33_ASAP7_75t_L      g20446(.A(new_n20702), .B(new_n20700), .Y(new_n20703));
  INVx1_ASAP7_75t_L         g20447(.A(new_n20703), .Y(new_n20704));
  AOI22xp33_ASAP7_75t_L     g20448(.A1(new_n11656), .A2(\b[60] ), .B1(new_n11654), .B2(new_n11234), .Y(new_n20705));
  OAI221xp5_ASAP7_75t_L     g20449(.A1(new_n12364), .A2(new_n10881), .B1(new_n10848), .B2(new_n13003), .C(new_n20705), .Y(new_n20706));
  XNOR2x2_ASAP7_75t_L       g20450(.A(\a[62] ), .B(new_n20706), .Y(new_n20707));
  NOR2xp33_ASAP7_75t_L      g20451(.A(new_n20707), .B(new_n20704), .Y(new_n20708));
  AND2x2_ASAP7_75t_L        g20452(.A(new_n20707), .B(new_n20704), .Y(new_n20709));
  NOR2xp33_ASAP7_75t_L      g20453(.A(new_n20708), .B(new_n20709), .Y(new_n20710));
  NAND2xp33_ASAP7_75t_L     g20454(.A(\b[63] ), .B(new_n10594), .Y(new_n20711));
  A2O1A1Ixp33_ASAP7_75t_L   g20455(.A1(new_n12607), .A2(new_n12603), .B(new_n10974), .C(new_n20711), .Y(new_n20712));
  AOI221xp5_ASAP7_75t_L     g20456(.A1(\b[61] ), .A2(new_n10973), .B1(\b[62] ), .B2(new_n10584), .C(new_n20712), .Y(new_n20713));
  XNOR2x2_ASAP7_75t_L       g20457(.A(new_n10588), .B(new_n20713), .Y(new_n20714));
  NAND2xp33_ASAP7_75t_L     g20458(.A(new_n20654), .B(new_n20661), .Y(new_n20715));
  NOR2xp33_ASAP7_75t_L      g20459(.A(new_n20714), .B(new_n20715), .Y(new_n20716));
  INVx1_ASAP7_75t_L         g20460(.A(new_n20716), .Y(new_n20717));
  NAND2xp33_ASAP7_75t_L     g20461(.A(new_n20714), .B(new_n20715), .Y(new_n20718));
  NAND3xp33_ASAP7_75t_L     g20462(.A(new_n20717), .B(new_n20710), .C(new_n20718), .Y(new_n20719));
  AO21x2_ASAP7_75t_L        g20463(.A1(new_n20718), .A2(new_n20717), .B(new_n20710), .Y(new_n20720));
  AND2x2_ASAP7_75t_L        g20464(.A(new_n20719), .B(new_n20720), .Y(new_n20721));
  O2A1O1Ixp33_ASAP7_75t_L   g20465(.A1(new_n20663), .A2(new_n20673), .B(new_n20672), .C(new_n20721), .Y(new_n20722));
  INVx1_ASAP7_75t_L         g20466(.A(new_n20722), .Y(new_n20723));
  NAND3xp33_ASAP7_75t_L     g20467(.A(new_n20676), .B(new_n20672), .C(new_n20721), .Y(new_n20724));
  AND2x2_ASAP7_75t_L        g20468(.A(new_n20723), .B(new_n20724), .Y(new_n20725));
  INVx1_ASAP7_75t_L         g20469(.A(new_n20725), .Y(new_n20726));
  A2O1A1O1Ixp25_ASAP7_75t_L g20470(.A1(new_n20631), .A2(new_n20687), .B(new_n20679), .C(new_n20680), .D(new_n20726), .Y(new_n20727));
  A2O1A1Ixp33_ASAP7_75t_L   g20471(.A1(new_n20687), .A2(new_n20631), .B(new_n20679), .C(new_n20680), .Y(new_n20728));
  NOR2xp33_ASAP7_75t_L      g20472(.A(new_n20725), .B(new_n20728), .Y(new_n20729));
  NOR2xp33_ASAP7_75t_L      g20473(.A(new_n20727), .B(new_n20729), .Y(\f[120] ));
  INVx1_ASAP7_75t_L         g20474(.A(new_n20702), .Y(new_n20731));
  NOR2xp33_ASAP7_75t_L      g20475(.A(new_n10488), .B(new_n12671), .Y(new_n20732));
  INVx1_ASAP7_75t_L         g20476(.A(new_n20697), .Y(new_n20733));
  A2O1A1O1Ixp25_ASAP7_75t_L g20477(.A1(new_n12669), .A2(\b[57] ), .B(new_n20690), .C(new_n9610), .D(new_n20733), .Y(new_n20734));
  A2O1A1Ixp33_ASAP7_75t_L   g20478(.A1(new_n12669), .A2(\b[58] ), .B(new_n20732), .C(new_n20734), .Y(new_n20735));
  O2A1O1Ixp33_ASAP7_75t_L   g20479(.A1(new_n12353), .A2(new_n12355), .B(\b[58] ), .C(new_n20732), .Y(new_n20736));
  INVx1_ASAP7_75t_L         g20480(.A(new_n20736), .Y(new_n20737));
  A2O1A1Ixp33_ASAP7_75t_L   g20481(.A1(new_n12669), .A2(\b[57] ), .B(new_n20690), .C(new_n9610), .Y(new_n20738));
  A2O1A1O1Ixp25_ASAP7_75t_L g20482(.A1(new_n20695), .A2(new_n20694), .B(new_n20604), .C(new_n20738), .D(new_n20737), .Y(new_n20739));
  INVx1_ASAP7_75t_L         g20483(.A(new_n20739), .Y(new_n20740));
  NAND2xp33_ASAP7_75t_L     g20484(.A(new_n20740), .B(new_n20735), .Y(new_n20741));
  NAND2xp33_ASAP7_75t_L     g20485(.A(\b[60] ), .B(new_n11647), .Y(new_n20742));
  OAI221xp5_ASAP7_75t_L     g20486(.A1(new_n12023), .A2(new_n11911), .B1(new_n12022), .B2(new_n11920), .C(new_n20742), .Y(new_n20743));
  AOI21xp33_ASAP7_75t_L     g20487(.A1(new_n12021), .A2(\b[59] ), .B(new_n20743), .Y(new_n20744));
  NAND2xp33_ASAP7_75t_L     g20488(.A(\a[62] ), .B(new_n20744), .Y(new_n20745));
  A2O1A1Ixp33_ASAP7_75t_L   g20489(.A1(\b[59] ), .A2(new_n12021), .B(new_n20743), .C(new_n11651), .Y(new_n20746));
  AND2x2_ASAP7_75t_L        g20490(.A(new_n20746), .B(new_n20745), .Y(new_n20747));
  NOR2xp33_ASAP7_75t_L      g20491(.A(new_n20741), .B(new_n20747), .Y(new_n20748));
  INVx1_ASAP7_75t_L         g20492(.A(new_n20748), .Y(new_n20749));
  NAND2xp33_ASAP7_75t_L     g20493(.A(new_n20741), .B(new_n20747), .Y(new_n20750));
  NAND2xp33_ASAP7_75t_L     g20494(.A(new_n20750), .B(new_n20749), .Y(new_n20751));
  O2A1O1Ixp33_ASAP7_75t_L   g20495(.A1(new_n20704), .A2(new_n20707), .B(new_n20731), .C(new_n20751), .Y(new_n20752));
  INVx1_ASAP7_75t_L         g20496(.A(new_n20752), .Y(new_n20753));
  INVx1_ASAP7_75t_L         g20497(.A(new_n20708), .Y(new_n20754));
  NAND3xp33_ASAP7_75t_L     g20498(.A(new_n20754), .B(new_n20731), .C(new_n20751), .Y(new_n20755));
  NAND2xp33_ASAP7_75t_L     g20499(.A(new_n20755), .B(new_n20753), .Y(new_n20756));
  A2O1A1Ixp33_ASAP7_75t_L   g20500(.A1(new_n12597), .A2(new_n12600), .B(new_n12628), .C(new_n10591), .Y(new_n20757));
  OAI221xp5_ASAP7_75t_L     g20501(.A1(new_n11335), .A2(new_n12599), .B1(new_n12273), .B2(new_n11330), .C(new_n20757), .Y(new_n20758));
  XNOR2x2_ASAP7_75t_L       g20502(.A(\a[59] ), .B(new_n20758), .Y(new_n20759));
  INVx1_ASAP7_75t_L         g20503(.A(new_n20759), .Y(new_n20760));
  XNOR2x2_ASAP7_75t_L       g20504(.A(new_n20760), .B(new_n20756), .Y(new_n20761));
  INVx1_ASAP7_75t_L         g20505(.A(new_n20761), .Y(new_n20762));
  NAND3xp33_ASAP7_75t_L     g20506(.A(new_n20762), .B(new_n20719), .C(new_n20717), .Y(new_n20763));
  O2A1O1Ixp33_ASAP7_75t_L   g20507(.A1(new_n20714), .A2(new_n20715), .B(new_n20719), .C(new_n20762), .Y(new_n20764));
  INVx1_ASAP7_75t_L         g20508(.A(new_n20764), .Y(new_n20765));
  AND2x2_ASAP7_75t_L        g20509(.A(new_n20763), .B(new_n20765), .Y(new_n20766));
  INVx1_ASAP7_75t_L         g20510(.A(new_n20766), .Y(new_n20767));
  A2O1A1O1Ixp25_ASAP7_75t_L g20511(.A1(new_n20680), .A2(new_n20683), .B(new_n20722), .C(new_n20724), .D(new_n20767), .Y(new_n20768));
  A2O1A1Ixp33_ASAP7_75t_L   g20512(.A1(new_n20683), .A2(new_n20680), .B(new_n20726), .C(new_n20724), .Y(new_n20769));
  NOR2xp33_ASAP7_75t_L      g20513(.A(new_n20766), .B(new_n20769), .Y(new_n20770));
  NOR2xp33_ASAP7_75t_L      g20514(.A(new_n20768), .B(new_n20770), .Y(\f[121] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20515(.A1(new_n20678), .A2(new_n20677), .B(new_n20684), .C(new_n20725), .Y(new_n20772));
  A2O1A1Ixp33_ASAP7_75t_L   g20516(.A1(new_n20772), .A2(new_n20724), .B(new_n20767), .C(new_n20765), .Y(new_n20773));
  AOI22xp33_ASAP7_75t_L     g20517(.A1(new_n11656), .A2(\b[62] ), .B1(new_n11654), .B2(new_n12280), .Y(new_n20774));
  OAI221xp5_ASAP7_75t_L     g20518(.A1(new_n12364), .A2(new_n11911), .B1(new_n11226), .B2(new_n13003), .C(new_n20774), .Y(new_n20775));
  XNOR2x2_ASAP7_75t_L       g20519(.A(\a[62] ), .B(new_n20775), .Y(new_n20776));
  A2O1A1Ixp33_ASAP7_75t_L   g20520(.A1(new_n12278), .A2(\b[61] ), .B(\b[62] ), .C(new_n10591), .Y(new_n20777));
  A2O1A1Ixp33_ASAP7_75t_L   g20521(.A1(new_n20777), .A2(new_n11330), .B(new_n12599), .C(\a[59] ), .Y(new_n20778));
  O2A1O1Ixp33_ASAP7_75t_L   g20522(.A1(new_n10974), .A2(new_n13934), .B(new_n11330), .C(new_n12599), .Y(new_n20779));
  NAND2xp33_ASAP7_75t_L     g20523(.A(new_n10588), .B(new_n20779), .Y(new_n20780));
  AND2x2_ASAP7_75t_L        g20524(.A(new_n20780), .B(new_n20778), .Y(new_n20781));
  NOR2xp33_ASAP7_75t_L      g20525(.A(new_n20781), .B(new_n20776), .Y(new_n20782));
  NAND2xp33_ASAP7_75t_L     g20526(.A(new_n20781), .B(new_n20776), .Y(new_n20783));
  INVx1_ASAP7_75t_L         g20527(.A(new_n20783), .Y(new_n20784));
  NOR2xp33_ASAP7_75t_L      g20528(.A(new_n20782), .B(new_n20784), .Y(new_n20785));
  A2O1A1O1Ixp25_ASAP7_75t_L g20529(.A1(new_n20692), .A2(new_n9610), .B(new_n20733), .C(new_n20736), .D(new_n20748), .Y(new_n20786));
  NOR2xp33_ASAP7_75t_L      g20530(.A(new_n10848), .B(new_n12671), .Y(new_n20787));
  A2O1A1Ixp33_ASAP7_75t_L   g20531(.A1(\b[59] ), .A2(new_n12669), .B(new_n20787), .C(new_n20736), .Y(new_n20788));
  O2A1O1Ixp33_ASAP7_75t_L   g20532(.A1(new_n12353), .A2(new_n12355), .B(\b[59] ), .C(new_n20787), .Y(new_n20789));
  A2O1A1Ixp33_ASAP7_75t_L   g20533(.A1(new_n12669), .A2(\b[58] ), .B(new_n20732), .C(new_n20789), .Y(new_n20790));
  NAND2xp33_ASAP7_75t_L     g20534(.A(new_n20790), .B(new_n20788), .Y(new_n20791));
  XNOR2x2_ASAP7_75t_L       g20535(.A(new_n20791), .B(new_n20786), .Y(new_n20792));
  XNOR2x2_ASAP7_75t_L       g20536(.A(new_n20785), .B(new_n20792), .Y(new_n20793));
  A2O1A1Ixp33_ASAP7_75t_L   g20537(.A1(new_n20754), .A2(new_n20731), .B(new_n20751), .C(new_n20759), .Y(new_n20794));
  NAND3xp33_ASAP7_75t_L     g20538(.A(new_n20793), .B(new_n20755), .C(new_n20794), .Y(new_n20795));
  INVx1_ASAP7_75t_L         g20539(.A(new_n20795), .Y(new_n20796));
  O2A1O1Ixp33_ASAP7_75t_L   g20540(.A1(new_n20752), .A2(new_n20760), .B(new_n20755), .C(new_n20793), .Y(new_n20797));
  NOR2xp33_ASAP7_75t_L      g20541(.A(new_n20797), .B(new_n20796), .Y(new_n20798));
  XOR2x2_ASAP7_75t_L        g20542(.A(new_n20798), .B(new_n20773), .Y(\f[122] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20543(.A1(new_n12669), .A2(\b[59] ), .B(new_n20787), .C(\a[59] ), .Y(new_n20800));
  AOI211xp5_ASAP7_75t_L     g20544(.A1(new_n12669), .A2(\b[59] ), .B(new_n20787), .C(\a[59] ), .Y(new_n20801));
  INVx1_ASAP7_75t_L         g20545(.A(new_n20801), .Y(new_n20802));
  NOR2xp33_ASAP7_75t_L      g20546(.A(new_n10881), .B(new_n12671), .Y(new_n20803));
  O2A1O1Ixp33_ASAP7_75t_L   g20547(.A1(new_n12353), .A2(new_n12355), .B(\b[60] ), .C(new_n20803), .Y(new_n20804));
  NAND3xp33_ASAP7_75t_L     g20548(.A(new_n20802), .B(new_n20800), .C(new_n20804), .Y(new_n20805));
  NAND2xp33_ASAP7_75t_L     g20549(.A(new_n20800), .B(new_n20802), .Y(new_n20806));
  A2O1A1Ixp33_ASAP7_75t_L   g20550(.A1(\b[60] ), .A2(new_n12669), .B(new_n20803), .C(new_n20806), .Y(new_n20807));
  AND2x2_ASAP7_75t_L        g20551(.A(new_n20805), .B(new_n20807), .Y(new_n20808));
  INVx1_ASAP7_75t_L         g20552(.A(new_n12603), .Y(new_n20809));
  NOR2xp33_ASAP7_75t_L      g20553(.A(new_n12599), .B(new_n12023), .Y(new_n20810));
  O2A1O1Ixp33_ASAP7_75t_L   g20554(.A1(new_n12606), .A2(new_n20809), .B(new_n11654), .C(new_n20810), .Y(new_n20811));
  OAI221xp5_ASAP7_75t_L     g20555(.A1(new_n12364), .A2(new_n12273), .B1(new_n11911), .B2(new_n13003), .C(new_n20811), .Y(new_n20812));
  NOR2xp33_ASAP7_75t_L      g20556(.A(new_n11651), .B(new_n20812), .Y(new_n20813));
  AND2x2_ASAP7_75t_L        g20557(.A(new_n11651), .B(new_n20812), .Y(new_n20814));
  NOR2xp33_ASAP7_75t_L      g20558(.A(new_n20813), .B(new_n20814), .Y(new_n20815));
  XOR2x2_ASAP7_75t_L        g20559(.A(new_n20808), .B(new_n20815), .Y(new_n20816));
  INVx1_ASAP7_75t_L         g20560(.A(new_n20786), .Y(new_n20817));
  A2O1A1O1Ixp25_ASAP7_75t_L g20561(.A1(new_n12669), .A2(\b[58] ), .B(new_n20732), .C(new_n20789), .D(new_n20817), .Y(new_n20818));
  A2O1A1O1Ixp25_ASAP7_75t_L g20562(.A1(new_n12669), .A2(\b[59] ), .B(new_n20787), .C(new_n20736), .D(new_n20818), .Y(new_n20819));
  XNOR2x2_ASAP7_75t_L       g20563(.A(new_n20816), .B(new_n20819), .Y(new_n20820));
  A2O1A1Ixp33_ASAP7_75t_L   g20564(.A1(new_n20778), .A2(new_n20780), .B(new_n20776), .C(new_n20792), .Y(new_n20821));
  NAND3xp33_ASAP7_75t_L     g20565(.A(new_n20820), .B(new_n20783), .C(new_n20821), .Y(new_n20822));
  AO21x2_ASAP7_75t_L        g20566(.A1(new_n20821), .A2(new_n20783), .B(new_n20820), .Y(new_n20823));
  AND2x2_ASAP7_75t_L        g20567(.A(new_n20822), .B(new_n20823), .Y(new_n20824));
  A2O1A1Ixp33_ASAP7_75t_L   g20568(.A1(new_n20773), .A2(new_n20798), .B(new_n20796), .C(new_n20824), .Y(new_n20825));
  A2O1A1O1Ixp25_ASAP7_75t_L g20569(.A1(new_n20766), .A2(new_n20769), .B(new_n20764), .C(new_n20798), .D(new_n20796), .Y(new_n20826));
  INVx1_ASAP7_75t_L         g20570(.A(new_n20824), .Y(new_n20827));
  NAND2xp33_ASAP7_75t_L     g20571(.A(new_n20827), .B(new_n20826), .Y(new_n20828));
  AND2x2_ASAP7_75t_L        g20572(.A(new_n20828), .B(new_n20825), .Y(\f[123] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20573(.A1(new_n20769), .A2(new_n20766), .B(new_n20764), .C(new_n20798), .Y(new_n20830));
  INVx1_ASAP7_75t_L         g20574(.A(new_n20819), .Y(new_n20831));
  NOR2xp33_ASAP7_75t_L      g20575(.A(new_n20816), .B(new_n20831), .Y(new_n20832));
  O2A1O1Ixp33_ASAP7_75t_L   g20576(.A1(new_n20813), .A2(new_n20814), .B(new_n20808), .C(new_n20832), .Y(new_n20833));
  NOR2xp33_ASAP7_75t_L      g20577(.A(new_n11226), .B(new_n12671), .Y(new_n20834));
  O2A1O1Ixp33_ASAP7_75t_L   g20578(.A1(new_n12353), .A2(new_n12355), .B(\b[61] ), .C(new_n20834), .Y(new_n20835));
  INVx1_ASAP7_75t_L         g20579(.A(new_n20835), .Y(new_n20836));
  A2O1A1Ixp33_ASAP7_75t_L   g20580(.A1(new_n12669), .A2(\b[59] ), .B(new_n20787), .C(new_n10588), .Y(new_n20837));
  A2O1A1O1Ixp25_ASAP7_75t_L g20581(.A1(new_n20800), .A2(new_n20802), .B(new_n20804), .C(new_n20837), .D(new_n20836), .Y(new_n20838));
  INVx1_ASAP7_75t_L         g20582(.A(new_n20838), .Y(new_n20839));
  INVx1_ASAP7_75t_L         g20583(.A(new_n20787), .Y(new_n20840));
  O2A1O1Ixp33_ASAP7_75t_L   g20584(.A1(new_n10881), .A2(new_n12356), .B(new_n20840), .C(\a[59] ), .Y(new_n20841));
  A2O1A1O1Ixp25_ASAP7_75t_L g20585(.A1(new_n12669), .A2(\b[60] ), .B(new_n20803), .C(new_n20806), .D(new_n20841), .Y(new_n20842));
  A2O1A1Ixp33_ASAP7_75t_L   g20586(.A1(new_n12669), .A2(\b[61] ), .B(new_n20834), .C(new_n20842), .Y(new_n20843));
  NAND2xp33_ASAP7_75t_L     g20587(.A(new_n20839), .B(new_n20843), .Y(new_n20844));
  OAI22xp33_ASAP7_75t_L     g20588(.A1(new_n13003), .A2(new_n12273), .B1(new_n12599), .B2(new_n12364), .Y(new_n20845));
  A2O1A1O1Ixp25_ASAP7_75t_L g20589(.A1(new_n12600), .A2(new_n12597), .B(new_n12628), .C(new_n11654), .D(new_n20845), .Y(new_n20846));
  NAND2xp33_ASAP7_75t_L     g20590(.A(\a[62] ), .B(new_n20846), .Y(new_n20847));
  A2O1A1Ixp33_ASAP7_75t_L   g20591(.A1(new_n19739), .A2(new_n11654), .B(new_n20845), .C(new_n11651), .Y(new_n20848));
  AO21x2_ASAP7_75t_L        g20592(.A1(new_n20847), .A2(new_n20848), .B(new_n20844), .Y(new_n20849));
  NAND3xp33_ASAP7_75t_L     g20593(.A(new_n20848), .B(new_n20847), .C(new_n20844), .Y(new_n20850));
  AND2x2_ASAP7_75t_L        g20594(.A(new_n20850), .B(new_n20849), .Y(new_n20851));
  INVx1_ASAP7_75t_L         g20595(.A(new_n20851), .Y(new_n20852));
  NOR2xp33_ASAP7_75t_L      g20596(.A(new_n20852), .B(new_n20833), .Y(new_n20853));
  INVx1_ASAP7_75t_L         g20597(.A(new_n20853), .Y(new_n20854));
  NAND2xp33_ASAP7_75t_L     g20598(.A(new_n20852), .B(new_n20833), .Y(new_n20855));
  AND2x2_ASAP7_75t_L        g20599(.A(new_n20855), .B(new_n20854), .Y(new_n20856));
  INVx1_ASAP7_75t_L         g20600(.A(new_n20856), .Y(new_n20857));
  A2O1A1O1Ixp25_ASAP7_75t_L g20601(.A1(new_n20795), .A2(new_n20830), .B(new_n20827), .C(new_n20822), .D(new_n20857), .Y(new_n20858));
  A2O1A1Ixp33_ASAP7_75t_L   g20602(.A1(new_n20830), .A2(new_n20795), .B(new_n20827), .C(new_n20822), .Y(new_n20859));
  NOR2xp33_ASAP7_75t_L      g20603(.A(new_n20856), .B(new_n20859), .Y(new_n20860));
  NOR2xp33_ASAP7_75t_L      g20604(.A(new_n20858), .B(new_n20860), .Y(\f[124] ));
  NAND2xp33_ASAP7_75t_L     g20605(.A(\b[61] ), .B(new_n12670), .Y(new_n20862));
  O2A1O1Ixp33_ASAP7_75t_L   g20606(.A1(new_n12356), .A2(new_n12273), .B(new_n20862), .C(new_n20836), .Y(new_n20863));
  INVx1_ASAP7_75t_L         g20607(.A(new_n20834), .Y(new_n20864));
  A2O1A1Ixp33_ASAP7_75t_L   g20608(.A1(new_n19241), .A2(new_n19242), .B(new_n12273), .C(new_n20862), .Y(new_n20865));
  O2A1O1Ixp33_ASAP7_75t_L   g20609(.A1(new_n11911), .A2(new_n12356), .B(new_n20864), .C(new_n20865), .Y(new_n20866));
  NOR2xp33_ASAP7_75t_L      g20610(.A(new_n20866), .B(new_n20863), .Y(new_n20867));
  O2A1O1Ixp33_ASAP7_75t_L   g20611(.A1(new_n11911), .A2(new_n12604), .B(new_n12273), .C(new_n12022), .Y(new_n20868));
  O2A1O1Ixp33_ASAP7_75t_L   g20612(.A1(new_n12021), .A2(new_n20868), .B(\b[63] ), .C(new_n11651), .Y(new_n20869));
  A2O1A1O1Ixp25_ASAP7_75t_L g20613(.A1(\b[61] ), .A2(new_n12278), .B(\b[62] ), .C(new_n11654), .D(new_n12021), .Y(new_n20870));
  NOR3xp33_ASAP7_75t_L      g20614(.A(new_n20870), .B(new_n12599), .C(\a[62] ), .Y(new_n20871));
  NOR2xp33_ASAP7_75t_L      g20615(.A(new_n20869), .B(new_n20871), .Y(new_n20872));
  XOR2x2_ASAP7_75t_L        g20616(.A(new_n20867), .B(new_n20872), .Y(new_n20873));
  O2A1O1Ixp33_ASAP7_75t_L   g20617(.A1(new_n20836), .A2(new_n20842), .B(new_n20849), .C(new_n20873), .Y(new_n20874));
  AND3x1_ASAP7_75t_L        g20618(.A(new_n20873), .B(new_n20849), .C(new_n20839), .Y(new_n20875));
  NOR2xp33_ASAP7_75t_L      g20619(.A(new_n20874), .B(new_n20875), .Y(new_n20876));
  INVx1_ASAP7_75t_L         g20620(.A(new_n20876), .Y(new_n20877));
  A2O1A1O1Ixp25_ASAP7_75t_L g20621(.A1(new_n20822), .A2(new_n20825), .B(new_n20857), .C(new_n20854), .D(new_n20877), .Y(new_n20878));
  A2O1A1Ixp33_ASAP7_75t_L   g20622(.A1(new_n20825), .A2(new_n20822), .B(new_n20857), .C(new_n20854), .Y(new_n20879));
  NOR2xp33_ASAP7_75t_L      g20623(.A(new_n20876), .B(new_n20879), .Y(new_n20880));
  NOR2xp33_ASAP7_75t_L      g20624(.A(new_n20878), .B(new_n20880), .Y(\f[125] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g20625(.A1(new_n20856), .A2(new_n20859), .B(new_n20853), .C(new_n20876), .D(new_n20874), .Y(new_n20882));
  O2A1O1Ixp33_ASAP7_75t_L   g20626(.A1(new_n20869), .A2(new_n20871), .B(new_n20867), .C(new_n20863), .Y(new_n20883));
  NOR2xp33_ASAP7_75t_L      g20627(.A(new_n12354), .B(new_n12599), .Y(new_n20884));
  INVx1_ASAP7_75t_L         g20628(.A(new_n20884), .Y(new_n20885));
  NOR3xp33_ASAP7_75t_L      g20629(.A(new_n11651), .B(new_n12354), .C(new_n12273), .Y(new_n20886));
  O2A1O1Ixp33_ASAP7_75t_L   g20630(.A1(new_n11651), .A2(\b[63] ), .B(new_n20885), .C(new_n20886), .Y(new_n20887));
  O2A1O1Ixp33_ASAP7_75t_L   g20631(.A1(new_n11911), .A2(new_n12356), .B(new_n20864), .C(new_n20887), .Y(new_n20888));
  AND2x2_ASAP7_75t_L        g20632(.A(new_n20887), .B(new_n20835), .Y(new_n20889));
  OR3x1_ASAP7_75t_L         g20633(.A(new_n20883), .B(new_n20888), .C(new_n20889), .Y(new_n20890));
  OAI21xp33_ASAP7_75t_L     g20634(.A1(new_n20888), .A2(new_n20889), .B(new_n20883), .Y(new_n20891));
  NAND2xp33_ASAP7_75t_L     g20635(.A(new_n20891), .B(new_n20890), .Y(new_n20892));
  XOR2x2_ASAP7_75t_L        g20636(.A(new_n20892), .B(new_n20882), .Y(\f[126] ));
  XNOR2x2_ASAP7_75t_L       g20637(.A(new_n20885), .B(new_n20888), .Y(new_n20894));
  OA211x2_ASAP7_75t_L       g20638(.A1(new_n20892), .A2(new_n20882), .B(new_n20890), .C(new_n20894), .Y(new_n20895));
  O2A1O1Ixp33_ASAP7_75t_L   g20639(.A1(new_n20892), .A2(new_n20882), .B(new_n20890), .C(new_n20894), .Y(new_n20896));
  NOR2xp33_ASAP7_75t_L      g20640(.A(new_n20896), .B(new_n20895), .Y(\f[127] ));
endmodule


