// Benchmark "top" written by ABC on Mon Dec 25 16:58:17 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386, new_n387, new_n388, new_n390, new_n391, new_n392, new_n393,
    new_n395, new_n396, new_n397, new_n398, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1369;
  NAND2xp33_ASAP7_75t_L     g000(.A(\b[0] ), .B(\a[0] ), .Y(new_n386));
  INVx1_ASAP7_75t_L         g001(.A(new_n386), .Y(new_n387));
  NOR2xp33_ASAP7_75t_L      g002(.A(\a[0] ), .B(\b[0] ), .Y(new_n388));
  NOR2xp33_ASAP7_75t_L      g003(.A(new_n388), .B(new_n387), .Y(\f[0] ));
  NOR2xp33_ASAP7_75t_L      g004(.A(\a[1] ), .B(\b[1] ), .Y(new_n390));
  NAND2xp33_ASAP7_75t_L     g005(.A(\b[1] ), .B(\a[1] ), .Y(new_n391));
  INVx1_ASAP7_75t_L         g006(.A(new_n391), .Y(new_n392));
  NOR2xp33_ASAP7_75t_L      g007(.A(new_n390), .B(new_n392), .Y(new_n393));
  XNOR2x2_ASAP7_75t_L       g008(.A(new_n386), .B(new_n393), .Y(\f[1] ));
  XNOR2x2_ASAP7_75t_L       g009(.A(\b[2] ), .B(\a[2] ), .Y(new_n395));
  OAI211xp5_ASAP7_75t_L     g010(.A1(new_n386), .A2(new_n390), .B(new_n395), .C(new_n391), .Y(new_n396));
  O2A1O1Ixp33_ASAP7_75t_L   g011(.A1(new_n386), .A2(new_n390), .B(new_n391), .C(new_n395), .Y(new_n397));
  INVx1_ASAP7_75t_L         g012(.A(new_n397), .Y(new_n398));
  AND2x2_ASAP7_75t_L        g013(.A(new_n396), .B(new_n398), .Y(\f[2] ));
  NAND2xp33_ASAP7_75t_L     g014(.A(\b[2] ), .B(\a[2] ), .Y(new_n400));
  NOR2xp33_ASAP7_75t_L      g015(.A(\a[3] ), .B(\b[3] ), .Y(new_n401));
  NAND2xp33_ASAP7_75t_L     g016(.A(\b[3] ), .B(\a[3] ), .Y(new_n402));
  INVx1_ASAP7_75t_L         g017(.A(new_n402), .Y(new_n403));
  OAI211xp5_ASAP7_75t_L     g018(.A1(new_n401), .A2(new_n403), .B(new_n398), .C(new_n400), .Y(new_n404));
  NOR2xp33_ASAP7_75t_L      g019(.A(new_n401), .B(new_n403), .Y(new_n405));
  A2O1A1Ixp33_ASAP7_75t_L   g020(.A1(\b[2] ), .A2(\a[2] ), .B(new_n397), .C(new_n405), .Y(new_n406));
  AND2x2_ASAP7_75t_L        g021(.A(new_n406), .B(new_n404), .Y(\f[3] ));
  NOR2xp33_ASAP7_75t_L      g022(.A(\a[4] ), .B(\b[4] ), .Y(new_n408));
  INVx1_ASAP7_75t_L         g023(.A(new_n408), .Y(new_n409));
  NAND2xp33_ASAP7_75t_L     g024(.A(\b[4] ), .B(\a[4] ), .Y(new_n410));
  A2O1A1Ixp33_ASAP7_75t_L   g025(.A1(new_n398), .A2(new_n400), .B(new_n401), .C(new_n402), .Y(new_n411));
  AOI21xp33_ASAP7_75t_L     g026(.A1(new_n410), .A2(new_n409), .B(new_n411), .Y(new_n412));
  NAND2xp33_ASAP7_75t_L     g027(.A(new_n410), .B(new_n409), .Y(new_n413));
  A2O1A1O1Ixp25_ASAP7_75t_L g028(.A1(new_n400), .A2(new_n398), .B(new_n401), .C(new_n402), .D(new_n413), .Y(new_n414));
  NOR2xp33_ASAP7_75t_L      g029(.A(new_n414), .B(new_n412), .Y(\f[4] ));
  NOR2xp33_ASAP7_75t_L      g030(.A(\a[5] ), .B(\b[5] ), .Y(new_n416));
  INVx1_ASAP7_75t_L         g031(.A(\a[5] ), .Y(new_n417));
  INVx1_ASAP7_75t_L         g032(.A(\b[5] ), .Y(new_n418));
  NOR2xp33_ASAP7_75t_L      g033(.A(new_n417), .B(new_n418), .Y(new_n419));
  NOR2xp33_ASAP7_75t_L      g034(.A(new_n416), .B(new_n419), .Y(new_n420));
  A2O1A1Ixp33_ASAP7_75t_L   g035(.A1(new_n406), .A2(new_n402), .B(new_n408), .C(new_n410), .Y(new_n421));
  NOR2xp33_ASAP7_75t_L      g036(.A(new_n420), .B(new_n421), .Y(new_n422));
  A2O1A1Ixp33_ASAP7_75t_L   g037(.A1(\b[4] ), .A2(\a[4] ), .B(new_n414), .C(new_n420), .Y(new_n423));
  INVx1_ASAP7_75t_L         g038(.A(new_n423), .Y(new_n424));
  NOR2xp33_ASAP7_75t_L      g039(.A(new_n422), .B(new_n424), .Y(\f[5] ));
  NOR2xp33_ASAP7_75t_L      g040(.A(\a[6] ), .B(\b[6] ), .Y(new_n426));
  AND2x2_ASAP7_75t_L        g041(.A(\a[6] ), .B(\b[6] ), .Y(new_n427));
  NOR2xp33_ASAP7_75t_L      g042(.A(new_n426), .B(new_n427), .Y(new_n428));
  INVx1_ASAP7_75t_L         g043(.A(new_n414), .Y(new_n429));
  INVx1_ASAP7_75t_L         g044(.A(new_n419), .Y(new_n430));
  A2O1A1Ixp33_ASAP7_75t_L   g045(.A1(new_n429), .A2(new_n410), .B(new_n416), .C(new_n430), .Y(new_n431));
  NOR2xp33_ASAP7_75t_L      g046(.A(new_n428), .B(new_n431), .Y(new_n432));
  INVx1_ASAP7_75t_L         g047(.A(new_n428), .Y(new_n433));
  A2O1A1O1Ixp25_ASAP7_75t_L g048(.A1(new_n410), .A2(new_n429), .B(new_n416), .C(new_n430), .D(new_n433), .Y(new_n434));
  NOR2xp33_ASAP7_75t_L      g049(.A(new_n434), .B(new_n432), .Y(\f[6] ));
  INVx1_ASAP7_75t_L         g050(.A(\a[7] ), .Y(new_n436));
  INVx1_ASAP7_75t_L         g051(.A(\b[7] ), .Y(new_n437));
  NAND2xp33_ASAP7_75t_L     g052(.A(new_n437), .B(new_n436), .Y(new_n438));
  NOR2xp33_ASAP7_75t_L      g053(.A(new_n436), .B(new_n437), .Y(new_n439));
  INVx1_ASAP7_75t_L         g054(.A(new_n439), .Y(new_n440));
  AND2x2_ASAP7_75t_L        g055(.A(new_n438), .B(new_n440), .Y(new_n441));
  A2O1A1O1Ixp25_ASAP7_75t_L g056(.A1(new_n420), .A2(new_n421), .B(new_n419), .C(new_n428), .D(new_n427), .Y(new_n442));
  XNOR2x2_ASAP7_75t_L       g057(.A(new_n441), .B(new_n442), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g058(.A(\a[8] ), .B(\b[8] ), .Y(new_n444));
  INVx1_ASAP7_75t_L         g059(.A(\a[8] ), .Y(new_n445));
  INVx1_ASAP7_75t_L         g060(.A(\b[8] ), .Y(new_n446));
  NOR2xp33_ASAP7_75t_L      g061(.A(new_n445), .B(new_n446), .Y(new_n447));
  NOR2xp33_ASAP7_75t_L      g062(.A(new_n444), .B(new_n447), .Y(new_n448));
  INVx1_ASAP7_75t_L         g063(.A(new_n448), .Y(new_n449));
  A2O1A1O1Ixp25_ASAP7_75t_L g064(.A1(new_n428), .A2(new_n431), .B(new_n427), .C(new_n438), .D(new_n439), .Y(new_n450));
  AND2x2_ASAP7_75t_L        g065(.A(new_n449), .B(new_n450), .Y(new_n451));
  A2O1A1Ixp33_ASAP7_75t_L   g066(.A1(new_n431), .A2(new_n428), .B(new_n427), .C(new_n441), .Y(new_n452));
  O2A1O1Ixp33_ASAP7_75t_L   g067(.A1(new_n436), .A2(new_n437), .B(new_n452), .C(new_n449), .Y(new_n453));
  NOR2xp33_ASAP7_75t_L      g068(.A(new_n453), .B(new_n451), .Y(\f[8] ));
  NOR2xp33_ASAP7_75t_L      g069(.A(\a[9] ), .B(\b[9] ), .Y(new_n455));
  INVx1_ASAP7_75t_L         g070(.A(\a[9] ), .Y(new_n456));
  INVx1_ASAP7_75t_L         g071(.A(\b[9] ), .Y(new_n457));
  NOR2xp33_ASAP7_75t_L      g072(.A(new_n456), .B(new_n457), .Y(new_n458));
  NOR2xp33_ASAP7_75t_L      g073(.A(new_n455), .B(new_n458), .Y(new_n459));
  INVx1_ASAP7_75t_L         g074(.A(new_n447), .Y(new_n460));
  A2O1A1Ixp33_ASAP7_75t_L   g075(.A1(new_n452), .A2(new_n440), .B(new_n444), .C(new_n460), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g076(.A(new_n459), .B(new_n461), .Y(new_n462));
  A2O1A1Ixp33_ASAP7_75t_L   g077(.A1(\b[8] ), .A2(\a[8] ), .B(new_n453), .C(new_n459), .Y(new_n463));
  INVx1_ASAP7_75t_L         g078(.A(new_n463), .Y(new_n464));
  NOR2xp33_ASAP7_75t_L      g079(.A(new_n462), .B(new_n464), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g080(.A(\a[10] ), .B(\b[10] ), .Y(new_n466));
  INVx1_ASAP7_75t_L         g081(.A(\a[10] ), .Y(new_n467));
  INVx1_ASAP7_75t_L         g082(.A(\b[10] ), .Y(new_n468));
  NOR2xp33_ASAP7_75t_L      g083(.A(new_n467), .B(new_n468), .Y(new_n469));
  NOR2xp33_ASAP7_75t_L      g084(.A(new_n466), .B(new_n469), .Y(new_n470));
  INVx1_ASAP7_75t_L         g085(.A(new_n453), .Y(new_n471));
  INVx1_ASAP7_75t_L         g086(.A(new_n458), .Y(new_n472));
  A2O1A1Ixp33_ASAP7_75t_L   g087(.A1(new_n471), .A2(new_n460), .B(new_n455), .C(new_n472), .Y(new_n473));
  NOR2xp33_ASAP7_75t_L      g088(.A(new_n470), .B(new_n473), .Y(new_n474));
  INVx1_ASAP7_75t_L         g089(.A(new_n470), .Y(new_n475));
  A2O1A1O1Ixp25_ASAP7_75t_L g090(.A1(new_n460), .A2(new_n471), .B(new_n455), .C(new_n472), .D(new_n475), .Y(new_n476));
  NOR2xp33_ASAP7_75t_L      g091(.A(new_n476), .B(new_n474), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g092(.A(\a[11] ), .B(\b[11] ), .Y(new_n478));
  INVx1_ASAP7_75t_L         g093(.A(\a[11] ), .Y(new_n479));
  INVx1_ASAP7_75t_L         g094(.A(\b[11] ), .Y(new_n480));
  NOR2xp33_ASAP7_75t_L      g095(.A(new_n479), .B(new_n480), .Y(new_n481));
  NOR2xp33_ASAP7_75t_L      g096(.A(new_n478), .B(new_n481), .Y(new_n482));
  INVx1_ASAP7_75t_L         g097(.A(new_n469), .Y(new_n483));
  A2O1A1Ixp33_ASAP7_75t_L   g098(.A1(new_n463), .A2(new_n472), .B(new_n466), .C(new_n483), .Y(new_n484));
  NOR2xp33_ASAP7_75t_L      g099(.A(new_n482), .B(new_n484), .Y(new_n485));
  A2O1A1Ixp33_ASAP7_75t_L   g100(.A1(new_n473), .A2(new_n470), .B(new_n469), .C(new_n482), .Y(new_n486));
  INVx1_ASAP7_75t_L         g101(.A(new_n486), .Y(new_n487));
  NOR2xp33_ASAP7_75t_L      g102(.A(new_n485), .B(new_n487), .Y(\f[11] ));
  NOR2xp33_ASAP7_75t_L      g103(.A(\a[12] ), .B(\b[12] ), .Y(new_n489));
  AND2x2_ASAP7_75t_L        g104(.A(\a[12] ), .B(\b[12] ), .Y(new_n490));
  NOR2xp33_ASAP7_75t_L      g105(.A(new_n489), .B(new_n490), .Y(new_n491));
  NOR3xp33_ASAP7_75t_L      g106(.A(new_n487), .B(new_n491), .C(new_n481), .Y(new_n492));
  INVx1_ASAP7_75t_L         g107(.A(new_n491), .Y(new_n493));
  O2A1O1Ixp33_ASAP7_75t_L   g108(.A1(new_n479), .A2(new_n480), .B(new_n486), .C(new_n493), .Y(new_n494));
  NOR2xp33_ASAP7_75t_L      g109(.A(new_n494), .B(new_n492), .Y(\f[12] ));
  NOR2xp33_ASAP7_75t_L      g110(.A(\a[13] ), .B(\b[13] ), .Y(new_n496));
  INVx1_ASAP7_75t_L         g111(.A(\a[13] ), .Y(new_n497));
  INVx1_ASAP7_75t_L         g112(.A(\b[13] ), .Y(new_n498));
  NOR2xp33_ASAP7_75t_L      g113(.A(new_n497), .B(new_n498), .Y(new_n499));
  NOR2xp33_ASAP7_75t_L      g114(.A(new_n496), .B(new_n499), .Y(new_n500));
  A2O1A1O1Ixp25_ASAP7_75t_L g115(.A1(new_n482), .A2(new_n484), .B(new_n481), .C(new_n491), .D(new_n490), .Y(new_n501));
  XNOR2x2_ASAP7_75t_L       g116(.A(new_n500), .B(new_n501), .Y(\f[13] ));
  NOR2xp33_ASAP7_75t_L      g117(.A(\a[14] ), .B(\b[14] ), .Y(new_n503));
  AND2x2_ASAP7_75t_L        g118(.A(\a[14] ), .B(\b[14] ), .Y(new_n504));
  NOR2xp33_ASAP7_75t_L      g119(.A(new_n503), .B(new_n504), .Y(new_n505));
  INVx1_ASAP7_75t_L         g120(.A(new_n505), .Y(new_n506));
  O2A1O1Ixp33_ASAP7_75t_L   g121(.A1(new_n490), .A2(new_n494), .B(new_n500), .C(new_n499), .Y(new_n507));
  AND2x2_ASAP7_75t_L        g122(.A(new_n506), .B(new_n507), .Y(new_n508));
  A2O1A1Ixp33_ASAP7_75t_L   g123(.A1(\b[12] ), .A2(\a[12] ), .B(new_n494), .C(new_n500), .Y(new_n509));
  O2A1O1Ixp33_ASAP7_75t_L   g124(.A1(new_n497), .A2(new_n498), .B(new_n509), .C(new_n506), .Y(new_n510));
  NOR2xp33_ASAP7_75t_L      g125(.A(new_n510), .B(new_n508), .Y(\f[14] ));
  NOR2xp33_ASAP7_75t_L      g126(.A(\a[15] ), .B(\b[15] ), .Y(new_n512));
  INVx1_ASAP7_75t_L         g127(.A(\a[15] ), .Y(new_n513));
  INVx1_ASAP7_75t_L         g128(.A(\b[15] ), .Y(new_n514));
  NOR2xp33_ASAP7_75t_L      g129(.A(new_n513), .B(new_n514), .Y(new_n515));
  NOR2xp33_ASAP7_75t_L      g130(.A(new_n512), .B(new_n515), .Y(new_n516));
  OR3x1_ASAP7_75t_L         g131(.A(new_n510), .B(new_n504), .C(new_n516), .Y(new_n517));
  A2O1A1Ixp33_ASAP7_75t_L   g132(.A1(\b[14] ), .A2(\a[14] ), .B(new_n510), .C(new_n516), .Y(new_n518));
  AND2x2_ASAP7_75t_L        g133(.A(new_n518), .B(new_n517), .Y(\f[15] ));
  NOR2xp33_ASAP7_75t_L      g134(.A(\a[16] ), .B(\b[16] ), .Y(new_n520));
  AND2x2_ASAP7_75t_L        g135(.A(\a[16] ), .B(\b[16] ), .Y(new_n521));
  NOR2xp33_ASAP7_75t_L      g136(.A(new_n520), .B(new_n521), .Y(new_n522));
  INVx1_ASAP7_75t_L         g137(.A(new_n522), .Y(new_n523));
  O2A1O1Ixp33_ASAP7_75t_L   g138(.A1(new_n504), .A2(new_n510), .B(new_n516), .C(new_n515), .Y(new_n524));
  AND2x2_ASAP7_75t_L        g139(.A(new_n523), .B(new_n524), .Y(new_n525));
  O2A1O1Ixp33_ASAP7_75t_L   g140(.A1(new_n513), .A2(new_n514), .B(new_n518), .C(new_n523), .Y(new_n526));
  NOR2xp33_ASAP7_75t_L      g141(.A(new_n526), .B(new_n525), .Y(\f[16] ));
  NOR2xp33_ASAP7_75t_L      g142(.A(\a[17] ), .B(\b[17] ), .Y(new_n528));
  INVx1_ASAP7_75t_L         g143(.A(\a[17] ), .Y(new_n529));
  INVx1_ASAP7_75t_L         g144(.A(\b[17] ), .Y(new_n530));
  NOR2xp33_ASAP7_75t_L      g145(.A(new_n529), .B(new_n530), .Y(new_n531));
  NOR2xp33_ASAP7_75t_L      g146(.A(new_n528), .B(new_n531), .Y(new_n532));
  OR3x1_ASAP7_75t_L         g147(.A(new_n526), .B(new_n521), .C(new_n532), .Y(new_n533));
  A2O1A1Ixp33_ASAP7_75t_L   g148(.A1(\b[16] ), .A2(\a[16] ), .B(new_n526), .C(new_n532), .Y(new_n534));
  AND2x2_ASAP7_75t_L        g149(.A(new_n534), .B(new_n533), .Y(\f[17] ));
  NOR2xp33_ASAP7_75t_L      g150(.A(\a[18] ), .B(\b[18] ), .Y(new_n536));
  AND2x2_ASAP7_75t_L        g151(.A(\a[18] ), .B(\b[18] ), .Y(new_n537));
  NOR2xp33_ASAP7_75t_L      g152(.A(new_n536), .B(new_n537), .Y(new_n538));
  INVx1_ASAP7_75t_L         g153(.A(new_n538), .Y(new_n539));
  O2A1O1Ixp33_ASAP7_75t_L   g154(.A1(new_n521), .A2(new_n526), .B(new_n532), .C(new_n531), .Y(new_n540));
  AND2x2_ASAP7_75t_L        g155(.A(new_n539), .B(new_n540), .Y(new_n541));
  O2A1O1Ixp33_ASAP7_75t_L   g156(.A1(new_n529), .A2(new_n530), .B(new_n534), .C(new_n539), .Y(new_n542));
  NOR2xp33_ASAP7_75t_L      g157(.A(new_n542), .B(new_n541), .Y(\f[18] ));
  NOR2xp33_ASAP7_75t_L      g158(.A(\a[19] ), .B(\b[19] ), .Y(new_n544));
  INVx1_ASAP7_75t_L         g159(.A(\a[19] ), .Y(new_n545));
  INVx1_ASAP7_75t_L         g160(.A(\b[19] ), .Y(new_n546));
  NOR2xp33_ASAP7_75t_L      g161(.A(new_n545), .B(new_n546), .Y(new_n547));
  NOR2xp33_ASAP7_75t_L      g162(.A(new_n544), .B(new_n547), .Y(new_n548));
  OR3x1_ASAP7_75t_L         g163(.A(new_n542), .B(new_n537), .C(new_n548), .Y(new_n549));
  A2O1A1Ixp33_ASAP7_75t_L   g164(.A1(\b[18] ), .A2(\a[18] ), .B(new_n542), .C(new_n548), .Y(new_n550));
  AND2x2_ASAP7_75t_L        g165(.A(new_n550), .B(new_n549), .Y(\f[19] ));
  NOR2xp33_ASAP7_75t_L      g166(.A(\a[20] ), .B(\b[20] ), .Y(new_n552));
  AND2x2_ASAP7_75t_L        g167(.A(\a[20] ), .B(\b[20] ), .Y(new_n553));
  NOR2xp33_ASAP7_75t_L      g168(.A(new_n552), .B(new_n553), .Y(new_n554));
  INVx1_ASAP7_75t_L         g169(.A(new_n554), .Y(new_n555));
  O2A1O1Ixp33_ASAP7_75t_L   g170(.A1(new_n537), .A2(new_n542), .B(new_n548), .C(new_n547), .Y(new_n556));
  AND2x2_ASAP7_75t_L        g171(.A(new_n555), .B(new_n556), .Y(new_n557));
  O2A1O1Ixp33_ASAP7_75t_L   g172(.A1(new_n545), .A2(new_n546), .B(new_n550), .C(new_n555), .Y(new_n558));
  NOR2xp33_ASAP7_75t_L      g173(.A(new_n558), .B(new_n557), .Y(\f[20] ));
  NOR2xp33_ASAP7_75t_L      g174(.A(\a[21] ), .B(\b[21] ), .Y(new_n560));
  INVx1_ASAP7_75t_L         g175(.A(\a[21] ), .Y(new_n561));
  INVx1_ASAP7_75t_L         g176(.A(\b[21] ), .Y(new_n562));
  NOR2xp33_ASAP7_75t_L      g177(.A(new_n561), .B(new_n562), .Y(new_n563));
  NOR2xp33_ASAP7_75t_L      g178(.A(new_n560), .B(new_n563), .Y(new_n564));
  OR3x1_ASAP7_75t_L         g179(.A(new_n558), .B(new_n553), .C(new_n564), .Y(new_n565));
  A2O1A1Ixp33_ASAP7_75t_L   g180(.A1(\b[20] ), .A2(\a[20] ), .B(new_n558), .C(new_n564), .Y(new_n566));
  AND2x2_ASAP7_75t_L        g181(.A(new_n566), .B(new_n565), .Y(\f[21] ));
  NOR2xp33_ASAP7_75t_L      g182(.A(\a[22] ), .B(\b[22] ), .Y(new_n568));
  AND2x2_ASAP7_75t_L        g183(.A(\a[22] ), .B(\b[22] ), .Y(new_n569));
  NOR2xp33_ASAP7_75t_L      g184(.A(new_n568), .B(new_n569), .Y(new_n570));
  INVx1_ASAP7_75t_L         g185(.A(new_n570), .Y(new_n571));
  O2A1O1Ixp33_ASAP7_75t_L   g186(.A1(new_n553), .A2(new_n558), .B(new_n564), .C(new_n563), .Y(new_n572));
  AND2x2_ASAP7_75t_L        g187(.A(new_n571), .B(new_n572), .Y(new_n573));
  O2A1O1Ixp33_ASAP7_75t_L   g188(.A1(new_n561), .A2(new_n562), .B(new_n566), .C(new_n571), .Y(new_n574));
  NOR2xp33_ASAP7_75t_L      g189(.A(new_n574), .B(new_n573), .Y(\f[22] ));
  NOR2xp33_ASAP7_75t_L      g190(.A(\a[23] ), .B(\b[23] ), .Y(new_n576));
  INVx1_ASAP7_75t_L         g191(.A(\a[23] ), .Y(new_n577));
  INVx1_ASAP7_75t_L         g192(.A(\b[23] ), .Y(new_n578));
  NOR2xp33_ASAP7_75t_L      g193(.A(new_n577), .B(new_n578), .Y(new_n579));
  NOR2xp33_ASAP7_75t_L      g194(.A(new_n576), .B(new_n579), .Y(new_n580));
  OR3x1_ASAP7_75t_L         g195(.A(new_n574), .B(new_n569), .C(new_n580), .Y(new_n581));
  A2O1A1Ixp33_ASAP7_75t_L   g196(.A1(\b[22] ), .A2(\a[22] ), .B(new_n574), .C(new_n580), .Y(new_n582));
  AND2x2_ASAP7_75t_L        g197(.A(new_n582), .B(new_n581), .Y(\f[23] ));
  NOR2xp33_ASAP7_75t_L      g198(.A(\a[24] ), .B(\b[24] ), .Y(new_n584));
  AND2x2_ASAP7_75t_L        g199(.A(\a[24] ), .B(\b[24] ), .Y(new_n585));
  NOR2xp33_ASAP7_75t_L      g200(.A(new_n584), .B(new_n585), .Y(new_n586));
  INVx1_ASAP7_75t_L         g201(.A(new_n586), .Y(new_n587));
  O2A1O1Ixp33_ASAP7_75t_L   g202(.A1(new_n569), .A2(new_n574), .B(new_n580), .C(new_n579), .Y(new_n588));
  AND2x2_ASAP7_75t_L        g203(.A(new_n587), .B(new_n588), .Y(new_n589));
  O2A1O1Ixp33_ASAP7_75t_L   g204(.A1(new_n577), .A2(new_n578), .B(new_n582), .C(new_n587), .Y(new_n590));
  NOR2xp33_ASAP7_75t_L      g205(.A(new_n590), .B(new_n589), .Y(\f[24] ));
  NOR2xp33_ASAP7_75t_L      g206(.A(\a[25] ), .B(\b[25] ), .Y(new_n592));
  INVx1_ASAP7_75t_L         g207(.A(\a[25] ), .Y(new_n593));
  INVx1_ASAP7_75t_L         g208(.A(\b[25] ), .Y(new_n594));
  NOR2xp33_ASAP7_75t_L      g209(.A(new_n593), .B(new_n594), .Y(new_n595));
  NOR2xp33_ASAP7_75t_L      g210(.A(new_n592), .B(new_n595), .Y(new_n596));
  OR3x1_ASAP7_75t_L         g211(.A(new_n590), .B(new_n585), .C(new_n596), .Y(new_n597));
  A2O1A1Ixp33_ASAP7_75t_L   g212(.A1(\b[24] ), .A2(\a[24] ), .B(new_n590), .C(new_n596), .Y(new_n598));
  AND2x2_ASAP7_75t_L        g213(.A(new_n598), .B(new_n597), .Y(\f[25] ));
  NOR2xp33_ASAP7_75t_L      g214(.A(\a[26] ), .B(\b[26] ), .Y(new_n600));
  AND2x2_ASAP7_75t_L        g215(.A(\a[26] ), .B(\b[26] ), .Y(new_n601));
  NOR2xp33_ASAP7_75t_L      g216(.A(new_n600), .B(new_n601), .Y(new_n602));
  INVx1_ASAP7_75t_L         g217(.A(new_n602), .Y(new_n603));
  O2A1O1Ixp33_ASAP7_75t_L   g218(.A1(new_n585), .A2(new_n590), .B(new_n596), .C(new_n595), .Y(new_n604));
  AND2x2_ASAP7_75t_L        g219(.A(new_n603), .B(new_n604), .Y(new_n605));
  O2A1O1Ixp33_ASAP7_75t_L   g220(.A1(new_n593), .A2(new_n594), .B(new_n598), .C(new_n603), .Y(new_n606));
  NOR2xp33_ASAP7_75t_L      g221(.A(new_n606), .B(new_n605), .Y(\f[26] ));
  NOR2xp33_ASAP7_75t_L      g222(.A(\a[27] ), .B(\b[27] ), .Y(new_n608));
  INVx1_ASAP7_75t_L         g223(.A(\a[27] ), .Y(new_n609));
  INVx1_ASAP7_75t_L         g224(.A(\b[27] ), .Y(new_n610));
  NOR2xp33_ASAP7_75t_L      g225(.A(new_n609), .B(new_n610), .Y(new_n611));
  NOR2xp33_ASAP7_75t_L      g226(.A(new_n608), .B(new_n611), .Y(new_n612));
  OR3x1_ASAP7_75t_L         g227(.A(new_n606), .B(new_n601), .C(new_n612), .Y(new_n613));
  A2O1A1Ixp33_ASAP7_75t_L   g228(.A1(\b[26] ), .A2(\a[26] ), .B(new_n606), .C(new_n612), .Y(new_n614));
  AND2x2_ASAP7_75t_L        g229(.A(new_n614), .B(new_n613), .Y(\f[27] ));
  NOR2xp33_ASAP7_75t_L      g230(.A(\a[28] ), .B(\b[28] ), .Y(new_n616));
  AND2x2_ASAP7_75t_L        g231(.A(\a[28] ), .B(\b[28] ), .Y(new_n617));
  NOR2xp33_ASAP7_75t_L      g232(.A(new_n616), .B(new_n617), .Y(new_n618));
  INVx1_ASAP7_75t_L         g233(.A(new_n618), .Y(new_n619));
  O2A1O1Ixp33_ASAP7_75t_L   g234(.A1(new_n601), .A2(new_n606), .B(new_n612), .C(new_n611), .Y(new_n620));
  AND2x2_ASAP7_75t_L        g235(.A(new_n619), .B(new_n620), .Y(new_n621));
  O2A1O1Ixp33_ASAP7_75t_L   g236(.A1(new_n609), .A2(new_n610), .B(new_n614), .C(new_n619), .Y(new_n622));
  NOR2xp33_ASAP7_75t_L      g237(.A(new_n622), .B(new_n621), .Y(\f[28] ));
  NOR2xp33_ASAP7_75t_L      g238(.A(\a[29] ), .B(\b[29] ), .Y(new_n624));
  INVx1_ASAP7_75t_L         g239(.A(\a[29] ), .Y(new_n625));
  INVx1_ASAP7_75t_L         g240(.A(\b[29] ), .Y(new_n626));
  NOR2xp33_ASAP7_75t_L      g241(.A(new_n625), .B(new_n626), .Y(new_n627));
  NOR2xp33_ASAP7_75t_L      g242(.A(new_n624), .B(new_n627), .Y(new_n628));
  OR3x1_ASAP7_75t_L         g243(.A(new_n622), .B(new_n617), .C(new_n628), .Y(new_n629));
  A2O1A1Ixp33_ASAP7_75t_L   g244(.A1(\b[28] ), .A2(\a[28] ), .B(new_n622), .C(new_n628), .Y(new_n630));
  AND2x2_ASAP7_75t_L        g245(.A(new_n630), .B(new_n629), .Y(\f[29] ));
  NOR2xp33_ASAP7_75t_L      g246(.A(\a[30] ), .B(\b[30] ), .Y(new_n632));
  AND2x2_ASAP7_75t_L        g247(.A(\a[30] ), .B(\b[30] ), .Y(new_n633));
  NOR2xp33_ASAP7_75t_L      g248(.A(new_n632), .B(new_n633), .Y(new_n634));
  INVx1_ASAP7_75t_L         g249(.A(new_n634), .Y(new_n635));
  O2A1O1Ixp33_ASAP7_75t_L   g250(.A1(new_n617), .A2(new_n622), .B(new_n628), .C(new_n627), .Y(new_n636));
  AND2x2_ASAP7_75t_L        g251(.A(new_n635), .B(new_n636), .Y(new_n637));
  O2A1O1Ixp33_ASAP7_75t_L   g252(.A1(new_n625), .A2(new_n626), .B(new_n630), .C(new_n635), .Y(new_n638));
  NOR2xp33_ASAP7_75t_L      g253(.A(new_n638), .B(new_n637), .Y(\f[30] ));
  NOR2xp33_ASAP7_75t_L      g254(.A(\a[31] ), .B(\b[31] ), .Y(new_n640));
  INVx1_ASAP7_75t_L         g255(.A(\a[31] ), .Y(new_n641));
  INVx1_ASAP7_75t_L         g256(.A(\b[31] ), .Y(new_n642));
  NOR2xp33_ASAP7_75t_L      g257(.A(new_n641), .B(new_n642), .Y(new_n643));
  NOR2xp33_ASAP7_75t_L      g258(.A(new_n640), .B(new_n643), .Y(new_n644));
  OR3x1_ASAP7_75t_L         g259(.A(new_n638), .B(new_n633), .C(new_n644), .Y(new_n645));
  A2O1A1Ixp33_ASAP7_75t_L   g260(.A1(\b[30] ), .A2(\a[30] ), .B(new_n638), .C(new_n644), .Y(new_n646));
  AND2x2_ASAP7_75t_L        g261(.A(new_n646), .B(new_n645), .Y(\f[31] ));
  NOR2xp33_ASAP7_75t_L      g262(.A(\a[32] ), .B(\b[32] ), .Y(new_n648));
  AND2x2_ASAP7_75t_L        g263(.A(\a[32] ), .B(\b[32] ), .Y(new_n649));
  NOR2xp33_ASAP7_75t_L      g264(.A(new_n648), .B(new_n649), .Y(new_n650));
  INVx1_ASAP7_75t_L         g265(.A(new_n650), .Y(new_n651));
  O2A1O1Ixp33_ASAP7_75t_L   g266(.A1(new_n633), .A2(new_n638), .B(new_n644), .C(new_n643), .Y(new_n652));
  AND2x2_ASAP7_75t_L        g267(.A(new_n651), .B(new_n652), .Y(new_n653));
  O2A1O1Ixp33_ASAP7_75t_L   g268(.A1(new_n641), .A2(new_n642), .B(new_n646), .C(new_n651), .Y(new_n654));
  NOR2xp33_ASAP7_75t_L      g269(.A(new_n654), .B(new_n653), .Y(\f[32] ));
  NOR2xp33_ASAP7_75t_L      g270(.A(\a[33] ), .B(\b[33] ), .Y(new_n656));
  INVx1_ASAP7_75t_L         g271(.A(\a[33] ), .Y(new_n657));
  INVx1_ASAP7_75t_L         g272(.A(\b[33] ), .Y(new_n658));
  NOR2xp33_ASAP7_75t_L      g273(.A(new_n657), .B(new_n658), .Y(new_n659));
  NOR2xp33_ASAP7_75t_L      g274(.A(new_n656), .B(new_n659), .Y(new_n660));
  OR3x1_ASAP7_75t_L         g275(.A(new_n654), .B(new_n649), .C(new_n660), .Y(new_n661));
  A2O1A1Ixp33_ASAP7_75t_L   g276(.A1(\b[32] ), .A2(\a[32] ), .B(new_n654), .C(new_n660), .Y(new_n662));
  AND2x2_ASAP7_75t_L        g277(.A(new_n662), .B(new_n661), .Y(\f[33] ));
  NOR2xp33_ASAP7_75t_L      g278(.A(\a[34] ), .B(\b[34] ), .Y(new_n664));
  AND2x2_ASAP7_75t_L        g279(.A(\a[34] ), .B(\b[34] ), .Y(new_n665));
  NOR2xp33_ASAP7_75t_L      g280(.A(new_n664), .B(new_n665), .Y(new_n666));
  INVx1_ASAP7_75t_L         g281(.A(new_n666), .Y(new_n667));
  O2A1O1Ixp33_ASAP7_75t_L   g282(.A1(new_n649), .A2(new_n654), .B(new_n660), .C(new_n659), .Y(new_n668));
  AND2x2_ASAP7_75t_L        g283(.A(new_n667), .B(new_n668), .Y(new_n669));
  O2A1O1Ixp33_ASAP7_75t_L   g284(.A1(new_n657), .A2(new_n658), .B(new_n662), .C(new_n667), .Y(new_n670));
  NOR2xp33_ASAP7_75t_L      g285(.A(new_n670), .B(new_n669), .Y(\f[34] ));
  NOR2xp33_ASAP7_75t_L      g286(.A(\a[35] ), .B(\b[35] ), .Y(new_n672));
  INVx1_ASAP7_75t_L         g287(.A(\a[35] ), .Y(new_n673));
  INVx1_ASAP7_75t_L         g288(.A(\b[35] ), .Y(new_n674));
  NOR2xp33_ASAP7_75t_L      g289(.A(new_n673), .B(new_n674), .Y(new_n675));
  NOR2xp33_ASAP7_75t_L      g290(.A(new_n672), .B(new_n675), .Y(new_n676));
  OR3x1_ASAP7_75t_L         g291(.A(new_n670), .B(new_n665), .C(new_n676), .Y(new_n677));
  A2O1A1Ixp33_ASAP7_75t_L   g292(.A1(\b[34] ), .A2(\a[34] ), .B(new_n670), .C(new_n676), .Y(new_n678));
  AND2x2_ASAP7_75t_L        g293(.A(new_n678), .B(new_n677), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g294(.A(\a[36] ), .B(\b[36] ), .Y(new_n680));
  AND2x2_ASAP7_75t_L        g295(.A(\a[36] ), .B(\b[36] ), .Y(new_n681));
  NOR2xp33_ASAP7_75t_L      g296(.A(new_n680), .B(new_n681), .Y(new_n682));
  INVx1_ASAP7_75t_L         g297(.A(new_n682), .Y(new_n683));
  O2A1O1Ixp33_ASAP7_75t_L   g298(.A1(new_n665), .A2(new_n670), .B(new_n676), .C(new_n675), .Y(new_n684));
  AND2x2_ASAP7_75t_L        g299(.A(new_n683), .B(new_n684), .Y(new_n685));
  O2A1O1Ixp33_ASAP7_75t_L   g300(.A1(new_n673), .A2(new_n674), .B(new_n678), .C(new_n683), .Y(new_n686));
  NOR2xp33_ASAP7_75t_L      g301(.A(new_n686), .B(new_n685), .Y(\f[36] ));
  INVx1_ASAP7_75t_L         g302(.A(\a[37] ), .Y(new_n688));
  INVx1_ASAP7_75t_L         g303(.A(\b[37] ), .Y(new_n689));
  NAND2xp33_ASAP7_75t_L     g304(.A(new_n689), .B(new_n688), .Y(new_n690));
  NOR2xp33_ASAP7_75t_L      g305(.A(new_n688), .B(new_n689), .Y(new_n691));
  INVx1_ASAP7_75t_L         g306(.A(new_n691), .Y(new_n692));
  AND2x2_ASAP7_75t_L        g307(.A(new_n690), .B(new_n692), .Y(new_n693));
  OR3x1_ASAP7_75t_L         g308(.A(new_n686), .B(new_n681), .C(new_n693), .Y(new_n694));
  A2O1A1Ixp33_ASAP7_75t_L   g309(.A1(\b[36] ), .A2(\a[36] ), .B(new_n686), .C(new_n693), .Y(new_n695));
  AND2x2_ASAP7_75t_L        g310(.A(new_n695), .B(new_n694), .Y(\f[37] ));
  NOR2xp33_ASAP7_75t_L      g311(.A(\a[38] ), .B(\b[38] ), .Y(new_n697));
  INVx1_ASAP7_75t_L         g312(.A(\a[38] ), .Y(new_n698));
  INVx1_ASAP7_75t_L         g313(.A(\b[38] ), .Y(new_n699));
  NOR2xp33_ASAP7_75t_L      g314(.A(new_n698), .B(new_n699), .Y(new_n700));
  NOR2xp33_ASAP7_75t_L      g315(.A(new_n697), .B(new_n700), .Y(new_n701));
  O2A1O1Ixp33_ASAP7_75t_L   g316(.A1(new_n681), .A2(new_n686), .B(new_n690), .C(new_n691), .Y(new_n702));
  XNOR2x2_ASAP7_75t_L       g317(.A(new_n701), .B(new_n702), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g318(.A(\a[39] ), .B(\b[39] ), .Y(new_n704));
  NAND2xp33_ASAP7_75t_L     g319(.A(\b[39] ), .B(\a[39] ), .Y(new_n705));
  INVx1_ASAP7_75t_L         g320(.A(new_n705), .Y(new_n706));
  NOR2xp33_ASAP7_75t_L      g321(.A(new_n704), .B(new_n706), .Y(new_n707));
  INVx1_ASAP7_75t_L         g322(.A(new_n700), .Y(new_n708));
  A2O1A1Ixp33_ASAP7_75t_L   g323(.A1(new_n695), .A2(new_n692), .B(new_n697), .C(new_n708), .Y(new_n709));
  NOR2xp33_ASAP7_75t_L      g324(.A(new_n707), .B(new_n709), .Y(new_n710));
  INVx1_ASAP7_75t_L         g325(.A(new_n707), .Y(new_n711));
  O2A1O1Ixp33_ASAP7_75t_L   g326(.A1(new_n697), .A2(new_n702), .B(new_n708), .C(new_n711), .Y(new_n712));
  NOR2xp33_ASAP7_75t_L      g327(.A(new_n712), .B(new_n710), .Y(\f[39] ));
  NOR2xp33_ASAP7_75t_L      g328(.A(\a[40] ), .B(\b[40] ), .Y(new_n714));
  INVx1_ASAP7_75t_L         g329(.A(\a[40] ), .Y(new_n715));
  INVx1_ASAP7_75t_L         g330(.A(\b[40] ), .Y(new_n716));
  NOR2xp33_ASAP7_75t_L      g331(.A(new_n715), .B(new_n716), .Y(new_n717));
  NOR2xp33_ASAP7_75t_L      g332(.A(new_n714), .B(new_n717), .Y(new_n718));
  OR3x1_ASAP7_75t_L         g333(.A(new_n712), .B(new_n706), .C(new_n718), .Y(new_n719));
  A2O1A1Ixp33_ASAP7_75t_L   g334(.A1(new_n709), .A2(new_n707), .B(new_n706), .C(new_n718), .Y(new_n720));
  AND2x2_ASAP7_75t_L        g335(.A(new_n720), .B(new_n719), .Y(\f[40] ));
  INVx1_ASAP7_75t_L         g336(.A(new_n717), .Y(new_n722));
  NOR2xp33_ASAP7_75t_L      g337(.A(\a[41] ), .B(\b[41] ), .Y(new_n723));
  NAND2xp33_ASAP7_75t_L     g338(.A(\b[41] ), .B(\a[41] ), .Y(new_n724));
  INVx1_ASAP7_75t_L         g339(.A(new_n724), .Y(new_n725));
  NOR2xp33_ASAP7_75t_L      g340(.A(new_n723), .B(new_n725), .Y(new_n726));
  INVx1_ASAP7_75t_L         g341(.A(new_n726), .Y(new_n727));
  AND3x1_ASAP7_75t_L        g342(.A(new_n720), .B(new_n727), .C(new_n722), .Y(new_n728));
  O2A1O1Ixp33_ASAP7_75t_L   g343(.A1(new_n715), .A2(new_n716), .B(new_n720), .C(new_n727), .Y(new_n729));
  NOR2xp33_ASAP7_75t_L      g344(.A(new_n729), .B(new_n728), .Y(\f[41] ));
  NOR2xp33_ASAP7_75t_L      g345(.A(\a[42] ), .B(\b[42] ), .Y(new_n731));
  AND2x2_ASAP7_75t_L        g346(.A(\a[42] ), .B(\b[42] ), .Y(new_n732));
  NOR2xp33_ASAP7_75t_L      g347(.A(new_n731), .B(new_n732), .Y(new_n733));
  A2O1A1Ixp33_ASAP7_75t_L   g348(.A1(new_n720), .A2(new_n722), .B(new_n723), .C(new_n724), .Y(new_n734));
  XOR2x2_ASAP7_75t_L        g349(.A(new_n733), .B(new_n734), .Y(\f[42] ));
  NOR2xp33_ASAP7_75t_L      g350(.A(\a[43] ), .B(\b[43] ), .Y(new_n736));
  INVx1_ASAP7_75t_L         g351(.A(\a[43] ), .Y(new_n737));
  INVx1_ASAP7_75t_L         g352(.A(\b[43] ), .Y(new_n738));
  NOR2xp33_ASAP7_75t_L      g353(.A(new_n737), .B(new_n738), .Y(new_n739));
  NOR2xp33_ASAP7_75t_L      g354(.A(new_n736), .B(new_n739), .Y(new_n740));
  O2A1O1Ixp33_ASAP7_75t_L   g355(.A1(new_n725), .A2(new_n729), .B(new_n733), .C(new_n732), .Y(new_n741));
  XNOR2x2_ASAP7_75t_L       g356(.A(new_n740), .B(new_n741), .Y(\f[43] ));
  INVx1_ASAP7_75t_L         g357(.A(new_n739), .Y(new_n743));
  A2O1A1Ixp33_ASAP7_75t_L   g358(.A1(new_n734), .A2(new_n733), .B(new_n732), .C(new_n740), .Y(new_n744));
  NOR2xp33_ASAP7_75t_L      g359(.A(\a[44] ), .B(\b[44] ), .Y(new_n745));
  NAND2xp33_ASAP7_75t_L     g360(.A(\b[44] ), .B(\a[44] ), .Y(new_n746));
  INVx1_ASAP7_75t_L         g361(.A(new_n746), .Y(new_n747));
  NOR2xp33_ASAP7_75t_L      g362(.A(new_n745), .B(new_n747), .Y(new_n748));
  INVx1_ASAP7_75t_L         g363(.A(new_n748), .Y(new_n749));
  AND3x1_ASAP7_75t_L        g364(.A(new_n744), .B(new_n749), .C(new_n743), .Y(new_n750));
  O2A1O1Ixp33_ASAP7_75t_L   g365(.A1(new_n737), .A2(new_n738), .B(new_n744), .C(new_n749), .Y(new_n751));
  NOR2xp33_ASAP7_75t_L      g366(.A(new_n751), .B(new_n750), .Y(\f[44] ));
  NOR2xp33_ASAP7_75t_L      g367(.A(\a[45] ), .B(\b[45] ), .Y(new_n753));
  AND2x2_ASAP7_75t_L        g368(.A(\a[45] ), .B(\b[45] ), .Y(new_n754));
  NOR2xp33_ASAP7_75t_L      g369(.A(new_n753), .B(new_n754), .Y(new_n755));
  A2O1A1Ixp33_ASAP7_75t_L   g370(.A1(new_n744), .A2(new_n743), .B(new_n745), .C(new_n746), .Y(new_n756));
  XOR2x2_ASAP7_75t_L        g371(.A(new_n755), .B(new_n756), .Y(\f[45] ));
  NOR2xp33_ASAP7_75t_L      g372(.A(\a[46] ), .B(\b[46] ), .Y(new_n758));
  INVx1_ASAP7_75t_L         g373(.A(\a[46] ), .Y(new_n759));
  INVx1_ASAP7_75t_L         g374(.A(\b[46] ), .Y(new_n760));
  NOR2xp33_ASAP7_75t_L      g375(.A(new_n759), .B(new_n760), .Y(new_n761));
  NOR2xp33_ASAP7_75t_L      g376(.A(new_n758), .B(new_n761), .Y(new_n762));
  O2A1O1Ixp33_ASAP7_75t_L   g377(.A1(new_n747), .A2(new_n751), .B(new_n755), .C(new_n754), .Y(new_n763));
  XNOR2x2_ASAP7_75t_L       g378(.A(new_n762), .B(new_n763), .Y(\f[46] ));
  INVx1_ASAP7_75t_L         g379(.A(new_n761), .Y(new_n765));
  A2O1A1Ixp33_ASAP7_75t_L   g380(.A1(new_n756), .A2(new_n755), .B(new_n754), .C(new_n762), .Y(new_n766));
  NOR2xp33_ASAP7_75t_L      g381(.A(\a[47] ), .B(\b[47] ), .Y(new_n767));
  NAND2xp33_ASAP7_75t_L     g382(.A(\b[47] ), .B(\a[47] ), .Y(new_n768));
  INVx1_ASAP7_75t_L         g383(.A(new_n768), .Y(new_n769));
  NOR2xp33_ASAP7_75t_L      g384(.A(new_n767), .B(new_n769), .Y(new_n770));
  INVx1_ASAP7_75t_L         g385(.A(new_n770), .Y(new_n771));
  AND3x1_ASAP7_75t_L        g386(.A(new_n766), .B(new_n771), .C(new_n765), .Y(new_n772));
  O2A1O1Ixp33_ASAP7_75t_L   g387(.A1(new_n759), .A2(new_n760), .B(new_n766), .C(new_n771), .Y(new_n773));
  NOR2xp33_ASAP7_75t_L      g388(.A(new_n773), .B(new_n772), .Y(\f[47] ));
  NOR2xp33_ASAP7_75t_L      g389(.A(\a[48] ), .B(\b[48] ), .Y(new_n775));
  AND2x2_ASAP7_75t_L        g390(.A(\a[48] ), .B(\b[48] ), .Y(new_n776));
  NOR2xp33_ASAP7_75t_L      g391(.A(new_n775), .B(new_n776), .Y(new_n777));
  A2O1A1Ixp33_ASAP7_75t_L   g392(.A1(new_n766), .A2(new_n765), .B(new_n767), .C(new_n768), .Y(new_n778));
  XOR2x2_ASAP7_75t_L        g393(.A(new_n777), .B(new_n778), .Y(\f[48] ));
  NOR2xp33_ASAP7_75t_L      g394(.A(\a[49] ), .B(\b[49] ), .Y(new_n780));
  INVx1_ASAP7_75t_L         g395(.A(\a[49] ), .Y(new_n781));
  INVx1_ASAP7_75t_L         g396(.A(\b[49] ), .Y(new_n782));
  NOR2xp33_ASAP7_75t_L      g397(.A(new_n781), .B(new_n782), .Y(new_n783));
  NOR2xp33_ASAP7_75t_L      g398(.A(new_n780), .B(new_n783), .Y(new_n784));
  O2A1O1Ixp33_ASAP7_75t_L   g399(.A1(new_n769), .A2(new_n773), .B(new_n777), .C(new_n776), .Y(new_n785));
  XNOR2x2_ASAP7_75t_L       g400(.A(new_n784), .B(new_n785), .Y(\f[49] ));
  INVx1_ASAP7_75t_L         g401(.A(new_n783), .Y(new_n787));
  A2O1A1Ixp33_ASAP7_75t_L   g402(.A1(new_n778), .A2(new_n777), .B(new_n776), .C(new_n784), .Y(new_n788));
  NOR2xp33_ASAP7_75t_L      g403(.A(\a[50] ), .B(\b[50] ), .Y(new_n789));
  NAND2xp33_ASAP7_75t_L     g404(.A(\b[50] ), .B(\a[50] ), .Y(new_n790));
  INVx1_ASAP7_75t_L         g405(.A(new_n790), .Y(new_n791));
  NOR2xp33_ASAP7_75t_L      g406(.A(new_n789), .B(new_n791), .Y(new_n792));
  INVx1_ASAP7_75t_L         g407(.A(new_n792), .Y(new_n793));
  AND3x1_ASAP7_75t_L        g408(.A(new_n788), .B(new_n793), .C(new_n787), .Y(new_n794));
  O2A1O1Ixp33_ASAP7_75t_L   g409(.A1(new_n781), .A2(new_n782), .B(new_n788), .C(new_n793), .Y(new_n795));
  NOR2xp33_ASAP7_75t_L      g410(.A(new_n795), .B(new_n794), .Y(\f[50] ));
  NOR2xp33_ASAP7_75t_L      g411(.A(\a[51] ), .B(\b[51] ), .Y(new_n797));
  AND2x2_ASAP7_75t_L        g412(.A(\a[51] ), .B(\b[51] ), .Y(new_n798));
  NOR2xp33_ASAP7_75t_L      g413(.A(new_n797), .B(new_n798), .Y(new_n799));
  A2O1A1Ixp33_ASAP7_75t_L   g414(.A1(new_n788), .A2(new_n787), .B(new_n789), .C(new_n790), .Y(new_n800));
  XOR2x2_ASAP7_75t_L        g415(.A(new_n799), .B(new_n800), .Y(\f[51] ));
  NOR2xp33_ASAP7_75t_L      g416(.A(\a[52] ), .B(\b[52] ), .Y(new_n802));
  INVx1_ASAP7_75t_L         g417(.A(\a[52] ), .Y(new_n803));
  INVx1_ASAP7_75t_L         g418(.A(\b[52] ), .Y(new_n804));
  NOR2xp33_ASAP7_75t_L      g419(.A(new_n803), .B(new_n804), .Y(new_n805));
  NOR2xp33_ASAP7_75t_L      g420(.A(new_n802), .B(new_n805), .Y(new_n806));
  O2A1O1Ixp33_ASAP7_75t_L   g421(.A1(new_n791), .A2(new_n795), .B(new_n799), .C(new_n798), .Y(new_n807));
  XNOR2x2_ASAP7_75t_L       g422(.A(new_n806), .B(new_n807), .Y(\f[52] ));
  INVx1_ASAP7_75t_L         g423(.A(new_n805), .Y(new_n809));
  A2O1A1Ixp33_ASAP7_75t_L   g424(.A1(new_n800), .A2(new_n799), .B(new_n798), .C(new_n806), .Y(new_n810));
  NOR2xp33_ASAP7_75t_L      g425(.A(\a[53] ), .B(\b[53] ), .Y(new_n811));
  NAND2xp33_ASAP7_75t_L     g426(.A(\b[53] ), .B(\a[53] ), .Y(new_n812));
  INVx1_ASAP7_75t_L         g427(.A(new_n812), .Y(new_n813));
  NOR2xp33_ASAP7_75t_L      g428(.A(new_n811), .B(new_n813), .Y(new_n814));
  INVx1_ASAP7_75t_L         g429(.A(new_n814), .Y(new_n815));
  AND3x1_ASAP7_75t_L        g430(.A(new_n810), .B(new_n815), .C(new_n809), .Y(new_n816));
  O2A1O1Ixp33_ASAP7_75t_L   g431(.A1(new_n803), .A2(new_n804), .B(new_n810), .C(new_n815), .Y(new_n817));
  NOR2xp33_ASAP7_75t_L      g432(.A(new_n817), .B(new_n816), .Y(\f[53] ));
  NOR2xp33_ASAP7_75t_L      g433(.A(\a[54] ), .B(\b[54] ), .Y(new_n819));
  AND2x2_ASAP7_75t_L        g434(.A(\a[54] ), .B(\b[54] ), .Y(new_n820));
  NOR2xp33_ASAP7_75t_L      g435(.A(new_n819), .B(new_n820), .Y(new_n821));
  A2O1A1Ixp33_ASAP7_75t_L   g436(.A1(new_n810), .A2(new_n809), .B(new_n811), .C(new_n812), .Y(new_n822));
  XOR2x2_ASAP7_75t_L        g437(.A(new_n821), .B(new_n822), .Y(\f[54] ));
  NOR2xp33_ASAP7_75t_L      g438(.A(\a[55] ), .B(\b[55] ), .Y(new_n824));
  INVx1_ASAP7_75t_L         g439(.A(\a[55] ), .Y(new_n825));
  INVx1_ASAP7_75t_L         g440(.A(\b[55] ), .Y(new_n826));
  NOR2xp33_ASAP7_75t_L      g441(.A(new_n825), .B(new_n826), .Y(new_n827));
  NOR2xp33_ASAP7_75t_L      g442(.A(new_n824), .B(new_n827), .Y(new_n828));
  O2A1O1Ixp33_ASAP7_75t_L   g443(.A1(new_n813), .A2(new_n817), .B(new_n821), .C(new_n820), .Y(new_n829));
  XNOR2x2_ASAP7_75t_L       g444(.A(new_n828), .B(new_n829), .Y(\f[55] ));
  INVx1_ASAP7_75t_L         g445(.A(new_n827), .Y(new_n831));
  A2O1A1Ixp33_ASAP7_75t_L   g446(.A1(new_n822), .A2(new_n821), .B(new_n820), .C(new_n828), .Y(new_n832));
  NOR2xp33_ASAP7_75t_L      g447(.A(\a[56] ), .B(\b[56] ), .Y(new_n833));
  NAND2xp33_ASAP7_75t_L     g448(.A(\b[56] ), .B(\a[56] ), .Y(new_n834));
  INVx1_ASAP7_75t_L         g449(.A(new_n834), .Y(new_n835));
  NOR2xp33_ASAP7_75t_L      g450(.A(new_n833), .B(new_n835), .Y(new_n836));
  INVx1_ASAP7_75t_L         g451(.A(new_n836), .Y(new_n837));
  AND3x1_ASAP7_75t_L        g452(.A(new_n832), .B(new_n837), .C(new_n831), .Y(new_n838));
  O2A1O1Ixp33_ASAP7_75t_L   g453(.A1(new_n825), .A2(new_n826), .B(new_n832), .C(new_n837), .Y(new_n839));
  NOR2xp33_ASAP7_75t_L      g454(.A(new_n839), .B(new_n838), .Y(\f[56] ));
  NOR2xp33_ASAP7_75t_L      g455(.A(\a[57] ), .B(\b[57] ), .Y(new_n841));
  AND2x2_ASAP7_75t_L        g456(.A(\a[57] ), .B(\b[57] ), .Y(new_n842));
  NOR2xp33_ASAP7_75t_L      g457(.A(new_n841), .B(new_n842), .Y(new_n843));
  A2O1A1Ixp33_ASAP7_75t_L   g458(.A1(new_n832), .A2(new_n831), .B(new_n833), .C(new_n834), .Y(new_n844));
  XOR2x2_ASAP7_75t_L        g459(.A(new_n843), .B(new_n844), .Y(\f[57] ));
  NOR2xp33_ASAP7_75t_L      g460(.A(\a[58] ), .B(\b[58] ), .Y(new_n846));
  INVx1_ASAP7_75t_L         g461(.A(\a[58] ), .Y(new_n847));
  INVx1_ASAP7_75t_L         g462(.A(\b[58] ), .Y(new_n848));
  NOR2xp33_ASAP7_75t_L      g463(.A(new_n847), .B(new_n848), .Y(new_n849));
  NOR2xp33_ASAP7_75t_L      g464(.A(new_n846), .B(new_n849), .Y(new_n850));
  O2A1O1Ixp33_ASAP7_75t_L   g465(.A1(new_n835), .A2(new_n839), .B(new_n843), .C(new_n842), .Y(new_n851));
  XNOR2x2_ASAP7_75t_L       g466(.A(new_n850), .B(new_n851), .Y(\f[58] ));
  INVx1_ASAP7_75t_L         g467(.A(new_n849), .Y(new_n853));
  A2O1A1Ixp33_ASAP7_75t_L   g468(.A1(new_n844), .A2(new_n843), .B(new_n842), .C(new_n850), .Y(new_n854));
  NOR2xp33_ASAP7_75t_L      g469(.A(\a[59] ), .B(\b[59] ), .Y(new_n855));
  NAND2xp33_ASAP7_75t_L     g470(.A(\b[59] ), .B(\a[59] ), .Y(new_n856));
  INVx1_ASAP7_75t_L         g471(.A(new_n856), .Y(new_n857));
  NOR2xp33_ASAP7_75t_L      g472(.A(new_n855), .B(new_n857), .Y(new_n858));
  INVx1_ASAP7_75t_L         g473(.A(new_n858), .Y(new_n859));
  AND3x1_ASAP7_75t_L        g474(.A(new_n854), .B(new_n859), .C(new_n853), .Y(new_n860));
  O2A1O1Ixp33_ASAP7_75t_L   g475(.A1(new_n847), .A2(new_n848), .B(new_n854), .C(new_n859), .Y(new_n861));
  NOR2xp33_ASAP7_75t_L      g476(.A(new_n861), .B(new_n860), .Y(\f[59] ));
  NOR2xp33_ASAP7_75t_L      g477(.A(\a[60] ), .B(\b[60] ), .Y(new_n863));
  AND2x2_ASAP7_75t_L        g478(.A(\a[60] ), .B(\b[60] ), .Y(new_n864));
  NOR2xp33_ASAP7_75t_L      g479(.A(new_n863), .B(new_n864), .Y(new_n865));
  A2O1A1Ixp33_ASAP7_75t_L   g480(.A1(new_n854), .A2(new_n853), .B(new_n855), .C(new_n856), .Y(new_n866));
  XOR2x2_ASAP7_75t_L        g481(.A(new_n865), .B(new_n866), .Y(\f[60] ));
  NOR2xp33_ASAP7_75t_L      g482(.A(\a[61] ), .B(\b[61] ), .Y(new_n868));
  INVx1_ASAP7_75t_L         g483(.A(\a[61] ), .Y(new_n869));
  INVx1_ASAP7_75t_L         g484(.A(\b[61] ), .Y(new_n870));
  NOR2xp33_ASAP7_75t_L      g485(.A(new_n869), .B(new_n870), .Y(new_n871));
  NOR2xp33_ASAP7_75t_L      g486(.A(new_n868), .B(new_n871), .Y(new_n872));
  O2A1O1Ixp33_ASAP7_75t_L   g487(.A1(new_n857), .A2(new_n861), .B(new_n865), .C(new_n864), .Y(new_n873));
  XNOR2x2_ASAP7_75t_L       g488(.A(new_n872), .B(new_n873), .Y(\f[61] ));
  INVx1_ASAP7_75t_L         g489(.A(new_n871), .Y(new_n875));
  A2O1A1Ixp33_ASAP7_75t_L   g490(.A1(new_n866), .A2(new_n865), .B(new_n864), .C(new_n872), .Y(new_n876));
  NOR2xp33_ASAP7_75t_L      g491(.A(\a[62] ), .B(\b[62] ), .Y(new_n877));
  NAND2xp33_ASAP7_75t_L     g492(.A(\b[62] ), .B(\a[62] ), .Y(new_n878));
  INVx1_ASAP7_75t_L         g493(.A(new_n878), .Y(new_n879));
  NOR2xp33_ASAP7_75t_L      g494(.A(new_n877), .B(new_n879), .Y(new_n880));
  INVx1_ASAP7_75t_L         g495(.A(new_n880), .Y(new_n881));
  AND3x1_ASAP7_75t_L        g496(.A(new_n876), .B(new_n881), .C(new_n875), .Y(new_n882));
  O2A1O1Ixp33_ASAP7_75t_L   g497(.A1(new_n869), .A2(new_n870), .B(new_n876), .C(new_n881), .Y(new_n883));
  NOR2xp33_ASAP7_75t_L      g498(.A(new_n883), .B(new_n882), .Y(\f[62] ));
  NOR2xp33_ASAP7_75t_L      g499(.A(\a[63] ), .B(\b[63] ), .Y(new_n885));
  AND2x2_ASAP7_75t_L        g500(.A(\a[63] ), .B(\b[63] ), .Y(new_n886));
  NOR2xp33_ASAP7_75t_L      g501(.A(new_n885), .B(new_n886), .Y(new_n887));
  A2O1A1Ixp33_ASAP7_75t_L   g502(.A1(new_n876), .A2(new_n875), .B(new_n877), .C(new_n878), .Y(new_n888));
  XOR2x2_ASAP7_75t_L        g503(.A(new_n887), .B(new_n888), .Y(\f[63] ));
  NOR2xp33_ASAP7_75t_L      g504(.A(\a[64] ), .B(\b[64] ), .Y(new_n890));
  INVx1_ASAP7_75t_L         g505(.A(\a[64] ), .Y(new_n891));
  INVx1_ASAP7_75t_L         g506(.A(\b[64] ), .Y(new_n892));
  NOR2xp33_ASAP7_75t_L      g507(.A(new_n891), .B(new_n892), .Y(new_n893));
  NOR2xp33_ASAP7_75t_L      g508(.A(new_n890), .B(new_n893), .Y(new_n894));
  O2A1O1Ixp33_ASAP7_75t_L   g509(.A1(new_n879), .A2(new_n883), .B(new_n887), .C(new_n886), .Y(new_n895));
  XNOR2x2_ASAP7_75t_L       g510(.A(new_n894), .B(new_n895), .Y(\f[64] ));
  INVx1_ASAP7_75t_L         g511(.A(new_n893), .Y(new_n897));
  A2O1A1Ixp33_ASAP7_75t_L   g512(.A1(new_n888), .A2(new_n887), .B(new_n886), .C(new_n894), .Y(new_n898));
  NOR2xp33_ASAP7_75t_L      g513(.A(\a[65] ), .B(\b[65] ), .Y(new_n899));
  NAND2xp33_ASAP7_75t_L     g514(.A(\b[65] ), .B(\a[65] ), .Y(new_n900));
  INVx1_ASAP7_75t_L         g515(.A(new_n900), .Y(new_n901));
  NOR2xp33_ASAP7_75t_L      g516(.A(new_n899), .B(new_n901), .Y(new_n902));
  INVx1_ASAP7_75t_L         g517(.A(new_n902), .Y(new_n903));
  AND3x1_ASAP7_75t_L        g518(.A(new_n898), .B(new_n903), .C(new_n897), .Y(new_n904));
  O2A1O1Ixp33_ASAP7_75t_L   g519(.A1(new_n891), .A2(new_n892), .B(new_n898), .C(new_n903), .Y(new_n905));
  NOR2xp33_ASAP7_75t_L      g520(.A(new_n905), .B(new_n904), .Y(\f[65] ));
  NOR2xp33_ASAP7_75t_L      g521(.A(\a[66] ), .B(\b[66] ), .Y(new_n907));
  AND2x2_ASAP7_75t_L        g522(.A(\a[66] ), .B(\b[66] ), .Y(new_n908));
  NOR2xp33_ASAP7_75t_L      g523(.A(new_n907), .B(new_n908), .Y(new_n909));
  A2O1A1Ixp33_ASAP7_75t_L   g524(.A1(new_n898), .A2(new_n897), .B(new_n899), .C(new_n900), .Y(new_n910));
  XOR2x2_ASAP7_75t_L        g525(.A(new_n909), .B(new_n910), .Y(\f[66] ));
  NOR2xp33_ASAP7_75t_L      g526(.A(\a[67] ), .B(\b[67] ), .Y(new_n912));
  INVx1_ASAP7_75t_L         g527(.A(\a[67] ), .Y(new_n913));
  INVx1_ASAP7_75t_L         g528(.A(\b[67] ), .Y(new_n914));
  NOR2xp33_ASAP7_75t_L      g529(.A(new_n913), .B(new_n914), .Y(new_n915));
  NOR2xp33_ASAP7_75t_L      g530(.A(new_n912), .B(new_n915), .Y(new_n916));
  O2A1O1Ixp33_ASAP7_75t_L   g531(.A1(new_n901), .A2(new_n905), .B(new_n909), .C(new_n908), .Y(new_n917));
  XNOR2x2_ASAP7_75t_L       g532(.A(new_n916), .B(new_n917), .Y(\f[67] ));
  INVx1_ASAP7_75t_L         g533(.A(new_n915), .Y(new_n919));
  A2O1A1Ixp33_ASAP7_75t_L   g534(.A1(new_n910), .A2(new_n909), .B(new_n908), .C(new_n916), .Y(new_n920));
  NOR2xp33_ASAP7_75t_L      g535(.A(\a[68] ), .B(\b[68] ), .Y(new_n921));
  NAND2xp33_ASAP7_75t_L     g536(.A(\b[68] ), .B(\a[68] ), .Y(new_n922));
  INVx1_ASAP7_75t_L         g537(.A(new_n922), .Y(new_n923));
  NOR2xp33_ASAP7_75t_L      g538(.A(new_n921), .B(new_n923), .Y(new_n924));
  INVx1_ASAP7_75t_L         g539(.A(new_n924), .Y(new_n925));
  AND3x1_ASAP7_75t_L        g540(.A(new_n920), .B(new_n925), .C(new_n919), .Y(new_n926));
  O2A1O1Ixp33_ASAP7_75t_L   g541(.A1(new_n913), .A2(new_n914), .B(new_n920), .C(new_n925), .Y(new_n927));
  NOR2xp33_ASAP7_75t_L      g542(.A(new_n927), .B(new_n926), .Y(\f[68] ));
  NOR2xp33_ASAP7_75t_L      g543(.A(\a[69] ), .B(\b[69] ), .Y(new_n929));
  AND2x2_ASAP7_75t_L        g544(.A(\a[69] ), .B(\b[69] ), .Y(new_n930));
  NOR2xp33_ASAP7_75t_L      g545(.A(new_n929), .B(new_n930), .Y(new_n931));
  A2O1A1Ixp33_ASAP7_75t_L   g546(.A1(new_n920), .A2(new_n919), .B(new_n921), .C(new_n922), .Y(new_n932));
  XOR2x2_ASAP7_75t_L        g547(.A(new_n931), .B(new_n932), .Y(\f[69] ));
  NOR2xp33_ASAP7_75t_L      g548(.A(\a[70] ), .B(\b[70] ), .Y(new_n934));
  INVx1_ASAP7_75t_L         g549(.A(\a[70] ), .Y(new_n935));
  INVx1_ASAP7_75t_L         g550(.A(\b[70] ), .Y(new_n936));
  NOR2xp33_ASAP7_75t_L      g551(.A(new_n935), .B(new_n936), .Y(new_n937));
  NOR2xp33_ASAP7_75t_L      g552(.A(new_n934), .B(new_n937), .Y(new_n938));
  O2A1O1Ixp33_ASAP7_75t_L   g553(.A1(new_n923), .A2(new_n927), .B(new_n931), .C(new_n930), .Y(new_n939));
  XNOR2x2_ASAP7_75t_L       g554(.A(new_n938), .B(new_n939), .Y(\f[70] ));
  INVx1_ASAP7_75t_L         g555(.A(new_n937), .Y(new_n941));
  A2O1A1Ixp33_ASAP7_75t_L   g556(.A1(new_n932), .A2(new_n931), .B(new_n930), .C(new_n938), .Y(new_n942));
  NOR2xp33_ASAP7_75t_L      g557(.A(\a[71] ), .B(\b[71] ), .Y(new_n943));
  NAND2xp33_ASAP7_75t_L     g558(.A(\b[71] ), .B(\a[71] ), .Y(new_n944));
  INVx1_ASAP7_75t_L         g559(.A(new_n944), .Y(new_n945));
  NOR2xp33_ASAP7_75t_L      g560(.A(new_n943), .B(new_n945), .Y(new_n946));
  INVx1_ASAP7_75t_L         g561(.A(new_n946), .Y(new_n947));
  AND3x1_ASAP7_75t_L        g562(.A(new_n942), .B(new_n947), .C(new_n941), .Y(new_n948));
  O2A1O1Ixp33_ASAP7_75t_L   g563(.A1(new_n935), .A2(new_n936), .B(new_n942), .C(new_n947), .Y(new_n949));
  NOR2xp33_ASAP7_75t_L      g564(.A(new_n949), .B(new_n948), .Y(\f[71] ));
  NOR2xp33_ASAP7_75t_L      g565(.A(\a[72] ), .B(\b[72] ), .Y(new_n951));
  AND2x2_ASAP7_75t_L        g566(.A(\a[72] ), .B(\b[72] ), .Y(new_n952));
  NOR2xp33_ASAP7_75t_L      g567(.A(new_n951), .B(new_n952), .Y(new_n953));
  A2O1A1Ixp33_ASAP7_75t_L   g568(.A1(new_n942), .A2(new_n941), .B(new_n943), .C(new_n944), .Y(new_n954));
  XOR2x2_ASAP7_75t_L        g569(.A(new_n953), .B(new_n954), .Y(\f[72] ));
  NOR2xp33_ASAP7_75t_L      g570(.A(\a[73] ), .B(\b[73] ), .Y(new_n956));
  INVx1_ASAP7_75t_L         g571(.A(\a[73] ), .Y(new_n957));
  INVx1_ASAP7_75t_L         g572(.A(\b[73] ), .Y(new_n958));
  NOR2xp33_ASAP7_75t_L      g573(.A(new_n957), .B(new_n958), .Y(new_n959));
  NOR2xp33_ASAP7_75t_L      g574(.A(new_n956), .B(new_n959), .Y(new_n960));
  O2A1O1Ixp33_ASAP7_75t_L   g575(.A1(new_n945), .A2(new_n949), .B(new_n953), .C(new_n952), .Y(new_n961));
  XNOR2x2_ASAP7_75t_L       g576(.A(new_n960), .B(new_n961), .Y(\f[73] ));
  INVx1_ASAP7_75t_L         g577(.A(new_n959), .Y(new_n963));
  A2O1A1Ixp33_ASAP7_75t_L   g578(.A1(new_n954), .A2(new_n953), .B(new_n952), .C(new_n960), .Y(new_n964));
  NOR2xp33_ASAP7_75t_L      g579(.A(\a[74] ), .B(\b[74] ), .Y(new_n965));
  NAND2xp33_ASAP7_75t_L     g580(.A(\b[74] ), .B(\a[74] ), .Y(new_n966));
  INVx1_ASAP7_75t_L         g581(.A(new_n966), .Y(new_n967));
  NOR2xp33_ASAP7_75t_L      g582(.A(new_n965), .B(new_n967), .Y(new_n968));
  INVx1_ASAP7_75t_L         g583(.A(new_n968), .Y(new_n969));
  AND3x1_ASAP7_75t_L        g584(.A(new_n964), .B(new_n969), .C(new_n963), .Y(new_n970));
  O2A1O1Ixp33_ASAP7_75t_L   g585(.A1(new_n957), .A2(new_n958), .B(new_n964), .C(new_n969), .Y(new_n971));
  NOR2xp33_ASAP7_75t_L      g586(.A(new_n971), .B(new_n970), .Y(\f[74] ));
  NOR2xp33_ASAP7_75t_L      g587(.A(\a[75] ), .B(\b[75] ), .Y(new_n973));
  AND2x2_ASAP7_75t_L        g588(.A(\a[75] ), .B(\b[75] ), .Y(new_n974));
  NOR2xp33_ASAP7_75t_L      g589(.A(new_n973), .B(new_n974), .Y(new_n975));
  A2O1A1Ixp33_ASAP7_75t_L   g590(.A1(new_n964), .A2(new_n963), .B(new_n965), .C(new_n966), .Y(new_n976));
  XOR2x2_ASAP7_75t_L        g591(.A(new_n975), .B(new_n976), .Y(\f[75] ));
  NOR2xp33_ASAP7_75t_L      g592(.A(\a[76] ), .B(\b[76] ), .Y(new_n978));
  INVx1_ASAP7_75t_L         g593(.A(\a[76] ), .Y(new_n979));
  INVx1_ASAP7_75t_L         g594(.A(\b[76] ), .Y(new_n980));
  NOR2xp33_ASAP7_75t_L      g595(.A(new_n979), .B(new_n980), .Y(new_n981));
  NOR2xp33_ASAP7_75t_L      g596(.A(new_n978), .B(new_n981), .Y(new_n982));
  O2A1O1Ixp33_ASAP7_75t_L   g597(.A1(new_n967), .A2(new_n971), .B(new_n975), .C(new_n974), .Y(new_n983));
  XNOR2x2_ASAP7_75t_L       g598(.A(new_n982), .B(new_n983), .Y(\f[76] ));
  INVx1_ASAP7_75t_L         g599(.A(new_n981), .Y(new_n985));
  A2O1A1Ixp33_ASAP7_75t_L   g600(.A1(new_n976), .A2(new_n975), .B(new_n974), .C(new_n982), .Y(new_n986));
  NOR2xp33_ASAP7_75t_L      g601(.A(\a[77] ), .B(\b[77] ), .Y(new_n987));
  NAND2xp33_ASAP7_75t_L     g602(.A(\b[77] ), .B(\a[77] ), .Y(new_n988));
  INVx1_ASAP7_75t_L         g603(.A(new_n988), .Y(new_n989));
  NOR2xp33_ASAP7_75t_L      g604(.A(new_n987), .B(new_n989), .Y(new_n990));
  INVx1_ASAP7_75t_L         g605(.A(new_n990), .Y(new_n991));
  AND3x1_ASAP7_75t_L        g606(.A(new_n986), .B(new_n991), .C(new_n985), .Y(new_n992));
  O2A1O1Ixp33_ASAP7_75t_L   g607(.A1(new_n979), .A2(new_n980), .B(new_n986), .C(new_n991), .Y(new_n993));
  NOR2xp33_ASAP7_75t_L      g608(.A(new_n993), .B(new_n992), .Y(\f[77] ));
  NOR2xp33_ASAP7_75t_L      g609(.A(\a[78] ), .B(\b[78] ), .Y(new_n995));
  AND2x2_ASAP7_75t_L        g610(.A(\a[78] ), .B(\b[78] ), .Y(new_n996));
  NOR2xp33_ASAP7_75t_L      g611(.A(new_n995), .B(new_n996), .Y(new_n997));
  A2O1A1Ixp33_ASAP7_75t_L   g612(.A1(new_n986), .A2(new_n985), .B(new_n987), .C(new_n988), .Y(new_n998));
  XOR2x2_ASAP7_75t_L        g613(.A(new_n997), .B(new_n998), .Y(\f[78] ));
  NOR2xp33_ASAP7_75t_L      g614(.A(\a[79] ), .B(\b[79] ), .Y(new_n1000));
  INVx1_ASAP7_75t_L         g615(.A(\a[79] ), .Y(new_n1001));
  INVx1_ASAP7_75t_L         g616(.A(\b[79] ), .Y(new_n1002));
  NOR2xp33_ASAP7_75t_L      g617(.A(new_n1001), .B(new_n1002), .Y(new_n1003));
  NOR2xp33_ASAP7_75t_L      g618(.A(new_n1000), .B(new_n1003), .Y(new_n1004));
  O2A1O1Ixp33_ASAP7_75t_L   g619(.A1(new_n989), .A2(new_n993), .B(new_n997), .C(new_n996), .Y(new_n1005));
  XNOR2x2_ASAP7_75t_L       g620(.A(new_n1004), .B(new_n1005), .Y(\f[79] ));
  INVx1_ASAP7_75t_L         g621(.A(new_n1003), .Y(new_n1007));
  A2O1A1Ixp33_ASAP7_75t_L   g622(.A1(new_n998), .A2(new_n997), .B(new_n996), .C(new_n1004), .Y(new_n1008));
  NOR2xp33_ASAP7_75t_L      g623(.A(\a[80] ), .B(\b[80] ), .Y(new_n1009));
  NAND2xp33_ASAP7_75t_L     g624(.A(\b[80] ), .B(\a[80] ), .Y(new_n1010));
  INVx1_ASAP7_75t_L         g625(.A(new_n1010), .Y(new_n1011));
  NOR2xp33_ASAP7_75t_L      g626(.A(new_n1009), .B(new_n1011), .Y(new_n1012));
  INVx1_ASAP7_75t_L         g627(.A(new_n1012), .Y(new_n1013));
  AND3x1_ASAP7_75t_L        g628(.A(new_n1008), .B(new_n1013), .C(new_n1007), .Y(new_n1014));
  O2A1O1Ixp33_ASAP7_75t_L   g629(.A1(new_n1001), .A2(new_n1002), .B(new_n1008), .C(new_n1013), .Y(new_n1015));
  NOR2xp33_ASAP7_75t_L      g630(.A(new_n1015), .B(new_n1014), .Y(\f[80] ));
  NOR2xp33_ASAP7_75t_L      g631(.A(\a[81] ), .B(\b[81] ), .Y(new_n1017));
  AND2x2_ASAP7_75t_L        g632(.A(\a[81] ), .B(\b[81] ), .Y(new_n1018));
  NOR2xp33_ASAP7_75t_L      g633(.A(new_n1017), .B(new_n1018), .Y(new_n1019));
  A2O1A1Ixp33_ASAP7_75t_L   g634(.A1(new_n1008), .A2(new_n1007), .B(new_n1009), .C(new_n1010), .Y(new_n1020));
  XOR2x2_ASAP7_75t_L        g635(.A(new_n1019), .B(new_n1020), .Y(\f[81] ));
  NOR2xp33_ASAP7_75t_L      g636(.A(\a[82] ), .B(\b[82] ), .Y(new_n1022));
  INVx1_ASAP7_75t_L         g637(.A(\a[82] ), .Y(new_n1023));
  INVx1_ASAP7_75t_L         g638(.A(\b[82] ), .Y(new_n1024));
  NOR2xp33_ASAP7_75t_L      g639(.A(new_n1023), .B(new_n1024), .Y(new_n1025));
  NOR2xp33_ASAP7_75t_L      g640(.A(new_n1022), .B(new_n1025), .Y(new_n1026));
  O2A1O1Ixp33_ASAP7_75t_L   g641(.A1(new_n1011), .A2(new_n1015), .B(new_n1019), .C(new_n1018), .Y(new_n1027));
  XNOR2x2_ASAP7_75t_L       g642(.A(new_n1026), .B(new_n1027), .Y(\f[82] ));
  INVx1_ASAP7_75t_L         g643(.A(new_n1025), .Y(new_n1029));
  A2O1A1Ixp33_ASAP7_75t_L   g644(.A1(new_n1020), .A2(new_n1019), .B(new_n1018), .C(new_n1026), .Y(new_n1030));
  NOR2xp33_ASAP7_75t_L      g645(.A(\a[83] ), .B(\b[83] ), .Y(new_n1031));
  NAND2xp33_ASAP7_75t_L     g646(.A(\b[83] ), .B(\a[83] ), .Y(new_n1032));
  INVx1_ASAP7_75t_L         g647(.A(new_n1032), .Y(new_n1033));
  NOR2xp33_ASAP7_75t_L      g648(.A(new_n1031), .B(new_n1033), .Y(new_n1034));
  INVx1_ASAP7_75t_L         g649(.A(new_n1034), .Y(new_n1035));
  AND3x1_ASAP7_75t_L        g650(.A(new_n1030), .B(new_n1035), .C(new_n1029), .Y(new_n1036));
  O2A1O1Ixp33_ASAP7_75t_L   g651(.A1(new_n1023), .A2(new_n1024), .B(new_n1030), .C(new_n1035), .Y(new_n1037));
  NOR2xp33_ASAP7_75t_L      g652(.A(new_n1037), .B(new_n1036), .Y(\f[83] ));
  NOR2xp33_ASAP7_75t_L      g653(.A(\a[84] ), .B(\b[84] ), .Y(new_n1039));
  AND2x2_ASAP7_75t_L        g654(.A(\a[84] ), .B(\b[84] ), .Y(new_n1040));
  NOR2xp33_ASAP7_75t_L      g655(.A(new_n1039), .B(new_n1040), .Y(new_n1041));
  A2O1A1Ixp33_ASAP7_75t_L   g656(.A1(new_n1030), .A2(new_n1029), .B(new_n1031), .C(new_n1032), .Y(new_n1042));
  XOR2x2_ASAP7_75t_L        g657(.A(new_n1041), .B(new_n1042), .Y(\f[84] ));
  NOR2xp33_ASAP7_75t_L      g658(.A(\a[85] ), .B(\b[85] ), .Y(new_n1044));
  INVx1_ASAP7_75t_L         g659(.A(\a[85] ), .Y(new_n1045));
  INVx1_ASAP7_75t_L         g660(.A(\b[85] ), .Y(new_n1046));
  NOR2xp33_ASAP7_75t_L      g661(.A(new_n1045), .B(new_n1046), .Y(new_n1047));
  NOR2xp33_ASAP7_75t_L      g662(.A(new_n1044), .B(new_n1047), .Y(new_n1048));
  O2A1O1Ixp33_ASAP7_75t_L   g663(.A1(new_n1033), .A2(new_n1037), .B(new_n1041), .C(new_n1040), .Y(new_n1049));
  XNOR2x2_ASAP7_75t_L       g664(.A(new_n1048), .B(new_n1049), .Y(\f[85] ));
  INVx1_ASAP7_75t_L         g665(.A(new_n1047), .Y(new_n1051));
  A2O1A1Ixp33_ASAP7_75t_L   g666(.A1(new_n1042), .A2(new_n1041), .B(new_n1040), .C(new_n1048), .Y(new_n1052));
  NOR2xp33_ASAP7_75t_L      g667(.A(\a[86] ), .B(\b[86] ), .Y(new_n1053));
  NAND2xp33_ASAP7_75t_L     g668(.A(\b[86] ), .B(\a[86] ), .Y(new_n1054));
  INVx1_ASAP7_75t_L         g669(.A(new_n1054), .Y(new_n1055));
  NOR2xp33_ASAP7_75t_L      g670(.A(new_n1053), .B(new_n1055), .Y(new_n1056));
  INVx1_ASAP7_75t_L         g671(.A(new_n1056), .Y(new_n1057));
  AND3x1_ASAP7_75t_L        g672(.A(new_n1052), .B(new_n1057), .C(new_n1051), .Y(new_n1058));
  O2A1O1Ixp33_ASAP7_75t_L   g673(.A1(new_n1045), .A2(new_n1046), .B(new_n1052), .C(new_n1057), .Y(new_n1059));
  NOR2xp33_ASAP7_75t_L      g674(.A(new_n1059), .B(new_n1058), .Y(\f[86] ));
  NOR2xp33_ASAP7_75t_L      g675(.A(\a[87] ), .B(\b[87] ), .Y(new_n1061));
  AND2x2_ASAP7_75t_L        g676(.A(\a[87] ), .B(\b[87] ), .Y(new_n1062));
  NOR2xp33_ASAP7_75t_L      g677(.A(new_n1061), .B(new_n1062), .Y(new_n1063));
  A2O1A1Ixp33_ASAP7_75t_L   g678(.A1(new_n1052), .A2(new_n1051), .B(new_n1053), .C(new_n1054), .Y(new_n1064));
  XOR2x2_ASAP7_75t_L        g679(.A(new_n1063), .B(new_n1064), .Y(\f[87] ));
  NOR2xp33_ASAP7_75t_L      g680(.A(\a[88] ), .B(\b[88] ), .Y(new_n1066));
  INVx1_ASAP7_75t_L         g681(.A(\a[88] ), .Y(new_n1067));
  INVx1_ASAP7_75t_L         g682(.A(\b[88] ), .Y(new_n1068));
  NOR2xp33_ASAP7_75t_L      g683(.A(new_n1067), .B(new_n1068), .Y(new_n1069));
  NOR2xp33_ASAP7_75t_L      g684(.A(new_n1066), .B(new_n1069), .Y(new_n1070));
  O2A1O1Ixp33_ASAP7_75t_L   g685(.A1(new_n1055), .A2(new_n1059), .B(new_n1063), .C(new_n1062), .Y(new_n1071));
  XNOR2x2_ASAP7_75t_L       g686(.A(new_n1070), .B(new_n1071), .Y(\f[88] ));
  INVx1_ASAP7_75t_L         g687(.A(new_n1069), .Y(new_n1073));
  A2O1A1Ixp33_ASAP7_75t_L   g688(.A1(new_n1064), .A2(new_n1063), .B(new_n1062), .C(new_n1070), .Y(new_n1074));
  NOR2xp33_ASAP7_75t_L      g689(.A(\a[89] ), .B(\b[89] ), .Y(new_n1075));
  NAND2xp33_ASAP7_75t_L     g690(.A(\b[89] ), .B(\a[89] ), .Y(new_n1076));
  INVx1_ASAP7_75t_L         g691(.A(new_n1076), .Y(new_n1077));
  NOR2xp33_ASAP7_75t_L      g692(.A(new_n1075), .B(new_n1077), .Y(new_n1078));
  INVx1_ASAP7_75t_L         g693(.A(new_n1078), .Y(new_n1079));
  AND3x1_ASAP7_75t_L        g694(.A(new_n1074), .B(new_n1079), .C(new_n1073), .Y(new_n1080));
  O2A1O1Ixp33_ASAP7_75t_L   g695(.A1(new_n1067), .A2(new_n1068), .B(new_n1074), .C(new_n1079), .Y(new_n1081));
  NOR2xp33_ASAP7_75t_L      g696(.A(new_n1081), .B(new_n1080), .Y(\f[89] ));
  NOR2xp33_ASAP7_75t_L      g697(.A(\a[90] ), .B(\b[90] ), .Y(new_n1083));
  AND2x2_ASAP7_75t_L        g698(.A(\a[90] ), .B(\b[90] ), .Y(new_n1084));
  NOR2xp33_ASAP7_75t_L      g699(.A(new_n1083), .B(new_n1084), .Y(new_n1085));
  A2O1A1Ixp33_ASAP7_75t_L   g700(.A1(new_n1074), .A2(new_n1073), .B(new_n1075), .C(new_n1076), .Y(new_n1086));
  XOR2x2_ASAP7_75t_L        g701(.A(new_n1085), .B(new_n1086), .Y(\f[90] ));
  NOR2xp33_ASAP7_75t_L      g702(.A(\a[91] ), .B(\b[91] ), .Y(new_n1088));
  INVx1_ASAP7_75t_L         g703(.A(\a[91] ), .Y(new_n1089));
  INVx1_ASAP7_75t_L         g704(.A(\b[91] ), .Y(new_n1090));
  NOR2xp33_ASAP7_75t_L      g705(.A(new_n1089), .B(new_n1090), .Y(new_n1091));
  NOR2xp33_ASAP7_75t_L      g706(.A(new_n1088), .B(new_n1091), .Y(new_n1092));
  O2A1O1Ixp33_ASAP7_75t_L   g707(.A1(new_n1077), .A2(new_n1081), .B(new_n1085), .C(new_n1084), .Y(new_n1093));
  XNOR2x2_ASAP7_75t_L       g708(.A(new_n1092), .B(new_n1093), .Y(\f[91] ));
  INVx1_ASAP7_75t_L         g709(.A(new_n1091), .Y(new_n1095));
  A2O1A1Ixp33_ASAP7_75t_L   g710(.A1(new_n1086), .A2(new_n1085), .B(new_n1084), .C(new_n1092), .Y(new_n1096));
  NOR2xp33_ASAP7_75t_L      g711(.A(\a[92] ), .B(\b[92] ), .Y(new_n1097));
  NAND2xp33_ASAP7_75t_L     g712(.A(\b[92] ), .B(\a[92] ), .Y(new_n1098));
  INVx1_ASAP7_75t_L         g713(.A(new_n1098), .Y(new_n1099));
  NOR2xp33_ASAP7_75t_L      g714(.A(new_n1097), .B(new_n1099), .Y(new_n1100));
  INVx1_ASAP7_75t_L         g715(.A(new_n1100), .Y(new_n1101));
  AND3x1_ASAP7_75t_L        g716(.A(new_n1096), .B(new_n1101), .C(new_n1095), .Y(new_n1102));
  O2A1O1Ixp33_ASAP7_75t_L   g717(.A1(new_n1089), .A2(new_n1090), .B(new_n1096), .C(new_n1101), .Y(new_n1103));
  NOR2xp33_ASAP7_75t_L      g718(.A(new_n1103), .B(new_n1102), .Y(\f[92] ));
  NOR2xp33_ASAP7_75t_L      g719(.A(\a[93] ), .B(\b[93] ), .Y(new_n1105));
  AND2x2_ASAP7_75t_L        g720(.A(\a[93] ), .B(\b[93] ), .Y(new_n1106));
  NOR2xp33_ASAP7_75t_L      g721(.A(new_n1105), .B(new_n1106), .Y(new_n1107));
  A2O1A1Ixp33_ASAP7_75t_L   g722(.A1(new_n1096), .A2(new_n1095), .B(new_n1097), .C(new_n1098), .Y(new_n1108));
  XOR2x2_ASAP7_75t_L        g723(.A(new_n1107), .B(new_n1108), .Y(\f[93] ));
  NOR2xp33_ASAP7_75t_L      g724(.A(\a[94] ), .B(\b[94] ), .Y(new_n1110));
  INVx1_ASAP7_75t_L         g725(.A(\a[94] ), .Y(new_n1111));
  INVx1_ASAP7_75t_L         g726(.A(\b[94] ), .Y(new_n1112));
  NOR2xp33_ASAP7_75t_L      g727(.A(new_n1111), .B(new_n1112), .Y(new_n1113));
  NOR2xp33_ASAP7_75t_L      g728(.A(new_n1110), .B(new_n1113), .Y(new_n1114));
  O2A1O1Ixp33_ASAP7_75t_L   g729(.A1(new_n1099), .A2(new_n1103), .B(new_n1107), .C(new_n1106), .Y(new_n1115));
  XNOR2x2_ASAP7_75t_L       g730(.A(new_n1114), .B(new_n1115), .Y(\f[94] ));
  INVx1_ASAP7_75t_L         g731(.A(new_n1113), .Y(new_n1117));
  A2O1A1Ixp33_ASAP7_75t_L   g732(.A1(new_n1108), .A2(new_n1107), .B(new_n1106), .C(new_n1114), .Y(new_n1118));
  NOR2xp33_ASAP7_75t_L      g733(.A(\a[95] ), .B(\b[95] ), .Y(new_n1119));
  NAND2xp33_ASAP7_75t_L     g734(.A(\b[95] ), .B(\a[95] ), .Y(new_n1120));
  INVx1_ASAP7_75t_L         g735(.A(new_n1120), .Y(new_n1121));
  NOR2xp33_ASAP7_75t_L      g736(.A(new_n1119), .B(new_n1121), .Y(new_n1122));
  INVx1_ASAP7_75t_L         g737(.A(new_n1122), .Y(new_n1123));
  AND3x1_ASAP7_75t_L        g738(.A(new_n1118), .B(new_n1123), .C(new_n1117), .Y(new_n1124));
  O2A1O1Ixp33_ASAP7_75t_L   g739(.A1(new_n1111), .A2(new_n1112), .B(new_n1118), .C(new_n1123), .Y(new_n1125));
  NOR2xp33_ASAP7_75t_L      g740(.A(new_n1125), .B(new_n1124), .Y(\f[95] ));
  NOR2xp33_ASAP7_75t_L      g741(.A(\a[96] ), .B(\b[96] ), .Y(new_n1127));
  AND2x2_ASAP7_75t_L        g742(.A(\a[96] ), .B(\b[96] ), .Y(new_n1128));
  NOR2xp33_ASAP7_75t_L      g743(.A(new_n1127), .B(new_n1128), .Y(new_n1129));
  A2O1A1Ixp33_ASAP7_75t_L   g744(.A1(new_n1118), .A2(new_n1117), .B(new_n1119), .C(new_n1120), .Y(new_n1130));
  XOR2x2_ASAP7_75t_L        g745(.A(new_n1129), .B(new_n1130), .Y(\f[96] ));
  NOR2xp33_ASAP7_75t_L      g746(.A(\a[97] ), .B(\b[97] ), .Y(new_n1132));
  INVx1_ASAP7_75t_L         g747(.A(\a[97] ), .Y(new_n1133));
  INVx1_ASAP7_75t_L         g748(.A(\b[97] ), .Y(new_n1134));
  NOR2xp33_ASAP7_75t_L      g749(.A(new_n1133), .B(new_n1134), .Y(new_n1135));
  NOR2xp33_ASAP7_75t_L      g750(.A(new_n1132), .B(new_n1135), .Y(new_n1136));
  O2A1O1Ixp33_ASAP7_75t_L   g751(.A1(new_n1121), .A2(new_n1125), .B(new_n1129), .C(new_n1128), .Y(new_n1137));
  XNOR2x2_ASAP7_75t_L       g752(.A(new_n1136), .B(new_n1137), .Y(\f[97] ));
  INVx1_ASAP7_75t_L         g753(.A(new_n1135), .Y(new_n1139));
  A2O1A1Ixp33_ASAP7_75t_L   g754(.A1(new_n1130), .A2(new_n1129), .B(new_n1128), .C(new_n1136), .Y(new_n1140));
  NOR2xp33_ASAP7_75t_L      g755(.A(\a[98] ), .B(\b[98] ), .Y(new_n1141));
  NAND2xp33_ASAP7_75t_L     g756(.A(\b[98] ), .B(\a[98] ), .Y(new_n1142));
  INVx1_ASAP7_75t_L         g757(.A(new_n1142), .Y(new_n1143));
  NOR2xp33_ASAP7_75t_L      g758(.A(new_n1141), .B(new_n1143), .Y(new_n1144));
  INVx1_ASAP7_75t_L         g759(.A(new_n1144), .Y(new_n1145));
  AND3x1_ASAP7_75t_L        g760(.A(new_n1140), .B(new_n1145), .C(new_n1139), .Y(new_n1146));
  O2A1O1Ixp33_ASAP7_75t_L   g761(.A1(new_n1133), .A2(new_n1134), .B(new_n1140), .C(new_n1145), .Y(new_n1147));
  NOR2xp33_ASAP7_75t_L      g762(.A(new_n1147), .B(new_n1146), .Y(\f[98] ));
  NOR2xp33_ASAP7_75t_L      g763(.A(\a[99] ), .B(\b[99] ), .Y(new_n1149));
  AND2x2_ASAP7_75t_L        g764(.A(\a[99] ), .B(\b[99] ), .Y(new_n1150));
  NOR2xp33_ASAP7_75t_L      g765(.A(new_n1149), .B(new_n1150), .Y(new_n1151));
  A2O1A1Ixp33_ASAP7_75t_L   g766(.A1(new_n1140), .A2(new_n1139), .B(new_n1141), .C(new_n1142), .Y(new_n1152));
  XOR2x2_ASAP7_75t_L        g767(.A(new_n1151), .B(new_n1152), .Y(\f[99] ));
  NOR2xp33_ASAP7_75t_L      g768(.A(\a[100] ), .B(\b[100] ), .Y(new_n1154));
  INVx1_ASAP7_75t_L         g769(.A(\a[100] ), .Y(new_n1155));
  INVx1_ASAP7_75t_L         g770(.A(\b[100] ), .Y(new_n1156));
  NOR2xp33_ASAP7_75t_L      g771(.A(new_n1155), .B(new_n1156), .Y(new_n1157));
  NOR2xp33_ASAP7_75t_L      g772(.A(new_n1154), .B(new_n1157), .Y(new_n1158));
  O2A1O1Ixp33_ASAP7_75t_L   g773(.A1(new_n1143), .A2(new_n1147), .B(new_n1151), .C(new_n1150), .Y(new_n1159));
  XNOR2x2_ASAP7_75t_L       g774(.A(new_n1158), .B(new_n1159), .Y(\f[100] ));
  INVx1_ASAP7_75t_L         g775(.A(new_n1157), .Y(new_n1161));
  A2O1A1Ixp33_ASAP7_75t_L   g776(.A1(new_n1152), .A2(new_n1151), .B(new_n1150), .C(new_n1158), .Y(new_n1162));
  NOR2xp33_ASAP7_75t_L      g777(.A(\a[101] ), .B(\b[101] ), .Y(new_n1163));
  NAND2xp33_ASAP7_75t_L     g778(.A(\b[101] ), .B(\a[101] ), .Y(new_n1164));
  INVx1_ASAP7_75t_L         g779(.A(new_n1164), .Y(new_n1165));
  NOR2xp33_ASAP7_75t_L      g780(.A(new_n1163), .B(new_n1165), .Y(new_n1166));
  INVx1_ASAP7_75t_L         g781(.A(new_n1166), .Y(new_n1167));
  AND3x1_ASAP7_75t_L        g782(.A(new_n1162), .B(new_n1167), .C(new_n1161), .Y(new_n1168));
  O2A1O1Ixp33_ASAP7_75t_L   g783(.A1(new_n1155), .A2(new_n1156), .B(new_n1162), .C(new_n1167), .Y(new_n1169));
  NOR2xp33_ASAP7_75t_L      g784(.A(new_n1169), .B(new_n1168), .Y(\f[101] ));
  NOR2xp33_ASAP7_75t_L      g785(.A(\a[102] ), .B(\b[102] ), .Y(new_n1171));
  AND2x2_ASAP7_75t_L        g786(.A(\a[102] ), .B(\b[102] ), .Y(new_n1172));
  NOR2xp33_ASAP7_75t_L      g787(.A(new_n1171), .B(new_n1172), .Y(new_n1173));
  A2O1A1Ixp33_ASAP7_75t_L   g788(.A1(new_n1162), .A2(new_n1161), .B(new_n1163), .C(new_n1164), .Y(new_n1174));
  XOR2x2_ASAP7_75t_L        g789(.A(new_n1173), .B(new_n1174), .Y(\f[102] ));
  NOR2xp33_ASAP7_75t_L      g790(.A(\a[103] ), .B(\b[103] ), .Y(new_n1176));
  INVx1_ASAP7_75t_L         g791(.A(\a[103] ), .Y(new_n1177));
  INVx1_ASAP7_75t_L         g792(.A(\b[103] ), .Y(new_n1178));
  NOR2xp33_ASAP7_75t_L      g793(.A(new_n1177), .B(new_n1178), .Y(new_n1179));
  NOR2xp33_ASAP7_75t_L      g794(.A(new_n1176), .B(new_n1179), .Y(new_n1180));
  O2A1O1Ixp33_ASAP7_75t_L   g795(.A1(new_n1165), .A2(new_n1169), .B(new_n1173), .C(new_n1172), .Y(new_n1181));
  XNOR2x2_ASAP7_75t_L       g796(.A(new_n1180), .B(new_n1181), .Y(\f[103] ));
  INVx1_ASAP7_75t_L         g797(.A(new_n1179), .Y(new_n1183));
  A2O1A1Ixp33_ASAP7_75t_L   g798(.A1(new_n1174), .A2(new_n1173), .B(new_n1172), .C(new_n1180), .Y(new_n1184));
  NOR2xp33_ASAP7_75t_L      g799(.A(\a[104] ), .B(\b[104] ), .Y(new_n1185));
  NAND2xp33_ASAP7_75t_L     g800(.A(\b[104] ), .B(\a[104] ), .Y(new_n1186));
  INVx1_ASAP7_75t_L         g801(.A(new_n1186), .Y(new_n1187));
  NOR2xp33_ASAP7_75t_L      g802(.A(new_n1185), .B(new_n1187), .Y(new_n1188));
  INVx1_ASAP7_75t_L         g803(.A(new_n1188), .Y(new_n1189));
  AND3x1_ASAP7_75t_L        g804(.A(new_n1184), .B(new_n1189), .C(new_n1183), .Y(new_n1190));
  O2A1O1Ixp33_ASAP7_75t_L   g805(.A1(new_n1177), .A2(new_n1178), .B(new_n1184), .C(new_n1189), .Y(new_n1191));
  NOR2xp33_ASAP7_75t_L      g806(.A(new_n1191), .B(new_n1190), .Y(\f[104] ));
  NOR2xp33_ASAP7_75t_L      g807(.A(\a[105] ), .B(\b[105] ), .Y(new_n1193));
  AND2x2_ASAP7_75t_L        g808(.A(\a[105] ), .B(\b[105] ), .Y(new_n1194));
  NOR2xp33_ASAP7_75t_L      g809(.A(new_n1193), .B(new_n1194), .Y(new_n1195));
  A2O1A1Ixp33_ASAP7_75t_L   g810(.A1(new_n1184), .A2(new_n1183), .B(new_n1185), .C(new_n1186), .Y(new_n1196));
  XOR2x2_ASAP7_75t_L        g811(.A(new_n1195), .B(new_n1196), .Y(\f[105] ));
  NOR2xp33_ASAP7_75t_L      g812(.A(\a[106] ), .B(\b[106] ), .Y(new_n1198));
  INVx1_ASAP7_75t_L         g813(.A(\a[106] ), .Y(new_n1199));
  INVx1_ASAP7_75t_L         g814(.A(\b[106] ), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g815(.A(new_n1199), .B(new_n1200), .Y(new_n1201));
  NOR2xp33_ASAP7_75t_L      g816(.A(new_n1198), .B(new_n1201), .Y(new_n1202));
  O2A1O1Ixp33_ASAP7_75t_L   g817(.A1(new_n1187), .A2(new_n1191), .B(new_n1195), .C(new_n1194), .Y(new_n1203));
  XNOR2x2_ASAP7_75t_L       g818(.A(new_n1202), .B(new_n1203), .Y(\f[106] ));
  INVx1_ASAP7_75t_L         g819(.A(new_n1201), .Y(new_n1205));
  A2O1A1Ixp33_ASAP7_75t_L   g820(.A1(new_n1196), .A2(new_n1195), .B(new_n1194), .C(new_n1202), .Y(new_n1206));
  NOR2xp33_ASAP7_75t_L      g821(.A(\a[107] ), .B(\b[107] ), .Y(new_n1207));
  NAND2xp33_ASAP7_75t_L     g822(.A(\b[107] ), .B(\a[107] ), .Y(new_n1208));
  INVx1_ASAP7_75t_L         g823(.A(new_n1208), .Y(new_n1209));
  NOR2xp33_ASAP7_75t_L      g824(.A(new_n1207), .B(new_n1209), .Y(new_n1210));
  INVx1_ASAP7_75t_L         g825(.A(new_n1210), .Y(new_n1211));
  AND3x1_ASAP7_75t_L        g826(.A(new_n1206), .B(new_n1211), .C(new_n1205), .Y(new_n1212));
  O2A1O1Ixp33_ASAP7_75t_L   g827(.A1(new_n1199), .A2(new_n1200), .B(new_n1206), .C(new_n1211), .Y(new_n1213));
  NOR2xp33_ASAP7_75t_L      g828(.A(new_n1213), .B(new_n1212), .Y(\f[107] ));
  NOR2xp33_ASAP7_75t_L      g829(.A(\a[108] ), .B(\b[108] ), .Y(new_n1215));
  AND2x2_ASAP7_75t_L        g830(.A(\a[108] ), .B(\b[108] ), .Y(new_n1216));
  NOR2xp33_ASAP7_75t_L      g831(.A(new_n1215), .B(new_n1216), .Y(new_n1217));
  A2O1A1Ixp33_ASAP7_75t_L   g832(.A1(new_n1206), .A2(new_n1205), .B(new_n1207), .C(new_n1208), .Y(new_n1218));
  XOR2x2_ASAP7_75t_L        g833(.A(new_n1217), .B(new_n1218), .Y(\f[108] ));
  NOR2xp33_ASAP7_75t_L      g834(.A(\a[109] ), .B(\b[109] ), .Y(new_n1220));
  INVx1_ASAP7_75t_L         g835(.A(\a[109] ), .Y(new_n1221));
  INVx1_ASAP7_75t_L         g836(.A(\b[109] ), .Y(new_n1222));
  NOR2xp33_ASAP7_75t_L      g837(.A(new_n1221), .B(new_n1222), .Y(new_n1223));
  NOR2xp33_ASAP7_75t_L      g838(.A(new_n1220), .B(new_n1223), .Y(new_n1224));
  O2A1O1Ixp33_ASAP7_75t_L   g839(.A1(new_n1209), .A2(new_n1213), .B(new_n1217), .C(new_n1216), .Y(new_n1225));
  XNOR2x2_ASAP7_75t_L       g840(.A(new_n1224), .B(new_n1225), .Y(\f[109] ));
  INVx1_ASAP7_75t_L         g841(.A(new_n1223), .Y(new_n1227));
  A2O1A1Ixp33_ASAP7_75t_L   g842(.A1(new_n1218), .A2(new_n1217), .B(new_n1216), .C(new_n1224), .Y(new_n1228));
  NOR2xp33_ASAP7_75t_L      g843(.A(\a[110] ), .B(\b[110] ), .Y(new_n1229));
  NAND2xp33_ASAP7_75t_L     g844(.A(\b[110] ), .B(\a[110] ), .Y(new_n1230));
  INVx1_ASAP7_75t_L         g845(.A(new_n1230), .Y(new_n1231));
  NOR2xp33_ASAP7_75t_L      g846(.A(new_n1229), .B(new_n1231), .Y(new_n1232));
  INVx1_ASAP7_75t_L         g847(.A(new_n1232), .Y(new_n1233));
  AND3x1_ASAP7_75t_L        g848(.A(new_n1228), .B(new_n1233), .C(new_n1227), .Y(new_n1234));
  O2A1O1Ixp33_ASAP7_75t_L   g849(.A1(new_n1221), .A2(new_n1222), .B(new_n1228), .C(new_n1233), .Y(new_n1235));
  NOR2xp33_ASAP7_75t_L      g850(.A(new_n1235), .B(new_n1234), .Y(\f[110] ));
  NOR2xp33_ASAP7_75t_L      g851(.A(\a[111] ), .B(\b[111] ), .Y(new_n1237));
  AND2x2_ASAP7_75t_L        g852(.A(\a[111] ), .B(\b[111] ), .Y(new_n1238));
  NOR2xp33_ASAP7_75t_L      g853(.A(new_n1237), .B(new_n1238), .Y(new_n1239));
  A2O1A1Ixp33_ASAP7_75t_L   g854(.A1(new_n1228), .A2(new_n1227), .B(new_n1229), .C(new_n1230), .Y(new_n1240));
  XOR2x2_ASAP7_75t_L        g855(.A(new_n1239), .B(new_n1240), .Y(\f[111] ));
  NOR2xp33_ASAP7_75t_L      g856(.A(\a[112] ), .B(\b[112] ), .Y(new_n1242));
  INVx1_ASAP7_75t_L         g857(.A(\a[112] ), .Y(new_n1243));
  INVx1_ASAP7_75t_L         g858(.A(\b[112] ), .Y(new_n1244));
  NOR2xp33_ASAP7_75t_L      g859(.A(new_n1243), .B(new_n1244), .Y(new_n1245));
  NOR2xp33_ASAP7_75t_L      g860(.A(new_n1242), .B(new_n1245), .Y(new_n1246));
  O2A1O1Ixp33_ASAP7_75t_L   g861(.A1(new_n1231), .A2(new_n1235), .B(new_n1239), .C(new_n1238), .Y(new_n1247));
  XNOR2x2_ASAP7_75t_L       g862(.A(new_n1246), .B(new_n1247), .Y(\f[112] ));
  INVx1_ASAP7_75t_L         g863(.A(new_n1245), .Y(new_n1249));
  A2O1A1Ixp33_ASAP7_75t_L   g864(.A1(new_n1240), .A2(new_n1239), .B(new_n1238), .C(new_n1246), .Y(new_n1250));
  NOR2xp33_ASAP7_75t_L      g865(.A(\a[113] ), .B(\b[113] ), .Y(new_n1251));
  NAND2xp33_ASAP7_75t_L     g866(.A(\b[113] ), .B(\a[113] ), .Y(new_n1252));
  INVx1_ASAP7_75t_L         g867(.A(new_n1252), .Y(new_n1253));
  NOR2xp33_ASAP7_75t_L      g868(.A(new_n1251), .B(new_n1253), .Y(new_n1254));
  INVx1_ASAP7_75t_L         g869(.A(new_n1254), .Y(new_n1255));
  AND3x1_ASAP7_75t_L        g870(.A(new_n1250), .B(new_n1255), .C(new_n1249), .Y(new_n1256));
  O2A1O1Ixp33_ASAP7_75t_L   g871(.A1(new_n1243), .A2(new_n1244), .B(new_n1250), .C(new_n1255), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g872(.A(new_n1257), .B(new_n1256), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g873(.A(\a[114] ), .B(\b[114] ), .Y(new_n1259));
  AND2x2_ASAP7_75t_L        g874(.A(\a[114] ), .B(\b[114] ), .Y(new_n1260));
  NOR2xp33_ASAP7_75t_L      g875(.A(new_n1259), .B(new_n1260), .Y(new_n1261));
  A2O1A1Ixp33_ASAP7_75t_L   g876(.A1(new_n1250), .A2(new_n1249), .B(new_n1251), .C(new_n1252), .Y(new_n1262));
  XOR2x2_ASAP7_75t_L        g877(.A(new_n1261), .B(new_n1262), .Y(\f[114] ));
  NOR2xp33_ASAP7_75t_L      g878(.A(\a[115] ), .B(\b[115] ), .Y(new_n1264));
  INVx1_ASAP7_75t_L         g879(.A(\a[115] ), .Y(new_n1265));
  INVx1_ASAP7_75t_L         g880(.A(\b[115] ), .Y(new_n1266));
  NOR2xp33_ASAP7_75t_L      g881(.A(new_n1265), .B(new_n1266), .Y(new_n1267));
  NOR2xp33_ASAP7_75t_L      g882(.A(new_n1264), .B(new_n1267), .Y(new_n1268));
  O2A1O1Ixp33_ASAP7_75t_L   g883(.A1(new_n1253), .A2(new_n1257), .B(new_n1261), .C(new_n1260), .Y(new_n1269));
  XNOR2x2_ASAP7_75t_L       g884(.A(new_n1268), .B(new_n1269), .Y(\f[115] ));
  INVx1_ASAP7_75t_L         g885(.A(new_n1267), .Y(new_n1271));
  A2O1A1Ixp33_ASAP7_75t_L   g886(.A1(new_n1262), .A2(new_n1261), .B(new_n1260), .C(new_n1268), .Y(new_n1272));
  NOR2xp33_ASAP7_75t_L      g887(.A(\a[116] ), .B(\b[116] ), .Y(new_n1273));
  NAND2xp33_ASAP7_75t_L     g888(.A(\b[116] ), .B(\a[116] ), .Y(new_n1274));
  INVx1_ASAP7_75t_L         g889(.A(new_n1274), .Y(new_n1275));
  NOR2xp33_ASAP7_75t_L      g890(.A(new_n1273), .B(new_n1275), .Y(new_n1276));
  INVx1_ASAP7_75t_L         g891(.A(new_n1276), .Y(new_n1277));
  AND3x1_ASAP7_75t_L        g892(.A(new_n1272), .B(new_n1277), .C(new_n1271), .Y(new_n1278));
  O2A1O1Ixp33_ASAP7_75t_L   g893(.A1(new_n1265), .A2(new_n1266), .B(new_n1272), .C(new_n1277), .Y(new_n1279));
  NOR2xp33_ASAP7_75t_L      g894(.A(new_n1279), .B(new_n1278), .Y(\f[116] ));
  NOR2xp33_ASAP7_75t_L      g895(.A(\a[117] ), .B(\b[117] ), .Y(new_n1281));
  AND2x2_ASAP7_75t_L        g896(.A(\a[117] ), .B(\b[117] ), .Y(new_n1282));
  NOR2xp33_ASAP7_75t_L      g897(.A(new_n1281), .B(new_n1282), .Y(new_n1283));
  A2O1A1Ixp33_ASAP7_75t_L   g898(.A1(new_n1272), .A2(new_n1271), .B(new_n1273), .C(new_n1274), .Y(new_n1284));
  XOR2x2_ASAP7_75t_L        g899(.A(new_n1283), .B(new_n1284), .Y(\f[117] ));
  NOR2xp33_ASAP7_75t_L      g900(.A(\a[118] ), .B(\b[118] ), .Y(new_n1286));
  INVx1_ASAP7_75t_L         g901(.A(\a[118] ), .Y(new_n1287));
  INVx1_ASAP7_75t_L         g902(.A(\b[118] ), .Y(new_n1288));
  NOR2xp33_ASAP7_75t_L      g903(.A(new_n1287), .B(new_n1288), .Y(new_n1289));
  NOR2xp33_ASAP7_75t_L      g904(.A(new_n1286), .B(new_n1289), .Y(new_n1290));
  O2A1O1Ixp33_ASAP7_75t_L   g905(.A1(new_n1275), .A2(new_n1279), .B(new_n1283), .C(new_n1282), .Y(new_n1291));
  XNOR2x2_ASAP7_75t_L       g906(.A(new_n1290), .B(new_n1291), .Y(\f[118] ));
  INVx1_ASAP7_75t_L         g907(.A(new_n1289), .Y(new_n1293));
  A2O1A1Ixp33_ASAP7_75t_L   g908(.A1(new_n1284), .A2(new_n1283), .B(new_n1282), .C(new_n1290), .Y(new_n1294));
  NOR2xp33_ASAP7_75t_L      g909(.A(\a[119] ), .B(\b[119] ), .Y(new_n1295));
  NAND2xp33_ASAP7_75t_L     g910(.A(\b[119] ), .B(\a[119] ), .Y(new_n1296));
  INVx1_ASAP7_75t_L         g911(.A(new_n1296), .Y(new_n1297));
  NOR2xp33_ASAP7_75t_L      g912(.A(new_n1295), .B(new_n1297), .Y(new_n1298));
  INVx1_ASAP7_75t_L         g913(.A(new_n1298), .Y(new_n1299));
  AND3x1_ASAP7_75t_L        g914(.A(new_n1294), .B(new_n1299), .C(new_n1293), .Y(new_n1300));
  O2A1O1Ixp33_ASAP7_75t_L   g915(.A1(new_n1287), .A2(new_n1288), .B(new_n1294), .C(new_n1299), .Y(new_n1301));
  NOR2xp33_ASAP7_75t_L      g916(.A(new_n1301), .B(new_n1300), .Y(\f[119] ));
  NOR2xp33_ASAP7_75t_L      g917(.A(\a[120] ), .B(\b[120] ), .Y(new_n1303));
  INVx1_ASAP7_75t_L         g918(.A(\a[120] ), .Y(new_n1304));
  INVx1_ASAP7_75t_L         g919(.A(\b[120] ), .Y(new_n1305));
  NOR2xp33_ASAP7_75t_L      g920(.A(new_n1304), .B(new_n1305), .Y(new_n1306));
  NOR2xp33_ASAP7_75t_L      g921(.A(new_n1303), .B(new_n1306), .Y(new_n1307));
  A2O1A1Ixp33_ASAP7_75t_L   g922(.A1(new_n1294), .A2(new_n1293), .B(new_n1295), .C(new_n1296), .Y(new_n1308));
  XOR2x2_ASAP7_75t_L        g923(.A(new_n1307), .B(new_n1308), .Y(\f[120] ));
  NOR2xp33_ASAP7_75t_L      g924(.A(\a[121] ), .B(\b[121] ), .Y(new_n1310));
  NAND2xp33_ASAP7_75t_L     g925(.A(\b[121] ), .B(\a[121] ), .Y(new_n1311));
  INVx1_ASAP7_75t_L         g926(.A(new_n1311), .Y(new_n1312));
  NOR2xp33_ASAP7_75t_L      g927(.A(new_n1310), .B(new_n1312), .Y(new_n1313));
  AOI211xp5_ASAP7_75t_L     g928(.A1(new_n1308), .A2(new_n1307), .B(new_n1313), .C(new_n1306), .Y(new_n1314));
  A2O1A1Ixp33_ASAP7_75t_L   g929(.A1(new_n1308), .A2(new_n1307), .B(new_n1306), .C(new_n1313), .Y(new_n1315));
  INVx1_ASAP7_75t_L         g930(.A(new_n1315), .Y(new_n1316));
  NOR2xp33_ASAP7_75t_L      g931(.A(new_n1314), .B(new_n1316), .Y(\f[121] ));
  NOR2xp33_ASAP7_75t_L      g932(.A(\a[122] ), .B(\b[122] ), .Y(new_n1318));
  INVx1_ASAP7_75t_L         g933(.A(\a[122] ), .Y(new_n1319));
  INVx1_ASAP7_75t_L         g934(.A(\b[122] ), .Y(new_n1320));
  NOR2xp33_ASAP7_75t_L      g935(.A(new_n1319), .B(new_n1320), .Y(new_n1321));
  NOR2xp33_ASAP7_75t_L      g936(.A(new_n1318), .B(new_n1321), .Y(new_n1322));
  A2O1A1O1Ixp25_ASAP7_75t_L g937(.A1(new_n1307), .A2(new_n1308), .B(new_n1306), .C(new_n1313), .D(new_n1312), .Y(new_n1323));
  XNOR2x2_ASAP7_75t_L       g938(.A(new_n1322), .B(new_n1323), .Y(\f[122] ));
  NOR2xp33_ASAP7_75t_L      g939(.A(\a[123] ), .B(\b[123] ), .Y(new_n1325));
  NAND2xp33_ASAP7_75t_L     g940(.A(\b[123] ), .B(\a[123] ), .Y(new_n1326));
  INVx1_ASAP7_75t_L         g941(.A(new_n1326), .Y(new_n1327));
  NOR2xp33_ASAP7_75t_L      g942(.A(new_n1325), .B(new_n1327), .Y(new_n1328));
  INVx1_ASAP7_75t_L         g943(.A(new_n1321), .Y(new_n1329));
  A2O1A1Ixp33_ASAP7_75t_L   g944(.A1(new_n1315), .A2(new_n1311), .B(new_n1318), .C(new_n1329), .Y(new_n1330));
  NOR2xp33_ASAP7_75t_L      g945(.A(new_n1328), .B(new_n1330), .Y(new_n1331));
  INVx1_ASAP7_75t_L         g946(.A(new_n1328), .Y(new_n1332));
  A2O1A1O1Ixp25_ASAP7_75t_L g947(.A1(new_n1311), .A2(new_n1315), .B(new_n1318), .C(new_n1329), .D(new_n1332), .Y(new_n1333));
  NOR2xp33_ASAP7_75t_L      g948(.A(new_n1333), .B(new_n1331), .Y(\f[123] ));
  NOR2xp33_ASAP7_75t_L      g949(.A(\a[124] ), .B(\b[124] ), .Y(new_n1335));
  INVx1_ASAP7_75t_L         g950(.A(\a[124] ), .Y(new_n1336));
  INVx1_ASAP7_75t_L         g951(.A(\b[124] ), .Y(new_n1337));
  NOR2xp33_ASAP7_75t_L      g952(.A(new_n1336), .B(new_n1337), .Y(new_n1338));
  NOR2xp33_ASAP7_75t_L      g953(.A(new_n1335), .B(new_n1338), .Y(new_n1339));
  A2O1A1Ixp33_ASAP7_75t_L   g954(.A1(\b[121] ), .A2(\a[121] ), .B(new_n1316), .C(new_n1322), .Y(new_n1340));
  A2O1A1Ixp33_ASAP7_75t_L   g955(.A1(new_n1340), .A2(new_n1329), .B(new_n1325), .C(new_n1326), .Y(new_n1341));
  XOR2x2_ASAP7_75t_L        g956(.A(new_n1339), .B(new_n1341), .Y(\f[124] ));
  INVx1_ASAP7_75t_L         g957(.A(new_n1338), .Y(new_n1343));
  A2O1A1Ixp33_ASAP7_75t_L   g958(.A1(new_n1330), .A2(new_n1328), .B(new_n1327), .C(new_n1339), .Y(new_n1344));
  NOR2xp33_ASAP7_75t_L      g959(.A(\a[125] ), .B(\b[125] ), .Y(new_n1345));
  NAND2xp33_ASAP7_75t_L     g960(.A(\b[125] ), .B(\a[125] ), .Y(new_n1346));
  INVx1_ASAP7_75t_L         g961(.A(new_n1346), .Y(new_n1347));
  NOR2xp33_ASAP7_75t_L      g962(.A(new_n1345), .B(new_n1347), .Y(new_n1348));
  INVx1_ASAP7_75t_L         g963(.A(new_n1348), .Y(new_n1349));
  AND3x1_ASAP7_75t_L        g964(.A(new_n1344), .B(new_n1349), .C(new_n1343), .Y(new_n1350));
  O2A1O1Ixp33_ASAP7_75t_L   g965(.A1(new_n1336), .A2(new_n1337), .B(new_n1344), .C(new_n1349), .Y(new_n1351));
  NOR2xp33_ASAP7_75t_L      g966(.A(new_n1351), .B(new_n1350), .Y(\f[125] ));
  NOR2xp33_ASAP7_75t_L      g967(.A(\a[126] ), .B(\b[126] ), .Y(new_n1353));
  NAND2xp33_ASAP7_75t_L     g968(.A(\b[126] ), .B(\a[126] ), .Y(new_n1354));
  INVx1_ASAP7_75t_L         g969(.A(new_n1354), .Y(new_n1355));
  NOR2xp33_ASAP7_75t_L      g970(.A(new_n1353), .B(new_n1355), .Y(new_n1356));
  A2O1A1Ixp33_ASAP7_75t_L   g971(.A1(new_n1344), .A2(new_n1343), .B(new_n1345), .C(new_n1346), .Y(new_n1357));
  XOR2x2_ASAP7_75t_L        g972(.A(new_n1356), .B(new_n1357), .Y(\f[126] ));
  NOR2xp33_ASAP7_75t_L      g973(.A(\a[127] ), .B(\b[127] ), .Y(new_n1359));
  NAND2xp33_ASAP7_75t_L     g974(.A(\b[127] ), .B(\a[127] ), .Y(new_n1360));
  INVx1_ASAP7_75t_L         g975(.A(new_n1360), .Y(new_n1361));
  NOR2xp33_ASAP7_75t_L      g976(.A(new_n1359), .B(new_n1361), .Y(new_n1362));
  A2O1A1Ixp33_ASAP7_75t_L   g977(.A1(new_n1341), .A2(new_n1339), .B(new_n1338), .C(new_n1348), .Y(new_n1363));
  A2O1A1Ixp33_ASAP7_75t_L   g978(.A1(new_n1363), .A2(new_n1346), .B(new_n1353), .C(new_n1354), .Y(new_n1364));
  NOR2xp33_ASAP7_75t_L      g979(.A(new_n1362), .B(new_n1364), .Y(new_n1365));
  INVx1_ASAP7_75t_L         g980(.A(new_n1362), .Y(new_n1366));
  A2O1A1O1Ixp25_ASAP7_75t_L g981(.A1(new_n1346), .A2(new_n1363), .B(new_n1353), .C(new_n1354), .D(new_n1366), .Y(new_n1367));
  NOR2xp33_ASAP7_75t_L      g982(.A(new_n1367), .B(new_n1365), .Y(\f[127] ));
  A2O1A1Ixp33_ASAP7_75t_L   g983(.A1(\b[125] ), .A2(\a[125] ), .B(new_n1351), .C(new_n1356), .Y(new_n1369));
  A2O1A1Ixp33_ASAP7_75t_L   g984(.A1(new_n1369), .A2(new_n1354), .B(new_n1359), .C(new_n1360), .Y(cOut));
endmodule


