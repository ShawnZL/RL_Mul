// Benchmark "top" written by ABC on Mon Dec 25 17:56:46 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1677, new_n1678,
    new_n1679, new_n1680, new_n1681, new_n1682, new_n1683, new_n1684,
    new_n1685, new_n1686, new_n1687, new_n1688, new_n1689, new_n1690,
    new_n1691, new_n1692, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1698, new_n1699, new_n1700, new_n1701, new_n1702,
    new_n1703, new_n1704, new_n1705, new_n1706, new_n1707, new_n1708,
    new_n1709, new_n1710, new_n1711, new_n1712, new_n1713, new_n1714,
    new_n1715, new_n1716, new_n1717, new_n1718, new_n1719, new_n1720,
    new_n1721, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1750,
    new_n1751, new_n1752, new_n1753, new_n1754, new_n1755, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2556, new_n2557, new_n2558, new_n2559, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572,
    new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703, new_n2704, new_n2705,
    new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2999, new_n3000, new_n3001,
    new_n3002, new_n3003, new_n3004, new_n3005, new_n3006, new_n3007,
    new_n3008, new_n3009, new_n3010, new_n3011, new_n3012, new_n3013,
    new_n3014, new_n3015, new_n3016, new_n3017, new_n3018, new_n3019,
    new_n3020, new_n3021, new_n3022, new_n3023, new_n3024, new_n3025,
    new_n3026, new_n3027, new_n3028, new_n3029, new_n3030, new_n3031,
    new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037,
    new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043,
    new_n3044, new_n3045, new_n3046, new_n3047, new_n3048, new_n3049,
    new_n3050, new_n3051, new_n3052, new_n3053, new_n3054, new_n3055,
    new_n3056, new_n3057, new_n3058, new_n3059, new_n3060, new_n3061,
    new_n3062, new_n3063, new_n3064, new_n3065, new_n3066, new_n3067,
    new_n3068, new_n3069, new_n3070, new_n3071, new_n3072, new_n3073,
    new_n3074, new_n3075, new_n3076, new_n3077, new_n3078, new_n3079,
    new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085,
    new_n3086, new_n3087, new_n3088, new_n3089, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125, new_n3126, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3799, new_n3800, new_n3801, new_n3802, new_n3803,
    new_n3804, new_n3805, new_n3806, new_n3807, new_n3808, new_n3809,
    new_n3810, new_n3811, new_n3812, new_n3813, new_n3814, new_n3815,
    new_n3816, new_n3817, new_n3818, new_n3819, new_n3820, new_n3821,
    new_n3822, new_n3823, new_n3824, new_n3825, new_n3826, new_n3827,
    new_n3828, new_n3829, new_n3830, new_n3831, new_n3832, new_n3833,
    new_n3834, new_n3835, new_n3836, new_n3837, new_n3838, new_n3839,
    new_n3840, new_n3841, new_n3842, new_n3843, new_n3844, new_n3845,
    new_n3846, new_n3847, new_n3848, new_n3849, new_n3850, new_n3851,
    new_n3852, new_n3853, new_n3854, new_n3855, new_n3856, new_n3857,
    new_n3858, new_n3859, new_n3860, new_n3861, new_n3862, new_n3863,
    new_n3864, new_n3865, new_n3866, new_n3867, new_n3868, new_n3869,
    new_n3870, new_n3871, new_n3872, new_n3873, new_n3874, new_n3875,
    new_n3876, new_n3877, new_n3878, new_n3879, new_n3880, new_n3881,
    new_n3882, new_n3883, new_n3884, new_n3885, new_n3886, new_n3887,
    new_n3888, new_n3889, new_n3890, new_n3891, new_n3892, new_n3893,
    new_n3894, new_n3895, new_n3896, new_n3897, new_n3898, new_n3899,
    new_n3900, new_n3901, new_n3902, new_n3903, new_n3904, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3930, new_n3931, new_n3932, new_n3933, new_n3934, new_n3935,
    new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941,
    new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947,
    new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953,
    new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959,
    new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965,
    new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971,
    new_n3972, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977,
    new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983,
    new_n3984, new_n3985, new_n3986, new_n3987, new_n3988, new_n3989,
    new_n3990, new_n3991, new_n3992, new_n3993, new_n3994, new_n3995,
    new_n3996, new_n3997, new_n3998, new_n3999, new_n4000, new_n4001,
    new_n4002, new_n4003, new_n4004, new_n4005, new_n4006, new_n4007,
    new_n4008, new_n4009, new_n4010, new_n4011, new_n4012, new_n4013,
    new_n4014, new_n4015, new_n4016, new_n4017, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4230, new_n4231,
    new_n4232, new_n4233, new_n4234, new_n4235, new_n4236, new_n4237,
    new_n4238, new_n4239, new_n4240, new_n4241, new_n4242, new_n4243,
    new_n4244, new_n4245, new_n4246, new_n4247, new_n4248, new_n4249,
    new_n4250, new_n4251, new_n4252, new_n4253, new_n4254, new_n4255,
    new_n4256, new_n4257, new_n4258, new_n4259, new_n4260, new_n4261,
    new_n4262, new_n4263, new_n4264, new_n4265, new_n4266, new_n4267,
    new_n4268, new_n4269, new_n4270, new_n4271, new_n4272, new_n4273,
    new_n4274, new_n4275, new_n4276, new_n4277, new_n4278, new_n4279,
    new_n4280, new_n4281, new_n4282, new_n4283, new_n4284, new_n4285,
    new_n4286, new_n4287, new_n4288, new_n4289, new_n4290, new_n4291,
    new_n4292, new_n4293, new_n4294, new_n4295, new_n4296, new_n4297,
    new_n4298, new_n4299, new_n4300, new_n4301, new_n4302, new_n4303,
    new_n4304, new_n4305, new_n4306, new_n4307, new_n4308, new_n4309,
    new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325, new_n4326, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374, new_n4375,
    new_n4376, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424, new_n4425, new_n4426, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646,
    new_n4647, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5096, new_n5097, new_n5098, new_n5099,
    new_n5100, new_n5101, new_n5102, new_n5103, new_n5104, new_n5105,
    new_n5106, new_n5107, new_n5108, new_n5109, new_n5110, new_n5111,
    new_n5112, new_n5113, new_n5114, new_n5115, new_n5116, new_n5117,
    new_n5118, new_n5119, new_n5120, new_n5121, new_n5122, new_n5123,
    new_n5124, new_n5125, new_n5126, new_n5127, new_n5128, new_n5129,
    new_n5130, new_n5131, new_n5132, new_n5133, new_n5134, new_n5135,
    new_n5136, new_n5137, new_n5138, new_n5139, new_n5140, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211, new_n5212, new_n5213,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219,
    new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225,
    new_n5226, new_n5227, new_n5228, new_n5229, new_n5230, new_n5231,
    new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237,
    new_n5238, new_n5239, new_n5240, new_n5241, new_n5242, new_n5243,
    new_n5244, new_n5245, new_n5246, new_n5247, new_n5248, new_n5249,
    new_n5250, new_n5251, new_n5252, new_n5253, new_n5254, new_n5255,
    new_n5256, new_n5257, new_n5258, new_n5259, new_n5260, new_n5261,
    new_n5262, new_n5263, new_n5264, new_n5265, new_n5266, new_n5267,
    new_n5268, new_n5269, new_n5270, new_n5271, new_n5272, new_n5273,
    new_n5274, new_n5275, new_n5276, new_n5277, new_n5278, new_n5279,
    new_n5280, new_n5281, new_n5282, new_n5283, new_n5284, new_n5285,
    new_n5286, new_n5287, new_n5288, new_n5289, new_n5290, new_n5291,
    new_n5292, new_n5293, new_n5294, new_n5295, new_n5296, new_n5297,
    new_n5298, new_n5299, new_n5300, new_n5301, new_n5302, new_n5303,
    new_n5304, new_n5305, new_n5306, new_n5307, new_n5308, new_n5309,
    new_n5310, new_n5311, new_n5312, new_n5313, new_n5314, new_n5315,
    new_n5316, new_n5317, new_n5318, new_n5319, new_n5320, new_n5321,
    new_n5322, new_n5323, new_n5324, new_n5325, new_n5326, new_n5327,
    new_n5328, new_n5329, new_n5330, new_n5331, new_n5332, new_n5333,
    new_n5334, new_n5336, new_n5337, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351, new_n5352,
    new_n5353, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5585, new_n5586, new_n5587,
    new_n5588, new_n5589, new_n5590, new_n5591, new_n5592, new_n5593,
    new_n5594, new_n5595, new_n5596, new_n5597, new_n5598, new_n5599,
    new_n5600, new_n5601, new_n5602, new_n5603, new_n5604, new_n5605,
    new_n5606, new_n5607, new_n5608, new_n5609, new_n5610, new_n5611,
    new_n5612, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696, new_n5697, new_n5698, new_n5699, new_n5700, new_n5701,
    new_n5702, new_n5703, new_n5704, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765, new_n5766, new_n5767,
    new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773,
    new_n5774, new_n5775, new_n5776, new_n5777, new_n5778, new_n5779,
    new_n5780, new_n5781, new_n5782, new_n5783, new_n5784, new_n5785,
    new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791,
    new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797,
    new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803,
    new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822, new_n5823, new_n5824, new_n5826, new_n5827, new_n5828,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5833, new_n5834,
    new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840,
    new_n5841, new_n5842, new_n5843, new_n5844, new_n5845, new_n5846,
    new_n5847, new_n5848, new_n5849, new_n5850, new_n5851, new_n5852,
    new_n5853, new_n5854, new_n5855, new_n5856, new_n5857, new_n5858,
    new_n5859, new_n5860, new_n5861, new_n5862, new_n5863, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936,
    new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942,
    new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948,
    new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038,
    new_n6039, new_n6040, new_n6041, new_n6042, new_n6043, new_n6044,
    new_n6045, new_n6046, new_n6047, new_n6048, new_n6049, new_n6050,
    new_n6051, new_n6052, new_n6053, new_n6054, new_n6055, new_n6056,
    new_n6057, new_n6058, new_n6059, new_n6060, new_n6061, new_n6062,
    new_n6063, new_n6064, new_n6065, new_n6066, new_n6067, new_n6068,
    new_n6069, new_n6070, new_n6071, new_n6072, new_n6073, new_n6074,
    new_n6075, new_n6076, new_n6077, new_n6078, new_n6079, new_n6080,
    new_n6082, new_n6083, new_n6084, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104, new_n6105,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189,
    new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255,
    new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273,
    new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309,
    new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6338, new_n6339, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376,
    new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382,
    new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430,
    new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556,
    new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587,
    new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611,
    new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653,
    new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7086, new_n7087,
    new_n7088, new_n7089, new_n7090, new_n7091, new_n7092, new_n7093,
    new_n7094, new_n7095, new_n7096, new_n7097, new_n7098, new_n7099,
    new_n7100, new_n7101, new_n7102, new_n7103, new_n7104, new_n7105,
    new_n7106, new_n7107, new_n7108, new_n7109, new_n7110, new_n7111,
    new_n7112, new_n7113, new_n7114, new_n7115, new_n7116, new_n7117,
    new_n7118, new_n7119, new_n7120, new_n7121, new_n7122, new_n7123,
    new_n7124, new_n7125, new_n7126, new_n7127, new_n7128, new_n7129,
    new_n7130, new_n7131, new_n7132, new_n7133, new_n7134, new_n7135,
    new_n7136, new_n7137, new_n7138, new_n7139, new_n7140, new_n7141,
    new_n7142, new_n7143, new_n7144, new_n7145, new_n7146, new_n7147,
    new_n7148, new_n7149, new_n7150, new_n7151, new_n7152, new_n7153,
    new_n7154, new_n7155, new_n7156, new_n7157, new_n7158, new_n7159,
    new_n7160, new_n7161, new_n7162, new_n7163, new_n7164, new_n7165,
    new_n7166, new_n7167, new_n7168, new_n7169, new_n7170, new_n7171,
    new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177,
    new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183,
    new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189,
    new_n7190, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195,
    new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201,
    new_n7202, new_n7203, new_n7204, new_n7205, new_n7206, new_n7207,
    new_n7208, new_n7209, new_n7210, new_n7211, new_n7212, new_n7213,
    new_n7214, new_n7215, new_n7216, new_n7217, new_n7218, new_n7219,
    new_n7220, new_n7221, new_n7222, new_n7223, new_n7224, new_n7225,
    new_n7226, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231,
    new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237,
    new_n7238, new_n7239, new_n7240, new_n7241, new_n7242, new_n7243,
    new_n7244, new_n7245, new_n7246, new_n7247, new_n7248, new_n7249,
    new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7334,
    new_n7335, new_n7336, new_n7337, new_n7338, new_n7339, new_n7340,
    new_n7341, new_n7342, new_n7343, new_n7344, new_n7345, new_n7346,
    new_n7347, new_n7348, new_n7349, new_n7350, new_n7351, new_n7352,
    new_n7353, new_n7354, new_n7355, new_n7356, new_n7357, new_n7358,
    new_n7359, new_n7360, new_n7361, new_n7362, new_n7363, new_n7364,
    new_n7365, new_n7366, new_n7367, new_n7368, new_n7369, new_n7370,
    new_n7371, new_n7372, new_n7373, new_n7374, new_n7375, new_n7376,
    new_n7377, new_n7378, new_n7379, new_n7380, new_n7381, new_n7382,
    new_n7383, new_n7384, new_n7385, new_n7386, new_n7387, new_n7388,
    new_n7389, new_n7390, new_n7391, new_n7392, new_n7393, new_n7394,
    new_n7395, new_n7396, new_n7397, new_n7398, new_n7399, new_n7400,
    new_n7401, new_n7402, new_n7403, new_n7404, new_n7405, new_n7406,
    new_n7407, new_n7408, new_n7409, new_n7410, new_n7411, new_n7412,
    new_n7413, new_n7414, new_n7415, new_n7416, new_n7417, new_n7418,
    new_n7419, new_n7420, new_n7421, new_n7422, new_n7423, new_n7424,
    new_n7425, new_n7426, new_n7427, new_n7428, new_n7429, new_n7430,
    new_n7431, new_n7432, new_n7433, new_n7434, new_n7435, new_n7436,
    new_n7437, new_n7438, new_n7439, new_n7440, new_n7441, new_n7442,
    new_n7443, new_n7444, new_n7445, new_n7446, new_n7447, new_n7448,
    new_n7449, new_n7450, new_n7451, new_n7452, new_n7453, new_n7454,
    new_n7455, new_n7456, new_n7457, new_n7458, new_n7459, new_n7460,
    new_n7461, new_n7462, new_n7463, new_n7464, new_n7465, new_n7466,
    new_n7467, new_n7468, new_n7469, new_n7470, new_n7471, new_n7472,
    new_n7473, new_n7474, new_n7475, new_n7476, new_n7477, new_n7478,
    new_n7479, new_n7480, new_n7481, new_n7482, new_n7483, new_n7484,
    new_n7485, new_n7486, new_n7487, new_n7488, new_n7489, new_n7490,
    new_n7491, new_n7492, new_n7493, new_n7494, new_n7495, new_n7496,
    new_n7497, new_n7498, new_n7499, new_n7500, new_n7501, new_n7502,
    new_n7503, new_n7504, new_n7505, new_n7506, new_n7507, new_n7508,
    new_n7509, new_n7510, new_n7511, new_n7512, new_n7513, new_n7514,
    new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592,
    new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598,
    new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604,
    new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610,
    new_n7611, new_n7613, new_n7614, new_n7615, new_n7616, new_n7617,
    new_n7618, new_n7619, new_n7620, new_n7621, new_n7622, new_n7623,
    new_n7624, new_n7625, new_n7626, new_n7627, new_n7628, new_n7629,
    new_n7630, new_n7631, new_n7632, new_n7633, new_n7634, new_n7635,
    new_n7636, new_n7637, new_n7638, new_n7639, new_n7640, new_n7641,
    new_n7642, new_n7643, new_n7644, new_n7645, new_n7646, new_n7647,
    new_n7648, new_n7649, new_n7650, new_n7651, new_n7652, new_n7653,
    new_n7654, new_n7655, new_n7656, new_n7657, new_n7658, new_n7659,
    new_n7660, new_n7661, new_n7662, new_n7663, new_n7664, new_n7665,
    new_n7666, new_n7667, new_n7668, new_n7669, new_n7670, new_n7671,
    new_n7672, new_n7673, new_n7674, new_n7675, new_n7676, new_n7677,
    new_n7678, new_n7679, new_n7680, new_n7681, new_n7682, new_n7683,
    new_n7684, new_n7685, new_n7686, new_n7687, new_n7688, new_n7689,
    new_n7690, new_n7691, new_n7692, new_n7693, new_n7694, new_n7695,
    new_n7696, new_n7697, new_n7698, new_n7699, new_n7700, new_n7701,
    new_n7702, new_n7703, new_n7704, new_n7705, new_n7706, new_n7707,
    new_n7708, new_n7709, new_n7710, new_n7711, new_n7712, new_n7713,
    new_n7714, new_n7715, new_n7716, new_n7717, new_n7718, new_n7719,
    new_n7720, new_n7721, new_n7722, new_n7723, new_n7724, new_n7725,
    new_n7726, new_n7727, new_n7728, new_n7729, new_n7730, new_n7731,
    new_n7732, new_n7733, new_n7734, new_n7735, new_n7736, new_n7737,
    new_n7738, new_n7739, new_n7740, new_n7741, new_n7742, new_n7743,
    new_n7744, new_n7745, new_n7746, new_n7747, new_n7748, new_n7749,
    new_n7750, new_n7751, new_n7752, new_n7753, new_n7754, new_n7755,
    new_n7756, new_n7757, new_n7758, new_n7759, new_n7760, new_n7761,
    new_n7762, new_n7763, new_n7764, new_n7765, new_n7766, new_n7767,
    new_n7768, new_n7769, new_n7770, new_n7771, new_n7772, new_n7773,
    new_n7774, new_n7775, new_n7776, new_n7777, new_n7778, new_n7779,
    new_n7780, new_n7781, new_n7782, new_n7783, new_n7784, new_n7785,
    new_n7786, new_n7787, new_n7788, new_n7789, new_n7790, new_n7791,
    new_n7792, new_n7793, new_n7794, new_n7795, new_n7796, new_n7797,
    new_n7798, new_n7799, new_n7800, new_n7801, new_n7802, new_n7803,
    new_n7804, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809,
    new_n7810, new_n7811, new_n7812, new_n7813, new_n7814, new_n7815,
    new_n7816, new_n7817, new_n7818, new_n7819, new_n7820, new_n7821,
    new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827,
    new_n7828, new_n7829, new_n7830, new_n7831, new_n7832, new_n7833,
    new_n7834, new_n7835, new_n7836, new_n7837, new_n7838, new_n7839,
    new_n7840, new_n7841, new_n7842, new_n7843, new_n7844, new_n7845,
    new_n7846, new_n7847, new_n7848, new_n7849, new_n7850, new_n7851,
    new_n7852, new_n7853, new_n7854, new_n7855, new_n7856, new_n7857,
    new_n7858, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863,
    new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869,
    new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875,
    new_n7876, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881,
    new_n7882, new_n7883, new_n7884, new_n7885, new_n7886, new_n7887,
    new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893,
    new_n7894, new_n7895, new_n7897, new_n7898, new_n7899, new_n7900,
    new_n7901, new_n7902, new_n7903, new_n7904, new_n7905, new_n7906,
    new_n7907, new_n7908, new_n7909, new_n7910, new_n7911, new_n7912,
    new_n7913, new_n7914, new_n7915, new_n7916, new_n7917, new_n7918,
    new_n7919, new_n7920, new_n7921, new_n7922, new_n7923, new_n7924,
    new_n7925, new_n7926, new_n7927, new_n7928, new_n7929, new_n7930,
    new_n7931, new_n7932, new_n7933, new_n7934, new_n7935, new_n7936,
    new_n7937, new_n7938, new_n7939, new_n7940, new_n7941, new_n7942,
    new_n7943, new_n7944, new_n7945, new_n7946, new_n7947, new_n7948,
    new_n7949, new_n7950, new_n7951, new_n7952, new_n7953, new_n7954,
    new_n7955, new_n7956, new_n7957, new_n7958, new_n7959, new_n7960,
    new_n7961, new_n7962, new_n7963, new_n7964, new_n7965, new_n7966,
    new_n7967, new_n7968, new_n7969, new_n7970, new_n7971, new_n7972,
    new_n7973, new_n7974, new_n7975, new_n7976, new_n7977, new_n7978,
    new_n7979, new_n7980, new_n7981, new_n7982, new_n7983, new_n7984,
    new_n7985, new_n7986, new_n7987, new_n7988, new_n7989, new_n7990,
    new_n7991, new_n7992, new_n7993, new_n7994, new_n7995, new_n7996,
    new_n7997, new_n7998, new_n7999, new_n8000, new_n8001, new_n8002,
    new_n8003, new_n8004, new_n8005, new_n8006, new_n8007, new_n8008,
    new_n8009, new_n8010, new_n8011, new_n8012, new_n8013, new_n8014,
    new_n8015, new_n8016, new_n8017, new_n8018, new_n8019, new_n8020,
    new_n8021, new_n8022, new_n8023, new_n8024, new_n8025, new_n8026,
    new_n8027, new_n8028, new_n8029, new_n8030, new_n8031, new_n8032,
    new_n8033, new_n8034, new_n8035, new_n8036, new_n8037, new_n8038,
    new_n8039, new_n8040, new_n8041, new_n8042, new_n8043, new_n8044,
    new_n8045, new_n8046, new_n8047, new_n8048, new_n8049, new_n8050,
    new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056,
    new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062,
    new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068,
    new_n8069, new_n8070, new_n8071, new_n8072, new_n8073, new_n8074,
    new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080,
    new_n8081, new_n8082, new_n8083, new_n8084, new_n8085, new_n8086,
    new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092,
    new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098,
    new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104,
    new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110,
    new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140,
    new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146,
    new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152,
    new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158,
    new_n8159, new_n8160, new_n8161, new_n8162, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285,
    new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303,
    new_n8304, new_n8305, new_n8306, new_n8307, new_n8308, new_n8309,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8460,
    new_n8461, new_n8462, new_n8463, new_n8464, new_n8465, new_n8466,
    new_n8467, new_n8468, new_n8469, new_n8470, new_n8471, new_n8472,
    new_n8473, new_n8474, new_n8475, new_n8476, new_n8477, new_n8478,
    new_n8479, new_n8480, new_n8481, new_n8482, new_n8483, new_n8484,
    new_n8485, new_n8486, new_n8487, new_n8488, new_n8489, new_n8490,
    new_n8491, new_n8492, new_n8493, new_n8494, new_n8495, new_n8496,
    new_n8497, new_n8498, new_n8499, new_n8500, new_n8501, new_n8502,
    new_n8503, new_n8504, new_n8505, new_n8506, new_n8507, new_n8508,
    new_n8509, new_n8510, new_n8511, new_n8512, new_n8513, new_n8514,
    new_n8515, new_n8516, new_n8517, new_n8518, new_n8519, new_n8520,
    new_n8521, new_n8522, new_n8523, new_n8524, new_n8525, new_n8526,
    new_n8527, new_n8528, new_n8529, new_n8530, new_n8531, new_n8532,
    new_n8533, new_n8534, new_n8535, new_n8536, new_n8537, new_n8538,
    new_n8539, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544,
    new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550,
    new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556,
    new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562,
    new_n8563, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568,
    new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574,
    new_n8575, new_n8576, new_n8577, new_n8578, new_n8579, new_n8580,
    new_n8581, new_n8582, new_n8583, new_n8584, new_n8585, new_n8586,
    new_n8587, new_n8588, new_n8589, new_n8590, new_n8591, new_n8592,
    new_n8593, new_n8594, new_n8595, new_n8596, new_n8597, new_n8598,
    new_n8599, new_n8600, new_n8601, new_n8602, new_n8603, new_n8604,
    new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610,
    new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616,
    new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622,
    new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628,
    new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634,
    new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8760, new_n8761,
    new_n8762, new_n8763, new_n8764, new_n8765, new_n8766, new_n8767,
    new_n8768, new_n8769, new_n8770, new_n8771, new_n8772, new_n8773,
    new_n8774, new_n8775, new_n8776, new_n8777, new_n8778, new_n8779,
    new_n8780, new_n8781, new_n8782, new_n8783, new_n8784, new_n8785,
    new_n8786, new_n8787, new_n8788, new_n8789, new_n8790, new_n8791,
    new_n8792, new_n8793, new_n8794, new_n8795, new_n8796, new_n8797,
    new_n8798, new_n8799, new_n8800, new_n8801, new_n8802, new_n8803,
    new_n8804, new_n8805, new_n8806, new_n8807, new_n8808, new_n8809,
    new_n8810, new_n8811, new_n8812, new_n8813, new_n8814, new_n8815,
    new_n8816, new_n8817, new_n8818, new_n8819, new_n8820, new_n8821,
    new_n8822, new_n8823, new_n8824, new_n8825, new_n8826, new_n8827,
    new_n8828, new_n8829, new_n8830, new_n8831, new_n8832, new_n8833,
    new_n8834, new_n8835, new_n8836, new_n8837, new_n8838, new_n8839,
    new_n8840, new_n8841, new_n8842, new_n8843, new_n8844, new_n8845,
    new_n8846, new_n8847, new_n8848, new_n8849, new_n8850, new_n8851,
    new_n8852, new_n8853, new_n8854, new_n8855, new_n8856, new_n8857,
    new_n8858, new_n8859, new_n8860, new_n8861, new_n8862, new_n8863,
    new_n8864, new_n8865, new_n8866, new_n8867, new_n8868, new_n8869,
    new_n8870, new_n8871, new_n8872, new_n8873, new_n8874, new_n8875,
    new_n8876, new_n8877, new_n8878, new_n8879, new_n8880, new_n8881,
    new_n8882, new_n8883, new_n8884, new_n8885, new_n8886, new_n8887,
    new_n8888, new_n8889, new_n8890, new_n8891, new_n8892, new_n8893,
    new_n8894, new_n8895, new_n8896, new_n8897, new_n8898, new_n8899,
    new_n8900, new_n8901, new_n8902, new_n8903, new_n8904, new_n8905,
    new_n8906, new_n8907, new_n8908, new_n8909, new_n8910, new_n8911,
    new_n8912, new_n8913, new_n8914, new_n8915, new_n8916, new_n8917,
    new_n8918, new_n8919, new_n8920, new_n8921, new_n8922, new_n8923,
    new_n8924, new_n8925, new_n8926, new_n8927, new_n8928, new_n8929,
    new_n8930, new_n8931, new_n8932, new_n8933, new_n8934, new_n8935,
    new_n8936, new_n8937, new_n8938, new_n8939, new_n8940, new_n8941,
    new_n8942, new_n8943, new_n8944, new_n8945, new_n8946, new_n8947,
    new_n8948, new_n8949, new_n8950, new_n8951, new_n8952, new_n8953,
    new_n8954, new_n8955, new_n8956, new_n8957, new_n8958, new_n8959,
    new_n8960, new_n8961, new_n8962, new_n8963, new_n8964, new_n8965,
    new_n8966, new_n8967, new_n8968, new_n8969, new_n8970, new_n8971,
    new_n8972, new_n8973, new_n8974, new_n8975, new_n8976, new_n8977,
    new_n8978, new_n8979, new_n8980, new_n8981, new_n8982, new_n8983,
    new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989,
    new_n8990, new_n8991, new_n8992, new_n8993, new_n8994, new_n8995,
    new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9001,
    new_n9002, new_n9003, new_n9004, new_n9005, new_n9006, new_n9007,
    new_n9008, new_n9009, new_n9010, new_n9011, new_n9012, new_n9013,
    new_n9014, new_n9015, new_n9016, new_n9017, new_n9018, new_n9019,
    new_n9020, new_n9021, new_n9022, new_n9023, new_n9024, new_n9025,
    new_n9026, new_n9027, new_n9028, new_n9029, new_n9030, new_n9031,
    new_n9032, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037,
    new_n9038, new_n9039, new_n9040, new_n9041, new_n9042, new_n9043,
    new_n9044, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9339,
    new_n9340, new_n9341, new_n9342, new_n9343, new_n9344, new_n9345,
    new_n9346, new_n9347, new_n9348, new_n9349, new_n9350, new_n9351,
    new_n9352, new_n9353, new_n9354, new_n9355, new_n9356, new_n9357,
    new_n9358, new_n9359, new_n9360, new_n9361, new_n9362, new_n9363,
    new_n9364, new_n9365, new_n9366, new_n9367, new_n9368, new_n9369,
    new_n9370, new_n9371, new_n9372, new_n9373, new_n9374, new_n9375,
    new_n9376, new_n9377, new_n9378, new_n9379, new_n9380, new_n9381,
    new_n9382, new_n9383, new_n9384, new_n9385, new_n9386, new_n9387,
    new_n9388, new_n9389, new_n9390, new_n9391, new_n9392, new_n9393,
    new_n9394, new_n9395, new_n9396, new_n9397, new_n9398, new_n9399,
    new_n9400, new_n9401, new_n9402, new_n9403, new_n9404, new_n9405,
    new_n9406, new_n9407, new_n9408, new_n9409, new_n9410, new_n9411,
    new_n9412, new_n9413, new_n9414, new_n9415, new_n9416, new_n9417,
    new_n9418, new_n9419, new_n9420, new_n9421, new_n9422, new_n9423,
    new_n9424, new_n9425, new_n9426, new_n9427, new_n9428, new_n9429,
    new_n9430, new_n9431, new_n9432, new_n9433, new_n9434, new_n9435,
    new_n9436, new_n9437, new_n9438, new_n9439, new_n9440, new_n9441,
    new_n9442, new_n9443, new_n9444, new_n9445, new_n9446, new_n9447,
    new_n9448, new_n9449, new_n9450, new_n9451, new_n9452, new_n9453,
    new_n9454, new_n9455, new_n9456, new_n9457, new_n9458, new_n9459,
    new_n9460, new_n9461, new_n9462, new_n9463, new_n9464, new_n9465,
    new_n9466, new_n9467, new_n9468, new_n9469, new_n9470, new_n9471,
    new_n9472, new_n9473, new_n9474, new_n9475, new_n9476, new_n9477,
    new_n9478, new_n9479, new_n9480, new_n9481, new_n9482, new_n9483,
    new_n9484, new_n9485, new_n9486, new_n9487, new_n9488, new_n9489,
    new_n9490, new_n9491, new_n9492, new_n9493, new_n9494, new_n9495,
    new_n9496, new_n9497, new_n9498, new_n9499, new_n9500, new_n9501,
    new_n9502, new_n9503, new_n9504, new_n9505, new_n9506, new_n9507,
    new_n9508, new_n9509, new_n9510, new_n9511, new_n9512, new_n9513,
    new_n9514, new_n9515, new_n9516, new_n9517, new_n9518, new_n9519,
    new_n9520, new_n9521, new_n9522, new_n9523, new_n9524, new_n9525,
    new_n9526, new_n9527, new_n9528, new_n9529, new_n9530, new_n9531,
    new_n9532, new_n9533, new_n9534, new_n9535, new_n9536, new_n9537,
    new_n9538, new_n9539, new_n9540, new_n9541, new_n9542, new_n9543,
    new_n9544, new_n9545, new_n9546, new_n9547, new_n9548, new_n9549,
    new_n9550, new_n9551, new_n9552, new_n9553, new_n9554, new_n9555,
    new_n9556, new_n9557, new_n9558, new_n9559, new_n9560, new_n9561,
    new_n9562, new_n9563, new_n9564, new_n9565, new_n9566, new_n9567,
    new_n9568, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622, new_n9623, new_n9624, new_n9625, new_n9626, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633,
    new_n9634, new_n9635, new_n9637, new_n9638, new_n9639, new_n9640,
    new_n9641, new_n9642, new_n9643, new_n9644, new_n9645, new_n9646,
    new_n9647, new_n9648, new_n9649, new_n9650, new_n9651, new_n9652,
    new_n9653, new_n9654, new_n9655, new_n9656, new_n9657, new_n9658,
    new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664,
    new_n9665, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670,
    new_n9671, new_n9672, new_n9673, new_n9674, new_n9675, new_n9676,
    new_n9677, new_n9678, new_n9679, new_n9680, new_n9681, new_n9682,
    new_n9683, new_n9684, new_n9685, new_n9686, new_n9687, new_n9688,
    new_n9689, new_n9690, new_n9691, new_n9692, new_n9693, new_n9694,
    new_n9695, new_n9696, new_n9697, new_n9698, new_n9699, new_n9700,
    new_n9701, new_n9702, new_n9703, new_n9704, new_n9705, new_n9706,
    new_n9707, new_n9708, new_n9709, new_n9710, new_n9711, new_n9712,
    new_n9713, new_n9714, new_n9715, new_n9716, new_n9717, new_n9718,
    new_n9719, new_n9720, new_n9721, new_n9722, new_n9723, new_n9724,
    new_n9725, new_n9726, new_n9727, new_n9728, new_n9729, new_n9730,
    new_n9731, new_n9732, new_n9733, new_n9734, new_n9735, new_n9736,
    new_n9737, new_n9738, new_n9739, new_n9740, new_n9741, new_n9742,
    new_n9743, new_n9744, new_n9745, new_n9746, new_n9747, new_n9748,
    new_n9749, new_n9750, new_n9751, new_n9752, new_n9753, new_n9754,
    new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760,
    new_n9761, new_n9762, new_n9763, new_n9764, new_n9765, new_n9766,
    new_n9767, new_n9768, new_n9769, new_n9770, new_n9771, new_n9772,
    new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778,
    new_n9779, new_n9780, new_n9781, new_n9782, new_n9783, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832,
    new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838,
    new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9867, new_n9868,
    new_n9869, new_n9870, new_n9871, new_n9872, new_n9873, new_n9874,
    new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880,
    new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886,
    new_n9887, new_n9888, new_n9889, new_n9890, new_n9891, new_n9892,
    new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898,
    new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904,
    new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910,
    new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916,
    new_n9917, new_n9918, new_n9919, new_n9920, new_n9921, new_n9922,
    new_n9923, new_n9924, new_n9925, new_n9926, new_n9927, new_n9928,
    new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934,
    new_n9935, new_n9936, new_n9937, new_n9938, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022, new_n10023, new_n10024, new_n10025,
    new_n10026, new_n10027, new_n10028, new_n10029, new_n10030, new_n10031,
    new_n10032, new_n10033, new_n10034, new_n10035, new_n10036, new_n10037,
    new_n10038, new_n10039, new_n10040, new_n10041, new_n10042, new_n10043,
    new_n10044, new_n10045, new_n10046, new_n10047, new_n10048, new_n10049,
    new_n10050, new_n10051, new_n10052, new_n10053, new_n10054, new_n10055,
    new_n10056, new_n10057, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127,
    new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133,
    new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139,
    new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145,
    new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151,
    new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163,
    new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236, new_n10237, new_n10238, new_n10239, new_n10240, new_n10241,
    new_n10242, new_n10243, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10572, new_n10573,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589, new_n10590, new_n10591,
    new_n10592, new_n10593, new_n10594, new_n10595, new_n10596, new_n10597,
    new_n10598, new_n10599, new_n10600, new_n10601, new_n10602, new_n10603,
    new_n10604, new_n10605, new_n10606, new_n10607, new_n10608, new_n10609,
    new_n10610, new_n10611, new_n10612, new_n10613, new_n10614, new_n10615,
    new_n10616, new_n10617, new_n10618, new_n10619, new_n10620, new_n10621,
    new_n10622, new_n10623, new_n10624, new_n10625, new_n10626, new_n10627,
    new_n10628, new_n10629, new_n10630, new_n10631, new_n10632, new_n10633,
    new_n10634, new_n10635, new_n10636, new_n10637, new_n10638, new_n10639,
    new_n10640, new_n10641, new_n10642, new_n10643, new_n10644, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693,
    new_n10694, new_n10695, new_n10696, new_n10697, new_n10698, new_n10699,
    new_n10700, new_n10701, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710, new_n10711,
    new_n10712, new_n10713, new_n10714, new_n10715, new_n10716, new_n10717,
    new_n10718, new_n10719, new_n10720, new_n10721, new_n10722, new_n10723,
    new_n10724, new_n10725, new_n10726, new_n10727, new_n10728, new_n10729,
    new_n10730, new_n10731, new_n10732, new_n10733, new_n10734, new_n10735,
    new_n10736, new_n10737, new_n10738, new_n10739, new_n10740, new_n10741,
    new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747,
    new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775, new_n10776, new_n10777,
    new_n10778, new_n10779, new_n10780, new_n10781, new_n10782, new_n10783,
    new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789,
    new_n10790, new_n10791, new_n10792, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817, new_n10818, new_n10819,
    new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825,
    new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831,
    new_n10832, new_n10833, new_n10834, new_n10835, new_n10836, new_n10837,
    new_n10838, new_n10839, new_n10840, new_n10841, new_n10842, new_n10843,
    new_n10844, new_n10845, new_n10846, new_n10847, new_n10848, new_n10849,
    new_n10850, new_n10851, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10875, new_n10876, new_n10877, new_n10878, new_n10879, new_n10880,
    new_n10881, new_n10882, new_n10883, new_n10884, new_n10885, new_n10886,
    new_n10887, new_n10888, new_n10889, new_n10890, new_n10891, new_n10892,
    new_n10893, new_n10894, new_n10895, new_n10896, new_n10897, new_n10898,
    new_n10899, new_n10900, new_n10901, new_n10902, new_n10903, new_n10904,
    new_n10905, new_n10906, new_n10907, new_n10908, new_n10909, new_n10910,
    new_n10911, new_n10912, new_n10913, new_n10914, new_n10915, new_n10916,
    new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922,
    new_n10923, new_n10924, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943, new_n10944, new_n10945, new_n10946,
    new_n10947, new_n10948, new_n10949, new_n10950, new_n10951, new_n10952,
    new_n10953, new_n10954, new_n10955, new_n10956, new_n10957, new_n10958,
    new_n10959, new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965, new_n10966, new_n10967, new_n10968, new_n10969, new_n10970,
    new_n10971, new_n10972, new_n10973, new_n10974, new_n10975, new_n10976,
    new_n10977, new_n10978, new_n10979, new_n10980, new_n10981, new_n10982,
    new_n10983, new_n10984, new_n10985, new_n10986, new_n10987, new_n10988,
    new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024,
    new_n11025, new_n11026, new_n11027, new_n11028, new_n11029, new_n11030,
    new_n11031, new_n11032, new_n11033, new_n11034, new_n11035, new_n11036,
    new_n11037, new_n11038, new_n11039, new_n11040, new_n11041, new_n11042,
    new_n11043, new_n11044, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056, new_n11057, new_n11058, new_n11059, new_n11060,
    new_n11061, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066,
    new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072,
    new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078,
    new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084,
    new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186,
    new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211,
    new_n11212, new_n11213, new_n11214, new_n11215, new_n11216, new_n11217,
    new_n11218, new_n11219, new_n11220, new_n11221, new_n11222, new_n11223,
    new_n11224, new_n11225, new_n11226, new_n11227, new_n11228, new_n11229,
    new_n11230, new_n11231, new_n11232, new_n11233, new_n11234, new_n11235,
    new_n11236, new_n11237, new_n11238, new_n11239, new_n11240, new_n11241,
    new_n11242, new_n11243, new_n11244, new_n11245, new_n11246, new_n11247,
    new_n11248, new_n11249, new_n11250, new_n11251, new_n11252, new_n11253,
    new_n11254, new_n11255, new_n11256, new_n11257, new_n11258, new_n11259,
    new_n11260, new_n11261, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266, new_n11267, new_n11268, new_n11269, new_n11270, new_n11271,
    new_n11272, new_n11273, new_n11274, new_n11275, new_n11276, new_n11277,
    new_n11278, new_n11279, new_n11280, new_n11281, new_n11282, new_n11283,
    new_n11284, new_n11285, new_n11286, new_n11287, new_n11288, new_n11289,
    new_n11290, new_n11291, new_n11292, new_n11293, new_n11294, new_n11295,
    new_n11296, new_n11297, new_n11298, new_n11299, new_n11300, new_n11301,
    new_n11302, new_n11303, new_n11304, new_n11305, new_n11306, new_n11307,
    new_n11308, new_n11309, new_n11310, new_n11311, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326, new_n11327, new_n11328, new_n11329, new_n11330, new_n11331,
    new_n11332, new_n11333, new_n11334, new_n11335, new_n11336, new_n11337,
    new_n11338, new_n11339, new_n11340, new_n11341, new_n11342, new_n11343,
    new_n11344, new_n11345, new_n11346, new_n11347, new_n11348, new_n11349,
    new_n11350, new_n11351, new_n11352, new_n11353, new_n11354, new_n11355,
    new_n11356, new_n11357, new_n11358, new_n11359, new_n11360, new_n11361,
    new_n11362, new_n11363, new_n11364, new_n11365, new_n11366, new_n11367,
    new_n11368, new_n11369, new_n11370, new_n11371, new_n11372, new_n11373,
    new_n11374, new_n11375, new_n11376, new_n11377, new_n11378, new_n11379,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386, new_n11387, new_n11388, new_n11389, new_n11390, new_n11391,
    new_n11392, new_n11393, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398, new_n11399, new_n11400, new_n11401, new_n11402, new_n11403,
    new_n11404, new_n11405, new_n11406, new_n11407, new_n11408, new_n11409,
    new_n11410, new_n11411, new_n11412, new_n11413, new_n11414, new_n11415,
    new_n11416, new_n11417, new_n11418, new_n11419, new_n11420, new_n11421,
    new_n11422, new_n11423, new_n11424, new_n11425, new_n11426, new_n11427,
    new_n11428, new_n11429, new_n11430, new_n11431, new_n11432, new_n11433,
    new_n11434, new_n11435, new_n11436, new_n11437, new_n11438, new_n11439,
    new_n11440, new_n11441, new_n11442, new_n11443, new_n11444, new_n11445,
    new_n11446, new_n11447, new_n11448, new_n11449, new_n11450, new_n11451,
    new_n11452, new_n11453, new_n11454, new_n11455, new_n11456, new_n11457,
    new_n11458, new_n11459, new_n11460, new_n11461, new_n11462, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470, new_n11471, new_n11472, new_n11473, new_n11474, new_n11475,
    new_n11476, new_n11477, new_n11478, new_n11479, new_n11480, new_n11481,
    new_n11482, new_n11483, new_n11484, new_n11485, new_n11486, new_n11487,
    new_n11488, new_n11489, new_n11490, new_n11491, new_n11492, new_n11493,
    new_n11494, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535, new_n11536,
    new_n11537, new_n11538, new_n11539, new_n11540, new_n11541, new_n11542,
    new_n11543, new_n11544, new_n11545, new_n11546, new_n11547, new_n11548,
    new_n11549, new_n11550, new_n11551, new_n11552, new_n11553, new_n11554,
    new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560,
    new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608,
    new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620,
    new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632,
    new_n11633, new_n11634, new_n11635, new_n11636, new_n11637, new_n11638,
    new_n11639, new_n11640, new_n11641, new_n11642, new_n11643, new_n11644,
    new_n11645, new_n11646, new_n11647, new_n11648, new_n11649, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662,
    new_n11663, new_n11664, new_n11665, new_n11666, new_n11667, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673, new_n11674,
    new_n11675, new_n11676, new_n11677, new_n11678, new_n11679, new_n11680,
    new_n11681, new_n11682, new_n11683, new_n11684, new_n11685, new_n11686,
    new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692,
    new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698,
    new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704,
    new_n11705, new_n11706, new_n11707, new_n11708, new_n11709, new_n11710,
    new_n11711, new_n11712, new_n11713, new_n11714, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755, new_n11756, new_n11757, new_n11758,
    new_n11759, new_n11760, new_n11761, new_n11762, new_n11763, new_n11764,
    new_n11765, new_n11766, new_n11767, new_n11768, new_n11769, new_n11770,
    new_n11771, new_n11772, new_n11773, new_n11774, new_n11775, new_n11776,
    new_n11777, new_n11778, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11790, new_n11791, new_n11792, new_n11793, new_n11794, new_n11795,
    new_n11796, new_n11797, new_n11798, new_n11799, new_n11800, new_n11801,
    new_n11802, new_n11803, new_n11804, new_n11805, new_n11806, new_n11807,
    new_n11808, new_n11809, new_n11810, new_n11811, new_n11812, new_n11813,
    new_n11814, new_n11815, new_n11816, new_n11817, new_n11818, new_n11819,
    new_n11820, new_n11821, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861,
    new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876, new_n11877, new_n11878, new_n11879,
    new_n11880, new_n11881, new_n11882, new_n11883, new_n11884, new_n11885,
    new_n11886, new_n11887, new_n11888, new_n11889, new_n11890, new_n11891,
    new_n11892, new_n11893, new_n11894, new_n11895, new_n11896, new_n11897,
    new_n11898, new_n11899, new_n11900, new_n11901, new_n11902, new_n11903,
    new_n11904, new_n11905, new_n11906, new_n11907, new_n11908, new_n11909,
    new_n11910, new_n11911, new_n11912, new_n11913, new_n11914, new_n11915,
    new_n11916, new_n11917, new_n11918, new_n11919, new_n11920, new_n11921,
    new_n11922, new_n11923, new_n11924, new_n11925, new_n11926, new_n11927,
    new_n11928, new_n11929, new_n11930, new_n11931, new_n11932, new_n11933,
    new_n11934, new_n11935, new_n11936, new_n11937, new_n11938, new_n11939,
    new_n11940, new_n11941, new_n11942, new_n11943, new_n11944, new_n11945,
    new_n11946, new_n11947, new_n11948, new_n11949, new_n11950, new_n11951,
    new_n11952, new_n11953, new_n11954, new_n11955, new_n11956, new_n11957,
    new_n11958, new_n11959, new_n11960, new_n11961, new_n11962, new_n11963,
    new_n11964, new_n11965, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980, new_n11981,
    new_n11982, new_n11983, new_n11984, new_n11985, new_n11986, new_n11987,
    new_n11988, new_n11989, new_n11990, new_n11991, new_n11992, new_n11993,
    new_n11994, new_n11995, new_n11996, new_n11997, new_n11998, new_n11999,
    new_n12000, new_n12001, new_n12002, new_n12003, new_n12004, new_n12005,
    new_n12006, new_n12007, new_n12008, new_n12009, new_n12010, new_n12011,
    new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017,
    new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047,
    new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053,
    new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059,
    new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065,
    new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072, new_n12073, new_n12074, new_n12075, new_n12076, new_n12077,
    new_n12078, new_n12079, new_n12080, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111, new_n12112, new_n12113, new_n12114,
    new_n12115, new_n12116, new_n12117, new_n12118, new_n12119, new_n12120,
    new_n12121, new_n12122, new_n12123, new_n12124, new_n12125, new_n12126,
    new_n12127, new_n12128, new_n12129, new_n12130, new_n12131, new_n12132,
    new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138,
    new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145, new_n12146, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152, new_n12153, new_n12154, new_n12155, new_n12156,
    new_n12157, new_n12158, new_n12159, new_n12160, new_n12161, new_n12162,
    new_n12163, new_n12164, new_n12165, new_n12166, new_n12167, new_n12168,
    new_n12169, new_n12170, new_n12171, new_n12172, new_n12173, new_n12174,
    new_n12175, new_n12176, new_n12177, new_n12178, new_n12179, new_n12180,
    new_n12181, new_n12182, new_n12183, new_n12184, new_n12185, new_n12186,
    new_n12187, new_n12188, new_n12189, new_n12190, new_n12191, new_n12192,
    new_n12193, new_n12194, new_n12195, new_n12196, new_n12197, new_n12198,
    new_n12199, new_n12200, new_n12201, new_n12202, new_n12203, new_n12204,
    new_n12205, new_n12206, new_n12207, new_n12208, new_n12209, new_n12210,
    new_n12211, new_n12212, new_n12213, new_n12214, new_n12215, new_n12216,
    new_n12217, new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223, new_n12224, new_n12225, new_n12226, new_n12227, new_n12228,
    new_n12229, new_n12230, new_n12231, new_n12232, new_n12233, new_n12234,
    new_n12235, new_n12236, new_n12237, new_n12238, new_n12239, new_n12240,
    new_n12241, new_n12242, new_n12243, new_n12244, new_n12245, new_n12246,
    new_n12247, new_n12248, new_n12249, new_n12250, new_n12251, new_n12252,
    new_n12253, new_n12254, new_n12255, new_n12256, new_n12257, new_n12258,
    new_n12259, new_n12260, new_n12261, new_n12262, new_n12263, new_n12264,
    new_n12265, new_n12266, new_n12267, new_n12268, new_n12269, new_n12270,
    new_n12271, new_n12272, new_n12273, new_n12274, new_n12275, new_n12276,
    new_n12277, new_n12278, new_n12279, new_n12280, new_n12281, new_n12282,
    new_n12283, new_n12284, new_n12285, new_n12286, new_n12287, new_n12288,
    new_n12289, new_n12290, new_n12291, new_n12292, new_n12293, new_n12294,
    new_n12295, new_n12296, new_n12297, new_n12298, new_n12299, new_n12300,
    new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324, new_n12325,
    new_n12326, new_n12327, new_n12328, new_n12329, new_n12330, new_n12331,
    new_n12332, new_n12333, new_n12334, new_n12335, new_n12336, new_n12337,
    new_n12338, new_n12339, new_n12340, new_n12341, new_n12342, new_n12343,
    new_n12344, new_n12345, new_n12346, new_n12347, new_n12348, new_n12349,
    new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355,
    new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361,
    new_n12362, new_n12363, new_n12364, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380, new_n12381, new_n12382, new_n12383, new_n12384, new_n12385,
    new_n12386, new_n12387, new_n12388, new_n12389, new_n12390, new_n12391,
    new_n12392, new_n12393, new_n12394, new_n12395, new_n12396, new_n12397,
    new_n12398, new_n12399, new_n12400, new_n12401, new_n12402, new_n12403,
    new_n12404, new_n12405, new_n12406, new_n12407, new_n12408, new_n12409,
    new_n12410, new_n12411, new_n12412, new_n12413, new_n12414, new_n12415,
    new_n12416, new_n12417, new_n12418, new_n12419, new_n12420, new_n12421,
    new_n12422, new_n12423, new_n12424, new_n12425, new_n12426, new_n12427,
    new_n12428, new_n12429, new_n12430, new_n12431, new_n12432, new_n12433,
    new_n12434, new_n12435, new_n12436, new_n12437, new_n12438, new_n12439,
    new_n12440, new_n12441, new_n12442, new_n12443, new_n12444, new_n12445,
    new_n12446, new_n12447, new_n12448, new_n12449, new_n12450, new_n12451,
    new_n12452, new_n12453, new_n12454, new_n12455, new_n12456, new_n12457,
    new_n12458, new_n12459, new_n12460, new_n12461, new_n12462, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467, new_n12468, new_n12469,
    new_n12470, new_n12471, new_n12472, new_n12473, new_n12474, new_n12475,
    new_n12476, new_n12477, new_n12478, new_n12479, new_n12480, new_n12481,
    new_n12482, new_n12483, new_n12484, new_n12485, new_n12486, new_n12487,
    new_n12488, new_n12489, new_n12490, new_n12491, new_n12492, new_n12493,
    new_n12494, new_n12495, new_n12496, new_n12497, new_n12498, new_n12499,
    new_n12500, new_n12501, new_n12502, new_n12503, new_n12504, new_n12505,
    new_n12506, new_n12507, new_n12508, new_n12509, new_n12510, new_n12511,
    new_n12512, new_n12513, new_n12514, new_n12515, new_n12516, new_n12517,
    new_n12518, new_n12519, new_n12520, new_n12521, new_n12522, new_n12523,
    new_n12524, new_n12525, new_n12526, new_n12527, new_n12528, new_n12529,
    new_n12530, new_n12531, new_n12532, new_n12533, new_n12534, new_n12535,
    new_n12536, new_n12537, new_n12538, new_n12539, new_n12540, new_n12541,
    new_n12542, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566,
    new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572,
    new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578,
    new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584,
    new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590,
    new_n12591, new_n12592, new_n12593, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607, new_n12608,
    new_n12609, new_n12610, new_n12611, new_n12612, new_n12613, new_n12614,
    new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702, new_n12703, new_n12704,
    new_n12705, new_n12706, new_n12707, new_n12708, new_n12709, new_n12710,
    new_n12711, new_n12712, new_n12713, new_n12714, new_n12715, new_n12716,
    new_n12717, new_n12718, new_n12719, new_n12720, new_n12721, new_n12722,
    new_n12723, new_n12724, new_n12725, new_n12726, new_n12727, new_n12728,
    new_n12729, new_n12730, new_n12731, new_n12732, new_n12733, new_n12734,
    new_n12735, new_n12736, new_n12737, new_n12738, new_n12739, new_n12740,
    new_n12741, new_n12742, new_n12743, new_n12744, new_n12745, new_n12746,
    new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752,
    new_n12753, new_n12754, new_n12755, new_n12756, new_n12757, new_n12758,
    new_n12759, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764,
    new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770,
    new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783, new_n12784, new_n12785, new_n12786, new_n12787, new_n12788,
    new_n12789, new_n12790, new_n12791, new_n12792, new_n12793, new_n12794,
    new_n12795, new_n12796, new_n12798, new_n12799, new_n12800, new_n12801,
    new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842, new_n12843,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860, new_n12861,
    new_n12862, new_n12863, new_n12864, new_n12865, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870, new_n12871, new_n12872, new_n12873,
    new_n12874, new_n12875, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897,
    new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903,
    new_n12904, new_n12905, new_n12906, new_n12907, new_n12908, new_n12909,
    new_n12910, new_n12911, new_n12912, new_n12913, new_n12914, new_n12915,
    new_n12916, new_n12917, new_n12918, new_n12919, new_n12920, new_n12921,
    new_n12922, new_n12923, new_n12924, new_n12925, new_n12926, new_n12927,
    new_n12928, new_n12929, new_n12930, new_n12931, new_n12932, new_n12933,
    new_n12934, new_n12935, new_n12936, new_n12937, new_n12938, new_n12939,
    new_n12940, new_n12941, new_n12942, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956, new_n12957,
    new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963,
    new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969,
    new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975,
    new_n12976, new_n12977, new_n12978, new_n12979, new_n12980, new_n12981,
    new_n12982, new_n12983, new_n12984, new_n12985, new_n12986, new_n12987,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992, new_n12993,
    new_n12994, new_n12995, new_n12996, new_n12997, new_n12998, new_n12999,
    new_n13000, new_n13001, new_n13002, new_n13003, new_n13004, new_n13005,
    new_n13006, new_n13007, new_n13008, new_n13009, new_n13010, new_n13011,
    new_n13012, new_n13013, new_n13014, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030,
    new_n13031, new_n13032, new_n13033, new_n13034, new_n13035, new_n13036,
    new_n13037, new_n13038, new_n13039, new_n13040, new_n13041, new_n13042,
    new_n13043, new_n13044, new_n13045, new_n13046, new_n13047, new_n13048,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053, new_n13054,
    new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126,
    new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132,
    new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138,
    new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144,
    new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150,
    new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156,
    new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162,
    new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13217,
    new_n13218, new_n13219, new_n13220, new_n13221, new_n13222, new_n13223,
    new_n13224, new_n13225, new_n13226, new_n13227, new_n13228, new_n13229,
    new_n13230, new_n13231, new_n13232, new_n13233, new_n13234, new_n13235,
    new_n13236, new_n13237, new_n13238, new_n13239, new_n13240, new_n13241,
    new_n13242, new_n13243, new_n13244, new_n13245, new_n13246, new_n13247,
    new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253,
    new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259,
    new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270, new_n13271,
    new_n13272, new_n13273, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283,
    new_n13284, new_n13285, new_n13286, new_n13287, new_n13288, new_n13289,
    new_n13290, new_n13291, new_n13292, new_n13293, new_n13294, new_n13295,
    new_n13296, new_n13297, new_n13298, new_n13299, new_n13300, new_n13301,
    new_n13302, new_n13303, new_n13304, new_n13305, new_n13306, new_n13307,
    new_n13308, new_n13309, new_n13310, new_n13311, new_n13312, new_n13313,
    new_n13314, new_n13315, new_n13316, new_n13317, new_n13318, new_n13319,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333, new_n13334, new_n13335, new_n13336, new_n13337,
    new_n13338, new_n13339, new_n13340, new_n13341, new_n13342, new_n13343,
    new_n13344, new_n13345, new_n13346, new_n13347, new_n13348, new_n13349,
    new_n13350, new_n13351, new_n13352, new_n13353, new_n13354, new_n13355,
    new_n13356, new_n13357, new_n13358, new_n13359, new_n13360, new_n13361,
    new_n13362, new_n13363, new_n13364, new_n13365, new_n13366, new_n13367,
    new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373,
    new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407, new_n13408, new_n13409,
    new_n13410, new_n13411, new_n13412, new_n13413, new_n13414, new_n13415,
    new_n13416, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506,
    new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512,
    new_n13513, new_n13514, new_n13515, new_n13516, new_n13517, new_n13518,
    new_n13519, new_n13520, new_n13521, new_n13522, new_n13523, new_n13524,
    new_n13525, new_n13526, new_n13527, new_n13528, new_n13529, new_n13530,
    new_n13531, new_n13532, new_n13533, new_n13534, new_n13535, new_n13536,
    new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13548,
    new_n13549, new_n13550, new_n13551, new_n13552, new_n13553, new_n13554,
    new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729,
    new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735,
    new_n13736, new_n13737, new_n13738, new_n13739, new_n13740, new_n13741,
    new_n13742, new_n13743, new_n13744, new_n13745, new_n13746, new_n13747,
    new_n13748, new_n13749, new_n13750, new_n13751, new_n13752, new_n13753,
    new_n13754, new_n13755, new_n13756, new_n13757, new_n13758, new_n13759,
    new_n13760, new_n13761, new_n13762, new_n13763, new_n13764, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775, new_n13776, new_n13777,
    new_n13778, new_n13779, new_n13780, new_n13781, new_n13782, new_n13783,
    new_n13784, new_n13785, new_n13786, new_n13787, new_n13788, new_n13789,
    new_n13790, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850,
    new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856,
    new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862,
    new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868,
    new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874,
    new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880,
    new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886,
    new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892,
    new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898,
    new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904,
    new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910,
    new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13919, new_n13920, new_n13921, new_n13922,
    new_n13923, new_n13924, new_n13925, new_n13926, new_n13927, new_n13928,
    new_n13929, new_n13930, new_n13931, new_n13932, new_n13933, new_n13934,
    new_n13935, new_n13936, new_n13937, new_n13938, new_n13939, new_n13940,
    new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946,
    new_n13947, new_n13948, new_n13949, new_n13950, new_n13951, new_n13952,
    new_n13953, new_n13954, new_n13955, new_n13956, new_n13957, new_n13958,
    new_n13959, new_n13960, new_n13961, new_n13962, new_n13963, new_n13964,
    new_n13965, new_n13966, new_n13967, new_n13968, new_n13969, new_n13970,
    new_n13971, new_n13972, new_n13973, new_n13974, new_n13975, new_n13976,
    new_n13977, new_n13978, new_n13979, new_n13980, new_n13981, new_n13982,
    new_n13983, new_n13984, new_n13985, new_n13986, new_n13987, new_n13988,
    new_n13989, new_n13990, new_n13991, new_n13992, new_n13993, new_n13994,
    new_n13995, new_n13996, new_n13997, new_n13998, new_n13999, new_n14000,
    new_n14002, new_n14003, new_n14004, new_n14005, new_n14006, new_n14007,
    new_n14008, new_n14009, new_n14010, new_n14011, new_n14012, new_n14013,
    new_n14014, new_n14015, new_n14016, new_n14017, new_n14018, new_n14019,
    new_n14020, new_n14021, new_n14022, new_n14023, new_n14024, new_n14025,
    new_n14026, new_n14027, new_n14028, new_n14029, new_n14030, new_n14031,
    new_n14032, new_n14033, new_n14034, new_n14035, new_n14036, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059, new_n14060, new_n14061,
    new_n14062, new_n14063, new_n14064, new_n14065, new_n14066, new_n14067,
    new_n14068, new_n14069, new_n14070, new_n14071, new_n14072, new_n14073,
    new_n14074, new_n14075, new_n14076, new_n14077, new_n14078, new_n14079,
    new_n14080, new_n14081, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090, new_n14091,
    new_n14092, new_n14093, new_n14094, new_n14095, new_n14096, new_n14097,
    new_n14098, new_n14099, new_n14100, new_n14101, new_n14102, new_n14103,
    new_n14104, new_n14105, new_n14106, new_n14107, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120, new_n14121,
    new_n14122, new_n14123, new_n14124, new_n14125, new_n14126, new_n14127,
    new_n14128, new_n14129, new_n14130, new_n14131, new_n14132, new_n14133,
    new_n14134, new_n14135, new_n14136, new_n14137, new_n14138, new_n14139,
    new_n14140, new_n14141, new_n14142, new_n14143, new_n14144, new_n14145,
    new_n14146, new_n14147, new_n14148, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14170,
    new_n14171, new_n14172, new_n14173, new_n14174, new_n14175, new_n14176,
    new_n14177, new_n14178, new_n14179, new_n14180, new_n14181, new_n14182,
    new_n14183, new_n14184, new_n14185, new_n14186, new_n14187, new_n14188,
    new_n14189, new_n14190, new_n14191, new_n14192, new_n14193, new_n14194,
    new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200,
    new_n14201, new_n14202, new_n14203, new_n14204, new_n14205, new_n14206,
    new_n14207, new_n14208, new_n14209, new_n14210, new_n14211, new_n14212,
    new_n14213, new_n14214, new_n14215, new_n14216, new_n14217, new_n14218,
    new_n14219, new_n14220, new_n14221, new_n14222, new_n14223, new_n14224,
    new_n14225, new_n14226, new_n14227, new_n14228, new_n14229, new_n14230,
    new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236,
    new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242,
    new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267, new_n14268, new_n14269, new_n14270, new_n14271, new_n14272,
    new_n14273, new_n14274, new_n14275, new_n14276, new_n14277, new_n14278,
    new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284,
    new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290,
    new_n14291, new_n14292, new_n14293, new_n14294, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310, new_n14311, new_n14312, new_n14313, new_n14314,
    new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320,
    new_n14321, new_n14322, new_n14323, new_n14324, new_n14325, new_n14326,
    new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332,
    new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342, new_n14343, new_n14344,
    new_n14345, new_n14346, new_n14347, new_n14348, new_n14349, new_n14350,
    new_n14351, new_n14352, new_n14353, new_n14354, new_n14355, new_n14357,
    new_n14358, new_n14359, new_n14360, new_n14361, new_n14362, new_n14363,
    new_n14364, new_n14365, new_n14366, new_n14367, new_n14368, new_n14369,
    new_n14370, new_n14371, new_n14372, new_n14373, new_n14374, new_n14375,
    new_n14376, new_n14377, new_n14378, new_n14379, new_n14380, new_n14381,
    new_n14382, new_n14383, new_n14384, new_n14385, new_n14386, new_n14387,
    new_n14388, new_n14389, new_n14390, new_n14391, new_n14392, new_n14393,
    new_n14394, new_n14395, new_n14396, new_n14397, new_n14398, new_n14399,
    new_n14400, new_n14401, new_n14402, new_n14403, new_n14404, new_n14405,
    new_n14406, new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412, new_n14413, new_n14414, new_n14415, new_n14416, new_n14417,
    new_n14418, new_n14419, new_n14420, new_n14421, new_n14422, new_n14423,
    new_n14424, new_n14425, new_n14426, new_n14427, new_n14428, new_n14429,
    new_n14430, new_n14431, new_n14432, new_n14433, new_n14434, new_n14435,
    new_n14436, new_n14437, new_n14438, new_n14439, new_n14440, new_n14441,
    new_n14442, new_n14443, new_n14444, new_n14445, new_n14446, new_n14447,
    new_n14448, new_n14449, new_n14450, new_n14451, new_n14452, new_n14453,
    new_n14454, new_n14455, new_n14456, new_n14457, new_n14458, new_n14459,
    new_n14460, new_n14461, new_n14462, new_n14463, new_n14464, new_n14465,
    new_n14466, new_n14467, new_n14468, new_n14469, new_n14470, new_n14471,
    new_n14472, new_n14473, new_n14474, new_n14475, new_n14476, new_n14477,
    new_n14478, new_n14479, new_n14480, new_n14481, new_n14482, new_n14483,
    new_n14484, new_n14485, new_n14486, new_n14487, new_n14488, new_n14489,
    new_n14490, new_n14491, new_n14492, new_n14493, new_n14494, new_n14495,
    new_n14496, new_n14497, new_n14498, new_n14499, new_n14500, new_n14501,
    new_n14502, new_n14503, new_n14504, new_n14505, new_n14506, new_n14507,
    new_n14508, new_n14509, new_n14510, new_n14511, new_n14512, new_n14513,
    new_n14514, new_n14515, new_n14516, new_n14517, new_n14518, new_n14519,
    new_n14520, new_n14521, new_n14522, new_n14523, new_n14524, new_n14525,
    new_n14526, new_n14527, new_n14528, new_n14529, new_n14530, new_n14531,
    new_n14532, new_n14533, new_n14534, new_n14535, new_n14536, new_n14537,
    new_n14538, new_n14539, new_n14540, new_n14541, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546, new_n14547, new_n14548, new_n14549,
    new_n14550, new_n14551, new_n14552, new_n14553, new_n14554, new_n14555,
    new_n14556, new_n14557, new_n14558, new_n14559, new_n14560, new_n14561,
    new_n14562, new_n14563, new_n14564, new_n14565, new_n14566, new_n14568,
    new_n14569, new_n14570, new_n14571, new_n14572, new_n14573, new_n14574,
    new_n14575, new_n14576, new_n14577, new_n14578, new_n14579, new_n14580,
    new_n14581, new_n14582, new_n14583, new_n14584, new_n14585, new_n14586,
    new_n14587, new_n14588, new_n14589, new_n14590, new_n14591, new_n14592,
    new_n14593, new_n14594, new_n14595, new_n14596, new_n14597, new_n14598,
    new_n14599, new_n14600, new_n14601, new_n14602, new_n14603, new_n14604,
    new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610,
    new_n14611, new_n14612, new_n14613, new_n14614, new_n14615, new_n14616,
    new_n14617, new_n14618, new_n14619, new_n14620, new_n14621, new_n14622,
    new_n14623, new_n14624, new_n14625, new_n14626, new_n14627, new_n14628,
    new_n14629, new_n14630, new_n14631, new_n14632, new_n14633, new_n14634,
    new_n14635, new_n14636, new_n14637, new_n14638, new_n14639, new_n14640,
    new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646,
    new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652,
    new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658,
    new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664,
    new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670,
    new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676,
    new_n14677, new_n14678, new_n14679, new_n14680, new_n14681, new_n14682,
    new_n14683, new_n14684, new_n14685, new_n14686, new_n14687, new_n14688,
    new_n14689, new_n14690, new_n14691, new_n14692, new_n14693, new_n14694,
    new_n14695, new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701, new_n14702, new_n14703, new_n14704, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14727, new_n14728, new_n14729, new_n14730, new_n14731,
    new_n14732, new_n14733, new_n14734, new_n14735, new_n14736, new_n14737,
    new_n14738, new_n14739, new_n14740, new_n14741, new_n14742, new_n14743,
    new_n14744, new_n14745, new_n14746, new_n14747, new_n14748, new_n14749,
    new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14755,
    new_n14756, new_n14757, new_n14758, new_n14759, new_n14760, new_n14761,
    new_n14762, new_n14763, new_n14764, new_n14765, new_n14766, new_n14767,
    new_n14768, new_n14769, new_n14770, new_n14771, new_n14772, new_n14773,
    new_n14774, new_n14775, new_n14776, new_n14777, new_n14778, new_n14779,
    new_n14780, new_n14781, new_n14782, new_n14783, new_n14784, new_n14785,
    new_n14786, new_n14787, new_n14788, new_n14789, new_n14790, new_n14791,
    new_n14792, new_n14793, new_n14794, new_n14795, new_n14796, new_n14797,
    new_n14798, new_n14799, new_n14800, new_n14801, new_n14802, new_n14803,
    new_n14804, new_n14805, new_n14806, new_n14807, new_n14808, new_n14809,
    new_n14810, new_n14811, new_n14812, new_n14813, new_n14814, new_n14815,
    new_n14816, new_n14817, new_n14818, new_n14819, new_n14820, new_n14821,
    new_n14822, new_n14823, new_n14824, new_n14825, new_n14826, new_n14827,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838, new_n14839,
    new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845,
    new_n14846, new_n14847, new_n14848, new_n14849, new_n14850, new_n14851,
    new_n14852, new_n14853, new_n14854, new_n14855, new_n14856, new_n14857,
    new_n14858, new_n14859, new_n14860, new_n14861, new_n14862, new_n14863,
    new_n14864, new_n14865, new_n14866, new_n14867, new_n14868, new_n14869,
    new_n14870, new_n14871, new_n14872, new_n14873, new_n14874, new_n14875,
    new_n14876, new_n14877, new_n14878, new_n14879, new_n14880, new_n14881,
    new_n14882, new_n14883, new_n14884, new_n14885, new_n14886, new_n14887,
    new_n14888, new_n14889, new_n14890, new_n14891, new_n14892, new_n14893,
    new_n14894, new_n14895, new_n14896, new_n14897, new_n14898, new_n14899,
    new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905,
    new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911,
    new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917,
    new_n14918, new_n14919, new_n14920, new_n14921, new_n14922, new_n14923,
    new_n14924, new_n14925, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931, new_n14932, new_n14933, new_n14934, new_n14935, new_n14936,
    new_n14937, new_n14938, new_n14939, new_n14940, new_n14941, new_n14942,
    new_n14943, new_n14944, new_n14945, new_n14946, new_n14947, new_n14948,
    new_n14949, new_n14950, new_n14951, new_n14952, new_n14953, new_n14954,
    new_n14955, new_n14956, new_n14957, new_n14958, new_n14959, new_n14960,
    new_n14961, new_n14962, new_n14963, new_n14964, new_n14965, new_n14966,
    new_n14967, new_n14968, new_n14969, new_n14970, new_n14971, new_n14972,
    new_n14973, new_n14974, new_n14975, new_n14976, new_n14977, new_n14978,
    new_n14979, new_n14980, new_n14981, new_n14982, new_n14983, new_n14984,
    new_n14985, new_n14986, new_n14987, new_n14988, new_n14989, new_n14990,
    new_n14991, new_n14992, new_n14993, new_n14994, new_n14995, new_n14996,
    new_n14997, new_n14998, new_n14999, new_n15000, new_n15001, new_n15002,
    new_n15003, new_n15004, new_n15005, new_n15006, new_n15007, new_n15008,
    new_n15009, new_n15010, new_n15011, new_n15012, new_n15013, new_n15014,
    new_n15015, new_n15016, new_n15017, new_n15018, new_n15019, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031, new_n15032,
    new_n15033, new_n15034, new_n15035, new_n15036, new_n15037, new_n15038,
    new_n15039, new_n15040, new_n15041, new_n15042, new_n15043, new_n15044,
    new_n15045, new_n15046, new_n15047, new_n15048, new_n15049, new_n15050,
    new_n15051, new_n15052, new_n15053, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077, new_n15078, new_n15079, new_n15080,
    new_n15081, new_n15082, new_n15083, new_n15084, new_n15085, new_n15086,
    new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094, new_n15095, new_n15096, new_n15097, new_n15098,
    new_n15099, new_n15100, new_n15101, new_n15103, new_n15104, new_n15105,
    new_n15106, new_n15107, new_n15108, new_n15109, new_n15110, new_n15111,
    new_n15112, new_n15113, new_n15114, new_n15115, new_n15116, new_n15117,
    new_n15118, new_n15119, new_n15120, new_n15121, new_n15122, new_n15123,
    new_n15124, new_n15125, new_n15126, new_n15127, new_n15128, new_n15129,
    new_n15130, new_n15131, new_n15132, new_n15133, new_n15134, new_n15135,
    new_n15136, new_n15137, new_n15138, new_n15139, new_n15140, new_n15141,
    new_n15142, new_n15143, new_n15144, new_n15145, new_n15146, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15160, new_n15161, new_n15162, new_n15163, new_n15164, new_n15165,
    new_n15166, new_n15167, new_n15168, new_n15169, new_n15170, new_n15171,
    new_n15172, new_n15173, new_n15174, new_n15175, new_n15176, new_n15177,
    new_n15178, new_n15179, new_n15180, new_n15181, new_n15182, new_n15183,
    new_n15184, new_n15185, new_n15186, new_n15187, new_n15188, new_n15189,
    new_n15190, new_n15191, new_n15192, new_n15193, new_n15194, new_n15195,
    new_n15196, new_n15197, new_n15198, new_n15199, new_n15200, new_n15201,
    new_n15202, new_n15203, new_n15204, new_n15205, new_n15206, new_n15207,
    new_n15208, new_n15209, new_n15210, new_n15211, new_n15212, new_n15213,
    new_n15214, new_n15215, new_n15216, new_n15217, new_n15218, new_n15219,
    new_n15220, new_n15221, new_n15222, new_n15223, new_n15224, new_n15225,
    new_n15226, new_n15227, new_n15228, new_n15229, new_n15230, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241, new_n15242, new_n15243,
    new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249,
    new_n15250, new_n15251, new_n15252, new_n15253, new_n15254, new_n15255,
    new_n15256, new_n15257, new_n15258, new_n15259, new_n15260, new_n15261,
    new_n15262, new_n15263, new_n15264, new_n15265, new_n15266, new_n15267,
    new_n15268, new_n15269, new_n15270, new_n15272, new_n15273, new_n15274,
    new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280,
    new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286,
    new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304,
    new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322,
    new_n15323, new_n15324, new_n15325, new_n15326, new_n15327, new_n15328,
    new_n15329, new_n15330, new_n15331, new_n15332, new_n15333, new_n15334,
    new_n15335, new_n15336, new_n15337, new_n15338, new_n15339, new_n15340,
    new_n15341, new_n15342, new_n15343, new_n15344, new_n15345, new_n15346,
    new_n15347, new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353, new_n15354, new_n15355, new_n15356, new_n15357, new_n15358,
    new_n15359, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366, new_n15367, new_n15368, new_n15369, new_n15370,
    new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376,
    new_n15377, new_n15378, new_n15379, new_n15380, new_n15381, new_n15382,
    new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388,
    new_n15389, new_n15390, new_n15391, new_n15392, new_n15393, new_n15394,
    new_n15395, new_n15396, new_n15397, new_n15398, new_n15399, new_n15400,
    new_n15401, new_n15402, new_n15403, new_n15404, new_n15405, new_n15406,
    new_n15407, new_n15408, new_n15409, new_n15410, new_n15411, new_n15412,
    new_n15413, new_n15414, new_n15415, new_n15416, new_n15417, new_n15418,
    new_n15419, new_n15420, new_n15421, new_n15422, new_n15423, new_n15424,
    new_n15425, new_n15426, new_n15427, new_n15428, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435, new_n15436,
    new_n15437, new_n15438, new_n15440, new_n15441, new_n15442, new_n15443,
    new_n15444, new_n15445, new_n15446, new_n15447, new_n15448, new_n15449,
    new_n15450, new_n15451, new_n15452, new_n15453, new_n15454, new_n15455,
    new_n15456, new_n15457, new_n15458, new_n15459, new_n15460, new_n15461,
    new_n15462, new_n15463, new_n15464, new_n15465, new_n15466, new_n15467,
    new_n15468, new_n15469, new_n15470, new_n15471, new_n15472, new_n15473,
    new_n15474, new_n15475, new_n15476, new_n15477, new_n15478, new_n15479,
    new_n15480, new_n15481, new_n15482, new_n15483, new_n15484, new_n15485,
    new_n15486, new_n15487, new_n15488, new_n15489, new_n15490, new_n15491,
    new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503,
    new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533,
    new_n15534, new_n15535, new_n15536, new_n15537, new_n15538, new_n15539,
    new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546, new_n15547, new_n15548, new_n15549, new_n15550, new_n15551,
    new_n15552, new_n15553, new_n15554, new_n15555, new_n15556, new_n15557,
    new_n15558, new_n15559, new_n15560, new_n15561, new_n15562, new_n15563,
    new_n15564, new_n15565, new_n15566, new_n15567, new_n15568, new_n15569,
    new_n15570, new_n15571, new_n15572, new_n15573, new_n15574, new_n15575,
    new_n15576, new_n15577, new_n15578, new_n15579, new_n15580, new_n15581,
    new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588, new_n15589, new_n15590, new_n15591, new_n15592, new_n15593,
    new_n15594, new_n15595, new_n15596, new_n15597, new_n15598, new_n15599,
    new_n15601, new_n15602, new_n15603, new_n15604, new_n15605, new_n15606,
    new_n15607, new_n15608, new_n15609, new_n15610, new_n15611, new_n15612,
    new_n15613, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635, new_n15636,
    new_n15637, new_n15638, new_n15639, new_n15640, new_n15641, new_n15642,
    new_n15643, new_n15644, new_n15645, new_n15646, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15757, new_n15758, new_n15760, new_n15761, new_n15762, new_n15763,
    new_n15764, new_n15765, new_n15766, new_n15767, new_n15768, new_n15769,
    new_n15770, new_n15771, new_n15772, new_n15773, new_n15774, new_n15775,
    new_n15776, new_n15777, new_n15778, new_n15779, new_n15780, new_n15781,
    new_n15782, new_n15783, new_n15784, new_n15785, new_n15786, new_n15787,
    new_n15788, new_n15789, new_n15790, new_n15791, new_n15792, new_n15793,
    new_n15794, new_n15795, new_n15796, new_n15797, new_n15798, new_n15799,
    new_n15800, new_n15801, new_n15802, new_n15803, new_n15804, new_n15805,
    new_n15806, new_n15807, new_n15808, new_n15809, new_n15810, new_n15811,
    new_n15812, new_n15813, new_n15814, new_n15815, new_n15816, new_n15817,
    new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823,
    new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829,
    new_n15830, new_n15831, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15842, new_n15843, new_n15844, new_n15845, new_n15846, new_n15847,
    new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853,
    new_n15854, new_n15855, new_n15856, new_n15857, new_n15858, new_n15859,
    new_n15860, new_n15861, new_n15862, new_n15863, new_n15864, new_n15865,
    new_n15866, new_n15867, new_n15868, new_n15869, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884, new_n15885, new_n15886, new_n15887, new_n15888, new_n15889,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917, new_n15918, new_n15919,
    new_n15920, new_n15921, new_n15922, new_n15923, new_n15924, new_n15925,
    new_n15926, new_n15927, new_n15928, new_n15930, new_n15931, new_n15932,
    new_n15933, new_n15934, new_n15935, new_n15936, new_n15937, new_n15938,
    new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944,
    new_n15945, new_n15946, new_n15947, new_n15948, new_n15949, new_n15950,
    new_n15951, new_n15952, new_n15953, new_n15954, new_n15955, new_n15956,
    new_n15957, new_n15958, new_n15959, new_n15960, new_n15961, new_n15962,
    new_n15963, new_n15964, new_n15965, new_n15966, new_n15967, new_n15968,
    new_n15969, new_n15970, new_n15971, new_n15972, new_n15973, new_n15974,
    new_n15975, new_n15976, new_n15977, new_n15978, new_n15979, new_n15980,
    new_n15981, new_n15982, new_n15983, new_n15984, new_n15985, new_n15986,
    new_n15987, new_n15988, new_n15989, new_n15990, new_n15991, new_n15992,
    new_n15993, new_n15994, new_n15995, new_n15996, new_n15997, new_n15998,
    new_n15999, new_n16000, new_n16001, new_n16002, new_n16003, new_n16004,
    new_n16005, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010,
    new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016,
    new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022,
    new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034,
    new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040,
    new_n16041, new_n16042, new_n16043, new_n16044, new_n16045, new_n16046,
    new_n16047, new_n16048, new_n16049, new_n16050, new_n16051, new_n16052,
    new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058,
    new_n16059, new_n16060, new_n16061, new_n16062, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068, new_n16069, new_n16070,
    new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076,
    new_n16077, new_n16078, new_n16079, new_n16080, new_n16081, new_n16082,
    new_n16083, new_n16084, new_n16085, new_n16086, new_n16088, new_n16089,
    new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095,
    new_n16096, new_n16097, new_n16098, new_n16099, new_n16100, new_n16101,
    new_n16102, new_n16103, new_n16104, new_n16105, new_n16106, new_n16107,
    new_n16108, new_n16109, new_n16110, new_n16111, new_n16112, new_n16113,
    new_n16114, new_n16115, new_n16116, new_n16117, new_n16118, new_n16119,
    new_n16120, new_n16121, new_n16122, new_n16123, new_n16124, new_n16125,
    new_n16126, new_n16127, new_n16128, new_n16129, new_n16130, new_n16131,
    new_n16132, new_n16133, new_n16134, new_n16135, new_n16136, new_n16137,
    new_n16138, new_n16139, new_n16140, new_n16141, new_n16142, new_n16143,
    new_n16144, new_n16145, new_n16146, new_n16147, new_n16148, new_n16149,
    new_n16150, new_n16151, new_n16152, new_n16153, new_n16154, new_n16155,
    new_n16156, new_n16157, new_n16158, new_n16159, new_n16160, new_n16161,
    new_n16162, new_n16163, new_n16164, new_n16165, new_n16166, new_n16167,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184, new_n16185,
    new_n16186, new_n16187, new_n16188, new_n16189, new_n16190, new_n16191,
    new_n16192, new_n16193, new_n16194, new_n16195, new_n16196, new_n16197,
    new_n16198, new_n16199, new_n16200, new_n16201, new_n16202, new_n16203,
    new_n16204, new_n16205, new_n16206, new_n16207, new_n16208, new_n16209,
    new_n16210, new_n16211, new_n16212, new_n16213, new_n16214, new_n16215,
    new_n16216, new_n16217, new_n16218, new_n16219, new_n16220, new_n16221,
    new_n16222, new_n16223, new_n16224, new_n16225, new_n16226, new_n16227,
    new_n16228, new_n16229, new_n16230, new_n16231, new_n16232, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16239, new_n16240,
    new_n16241, new_n16242, new_n16243, new_n16244, new_n16245, new_n16246,
    new_n16247, new_n16248, new_n16249, new_n16250, new_n16251, new_n16252,
    new_n16253, new_n16254, new_n16255, new_n16256, new_n16257, new_n16258,
    new_n16259, new_n16260, new_n16261, new_n16262, new_n16263, new_n16264,
    new_n16265, new_n16266, new_n16267, new_n16268, new_n16269, new_n16270,
    new_n16271, new_n16272, new_n16273, new_n16274, new_n16275, new_n16276,
    new_n16277, new_n16278, new_n16279, new_n16280, new_n16281, new_n16282,
    new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288,
    new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294,
    new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300,
    new_n16301, new_n16302, new_n16303, new_n16304, new_n16305, new_n16306,
    new_n16307, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312,
    new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318,
    new_n16319, new_n16320, new_n16321, new_n16322, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327, new_n16328, new_n16329, new_n16330,
    new_n16331, new_n16332, new_n16333, new_n16334, new_n16335, new_n16336,
    new_n16337, new_n16338, new_n16339, new_n16340, new_n16341, new_n16342,
    new_n16343, new_n16344, new_n16345, new_n16346, new_n16347, new_n16348,
    new_n16349, new_n16350, new_n16351, new_n16352, new_n16353, new_n16354,
    new_n16355, new_n16356, new_n16357, new_n16358, new_n16359, new_n16360,
    new_n16361, new_n16362, new_n16363, new_n16364, new_n16365, new_n16366,
    new_n16367, new_n16368, new_n16369, new_n16370, new_n16371, new_n16372,
    new_n16373, new_n16374, new_n16375, new_n16376, new_n16377, new_n16378,
    new_n16379, new_n16380, new_n16381, new_n16382, new_n16383, new_n16384,
    new_n16385, new_n16386, new_n16387, new_n16388, new_n16389, new_n16390,
    new_n16391, new_n16392, new_n16393, new_n16394, new_n16396, new_n16397,
    new_n16398, new_n16399, new_n16400, new_n16401, new_n16402, new_n16403,
    new_n16404, new_n16405, new_n16406, new_n16407, new_n16408, new_n16409,
    new_n16410, new_n16411, new_n16412, new_n16413, new_n16414, new_n16415,
    new_n16416, new_n16417, new_n16418, new_n16419, new_n16420, new_n16421,
    new_n16422, new_n16423, new_n16424, new_n16425, new_n16426, new_n16427,
    new_n16428, new_n16429, new_n16430, new_n16431, new_n16432, new_n16433,
    new_n16434, new_n16435, new_n16436, new_n16437, new_n16438, new_n16439,
    new_n16440, new_n16441, new_n16442, new_n16443, new_n16444, new_n16445,
    new_n16446, new_n16447, new_n16448, new_n16449, new_n16450, new_n16451,
    new_n16452, new_n16453, new_n16454, new_n16455, new_n16456, new_n16457,
    new_n16458, new_n16459, new_n16460, new_n16461, new_n16462, new_n16463,
    new_n16464, new_n16465, new_n16466, new_n16467, new_n16468, new_n16469,
    new_n16470, new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476, new_n16477, new_n16478, new_n16479, new_n16480, new_n16481,
    new_n16482, new_n16483, new_n16484, new_n16485, new_n16486, new_n16487,
    new_n16488, new_n16489, new_n16490, new_n16491, new_n16492, new_n16493,
    new_n16494, new_n16495, new_n16496, new_n16497, new_n16498, new_n16499,
    new_n16500, new_n16501, new_n16502, new_n16503, new_n16504, new_n16505,
    new_n16506, new_n16507, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516, new_n16517,
    new_n16518, new_n16519, new_n16520, new_n16521, new_n16522, new_n16523,
    new_n16524, new_n16525, new_n16526, new_n16527, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544, new_n16546, new_n16547, new_n16548,
    new_n16549, new_n16550, new_n16551, new_n16552, new_n16553, new_n16554,
    new_n16555, new_n16556, new_n16557, new_n16558, new_n16559, new_n16560,
    new_n16561, new_n16562, new_n16563, new_n16564, new_n16565, new_n16566,
    new_n16567, new_n16568, new_n16569, new_n16570, new_n16571, new_n16572,
    new_n16573, new_n16574, new_n16575, new_n16576, new_n16577, new_n16578,
    new_n16579, new_n16580, new_n16581, new_n16582, new_n16583, new_n16584,
    new_n16585, new_n16586, new_n16587, new_n16588, new_n16589, new_n16590,
    new_n16591, new_n16592, new_n16593, new_n16594, new_n16595, new_n16596,
    new_n16597, new_n16598, new_n16599, new_n16600, new_n16601, new_n16602,
    new_n16603, new_n16604, new_n16605, new_n16606, new_n16607, new_n16608,
    new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617, new_n16618, new_n16619, new_n16620,
    new_n16621, new_n16622, new_n16623, new_n16624, new_n16625, new_n16626,
    new_n16627, new_n16628, new_n16629, new_n16630, new_n16631, new_n16632,
    new_n16633, new_n16634, new_n16635, new_n16636, new_n16637, new_n16638,
    new_n16639, new_n16640, new_n16641, new_n16642, new_n16643, new_n16644,
    new_n16645, new_n16646, new_n16647, new_n16648, new_n16649, new_n16650,
    new_n16651, new_n16652, new_n16653, new_n16654, new_n16655, new_n16656,
    new_n16657, new_n16658, new_n16659, new_n16660, new_n16661, new_n16662,
    new_n16663, new_n16664, new_n16665, new_n16666, new_n16667, new_n16668,
    new_n16669, new_n16670, new_n16671, new_n16672, new_n16673, new_n16674,
    new_n16675, new_n16676, new_n16677, new_n16678, new_n16679, new_n16680,
    new_n16681, new_n16682, new_n16683, new_n16684, new_n16685, new_n16686,
    new_n16687, new_n16688, new_n16689, new_n16690, new_n16691, new_n16693,
    new_n16694, new_n16695, new_n16696, new_n16697, new_n16698, new_n16699,
    new_n16700, new_n16701, new_n16702, new_n16703, new_n16704, new_n16705,
    new_n16706, new_n16707, new_n16708, new_n16709, new_n16710, new_n16711,
    new_n16712, new_n16713, new_n16714, new_n16715, new_n16716, new_n16717,
    new_n16718, new_n16719, new_n16720, new_n16721, new_n16722, new_n16723,
    new_n16724, new_n16725, new_n16726, new_n16727, new_n16728, new_n16729,
    new_n16730, new_n16731, new_n16732, new_n16733, new_n16734, new_n16735,
    new_n16736, new_n16737, new_n16738, new_n16739, new_n16740, new_n16741,
    new_n16742, new_n16743, new_n16744, new_n16745, new_n16746, new_n16747,
    new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753,
    new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759,
    new_n16760, new_n16761, new_n16762, new_n16763, new_n16764, new_n16765,
    new_n16766, new_n16767, new_n16768, new_n16769, new_n16770, new_n16771,
    new_n16772, new_n16773, new_n16774, new_n16775, new_n16776, new_n16777,
    new_n16778, new_n16779, new_n16780, new_n16781, new_n16782, new_n16783,
    new_n16784, new_n16785, new_n16786, new_n16787, new_n16788, new_n16789,
    new_n16790, new_n16791, new_n16792, new_n16793, new_n16794, new_n16795,
    new_n16796, new_n16797, new_n16798, new_n16799, new_n16800, new_n16801,
    new_n16802, new_n16803, new_n16804, new_n16805, new_n16806, new_n16807,
    new_n16808, new_n16809, new_n16810, new_n16811, new_n16812, new_n16813,
    new_n16814, new_n16815, new_n16816, new_n16817, new_n16818, new_n16819,
    new_n16820, new_n16821, new_n16822, new_n16823, new_n16824, new_n16825,
    new_n16826, new_n16827, new_n16828, new_n16829, new_n16830, new_n16831,
    new_n16832, new_n16833, new_n16834, new_n16835, new_n16837, new_n16838,
    new_n16839, new_n16840, new_n16841, new_n16842, new_n16843, new_n16844,
    new_n16845, new_n16846, new_n16847, new_n16848, new_n16849, new_n16850,
    new_n16851, new_n16852, new_n16853, new_n16854, new_n16855, new_n16856,
    new_n16857, new_n16858, new_n16859, new_n16860, new_n16861, new_n16862,
    new_n16863, new_n16864, new_n16865, new_n16866, new_n16867, new_n16868,
    new_n16869, new_n16870, new_n16871, new_n16872, new_n16873, new_n16874,
    new_n16875, new_n16876, new_n16877, new_n16878, new_n16879, new_n16880,
    new_n16881, new_n16882, new_n16883, new_n16884, new_n16885, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905, new_n16906, new_n16907, new_n16908, new_n16909, new_n16910,
    new_n16911, new_n16912, new_n16913, new_n16914, new_n16915, new_n16916,
    new_n16917, new_n16918, new_n16919, new_n16920, new_n16921, new_n16922,
    new_n16923, new_n16924, new_n16925, new_n16926, new_n16927, new_n16928,
    new_n16929, new_n16930, new_n16931, new_n16932, new_n16933, new_n16934,
    new_n16935, new_n16936, new_n16937, new_n16938, new_n16939, new_n16940,
    new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946,
    new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952,
    new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958,
    new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964,
    new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970,
    new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976,
    new_n16977, new_n16978, new_n16979, new_n16980, new_n16982, new_n16983,
    new_n16984, new_n16985, new_n16986, new_n16987, new_n16988, new_n16989,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994, new_n16995,
    new_n16996, new_n16997, new_n16998, new_n16999, new_n17000, new_n17001,
    new_n17002, new_n17003, new_n17004, new_n17005, new_n17006, new_n17007,
    new_n17008, new_n17009, new_n17010, new_n17011, new_n17012, new_n17013,
    new_n17014, new_n17015, new_n17016, new_n17017, new_n17018, new_n17019,
    new_n17020, new_n17021, new_n17022, new_n17023, new_n17024, new_n17025,
    new_n17026, new_n17027, new_n17028, new_n17029, new_n17030, new_n17031,
    new_n17032, new_n17033, new_n17034, new_n17035, new_n17036, new_n17037,
    new_n17038, new_n17039, new_n17040, new_n17041, new_n17042, new_n17043,
    new_n17044, new_n17045, new_n17046, new_n17047, new_n17048, new_n17049,
    new_n17050, new_n17051, new_n17052, new_n17053, new_n17054, new_n17055,
    new_n17056, new_n17057, new_n17058, new_n17059, new_n17060, new_n17061,
    new_n17062, new_n17063, new_n17064, new_n17065, new_n17066, new_n17067,
    new_n17068, new_n17069, new_n17070, new_n17071, new_n17072, new_n17073,
    new_n17074, new_n17075, new_n17076, new_n17077, new_n17078, new_n17079,
    new_n17080, new_n17081, new_n17082, new_n17083, new_n17084, new_n17085,
    new_n17086, new_n17087, new_n17088, new_n17089, new_n17090, new_n17091,
    new_n17092, new_n17093, new_n17094, new_n17095, new_n17096, new_n17097,
    new_n17098, new_n17099, new_n17100, new_n17101, new_n17102, new_n17103,
    new_n17104, new_n17105, new_n17106, new_n17107, new_n17108, new_n17109,
    new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17116,
    new_n17117, new_n17118, new_n17119, new_n17120, new_n17121, new_n17122,
    new_n17123, new_n17124, new_n17125, new_n17126, new_n17127, new_n17128,
    new_n17129, new_n17130, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138, new_n17139, new_n17140,
    new_n17141, new_n17142, new_n17143, new_n17144, new_n17145, new_n17146,
    new_n17147, new_n17148, new_n17149, new_n17150, new_n17151, new_n17152,
    new_n17153, new_n17154, new_n17155, new_n17156, new_n17157, new_n17158,
    new_n17159, new_n17160, new_n17161, new_n17162, new_n17163, new_n17164,
    new_n17165, new_n17166, new_n17167, new_n17168, new_n17169, new_n17170,
    new_n17171, new_n17172, new_n17173, new_n17174, new_n17175, new_n17176,
    new_n17177, new_n17178, new_n17179, new_n17180, new_n17181, new_n17182,
    new_n17183, new_n17184, new_n17185, new_n17186, new_n17187, new_n17188,
    new_n17189, new_n17190, new_n17191, new_n17192, new_n17193, new_n17194,
    new_n17195, new_n17196, new_n17197, new_n17198, new_n17199, new_n17200,
    new_n17201, new_n17202, new_n17203, new_n17204, new_n17205, new_n17206,
    new_n17207, new_n17208, new_n17209, new_n17210, new_n17211, new_n17212,
    new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218,
    new_n17219, new_n17220, new_n17221, new_n17222, new_n17223, new_n17224,
    new_n17225, new_n17226, new_n17227, new_n17228, new_n17229, new_n17230,
    new_n17231, new_n17232, new_n17233, new_n17234, new_n17235, new_n17236,
    new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243, new_n17244, new_n17245, new_n17246, new_n17247, new_n17248,
    new_n17249, new_n17250, new_n17251, new_n17252, new_n17253, new_n17254,
    new_n17255, new_n17256, new_n17258, new_n17259, new_n17260, new_n17261,
    new_n17262, new_n17263, new_n17264, new_n17265, new_n17266, new_n17267,
    new_n17268, new_n17269, new_n17270, new_n17271, new_n17272, new_n17273,
    new_n17274, new_n17275, new_n17276, new_n17277, new_n17278, new_n17279,
    new_n17280, new_n17281, new_n17282, new_n17283, new_n17284, new_n17285,
    new_n17286, new_n17287, new_n17288, new_n17289, new_n17290, new_n17291,
    new_n17292, new_n17293, new_n17294, new_n17295, new_n17296, new_n17297,
    new_n17298, new_n17299, new_n17300, new_n17301, new_n17302, new_n17303,
    new_n17304, new_n17305, new_n17306, new_n17307, new_n17308, new_n17309,
    new_n17310, new_n17311, new_n17312, new_n17313, new_n17314, new_n17315,
    new_n17316, new_n17317, new_n17318, new_n17319, new_n17320, new_n17321,
    new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327,
    new_n17328, new_n17329, new_n17330, new_n17331, new_n17332, new_n17333,
    new_n17334, new_n17335, new_n17336, new_n17337, new_n17338, new_n17339,
    new_n17340, new_n17341, new_n17342, new_n17343, new_n17344, new_n17345,
    new_n17346, new_n17347, new_n17348, new_n17349, new_n17350, new_n17351,
    new_n17352, new_n17353, new_n17354, new_n17355, new_n17356, new_n17357,
    new_n17358, new_n17359, new_n17360, new_n17361, new_n17362, new_n17363,
    new_n17364, new_n17365, new_n17366, new_n17367, new_n17368, new_n17369,
    new_n17370, new_n17371, new_n17372, new_n17373, new_n17374, new_n17375,
    new_n17376, new_n17377, new_n17378, new_n17379, new_n17380, new_n17381,
    new_n17382, new_n17383, new_n17384, new_n17385, new_n17387, new_n17388,
    new_n17389, new_n17390, new_n17391, new_n17392, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421, new_n17422, new_n17423, new_n17424,
    new_n17425, new_n17426, new_n17427, new_n17428, new_n17429, new_n17430,
    new_n17431, new_n17432, new_n17433, new_n17434, new_n17435, new_n17436,
    new_n17437, new_n17438, new_n17439, new_n17440, new_n17441, new_n17442,
    new_n17443, new_n17444, new_n17445, new_n17446, new_n17447, new_n17448,
    new_n17449, new_n17450, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458, new_n17459, new_n17460,
    new_n17461, new_n17462, new_n17463, new_n17464, new_n17465, new_n17466,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490,
    new_n17491, new_n17492, new_n17493, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508,
    new_n17509, new_n17510, new_n17511, new_n17512, new_n17514, new_n17515,
    new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521,
    new_n17522, new_n17523, new_n17524, new_n17525, new_n17526, new_n17527,
    new_n17528, new_n17529, new_n17530, new_n17531, new_n17532, new_n17533,
    new_n17534, new_n17535, new_n17536, new_n17537, new_n17538, new_n17539,
    new_n17540, new_n17541, new_n17542, new_n17543, new_n17544, new_n17545,
    new_n17546, new_n17547, new_n17548, new_n17549, new_n17550, new_n17551,
    new_n17552, new_n17553, new_n17554, new_n17555, new_n17556, new_n17557,
    new_n17558, new_n17559, new_n17560, new_n17561, new_n17562, new_n17563,
    new_n17564, new_n17565, new_n17566, new_n17567, new_n17568, new_n17569,
    new_n17570, new_n17571, new_n17572, new_n17573, new_n17574, new_n17575,
    new_n17576, new_n17577, new_n17578, new_n17579, new_n17580, new_n17581,
    new_n17582, new_n17583, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592, new_n17593,
    new_n17594, new_n17595, new_n17596, new_n17597, new_n17598, new_n17599,
    new_n17600, new_n17601, new_n17602, new_n17603, new_n17604, new_n17605,
    new_n17606, new_n17607, new_n17608, new_n17609, new_n17610, new_n17611,
    new_n17612, new_n17613, new_n17614, new_n17615, new_n17616, new_n17617,
    new_n17618, new_n17619, new_n17620, new_n17621, new_n17622, new_n17623,
    new_n17624, new_n17625, new_n17626, new_n17627, new_n17628, new_n17629,
    new_n17630, new_n17631, new_n17632, new_n17633, new_n17634, new_n17635,
    new_n17636, new_n17637, new_n17638, new_n17639, new_n17640, new_n17641,
    new_n17642, new_n17643, new_n17644, new_n17645, new_n17646, new_n17647,
    new_n17648, new_n17649, new_n17651, new_n17652, new_n17653, new_n17654,
    new_n17655, new_n17656, new_n17657, new_n17658, new_n17659, new_n17660,
    new_n17661, new_n17662, new_n17663, new_n17664, new_n17665, new_n17666,
    new_n17667, new_n17668, new_n17669, new_n17670, new_n17671, new_n17672,
    new_n17673, new_n17674, new_n17675, new_n17676, new_n17677, new_n17678,
    new_n17679, new_n17680, new_n17681, new_n17682, new_n17683, new_n17684,
    new_n17685, new_n17686, new_n17687, new_n17688, new_n17689, new_n17690,
    new_n17691, new_n17692, new_n17693, new_n17694, new_n17695, new_n17696,
    new_n17697, new_n17698, new_n17699, new_n17700, new_n17701, new_n17702,
    new_n17703, new_n17704, new_n17705, new_n17706, new_n17707, new_n17708,
    new_n17709, new_n17710, new_n17711, new_n17712, new_n17713, new_n17714,
    new_n17715, new_n17716, new_n17717, new_n17718, new_n17719, new_n17720,
    new_n17721, new_n17722, new_n17723, new_n17724, new_n17725, new_n17726,
    new_n17727, new_n17728, new_n17729, new_n17730, new_n17731, new_n17732,
    new_n17733, new_n17734, new_n17735, new_n17736, new_n17737, new_n17738,
    new_n17739, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744,
    new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17777, new_n17778, new_n17779, new_n17780, new_n17781,
    new_n17782, new_n17783, new_n17784, new_n17785, new_n17786, new_n17787,
    new_n17788, new_n17789, new_n17790, new_n17791, new_n17792, new_n17793,
    new_n17794, new_n17795, new_n17796, new_n17797, new_n17798, new_n17799,
    new_n17800, new_n17801, new_n17802, new_n17803, new_n17804, new_n17805,
    new_n17806, new_n17807, new_n17808, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820, new_n17821, new_n17822, new_n17823,
    new_n17824, new_n17825, new_n17826, new_n17827, new_n17828, new_n17829,
    new_n17830, new_n17831, new_n17832, new_n17833, new_n17834, new_n17835,
    new_n17836, new_n17837, new_n17838, new_n17839, new_n17840, new_n17841,
    new_n17842, new_n17843, new_n17844, new_n17845, new_n17846, new_n17847,
    new_n17848, new_n17849, new_n17850, new_n17851, new_n17852, new_n17853,
    new_n17854, new_n17855, new_n17856, new_n17857, new_n17858, new_n17859,
    new_n17860, new_n17861, new_n17862, new_n17863, new_n17864, new_n17865,
    new_n17866, new_n17867, new_n17868, new_n17869, new_n17870, new_n17871,
    new_n17872, new_n17873, new_n17874, new_n17875, new_n17876, new_n17877,
    new_n17878, new_n17879, new_n17880, new_n17881, new_n17882, new_n17883,
    new_n17884, new_n17885, new_n17886, new_n17887, new_n17888, new_n17889,
    new_n17890, new_n17891, new_n17893, new_n17894, new_n17895, new_n17896,
    new_n17897, new_n17898, new_n17899, new_n17900, new_n17901, new_n17902,
    new_n17903, new_n17904, new_n17905, new_n17906, new_n17907, new_n17908,
    new_n17909, new_n17910, new_n17911, new_n17912, new_n17913, new_n17914,
    new_n17915, new_n17916, new_n17917, new_n17918, new_n17919, new_n17920,
    new_n17921, new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17927, new_n17928, new_n17929, new_n17930, new_n17931, new_n17932,
    new_n17933, new_n17934, new_n17935, new_n17936, new_n17937, new_n17938,
    new_n17939, new_n17940, new_n17941, new_n17942, new_n17943, new_n17944,
    new_n17945, new_n17946, new_n17947, new_n17948, new_n17949, new_n17950,
    new_n17951, new_n17952, new_n17953, new_n17954, new_n17955, new_n17956,
    new_n17957, new_n17958, new_n17959, new_n17960, new_n17961, new_n17962,
    new_n17963, new_n17964, new_n17965, new_n17966, new_n17967, new_n17968,
    new_n17969, new_n17970, new_n17971, new_n17972, new_n17973, new_n17974,
    new_n17975, new_n17976, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17995, new_n17996, new_n17997, new_n17998,
    new_n17999, new_n18000, new_n18001, new_n18002, new_n18003, new_n18004,
    new_n18005, new_n18006, new_n18007, new_n18008, new_n18009, new_n18010,
    new_n18011, new_n18012, new_n18013, new_n18014, new_n18015, new_n18016,
    new_n18017, new_n18018, new_n18019, new_n18020, new_n18021, new_n18023,
    new_n18024, new_n18025, new_n18026, new_n18027, new_n18028, new_n18029,
    new_n18030, new_n18031, new_n18032, new_n18033, new_n18034, new_n18035,
    new_n18036, new_n18037, new_n18038, new_n18039, new_n18040, new_n18041,
    new_n18042, new_n18043, new_n18044, new_n18045, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053,
    new_n18054, new_n18055, new_n18056, new_n18057, new_n18058, new_n18059,
    new_n18060, new_n18061, new_n18062, new_n18063, new_n18064, new_n18065,
    new_n18066, new_n18067, new_n18068, new_n18069, new_n18070, new_n18071,
    new_n18072, new_n18073, new_n18074, new_n18075, new_n18076, new_n18077,
    new_n18078, new_n18079, new_n18080, new_n18081, new_n18082, new_n18083,
    new_n18084, new_n18085, new_n18086, new_n18087, new_n18088, new_n18089,
    new_n18090, new_n18091, new_n18092, new_n18093, new_n18094, new_n18095,
    new_n18096, new_n18097, new_n18098, new_n18099, new_n18100, new_n18101,
    new_n18102, new_n18103, new_n18104, new_n18105, new_n18106, new_n18107,
    new_n18108, new_n18109, new_n18110, new_n18111, new_n18112, new_n18113,
    new_n18114, new_n18115, new_n18116, new_n18117, new_n18118, new_n18119,
    new_n18120, new_n18121, new_n18122, new_n18123, new_n18124, new_n18125,
    new_n18126, new_n18127, new_n18128, new_n18129, new_n18130, new_n18131,
    new_n18132, new_n18133, new_n18134, new_n18135, new_n18136, new_n18137,
    new_n18138, new_n18140, new_n18141, new_n18142, new_n18143, new_n18144,
    new_n18145, new_n18146, new_n18147, new_n18148, new_n18149, new_n18150,
    new_n18151, new_n18152, new_n18153, new_n18154, new_n18155, new_n18156,
    new_n18157, new_n18158, new_n18159, new_n18160, new_n18161, new_n18162,
    new_n18163, new_n18164, new_n18165, new_n18166, new_n18167, new_n18168,
    new_n18169, new_n18170, new_n18171, new_n18172, new_n18173, new_n18174,
    new_n18175, new_n18176, new_n18177, new_n18178, new_n18179, new_n18180,
    new_n18181, new_n18182, new_n18183, new_n18184, new_n18185, new_n18186,
    new_n18187, new_n18188, new_n18189, new_n18190, new_n18191, new_n18192,
    new_n18193, new_n18194, new_n18195, new_n18196, new_n18197, new_n18198,
    new_n18199, new_n18200, new_n18201, new_n18202, new_n18203, new_n18204,
    new_n18205, new_n18206, new_n18207, new_n18208, new_n18209, new_n18210,
    new_n18211, new_n18212, new_n18213, new_n18214, new_n18215, new_n18216,
    new_n18217, new_n18218, new_n18219, new_n18220, new_n18221, new_n18222,
    new_n18223, new_n18224, new_n18225, new_n18226, new_n18227, new_n18228,
    new_n18229, new_n18230, new_n18231, new_n18232, new_n18233, new_n18234,
    new_n18235, new_n18236, new_n18237, new_n18238, new_n18239, new_n18240,
    new_n18241, new_n18242, new_n18243, new_n18244, new_n18245, new_n18246,
    new_n18247, new_n18248, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254, new_n18255, new_n18256, new_n18257, new_n18258, new_n18259,
    new_n18260, new_n18261, new_n18262, new_n18263, new_n18264, new_n18265,
    new_n18266, new_n18267, new_n18268, new_n18269, new_n18270, new_n18271,
    new_n18272, new_n18273, new_n18274, new_n18275, new_n18276, new_n18277,
    new_n18278, new_n18279, new_n18280, new_n18281, new_n18282, new_n18283,
    new_n18284, new_n18285, new_n18286, new_n18287, new_n18288, new_n18289,
    new_n18290, new_n18291, new_n18292, new_n18293, new_n18294, new_n18295,
    new_n18296, new_n18297, new_n18298, new_n18299, new_n18300, new_n18301,
    new_n18302, new_n18303, new_n18304, new_n18305, new_n18306, new_n18307,
    new_n18308, new_n18309, new_n18310, new_n18311, new_n18312, new_n18313,
    new_n18314, new_n18315, new_n18316, new_n18317, new_n18318, new_n18319,
    new_n18320, new_n18321, new_n18322, new_n18323, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332, new_n18333, new_n18334, new_n18335, new_n18336, new_n18337,
    new_n18338, new_n18339, new_n18340, new_n18341, new_n18342, new_n18343,
    new_n18344, new_n18345, new_n18346, new_n18347, new_n18348, new_n18349,
    new_n18350, new_n18351, new_n18352, new_n18353, new_n18354, new_n18355,
    new_n18356, new_n18357, new_n18358, new_n18359, new_n18360, new_n18361,
    new_n18362, new_n18363, new_n18364, new_n18366, new_n18367, new_n18368,
    new_n18369, new_n18370, new_n18371, new_n18372, new_n18373, new_n18374,
    new_n18375, new_n18376, new_n18377, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392,
    new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18398,
    new_n18399, new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405, new_n18406, new_n18407, new_n18408, new_n18409, new_n18410,
    new_n18411, new_n18412, new_n18413, new_n18414, new_n18415, new_n18416,
    new_n18417, new_n18418, new_n18419, new_n18420, new_n18421, new_n18422,
    new_n18423, new_n18424, new_n18425, new_n18426, new_n18427, new_n18428,
    new_n18429, new_n18430, new_n18431, new_n18432, new_n18433, new_n18434,
    new_n18435, new_n18436, new_n18437, new_n18438, new_n18439, new_n18440,
    new_n18441, new_n18442, new_n18443, new_n18444, new_n18445, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18452,
    new_n18453, new_n18454, new_n18455, new_n18456, new_n18457, new_n18458,
    new_n18459, new_n18460, new_n18461, new_n18462, new_n18463, new_n18464,
    new_n18465, new_n18467, new_n18468, new_n18469, new_n18470, new_n18471,
    new_n18472, new_n18473, new_n18474, new_n18475, new_n18476, new_n18477,
    new_n18478, new_n18479, new_n18480, new_n18481, new_n18482, new_n18483,
    new_n18484, new_n18485, new_n18486, new_n18487, new_n18488, new_n18489,
    new_n18490, new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496, new_n18497, new_n18498, new_n18499, new_n18500, new_n18501,
    new_n18502, new_n18503, new_n18504, new_n18505, new_n18506, new_n18507,
    new_n18508, new_n18509, new_n18510, new_n18511, new_n18512, new_n18513,
    new_n18514, new_n18515, new_n18516, new_n18517, new_n18518, new_n18519,
    new_n18520, new_n18521, new_n18522, new_n18523, new_n18524, new_n18525,
    new_n18526, new_n18527, new_n18528, new_n18529, new_n18530, new_n18531,
    new_n18532, new_n18533, new_n18534, new_n18535, new_n18536, new_n18537,
    new_n18538, new_n18539, new_n18540, new_n18541, new_n18542, new_n18543,
    new_n18544, new_n18545, new_n18546, new_n18547, new_n18548, new_n18549,
    new_n18550, new_n18551, new_n18552, new_n18553, new_n18554, new_n18555,
    new_n18556, new_n18558, new_n18559, new_n18560, new_n18561, new_n18562,
    new_n18563, new_n18564, new_n18565, new_n18566, new_n18567, new_n18568,
    new_n18569, new_n18570, new_n18571, new_n18572, new_n18573, new_n18574,
    new_n18575, new_n18576, new_n18577, new_n18578, new_n18579, new_n18580,
    new_n18581, new_n18582, new_n18583, new_n18584, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18591, new_n18592,
    new_n18593, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598,
    new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604,
    new_n18605, new_n18606, new_n18607, new_n18608, new_n18609, new_n18610,
    new_n18611, new_n18612, new_n18613, new_n18614, new_n18615, new_n18616,
    new_n18617, new_n18618, new_n18619, new_n18620, new_n18621, new_n18622,
    new_n18623, new_n18624, new_n18625, new_n18626, new_n18627, new_n18628,
    new_n18629, new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635, new_n18636, new_n18637, new_n18638, new_n18639, new_n18640,
    new_n18641, new_n18642, new_n18643, new_n18644, new_n18645, new_n18646,
    new_n18647, new_n18648, new_n18649, new_n18650, new_n18651, new_n18652,
    new_n18653, new_n18654, new_n18656, new_n18657, new_n18658, new_n18659,
    new_n18660, new_n18661, new_n18662, new_n18663, new_n18664, new_n18665,
    new_n18666, new_n18667, new_n18668, new_n18669, new_n18670, new_n18671,
    new_n18672, new_n18673, new_n18674, new_n18675, new_n18676, new_n18677,
    new_n18678, new_n18679, new_n18680, new_n18681, new_n18682, new_n18683,
    new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18690, new_n18691, new_n18692, new_n18693, new_n18694, new_n18695,
    new_n18696, new_n18697, new_n18698, new_n18699, new_n18700, new_n18701,
    new_n18702, new_n18703, new_n18704, new_n18705, new_n18706, new_n18707,
    new_n18708, new_n18709, new_n18710, new_n18711, new_n18712, new_n18713,
    new_n18714, new_n18715, new_n18716, new_n18717, new_n18718, new_n18719,
    new_n18720, new_n18721, new_n18722, new_n18723, new_n18724, new_n18725,
    new_n18726, new_n18727, new_n18728, new_n18729, new_n18730, new_n18731,
    new_n18732, new_n18733, new_n18734, new_n18735, new_n18736, new_n18737,
    new_n18738, new_n18739, new_n18740, new_n18741, new_n18742, new_n18743,
    new_n18744, new_n18745, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843, new_n18844, new_n18845, new_n18846, new_n18847,
    new_n18848, new_n18849, new_n18850, new_n18851, new_n18852, new_n18853,
    new_n18854, new_n18855, new_n18856, new_n18857, new_n18858, new_n18859,
    new_n18860, new_n18861, new_n18862, new_n18863, new_n18864, new_n18865,
    new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871,
    new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877,
    new_n18878, new_n18879, new_n18880, new_n18881, new_n18882, new_n18883,
    new_n18884, new_n18885, new_n18886, new_n18887, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900, new_n18901,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906, new_n18907,
    new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18914,
    new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962,
    new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968,
    new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18992, new_n18993,
    new_n18994, new_n18995, new_n18996, new_n18997, new_n18998, new_n18999,
    new_n19000, new_n19001, new_n19002, new_n19003, new_n19004, new_n19005,
    new_n19006, new_n19007, new_n19008, new_n19009, new_n19010, new_n19011,
    new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017,
    new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023,
    new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033, new_n19034, new_n19035,
    new_n19036, new_n19037, new_n19038, new_n19039, new_n19040, new_n19041,
    new_n19042, new_n19043, new_n19044, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19073, new_n19074, new_n19075, new_n19076, new_n19077, new_n19078,
    new_n19079, new_n19080, new_n19081, new_n19082, new_n19083, new_n19084,
    new_n19085, new_n19086, new_n19087, new_n19088, new_n19089, new_n19090,
    new_n19091, new_n19092, new_n19093, new_n19094, new_n19095, new_n19096,
    new_n19097, new_n19098, new_n19099, new_n19100, new_n19101, new_n19102,
    new_n19103, new_n19104, new_n19105, new_n19106, new_n19107, new_n19108,
    new_n19109, new_n19110, new_n19111, new_n19112, new_n19113, new_n19114,
    new_n19115, new_n19116, new_n19117, new_n19118, new_n19119, new_n19120,
    new_n19121, new_n19122, new_n19123, new_n19124, new_n19125, new_n19126,
    new_n19127, new_n19128, new_n19129, new_n19130, new_n19131, new_n19132,
    new_n19133, new_n19134, new_n19135, new_n19136, new_n19137, new_n19138,
    new_n19139, new_n19140, new_n19141, new_n19142, new_n19143, new_n19144,
    new_n19145, new_n19147, new_n19148, new_n19149, new_n19150, new_n19151,
    new_n19152, new_n19153, new_n19154, new_n19155, new_n19156, new_n19157,
    new_n19158, new_n19159, new_n19160, new_n19161, new_n19162, new_n19163,
    new_n19164, new_n19165, new_n19166, new_n19167, new_n19168, new_n19169,
    new_n19170, new_n19171, new_n19172, new_n19173, new_n19174, new_n19175,
    new_n19176, new_n19177, new_n19178, new_n19179, new_n19180, new_n19181,
    new_n19182, new_n19183, new_n19184, new_n19185, new_n19186, new_n19187,
    new_n19188, new_n19189, new_n19190, new_n19191, new_n19192, new_n19193,
    new_n19194, new_n19195, new_n19196, new_n19197, new_n19198, new_n19199,
    new_n19200, new_n19201, new_n19202, new_n19203, new_n19204, new_n19205,
    new_n19206, new_n19207, new_n19208, new_n19209, new_n19210, new_n19211,
    new_n19212, new_n19213, new_n19214, new_n19215, new_n19216, new_n19217,
    new_n19218, new_n19220, new_n19221, new_n19222, new_n19223, new_n19224,
    new_n19225, new_n19226, new_n19227, new_n19228, new_n19229, new_n19230,
    new_n19231, new_n19232, new_n19233, new_n19234, new_n19235, new_n19236,
    new_n19237, new_n19238, new_n19239, new_n19240, new_n19241, new_n19242,
    new_n19243, new_n19244, new_n19245, new_n19246, new_n19247, new_n19248,
    new_n19249, new_n19250, new_n19251, new_n19252, new_n19253, new_n19254,
    new_n19255, new_n19256, new_n19257, new_n19258, new_n19259, new_n19260,
    new_n19261, new_n19262, new_n19263, new_n19264, new_n19265, new_n19266,
    new_n19267, new_n19268, new_n19269, new_n19270, new_n19271, new_n19272,
    new_n19273, new_n19274, new_n19275, new_n19276, new_n19277, new_n19278,
    new_n19279, new_n19280, new_n19281, new_n19283, new_n19284, new_n19285,
    new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291,
    new_n19292, new_n19293, new_n19294, new_n19295, new_n19296, new_n19297,
    new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303,
    new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309,
    new_n19310, new_n19311, new_n19312, new_n19313, new_n19314, new_n19315,
    new_n19316, new_n19317, new_n19318, new_n19319, new_n19320, new_n19321,
    new_n19322, new_n19323, new_n19324, new_n19325, new_n19326, new_n19327,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332, new_n19333,
    new_n19334, new_n19335, new_n19336, new_n19337, new_n19338, new_n19339,
    new_n19340, new_n19341, new_n19342, new_n19343, new_n19344, new_n19345,
    new_n19346, new_n19348, new_n19349, new_n19350, new_n19351, new_n19352,
    new_n19353, new_n19354, new_n19355, new_n19356, new_n19357, new_n19358,
    new_n19359, new_n19360, new_n19361, new_n19362, new_n19363, new_n19364,
    new_n19365, new_n19366, new_n19367, new_n19368, new_n19369, new_n19370,
    new_n19371, new_n19372, new_n19373, new_n19374, new_n19375, new_n19376,
    new_n19377, new_n19378, new_n19379, new_n19380, new_n19381, new_n19382,
    new_n19383, new_n19384, new_n19385, new_n19386, new_n19387, new_n19388,
    new_n19389, new_n19390, new_n19391, new_n19392, new_n19393, new_n19394,
    new_n19395, new_n19396, new_n19397, new_n19398, new_n19399, new_n19401,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414, new_n19415, new_n19416, new_n19417, new_n19418, new_n19419,
    new_n19420, new_n19421, new_n19422, new_n19423, new_n19424, new_n19425,
    new_n19426, new_n19427, new_n19428, new_n19429, new_n19430, new_n19431,
    new_n19432, new_n19433, new_n19434, new_n19435, new_n19436, new_n19437,
    new_n19438, new_n19439, new_n19440, new_n19441, new_n19442, new_n19443,
    new_n19444, new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450, new_n19451, new_n19452, new_n19453, new_n19454, new_n19455,
    new_n19457, new_n19458, new_n19459, new_n19460, new_n19461, new_n19462,
    new_n19463, new_n19464, new_n19465, new_n19466, new_n19467, new_n19468,
    new_n19469, new_n19470, new_n19471, new_n19472, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477, new_n19478, new_n19479, new_n19480,
    new_n19481, new_n19482, new_n19483, new_n19484, new_n19485, new_n19486,
    new_n19487, new_n19488, new_n19489, new_n19490, new_n19491, new_n19492,
    new_n19493, new_n19494, new_n19495, new_n19496, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19506, new_n19507, new_n19508, new_n19509, new_n19510, new_n19511,
    new_n19512, new_n19513, new_n19514, new_n19515, new_n19516, new_n19517,
    new_n19518, new_n19519, new_n19520, new_n19521, new_n19522, new_n19523,
    new_n19524, new_n19525, new_n19526, new_n19527, new_n19528, new_n19529,
    new_n19530, new_n19531, new_n19532, new_n19533, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539, new_n19540, new_n19541,
    new_n19542, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547,
    new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553,
    new_n19554, new_n19555, new_n19557, new_n19558, new_n19559, new_n19560,
    new_n19561, new_n19562, new_n19563, new_n19564, new_n19565, new_n19566,
    new_n19567, new_n19568, new_n19569, new_n19570, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575, new_n19576, new_n19577, new_n19578,
    new_n19579, new_n19580, new_n19581, new_n19582, new_n19583, new_n19584,
    new_n19585, new_n19586, new_n19587, new_n19588, new_n19589, new_n19590,
    new_n19591, new_n19592, new_n19593, new_n19594, new_n19595, new_n19596,
    new_n19597, new_n19598, new_n19600, new_n19601, new_n19602, new_n19603,
    new_n19604, new_n19605, new_n19606, new_n19607, new_n19608, new_n19609,
    new_n19610, new_n19611, new_n19612, new_n19613, new_n19614, new_n19615,
    new_n19616, new_n19617, new_n19618, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623, new_n19624, new_n19625, new_n19626, new_n19627,
    new_n19628, new_n19629, new_n19630, new_n19631, new_n19632, new_n19633,
    new_n19634, new_n19635, new_n19636, new_n19637, new_n19638, new_n19639,
    new_n19640, new_n19641, new_n19642, new_n19643, new_n19645, new_n19646,
    new_n19647, new_n19648, new_n19649, new_n19650, new_n19651, new_n19652,
    new_n19653, new_n19654, new_n19655, new_n19656, new_n19657, new_n19658,
    new_n19659, new_n19660, new_n19661, new_n19662, new_n19663, new_n19664,
    new_n19665, new_n19666, new_n19667, new_n19668, new_n19669, new_n19670,
    new_n19671, new_n19672, new_n19674, new_n19675, new_n19676, new_n19677,
    new_n19678, new_n19679, new_n19680, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700, new_n19701,
    new_n19702, new_n19703, new_n19704, new_n19705, new_n19707, new_n19708,
    new_n19709, new_n19710, new_n19711, new_n19712, new_n19713, new_n19714,
    new_n19715, new_n19716, new_n19717, new_n19718, new_n19719, new_n19720,
    new_n19721, new_n19722, new_n19723, new_n19724, new_n19725, new_n19726,
    new_n19727, new_n19728, new_n19729, new_n19730, new_n19731, new_n19732,
    new_n19733, new_n19734, new_n19735, new_n19736, new_n19737, new_n19738,
    new_n19739, new_n19740, new_n19741, new_n19743, new_n19744, new_n19745,
    new_n19746, new_n19747, new_n19748, new_n19749, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756, new_n19757,
    new_n19758, new_n19759, new_n19760, new_n19761, new_n19762, new_n19763,
    new_n19764, new_n19766, new_n19767, new_n19768, new_n19769, new_n19770,
    new_n19771, new_n19772, new_n19773, new_n19774, new_n19775, new_n19776,
    new_n19777, new_n19778, new_n19779, new_n19780, new_n19781, new_n19782,
    new_n19784, new_n19785, new_n19786, new_n19787, new_n19788, new_n19789,
    new_n19790, new_n19791, new_n19792;
  INVx1_ASAP7_75t_L         g00000(.A(\a[0] ), .Y(new_n257));
  INVx1_ASAP7_75t_L         g00001(.A(\b[0] ), .Y(new_n258));
  NOR2xp33_ASAP7_75t_L      g00002(.A(new_n257), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00003(.A(\a[2] ), .B(\f[0] ), .Y(new_n260));
  INVx1_ASAP7_75t_L         g00004(.A(\b[1] ), .Y(new_n261));
  INVx1_ASAP7_75t_L         g00005(.A(\a[2] ), .Y(new_n262));
  NOR2xp33_ASAP7_75t_L      g00006(.A(\a[1] ), .B(new_n262), .Y(new_n263));
  INVx1_ASAP7_75t_L         g00007(.A(\a[1] ), .Y(new_n264));
  NOR2xp33_ASAP7_75t_L      g00008(.A(\a[2] ), .B(new_n264), .Y(new_n265));
  NOR2xp33_ASAP7_75t_L      g00009(.A(new_n263), .B(new_n265), .Y(new_n266));
  NOR2xp33_ASAP7_75t_L      g00010(.A(new_n257), .B(new_n266), .Y(new_n267));
  INVx1_ASAP7_75t_L         g00011(.A(new_n267), .Y(new_n268));
  XOR2x2_ASAP7_75t_L        g00012(.A(\b[1] ), .B(\b[0] ), .Y(new_n269));
  INVx1_ASAP7_75t_L         g00013(.A(new_n269), .Y(new_n270));
  NAND2xp33_ASAP7_75t_L     g00014(.A(\a[0] ), .B(new_n266), .Y(new_n271));
  NOR2xp33_ASAP7_75t_L      g00015(.A(\a[0] ), .B(new_n264), .Y(new_n272));
  NAND2xp33_ASAP7_75t_L     g00016(.A(\b[0] ), .B(new_n272), .Y(new_n273));
  OAI221xp5_ASAP7_75t_L     g00017(.A1(new_n271), .A2(new_n261), .B1(new_n270), .B2(new_n268), .C(new_n273), .Y(new_n274));
  XNOR2x2_ASAP7_75t_L       g00018(.A(new_n260), .B(new_n274), .Y(\f[1] ));
  INVx1_ASAP7_75t_L         g00019(.A(\b[2] ), .Y(new_n276));
  NAND3xp33_ASAP7_75t_L     g00020(.A(new_n276), .B(\b[1] ), .C(\b[0] ), .Y(new_n277));
  NAND2xp33_ASAP7_75t_L     g00021(.A(\b[1] ), .B(\b[0] ), .Y(new_n278));
  OAI21xp33_ASAP7_75t_L     g00022(.A1(\b[1] ), .A2(new_n276), .B(new_n278), .Y(new_n279));
  A2O1A1Ixp33_ASAP7_75t_L   g00023(.A1(\b[1] ), .A2(new_n276), .B(new_n279), .C(new_n277), .Y(new_n280));
  INVx1_ASAP7_75t_L         g00024(.A(new_n280), .Y(new_n281));
  NOR3xp33_ASAP7_75t_L      g00025(.A(new_n262), .B(\a[1] ), .C(\a[0] ), .Y(new_n282));
  INVx1_ASAP7_75t_L         g00026(.A(new_n282), .Y(new_n283));
  OAI22xp33_ASAP7_75t_L     g00027(.A1(new_n271), .A2(new_n276), .B1(new_n258), .B2(new_n283), .Y(new_n284));
  AOI221xp5_ASAP7_75t_L     g00028(.A1(new_n267), .A2(new_n281), .B1(new_n272), .B2(\b[1] ), .C(new_n284), .Y(new_n285));
  INVx1_ASAP7_75t_L         g00029(.A(new_n285), .Y(new_n286));
  O2A1O1Ixp33_ASAP7_75t_L   g00030(.A1(\f[0] ), .A2(new_n274), .B(\a[2] ), .C(new_n286), .Y(new_n287));
  A2O1A1Ixp33_ASAP7_75t_L   g00031(.A1(\a[0] ), .A2(\b[0] ), .B(new_n274), .C(\a[2] ), .Y(new_n288));
  NOR2xp33_ASAP7_75t_L      g00032(.A(new_n285), .B(new_n288), .Y(new_n289));
  NOR2xp33_ASAP7_75t_L      g00033(.A(new_n289), .B(new_n287), .Y(\f[2] ));
  INVx1_ASAP7_75t_L         g00034(.A(new_n272), .Y(new_n291));
  NOR2xp33_ASAP7_75t_L      g00035(.A(\b[2] ), .B(new_n278), .Y(new_n292));
  NOR2xp33_ASAP7_75t_L      g00036(.A(\b[2] ), .B(\b[3] ), .Y(new_n293));
  NAND2xp33_ASAP7_75t_L     g00037(.A(\b[3] ), .B(\b[2] ), .Y(new_n294));
  INVx1_ASAP7_75t_L         g00038(.A(new_n294), .Y(new_n295));
  NOR2xp33_ASAP7_75t_L      g00039(.A(new_n293), .B(new_n295), .Y(new_n296));
  A2O1A1Ixp33_ASAP7_75t_L   g00040(.A1(\b[2] ), .A2(\b[1] ), .B(new_n292), .C(new_n296), .Y(new_n297));
  INVx1_ASAP7_75t_L         g00041(.A(\b[3] ), .Y(new_n298));
  NAND2xp33_ASAP7_75t_L     g00042(.A(new_n298), .B(new_n276), .Y(new_n299));
  NAND2xp33_ASAP7_75t_L     g00043(.A(new_n294), .B(new_n299), .Y(new_n300));
  A2O1A1Ixp33_ASAP7_75t_L   g00044(.A1(new_n276), .A2(new_n258), .B(new_n261), .C(new_n300), .Y(new_n301));
  NAND2xp33_ASAP7_75t_L     g00045(.A(new_n301), .B(new_n297), .Y(new_n302));
  INVx1_ASAP7_75t_L         g00046(.A(new_n271), .Y(new_n303));
  AOI22xp33_ASAP7_75t_L     g00047(.A1(\b[1] ), .A2(new_n282), .B1(\b[3] ), .B2(new_n303), .Y(new_n304));
  OAI221xp5_ASAP7_75t_L     g00048(.A1(new_n291), .A2(new_n276), .B1(new_n268), .B2(new_n302), .C(new_n304), .Y(new_n305));
  XNOR2x2_ASAP7_75t_L       g00049(.A(\a[2] ), .B(new_n305), .Y(new_n306));
  INVx1_ASAP7_75t_L         g00050(.A(new_n306), .Y(new_n307));
  INVx1_ASAP7_75t_L         g00051(.A(\a[3] ), .Y(new_n308));
  NAND2xp33_ASAP7_75t_L     g00052(.A(\a[2] ), .B(new_n308), .Y(new_n309));
  NAND2xp33_ASAP7_75t_L     g00053(.A(\a[3] ), .B(new_n262), .Y(new_n310));
  NAND2xp33_ASAP7_75t_L     g00054(.A(new_n310), .B(new_n309), .Y(new_n311));
  NAND2xp33_ASAP7_75t_L     g00055(.A(\b[0] ), .B(new_n311), .Y(new_n312));
  INVx1_ASAP7_75t_L         g00056(.A(new_n312), .Y(new_n313));
  NAND2xp33_ASAP7_75t_L     g00057(.A(new_n313), .B(new_n307), .Y(new_n314));
  A2O1A1Ixp33_ASAP7_75t_L   g00058(.A1(new_n309), .A2(new_n310), .B(new_n258), .C(new_n306), .Y(new_n315));
  NAND2xp33_ASAP7_75t_L     g00059(.A(new_n315), .B(new_n314), .Y(new_n316));
  NOR3xp33_ASAP7_75t_L      g00060(.A(new_n274), .B(\f[0] ), .C(new_n262), .Y(new_n317));
  NAND2xp33_ASAP7_75t_L     g00061(.A(new_n285), .B(new_n317), .Y(new_n318));
  XOR2x2_ASAP7_75t_L        g00062(.A(new_n318), .B(new_n316), .Y(\f[3] ));
  OAI21xp33_ASAP7_75t_L     g00063(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n320));
  OAI21xp33_ASAP7_75t_L     g00064(.A1(new_n293), .A2(new_n320), .B(new_n294), .Y(new_n321));
  INVx1_ASAP7_75t_L         g00065(.A(new_n321), .Y(new_n322));
  NOR2xp33_ASAP7_75t_L      g00066(.A(\b[3] ), .B(\b[4] ), .Y(new_n323));
  INVx1_ASAP7_75t_L         g00067(.A(\b[4] ), .Y(new_n324));
  NOR2xp33_ASAP7_75t_L      g00068(.A(new_n298), .B(new_n324), .Y(new_n325));
  NOR3xp33_ASAP7_75t_L      g00069(.A(new_n322), .B(new_n323), .C(new_n325), .Y(new_n326));
  NOR2xp33_ASAP7_75t_L      g00070(.A(new_n323), .B(new_n325), .Y(new_n327));
  NOR2xp33_ASAP7_75t_L      g00071(.A(new_n321), .B(new_n327), .Y(new_n328));
  NOR2xp33_ASAP7_75t_L      g00072(.A(new_n328), .B(new_n326), .Y(new_n329));
  INVx1_ASAP7_75t_L         g00073(.A(new_n329), .Y(new_n330));
  AOI22xp33_ASAP7_75t_L     g00074(.A1(\b[2] ), .A2(new_n282), .B1(\b[4] ), .B2(new_n303), .Y(new_n331));
  OAI221xp5_ASAP7_75t_L     g00075(.A1(new_n291), .A2(new_n298), .B1(new_n268), .B2(new_n330), .C(new_n331), .Y(new_n332));
  XNOR2x2_ASAP7_75t_L       g00076(.A(new_n262), .B(new_n332), .Y(new_n333));
  NAND2xp33_ASAP7_75t_L     g00077(.A(\a[5] ), .B(new_n313), .Y(new_n334));
  INVx1_ASAP7_75t_L         g00078(.A(new_n311), .Y(new_n335));
  INVx1_ASAP7_75t_L         g00079(.A(\a[4] ), .Y(new_n336));
  NAND2xp33_ASAP7_75t_L     g00080(.A(\a[5] ), .B(new_n336), .Y(new_n337));
  INVx1_ASAP7_75t_L         g00081(.A(\a[5] ), .Y(new_n338));
  NAND2xp33_ASAP7_75t_L     g00082(.A(\a[4] ), .B(new_n338), .Y(new_n339));
  AND2x2_ASAP7_75t_L        g00083(.A(new_n337), .B(new_n339), .Y(new_n340));
  NOR2xp33_ASAP7_75t_L      g00084(.A(new_n340), .B(new_n335), .Y(new_n341));
  NAND2xp33_ASAP7_75t_L     g00085(.A(new_n269), .B(new_n341), .Y(new_n342));
  NAND2xp33_ASAP7_75t_L     g00086(.A(new_n311), .B(new_n340), .Y(new_n343));
  INVx1_ASAP7_75t_L         g00087(.A(new_n343), .Y(new_n344));
  NAND2xp33_ASAP7_75t_L     g00088(.A(\b[1] ), .B(new_n344), .Y(new_n345));
  XNOR2x2_ASAP7_75t_L       g00089(.A(\a[4] ), .B(\a[3] ), .Y(new_n346));
  NOR2xp33_ASAP7_75t_L      g00090(.A(new_n346), .B(new_n311), .Y(new_n347));
  NAND2xp33_ASAP7_75t_L     g00091(.A(\b[0] ), .B(new_n347), .Y(new_n348));
  NAND3xp33_ASAP7_75t_L     g00092(.A(new_n345), .B(new_n342), .C(new_n348), .Y(new_n349));
  XNOR2x2_ASAP7_75t_L       g00093(.A(new_n334), .B(new_n349), .Y(new_n350));
  XNOR2x2_ASAP7_75t_L       g00094(.A(new_n350), .B(new_n333), .Y(new_n351));
  MAJIxp5_ASAP7_75t_L       g00095(.A(new_n306), .B(new_n312), .C(new_n318), .Y(new_n352));
  XNOR2x2_ASAP7_75t_L       g00096(.A(new_n352), .B(new_n351), .Y(\f[4] ));
  INVx1_ASAP7_75t_L         g00097(.A(\b[5] ), .Y(new_n354));
  XOR2x2_ASAP7_75t_L        g00098(.A(\b[5] ), .B(\b[4] ), .Y(new_n355));
  A2O1A1Ixp33_ASAP7_75t_L   g00099(.A1(new_n327), .A2(new_n321), .B(new_n325), .C(new_n355), .Y(new_n356));
  INVx1_ASAP7_75t_L         g00100(.A(new_n356), .Y(new_n357));
  AOI211xp5_ASAP7_75t_L     g00101(.A1(new_n327), .A2(new_n321), .B(new_n355), .C(new_n325), .Y(new_n358));
  NOR2xp33_ASAP7_75t_L      g00102(.A(new_n358), .B(new_n357), .Y(new_n359));
  NAND2xp33_ASAP7_75t_L     g00103(.A(new_n267), .B(new_n359), .Y(new_n360));
  OAI221xp5_ASAP7_75t_L     g00104(.A1(new_n271), .A2(new_n354), .B1(new_n298), .B2(new_n283), .C(new_n360), .Y(new_n361));
  AOI21xp33_ASAP7_75t_L     g00105(.A1(new_n272), .A2(\b[4] ), .B(new_n361), .Y(new_n362));
  NAND2xp33_ASAP7_75t_L     g00106(.A(\a[2] ), .B(new_n362), .Y(new_n363));
  A2O1A1Ixp33_ASAP7_75t_L   g00107(.A1(\b[4] ), .A2(new_n272), .B(new_n361), .C(new_n262), .Y(new_n364));
  AND2x2_ASAP7_75t_L        g00108(.A(new_n364), .B(new_n363), .Y(new_n365));
  INVx1_ASAP7_75t_L         g00109(.A(new_n341), .Y(new_n366));
  A2O1A1Ixp33_ASAP7_75t_L   g00110(.A1(\b[0] ), .A2(new_n311), .B(new_n349), .C(\a[5] ), .Y(new_n367));
  NOR2xp33_ASAP7_75t_L      g00111(.A(new_n276), .B(new_n343), .Y(new_n368));
  NAND2xp33_ASAP7_75t_L     g00112(.A(new_n339), .B(new_n337), .Y(new_n369));
  AND3x1_ASAP7_75t_L        g00113(.A(new_n335), .B(new_n346), .C(new_n369), .Y(new_n370));
  AOI221xp5_ASAP7_75t_L     g00114(.A1(new_n347), .A2(\b[1] ), .B1(new_n370), .B2(\b[0] ), .C(new_n368), .Y(new_n371));
  O2A1O1Ixp33_ASAP7_75t_L   g00115(.A1(new_n366), .A2(new_n280), .B(new_n371), .C(new_n367), .Y(new_n372));
  A2O1A1Ixp33_ASAP7_75t_L   g00116(.A1(new_n309), .A2(new_n310), .B(new_n258), .C(\a[5] ), .Y(new_n373));
  OAI21xp33_ASAP7_75t_L     g00117(.A1(new_n280), .A2(new_n366), .B(new_n371), .Y(new_n374));
  O2A1O1Ixp33_ASAP7_75t_L   g00118(.A1(new_n349), .A2(new_n373), .B(\a[5] ), .C(new_n374), .Y(new_n375));
  OR2x4_ASAP7_75t_L         g00119(.A(new_n375), .B(new_n372), .Y(new_n376));
  XNOR2x2_ASAP7_75t_L       g00120(.A(new_n376), .B(new_n365), .Y(new_n377));
  MAJIxp5_ASAP7_75t_L       g00121(.A(new_n352), .B(new_n350), .C(new_n333), .Y(new_n378));
  XOR2x2_ASAP7_75t_L        g00122(.A(new_n378), .B(new_n377), .Y(\f[5] ));
  MAJIxp5_ASAP7_75t_L       g00123(.A(new_n365), .B(new_n376), .C(new_n378), .Y(new_n380));
  INVx1_ASAP7_75t_L         g00124(.A(new_n380), .Y(new_n381));
  NOR2xp33_ASAP7_75t_L      g00125(.A(\b[5] ), .B(\b[6] ), .Y(new_n382));
  NAND2xp33_ASAP7_75t_L     g00126(.A(\b[6] ), .B(\b[5] ), .Y(new_n383));
  INVx1_ASAP7_75t_L         g00127(.A(new_n383), .Y(new_n384));
  NOR2xp33_ASAP7_75t_L      g00128(.A(new_n382), .B(new_n384), .Y(new_n385));
  INVx1_ASAP7_75t_L         g00129(.A(new_n385), .Y(new_n386));
  O2A1O1Ixp33_ASAP7_75t_L   g00130(.A1(new_n324), .A2(new_n354), .B(new_n356), .C(new_n386), .Y(new_n387));
  NAND2xp33_ASAP7_75t_L     g00131(.A(\b[5] ), .B(\b[4] ), .Y(new_n388));
  AND3x1_ASAP7_75t_L        g00132(.A(new_n356), .B(new_n386), .C(new_n388), .Y(new_n389));
  OR2x4_ASAP7_75t_L         g00133(.A(new_n387), .B(new_n389), .Y(new_n390));
  AOI22xp33_ASAP7_75t_L     g00134(.A1(\b[4] ), .A2(new_n282), .B1(\b[6] ), .B2(new_n303), .Y(new_n391));
  OAI221xp5_ASAP7_75t_L     g00135(.A1(new_n291), .A2(new_n354), .B1(new_n268), .B2(new_n390), .C(new_n391), .Y(new_n392));
  XNOR2x2_ASAP7_75t_L       g00136(.A(\a[2] ), .B(new_n392), .Y(new_n393));
  INVx1_ASAP7_75t_L         g00137(.A(\a[6] ), .Y(new_n394));
  NAND2xp33_ASAP7_75t_L     g00138(.A(\a[5] ), .B(new_n394), .Y(new_n395));
  NAND2xp33_ASAP7_75t_L     g00139(.A(\a[6] ), .B(new_n338), .Y(new_n396));
  NOR3xp33_ASAP7_75t_L      g00140(.A(new_n374), .B(new_n373), .C(new_n349), .Y(new_n397));
  A2O1A1Ixp33_ASAP7_75t_L   g00141(.A1(new_n395), .A2(new_n396), .B(new_n258), .C(new_n397), .Y(new_n398));
  NAND2xp33_ASAP7_75t_L     g00142(.A(new_n396), .B(new_n395), .Y(new_n399));
  NAND2xp33_ASAP7_75t_L     g00143(.A(\b[0] ), .B(new_n399), .Y(new_n400));
  INVx1_ASAP7_75t_L         g00144(.A(new_n400), .Y(new_n401));
  OAI31xp33_ASAP7_75t_L     g00145(.A1(new_n374), .A2(new_n349), .A3(new_n373), .B(new_n401), .Y(new_n402));
  NAND2xp33_ASAP7_75t_L     g00146(.A(new_n402), .B(new_n398), .Y(new_n403));
  O2A1O1Ixp33_ASAP7_75t_L   g00147(.A1(new_n261), .A2(new_n276), .B(new_n277), .C(new_n300), .Y(new_n404));
  O2A1O1Ixp33_ASAP7_75t_L   g00148(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n296), .Y(new_n405));
  NOR2xp33_ASAP7_75t_L      g00149(.A(new_n404), .B(new_n405), .Y(new_n406));
  NAND3xp33_ASAP7_75t_L     g00150(.A(new_n335), .B(new_n369), .C(new_n346), .Y(new_n407));
  OAI22xp33_ASAP7_75t_L     g00151(.A1(new_n407), .A2(new_n261), .B1(new_n298), .B2(new_n343), .Y(new_n408));
  AOI221xp5_ASAP7_75t_L     g00152(.A1(\b[2] ), .A2(new_n347), .B1(new_n406), .B2(new_n341), .C(new_n408), .Y(new_n409));
  XNOR2x2_ASAP7_75t_L       g00153(.A(\a[5] ), .B(new_n409), .Y(new_n410));
  XNOR2x2_ASAP7_75t_L       g00154(.A(new_n410), .B(new_n403), .Y(new_n411));
  XNOR2x2_ASAP7_75t_L       g00155(.A(new_n393), .B(new_n411), .Y(new_n412));
  NOR2xp33_ASAP7_75t_L      g00156(.A(new_n381), .B(new_n412), .Y(new_n413));
  AND2x2_ASAP7_75t_L        g00157(.A(new_n381), .B(new_n412), .Y(new_n414));
  NOR2xp33_ASAP7_75t_L      g00158(.A(new_n413), .B(new_n414), .Y(\f[6] ));
  NOR2xp33_ASAP7_75t_L      g00159(.A(new_n393), .B(new_n411), .Y(new_n416));
  NOR2xp33_ASAP7_75t_L      g00160(.A(new_n416), .B(new_n413), .Y(new_n417));
  INVx1_ASAP7_75t_L         g00161(.A(\b[6] ), .Y(new_n418));
  A2O1A1Ixp33_ASAP7_75t_L   g00162(.A1(new_n356), .A2(new_n388), .B(new_n382), .C(new_n383), .Y(new_n419));
  INVx1_ASAP7_75t_L         g00163(.A(\b[7] ), .Y(new_n420));
  NAND2xp33_ASAP7_75t_L     g00164(.A(new_n420), .B(new_n418), .Y(new_n421));
  NAND2xp33_ASAP7_75t_L     g00165(.A(\b[7] ), .B(\b[6] ), .Y(new_n422));
  NAND2xp33_ASAP7_75t_L     g00166(.A(new_n422), .B(new_n421), .Y(new_n423));
  INVx1_ASAP7_75t_L         g00167(.A(new_n423), .Y(new_n424));
  XNOR2x2_ASAP7_75t_L       g00168(.A(new_n424), .B(new_n419), .Y(new_n425));
  AOI22xp33_ASAP7_75t_L     g00169(.A1(\b[5] ), .A2(new_n282), .B1(\b[7] ), .B2(new_n303), .Y(new_n426));
  OAI221xp5_ASAP7_75t_L     g00170(.A1(new_n291), .A2(new_n418), .B1(new_n268), .B2(new_n425), .C(new_n426), .Y(new_n427));
  XNOR2x2_ASAP7_75t_L       g00171(.A(\a[2] ), .B(new_n427), .Y(new_n428));
  INVx1_ASAP7_75t_L         g00172(.A(new_n347), .Y(new_n429));
  NOR2xp33_ASAP7_75t_L      g00173(.A(new_n298), .B(new_n429), .Y(new_n430));
  NAND2xp33_ASAP7_75t_L     g00174(.A(\b[2] ), .B(new_n370), .Y(new_n431));
  OAI221xp5_ASAP7_75t_L     g00175(.A1(new_n343), .A2(new_n324), .B1(new_n366), .B2(new_n330), .C(new_n431), .Y(new_n432));
  NOR3xp33_ASAP7_75t_L      g00176(.A(new_n432), .B(new_n430), .C(new_n338), .Y(new_n433));
  OA21x2_ASAP7_75t_L        g00177(.A1(new_n430), .A2(new_n432), .B(new_n338), .Y(new_n434));
  INVx1_ASAP7_75t_L         g00178(.A(\a[8] ), .Y(new_n435));
  NOR2xp33_ASAP7_75t_L      g00179(.A(new_n435), .B(new_n400), .Y(new_n436));
  AND2x2_ASAP7_75t_L        g00180(.A(new_n395), .B(new_n396), .Y(new_n437));
  INVx1_ASAP7_75t_L         g00181(.A(\a[7] ), .Y(new_n438));
  NAND2xp33_ASAP7_75t_L     g00182(.A(\a[8] ), .B(new_n438), .Y(new_n439));
  NAND2xp33_ASAP7_75t_L     g00183(.A(\a[7] ), .B(new_n435), .Y(new_n440));
  AOI21xp33_ASAP7_75t_L     g00184(.A1(new_n440), .A2(new_n439), .B(new_n437), .Y(new_n441));
  NAND2xp33_ASAP7_75t_L     g00185(.A(new_n269), .B(new_n441), .Y(new_n442));
  NAND2xp33_ASAP7_75t_L     g00186(.A(new_n440), .B(new_n439), .Y(new_n443));
  NOR2xp33_ASAP7_75t_L      g00187(.A(new_n443), .B(new_n437), .Y(new_n444));
  NAND2xp33_ASAP7_75t_L     g00188(.A(\b[1] ), .B(new_n444), .Y(new_n445));
  XNOR2x2_ASAP7_75t_L       g00189(.A(\a[7] ), .B(\a[6] ), .Y(new_n446));
  NOR2xp33_ASAP7_75t_L      g00190(.A(new_n446), .B(new_n399), .Y(new_n447));
  NAND2xp33_ASAP7_75t_L     g00191(.A(\b[0] ), .B(new_n447), .Y(new_n448));
  NAND3xp33_ASAP7_75t_L     g00192(.A(new_n442), .B(new_n445), .C(new_n448), .Y(new_n449));
  XNOR2x2_ASAP7_75t_L       g00193(.A(new_n436), .B(new_n449), .Y(new_n450));
  OR3x1_ASAP7_75t_L         g00194(.A(new_n434), .B(new_n433), .C(new_n450), .Y(new_n451));
  OAI21xp33_ASAP7_75t_L     g00195(.A1(new_n433), .A2(new_n434), .B(new_n450), .Y(new_n452));
  MAJIxp5_ASAP7_75t_L       g00196(.A(new_n410), .B(new_n401), .C(new_n397), .Y(new_n453));
  AOI21xp33_ASAP7_75t_L     g00197(.A1(new_n451), .A2(new_n452), .B(new_n453), .Y(new_n454));
  AND3x1_ASAP7_75t_L        g00198(.A(new_n451), .B(new_n453), .C(new_n452), .Y(new_n455));
  NOR3xp33_ASAP7_75t_L      g00199(.A(new_n455), .B(new_n454), .C(new_n428), .Y(new_n456));
  INVx1_ASAP7_75t_L         g00200(.A(new_n456), .Y(new_n457));
  OAI21xp33_ASAP7_75t_L     g00201(.A1(new_n454), .A2(new_n455), .B(new_n428), .Y(new_n458));
  NAND2xp33_ASAP7_75t_L     g00202(.A(new_n458), .B(new_n457), .Y(new_n459));
  XOR2x2_ASAP7_75t_L        g00203(.A(new_n459), .B(new_n417), .Y(\f[7] ));
  NAND2xp33_ASAP7_75t_L     g00204(.A(\b[4] ), .B(new_n347), .Y(new_n461));
  NAND2xp33_ASAP7_75t_L     g00205(.A(\b[5] ), .B(new_n344), .Y(new_n462));
  AOI22xp33_ASAP7_75t_L     g00206(.A1(\b[3] ), .A2(new_n370), .B1(new_n341), .B2(new_n359), .Y(new_n463));
  NAND4xp25_ASAP7_75t_L     g00207(.A(new_n463), .B(\a[5] ), .C(new_n461), .D(new_n462), .Y(new_n464));
  NAND2xp33_ASAP7_75t_L     g00208(.A(new_n462), .B(new_n463), .Y(new_n465));
  A2O1A1Ixp33_ASAP7_75t_L   g00209(.A1(\b[4] ), .A2(new_n347), .B(new_n465), .C(new_n338), .Y(new_n466));
  NAND2xp33_ASAP7_75t_L     g00210(.A(new_n464), .B(new_n466), .Y(new_n467));
  INVx1_ASAP7_75t_L         g00211(.A(new_n447), .Y(new_n468));
  NAND2xp33_ASAP7_75t_L     g00212(.A(new_n443), .B(new_n399), .Y(new_n469));
  NOR2xp33_ASAP7_75t_L      g00213(.A(new_n280), .B(new_n469), .Y(new_n470));
  AND3x1_ASAP7_75t_L        g00214(.A(new_n437), .B(new_n446), .C(new_n443), .Y(new_n471));
  AOI221xp5_ASAP7_75t_L     g00215(.A1(new_n444), .A2(\b[2] ), .B1(new_n471), .B2(\b[0] ), .C(new_n470), .Y(new_n472));
  OAI21xp33_ASAP7_75t_L     g00216(.A1(new_n261), .A2(new_n468), .B(new_n472), .Y(new_n473));
  O2A1O1Ixp33_ASAP7_75t_L   g00217(.A1(new_n401), .A2(new_n449), .B(\a[8] ), .C(new_n473), .Y(new_n474));
  A2O1A1Ixp33_ASAP7_75t_L   g00218(.A1(\b[0] ), .A2(new_n399), .B(new_n449), .C(\a[8] ), .Y(new_n475));
  O2A1O1Ixp33_ASAP7_75t_L   g00219(.A1(new_n468), .A2(new_n261), .B(new_n472), .C(new_n475), .Y(new_n476));
  NOR2xp33_ASAP7_75t_L      g00220(.A(new_n474), .B(new_n476), .Y(new_n477));
  INVx1_ASAP7_75t_L         g00221(.A(new_n477), .Y(new_n478));
  NOR2xp33_ASAP7_75t_L      g00222(.A(new_n467), .B(new_n478), .Y(new_n479));
  AOI21xp33_ASAP7_75t_L     g00223(.A1(new_n464), .A2(new_n466), .B(new_n477), .Y(new_n480));
  NOR2xp33_ASAP7_75t_L      g00224(.A(new_n433), .B(new_n434), .Y(new_n481));
  MAJIxp5_ASAP7_75t_L       g00225(.A(new_n453), .B(new_n450), .C(new_n481), .Y(new_n482));
  NOR3xp33_ASAP7_75t_L      g00226(.A(new_n482), .B(new_n480), .C(new_n479), .Y(new_n483));
  OA21x2_ASAP7_75t_L        g00227(.A1(new_n480), .A2(new_n479), .B(new_n482), .Y(new_n484));
  OR2x4_ASAP7_75t_L         g00228(.A(new_n483), .B(new_n484), .Y(new_n485));
  INVx1_ASAP7_75t_L         g00229(.A(new_n422), .Y(new_n486));
  NOR2xp33_ASAP7_75t_L      g00230(.A(\b[7] ), .B(\b[8] ), .Y(new_n487));
  INVx1_ASAP7_75t_L         g00231(.A(\b[8] ), .Y(new_n488));
  NOR2xp33_ASAP7_75t_L      g00232(.A(new_n420), .B(new_n488), .Y(new_n489));
  NOR2xp33_ASAP7_75t_L      g00233(.A(new_n487), .B(new_n489), .Y(new_n490));
  A2O1A1Ixp33_ASAP7_75t_L   g00234(.A1(new_n419), .A2(new_n424), .B(new_n486), .C(new_n490), .Y(new_n491));
  A2O1A1O1Ixp25_ASAP7_75t_L g00235(.A1(new_n388), .A2(new_n356), .B(new_n382), .C(new_n383), .D(new_n423), .Y(new_n492));
  OR3x1_ASAP7_75t_L         g00236(.A(new_n492), .B(new_n486), .C(new_n490), .Y(new_n493));
  NAND2xp33_ASAP7_75t_L     g00237(.A(new_n491), .B(new_n493), .Y(new_n494));
  AOI22xp33_ASAP7_75t_L     g00238(.A1(\b[6] ), .A2(new_n282), .B1(\b[8] ), .B2(new_n303), .Y(new_n495));
  OAI221xp5_ASAP7_75t_L     g00239(.A1(new_n291), .A2(new_n420), .B1(new_n268), .B2(new_n494), .C(new_n495), .Y(new_n496));
  XNOR2x2_ASAP7_75t_L       g00240(.A(\a[2] ), .B(new_n496), .Y(new_n497));
  XNOR2x2_ASAP7_75t_L       g00241(.A(new_n497), .B(new_n485), .Y(new_n498));
  O2A1O1Ixp33_ASAP7_75t_L   g00242(.A1(new_n459), .A2(new_n417), .B(new_n457), .C(new_n498), .Y(new_n499));
  NAND2xp33_ASAP7_75t_L     g00243(.A(new_n393), .B(new_n411), .Y(new_n500));
  A2O1A1O1Ixp25_ASAP7_75t_L g00244(.A1(new_n380), .A2(new_n500), .B(new_n416), .C(new_n458), .D(new_n456), .Y(new_n501));
  AND2x2_ASAP7_75t_L        g00245(.A(new_n501), .B(new_n498), .Y(new_n502));
  NOR2xp33_ASAP7_75t_L      g00246(.A(new_n502), .B(new_n499), .Y(\f[8] ));
  NAND5xp2_ASAP7_75t_L      g00247(.A(\a[8] ), .B(new_n442), .C(new_n445), .D(new_n448), .E(new_n400), .Y(new_n504));
  INVx1_ASAP7_75t_L         g00248(.A(\a[9] ), .Y(new_n505));
  NAND2xp33_ASAP7_75t_L     g00249(.A(\a[8] ), .B(new_n505), .Y(new_n506));
  NAND2xp33_ASAP7_75t_L     g00250(.A(\a[9] ), .B(new_n435), .Y(new_n507));
  AND2x2_ASAP7_75t_L        g00251(.A(new_n506), .B(new_n507), .Y(new_n508));
  NOR2xp33_ASAP7_75t_L      g00252(.A(new_n258), .B(new_n508), .Y(new_n509));
  OAI21xp33_ASAP7_75t_L     g00253(.A1(new_n504), .A2(new_n473), .B(new_n509), .Y(new_n510));
  INVx1_ASAP7_75t_L         g00254(.A(new_n504), .Y(new_n511));
  NAND2xp33_ASAP7_75t_L     g00255(.A(\b[1] ), .B(new_n447), .Y(new_n512));
  INVx1_ASAP7_75t_L         g00256(.A(new_n509), .Y(new_n513));
  NAND4xp25_ASAP7_75t_L     g00257(.A(new_n511), .B(new_n513), .C(new_n472), .D(new_n512), .Y(new_n514));
  NAND3xp33_ASAP7_75t_L     g00258(.A(new_n399), .B(new_n439), .C(new_n440), .Y(new_n515));
  NAND3xp33_ASAP7_75t_L     g00259(.A(new_n437), .B(new_n443), .C(new_n446), .Y(new_n516));
  OAI22xp33_ASAP7_75t_L     g00260(.A1(new_n516), .A2(new_n261), .B1(new_n298), .B2(new_n515), .Y(new_n517));
  AOI221xp5_ASAP7_75t_L     g00261(.A1(\b[2] ), .A2(new_n447), .B1(new_n406), .B2(new_n441), .C(new_n517), .Y(new_n518));
  XNOR2x2_ASAP7_75t_L       g00262(.A(new_n435), .B(new_n518), .Y(new_n519));
  AOI21xp33_ASAP7_75t_L     g00263(.A1(new_n514), .A2(new_n510), .B(new_n519), .Y(new_n520));
  INVx1_ASAP7_75t_L         g00264(.A(new_n520), .Y(new_n521));
  NAND3xp33_ASAP7_75t_L     g00265(.A(new_n519), .B(new_n514), .C(new_n510), .Y(new_n522));
  NOR2xp33_ASAP7_75t_L      g00266(.A(new_n354), .B(new_n429), .Y(new_n523));
  INVx1_ASAP7_75t_L         g00267(.A(new_n523), .Y(new_n524));
  NAND2xp33_ASAP7_75t_L     g00268(.A(\b[6] ), .B(new_n344), .Y(new_n525));
  NOR2xp33_ASAP7_75t_L      g00269(.A(new_n387), .B(new_n389), .Y(new_n526));
  AOI22xp33_ASAP7_75t_L     g00270(.A1(new_n370), .A2(\b[4] ), .B1(new_n341), .B2(new_n526), .Y(new_n527));
  AND4x1_ASAP7_75t_L        g00271(.A(new_n527), .B(new_n525), .C(new_n524), .D(\a[5] ), .Y(new_n528));
  AOI31xp33_ASAP7_75t_L     g00272(.A1(new_n527), .A2(new_n525), .A3(new_n524), .B(\a[5] ), .Y(new_n529));
  NOR2xp33_ASAP7_75t_L      g00273(.A(new_n529), .B(new_n528), .Y(new_n530));
  NAND3xp33_ASAP7_75t_L     g00274(.A(new_n521), .B(new_n522), .C(new_n530), .Y(new_n531));
  AO21x2_ASAP7_75t_L        g00275(.A1(new_n522), .A2(new_n521), .B(new_n530), .Y(new_n532));
  AND2x2_ASAP7_75t_L        g00276(.A(new_n531), .B(new_n532), .Y(new_n533));
  AOI21xp33_ASAP7_75t_L     g00277(.A1(new_n466), .A2(new_n464), .B(new_n478), .Y(new_n534));
  O2A1O1Ixp33_ASAP7_75t_L   g00278(.A1(new_n480), .A2(new_n479), .B(new_n482), .C(new_n534), .Y(new_n535));
  NAND2xp33_ASAP7_75t_L     g00279(.A(new_n535), .B(new_n533), .Y(new_n536));
  NAND2xp33_ASAP7_75t_L     g00280(.A(new_n531), .B(new_n532), .Y(new_n537));
  A2O1A1Ixp33_ASAP7_75t_L   g00281(.A1(new_n477), .A2(new_n467), .B(new_n484), .C(new_n537), .Y(new_n538));
  NOR2xp33_ASAP7_75t_L      g00282(.A(\b[8] ), .B(\b[9] ), .Y(new_n539));
  INVx1_ASAP7_75t_L         g00283(.A(\b[9] ), .Y(new_n540));
  NOR2xp33_ASAP7_75t_L      g00284(.A(new_n488), .B(new_n540), .Y(new_n541));
  NOR2xp33_ASAP7_75t_L      g00285(.A(new_n539), .B(new_n541), .Y(new_n542));
  INVx1_ASAP7_75t_L         g00286(.A(new_n542), .Y(new_n543));
  O2A1O1Ixp33_ASAP7_75t_L   g00287(.A1(new_n420), .A2(new_n488), .B(new_n491), .C(new_n543), .Y(new_n544));
  INVx1_ASAP7_75t_L         g00288(.A(new_n544), .Y(new_n545));
  A2O1A1O1Ixp25_ASAP7_75t_L g00289(.A1(new_n424), .A2(new_n419), .B(new_n486), .C(new_n490), .D(new_n489), .Y(new_n546));
  NAND2xp33_ASAP7_75t_L     g00290(.A(new_n543), .B(new_n546), .Y(new_n547));
  NAND2xp33_ASAP7_75t_L     g00291(.A(new_n547), .B(new_n545), .Y(new_n548));
  AOI22xp33_ASAP7_75t_L     g00292(.A1(\b[7] ), .A2(new_n282), .B1(\b[9] ), .B2(new_n303), .Y(new_n549));
  OAI221xp5_ASAP7_75t_L     g00293(.A1(new_n291), .A2(new_n488), .B1(new_n268), .B2(new_n548), .C(new_n549), .Y(new_n550));
  XNOR2x2_ASAP7_75t_L       g00294(.A(\a[2] ), .B(new_n550), .Y(new_n551));
  NAND3xp33_ASAP7_75t_L     g00295(.A(new_n536), .B(new_n538), .C(new_n551), .Y(new_n552));
  NOR3xp33_ASAP7_75t_L      g00296(.A(new_n537), .B(new_n484), .C(new_n534), .Y(new_n553));
  NOR2xp33_ASAP7_75t_L      g00297(.A(new_n535), .B(new_n533), .Y(new_n554));
  INVx1_ASAP7_75t_L         g00298(.A(new_n551), .Y(new_n555));
  OAI21xp33_ASAP7_75t_L     g00299(.A1(new_n553), .A2(new_n554), .B(new_n555), .Y(new_n556));
  NAND2xp33_ASAP7_75t_L     g00300(.A(new_n552), .B(new_n556), .Y(new_n557));
  MAJIxp5_ASAP7_75t_L       g00301(.A(new_n501), .B(new_n485), .C(new_n497), .Y(new_n558));
  XOR2x2_ASAP7_75t_L        g00302(.A(new_n557), .B(new_n558), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g00303(.A(new_n497), .B(new_n485), .Y(new_n560));
  NOR3xp33_ASAP7_75t_L      g00304(.A(new_n554), .B(new_n553), .C(new_n551), .Y(new_n561));
  O2A1O1Ixp33_ASAP7_75t_L   g00305(.A1(new_n560), .A2(new_n499), .B(new_n557), .C(new_n561), .Y(new_n562));
  NOR3xp33_ASAP7_75t_L      g00306(.A(new_n473), .B(new_n513), .C(new_n504), .Y(new_n563));
  NAND2xp33_ASAP7_75t_L     g00307(.A(\b[3] ), .B(new_n447), .Y(new_n564));
  AOI22xp33_ASAP7_75t_L     g00308(.A1(new_n444), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n471), .Y(new_n565));
  OA211x2_ASAP7_75t_L       g00309(.A1(new_n469), .A2(new_n330), .B(new_n565), .C(new_n564), .Y(new_n566));
  NAND2xp33_ASAP7_75t_L     g00310(.A(\a[8] ), .B(new_n566), .Y(new_n567));
  OAI211xp5_ASAP7_75t_L     g00311(.A1(new_n469), .A2(new_n330), .B(new_n564), .C(new_n565), .Y(new_n568));
  NAND2xp33_ASAP7_75t_L     g00312(.A(new_n435), .B(new_n568), .Y(new_n569));
  NAND2xp33_ASAP7_75t_L     g00313(.A(\a[11] ), .B(new_n509), .Y(new_n570));
  NAND2xp33_ASAP7_75t_L     g00314(.A(new_n507), .B(new_n506), .Y(new_n571));
  INVx1_ASAP7_75t_L         g00315(.A(\a[10] ), .Y(new_n572));
  NAND2xp33_ASAP7_75t_L     g00316(.A(\a[11] ), .B(new_n572), .Y(new_n573));
  INVx1_ASAP7_75t_L         g00317(.A(\a[11] ), .Y(new_n574));
  NAND2xp33_ASAP7_75t_L     g00318(.A(\a[10] ), .B(new_n574), .Y(new_n575));
  NAND2xp33_ASAP7_75t_L     g00319(.A(new_n575), .B(new_n573), .Y(new_n576));
  NAND2xp33_ASAP7_75t_L     g00320(.A(new_n576), .B(new_n571), .Y(new_n577));
  INVx1_ASAP7_75t_L         g00321(.A(new_n577), .Y(new_n578));
  NAND2xp33_ASAP7_75t_L     g00322(.A(new_n269), .B(new_n578), .Y(new_n579));
  NAND3xp33_ASAP7_75t_L     g00323(.A(new_n571), .B(new_n573), .C(new_n575), .Y(new_n580));
  INVx1_ASAP7_75t_L         g00324(.A(new_n580), .Y(new_n581));
  NAND2xp33_ASAP7_75t_L     g00325(.A(\b[1] ), .B(new_n581), .Y(new_n582));
  XNOR2x2_ASAP7_75t_L       g00326(.A(\a[10] ), .B(\a[9] ), .Y(new_n583));
  NOR2xp33_ASAP7_75t_L      g00327(.A(new_n583), .B(new_n571), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(\b[0] ), .B(new_n584), .Y(new_n585));
  NAND3xp33_ASAP7_75t_L     g00329(.A(new_n582), .B(new_n579), .C(new_n585), .Y(new_n586));
  XOR2x2_ASAP7_75t_L        g00330(.A(new_n570), .B(new_n586), .Y(new_n587));
  NAND3xp33_ASAP7_75t_L     g00331(.A(new_n567), .B(new_n587), .C(new_n569), .Y(new_n588));
  NOR2xp33_ASAP7_75t_L      g00332(.A(new_n435), .B(new_n568), .Y(new_n589));
  NOR2xp33_ASAP7_75t_L      g00333(.A(\a[8] ), .B(new_n566), .Y(new_n590));
  XNOR2x2_ASAP7_75t_L       g00334(.A(new_n570), .B(new_n586), .Y(new_n591));
  OAI21xp33_ASAP7_75t_L     g00335(.A1(new_n589), .A2(new_n590), .B(new_n591), .Y(new_n592));
  OAI211xp5_ASAP7_75t_L     g00336(.A1(new_n563), .A2(new_n520), .B(new_n588), .C(new_n592), .Y(new_n593));
  NOR2xp33_ASAP7_75t_L      g00337(.A(new_n504), .B(new_n473), .Y(new_n594));
  XNOR2x2_ASAP7_75t_L       g00338(.A(\a[8] ), .B(new_n518), .Y(new_n595));
  MAJIxp5_ASAP7_75t_L       g00339(.A(new_n595), .B(new_n509), .C(new_n594), .Y(new_n596));
  NOR3xp33_ASAP7_75t_L      g00340(.A(new_n590), .B(new_n591), .C(new_n589), .Y(new_n597));
  AOI21xp33_ASAP7_75t_L     g00341(.A1(new_n567), .A2(new_n569), .B(new_n587), .Y(new_n598));
  OAI21xp33_ASAP7_75t_L     g00342(.A1(new_n598), .A2(new_n597), .B(new_n596), .Y(new_n599));
  NAND2xp33_ASAP7_75t_L     g00343(.A(\b[7] ), .B(new_n344), .Y(new_n600));
  OAI221xp5_ASAP7_75t_L     g00344(.A1(new_n407), .A2(new_n354), .B1(new_n366), .B2(new_n425), .C(new_n600), .Y(new_n601));
  AOI21xp33_ASAP7_75t_L     g00345(.A1(new_n347), .A2(\b[6] ), .B(new_n601), .Y(new_n602));
  NAND2xp33_ASAP7_75t_L     g00346(.A(\a[5] ), .B(new_n602), .Y(new_n603));
  A2O1A1Ixp33_ASAP7_75t_L   g00347(.A1(\b[6] ), .A2(new_n347), .B(new_n601), .C(new_n338), .Y(new_n604));
  NAND4xp25_ASAP7_75t_L     g00348(.A(new_n593), .B(new_n604), .C(new_n603), .D(new_n599), .Y(new_n605));
  NAND2xp33_ASAP7_75t_L     g00349(.A(new_n599), .B(new_n593), .Y(new_n606));
  NAND2xp33_ASAP7_75t_L     g00350(.A(new_n604), .B(new_n603), .Y(new_n607));
  NAND2xp33_ASAP7_75t_L     g00351(.A(new_n607), .B(new_n606), .Y(new_n608));
  NAND2xp33_ASAP7_75t_L     g00352(.A(new_n605), .B(new_n608), .Y(new_n609));
  OAI211xp5_ASAP7_75t_L     g00353(.A1(new_n528), .A2(new_n529), .B(new_n521), .C(new_n522), .Y(new_n610));
  A2O1A1Ixp33_ASAP7_75t_L   g00354(.A1(new_n532), .A2(new_n531), .B(new_n535), .C(new_n610), .Y(new_n611));
  NOR2xp33_ASAP7_75t_L      g00355(.A(new_n611), .B(new_n609), .Y(new_n612));
  AOI22xp33_ASAP7_75t_L     g00356(.A1(new_n605), .A2(new_n608), .B1(new_n610), .B2(new_n538), .Y(new_n613));
  INVx1_ASAP7_75t_L         g00357(.A(new_n489), .Y(new_n614));
  INVx1_ASAP7_75t_L         g00358(.A(new_n541), .Y(new_n615));
  NOR2xp33_ASAP7_75t_L      g00359(.A(\b[9] ), .B(\b[10] ), .Y(new_n616));
  INVx1_ASAP7_75t_L         g00360(.A(\b[10] ), .Y(new_n617));
  NOR2xp33_ASAP7_75t_L      g00361(.A(new_n540), .B(new_n617), .Y(new_n618));
  NOR2xp33_ASAP7_75t_L      g00362(.A(new_n616), .B(new_n618), .Y(new_n619));
  INVx1_ASAP7_75t_L         g00363(.A(new_n619), .Y(new_n620));
  A2O1A1O1Ixp25_ASAP7_75t_L g00364(.A1(new_n614), .A2(new_n491), .B(new_n539), .C(new_n615), .D(new_n620), .Y(new_n621));
  INVx1_ASAP7_75t_L         g00365(.A(new_n621), .Y(new_n622));
  OAI211xp5_ASAP7_75t_L     g00366(.A1(new_n543), .A2(new_n546), .B(new_n615), .C(new_n620), .Y(new_n623));
  NAND2xp33_ASAP7_75t_L     g00367(.A(new_n623), .B(new_n622), .Y(new_n624));
  AOI22xp33_ASAP7_75t_L     g00368(.A1(\b[8] ), .A2(new_n282), .B1(\b[10] ), .B2(new_n303), .Y(new_n625));
  OAI221xp5_ASAP7_75t_L     g00369(.A1(new_n291), .A2(new_n540), .B1(new_n268), .B2(new_n624), .C(new_n625), .Y(new_n626));
  XNOR2x2_ASAP7_75t_L       g00370(.A(\a[2] ), .B(new_n626), .Y(new_n627));
  OAI21xp33_ASAP7_75t_L     g00371(.A1(new_n612), .A2(new_n613), .B(new_n627), .Y(new_n628));
  NOR3xp33_ASAP7_75t_L      g00372(.A(new_n613), .B(new_n627), .C(new_n612), .Y(new_n629));
  INVx1_ASAP7_75t_L         g00373(.A(new_n629), .Y(new_n630));
  NAND2xp33_ASAP7_75t_L     g00374(.A(new_n628), .B(new_n630), .Y(new_n631));
  XOR2x2_ASAP7_75t_L        g00375(.A(new_n631), .B(new_n562), .Y(\f[10] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g00376(.A1(new_n557), .A2(new_n558), .B(new_n561), .C(new_n628), .D(new_n629), .Y(new_n633));
  AOI21xp33_ASAP7_75t_L     g00377(.A1(new_n604), .A2(new_n603), .B(new_n606), .Y(new_n634));
  NAND2xp33_ASAP7_75t_L     g00378(.A(\b[8] ), .B(new_n344), .Y(new_n635));
  OAI221xp5_ASAP7_75t_L     g00379(.A1(new_n407), .A2(new_n418), .B1(new_n366), .B2(new_n494), .C(new_n635), .Y(new_n636));
  AOI211xp5_ASAP7_75t_L     g00380(.A1(\b[7] ), .A2(new_n347), .B(new_n338), .C(new_n636), .Y(new_n637));
  A2O1A1Ixp33_ASAP7_75t_L   g00381(.A1(\b[7] ), .A2(new_n347), .B(new_n636), .C(new_n338), .Y(new_n638));
  INVx1_ASAP7_75t_L         g00382(.A(new_n638), .Y(new_n639));
  NAND2xp33_ASAP7_75t_L     g00383(.A(new_n510), .B(new_n514), .Y(new_n640));
  A2O1A1O1Ixp25_ASAP7_75t_L g00384(.A1(new_n595), .A2(new_n640), .B(new_n563), .C(new_n588), .D(new_n598), .Y(new_n641));
  NAND2xp33_ASAP7_75t_L     g00385(.A(\b[4] ), .B(new_n447), .Y(new_n642));
  INVx1_ASAP7_75t_L         g00386(.A(new_n642), .Y(new_n643));
  NOR3xp33_ASAP7_75t_L      g00387(.A(new_n357), .B(new_n358), .C(new_n469), .Y(new_n644));
  OAI22xp33_ASAP7_75t_L     g00388(.A1(new_n516), .A2(new_n298), .B1(new_n354), .B2(new_n515), .Y(new_n645));
  NOR4xp25_ASAP7_75t_L      g00389(.A(new_n644), .B(new_n435), .C(new_n645), .D(new_n643), .Y(new_n646));
  INVx1_ASAP7_75t_L         g00390(.A(new_n646), .Y(new_n647));
  OAI31xp33_ASAP7_75t_L     g00391(.A1(new_n644), .A2(new_n643), .A3(new_n645), .B(new_n435), .Y(new_n648));
  NAND2xp33_ASAP7_75t_L     g00392(.A(\b[1] ), .B(new_n584), .Y(new_n649));
  NOR2xp33_ASAP7_75t_L      g00393(.A(new_n280), .B(new_n577), .Y(new_n650));
  AND3x1_ASAP7_75t_L        g00394(.A(new_n508), .B(new_n583), .C(new_n576), .Y(new_n651));
  AOI221xp5_ASAP7_75t_L     g00395(.A1(new_n651), .A2(\b[0] ), .B1(\b[2] ), .B2(new_n581), .C(new_n650), .Y(new_n652));
  NAND2xp33_ASAP7_75t_L     g00396(.A(new_n649), .B(new_n652), .Y(new_n653));
  O2A1O1Ixp33_ASAP7_75t_L   g00397(.A1(new_n509), .A2(new_n586), .B(\a[11] ), .C(new_n653), .Y(new_n654));
  INVx1_ASAP7_75t_L         g00398(.A(new_n654), .Y(new_n655));
  NAND5xp2_ASAP7_75t_L      g00399(.A(\a[11] ), .B(new_n582), .C(new_n579), .D(new_n585), .E(new_n513), .Y(new_n656));
  NAND3xp33_ASAP7_75t_L     g00400(.A(new_n653), .B(new_n656), .C(\a[11] ), .Y(new_n657));
  NAND4xp25_ASAP7_75t_L     g00401(.A(new_n657), .B(new_n647), .C(new_n648), .D(new_n655), .Y(new_n658));
  NAND2xp33_ASAP7_75t_L     g00402(.A(new_n648), .B(new_n647), .Y(new_n659));
  INVx1_ASAP7_75t_L         g00403(.A(new_n657), .Y(new_n660));
  OAI21xp33_ASAP7_75t_L     g00404(.A1(new_n654), .A2(new_n660), .B(new_n659), .Y(new_n661));
  AOI21xp33_ASAP7_75t_L     g00405(.A1(new_n661), .A2(new_n658), .B(new_n641), .Y(new_n662));
  OAI21xp33_ASAP7_75t_L     g00406(.A1(new_n597), .A2(new_n596), .B(new_n592), .Y(new_n663));
  NAND2xp33_ASAP7_75t_L     g00407(.A(new_n661), .B(new_n658), .Y(new_n664));
  NOR2xp33_ASAP7_75t_L      g00408(.A(new_n663), .B(new_n664), .Y(new_n665));
  OAI22xp33_ASAP7_75t_L     g00409(.A1(new_n665), .A2(new_n662), .B1(new_n639), .B2(new_n637), .Y(new_n666));
  INVx1_ASAP7_75t_L         g00410(.A(new_n637), .Y(new_n667));
  NAND2xp33_ASAP7_75t_L     g00411(.A(new_n663), .B(new_n664), .Y(new_n668));
  NAND3xp33_ASAP7_75t_L     g00412(.A(new_n641), .B(new_n658), .C(new_n661), .Y(new_n669));
  NAND4xp25_ASAP7_75t_L     g00413(.A(new_n669), .B(new_n668), .C(new_n667), .D(new_n638), .Y(new_n670));
  NAND2xp33_ASAP7_75t_L     g00414(.A(new_n670), .B(new_n666), .Y(new_n671));
  INVx1_ASAP7_75t_L         g00415(.A(new_n671), .Y(new_n672));
  A2O1A1Ixp33_ASAP7_75t_L   g00416(.A1(new_n611), .A2(new_n609), .B(new_n634), .C(new_n672), .Y(new_n673));
  AOI21xp33_ASAP7_75t_L     g00417(.A1(new_n609), .A2(new_n611), .B(new_n634), .Y(new_n674));
  NAND2xp33_ASAP7_75t_L     g00418(.A(new_n671), .B(new_n674), .Y(new_n675));
  NAND2xp33_ASAP7_75t_L     g00419(.A(new_n675), .B(new_n673), .Y(new_n676));
  A2O1A1Ixp33_ASAP7_75t_L   g00420(.A1(new_n491), .A2(new_n614), .B(new_n539), .C(new_n615), .Y(new_n677));
  NOR2xp33_ASAP7_75t_L      g00421(.A(\b[10] ), .B(\b[11] ), .Y(new_n678));
  INVx1_ASAP7_75t_L         g00422(.A(\b[11] ), .Y(new_n679));
  NOR2xp33_ASAP7_75t_L      g00423(.A(new_n617), .B(new_n679), .Y(new_n680));
  NOR2xp33_ASAP7_75t_L      g00424(.A(new_n678), .B(new_n680), .Y(new_n681));
  A2O1A1Ixp33_ASAP7_75t_L   g00425(.A1(new_n677), .A2(new_n619), .B(new_n618), .C(new_n681), .Y(new_n682));
  O2A1O1Ixp33_ASAP7_75t_L   g00426(.A1(new_n541), .A2(new_n544), .B(new_n619), .C(new_n618), .Y(new_n683));
  OAI21xp33_ASAP7_75t_L     g00427(.A1(new_n678), .A2(new_n680), .B(new_n683), .Y(new_n684));
  NAND2xp33_ASAP7_75t_L     g00428(.A(new_n682), .B(new_n684), .Y(new_n685));
  AOI22xp33_ASAP7_75t_L     g00429(.A1(\b[9] ), .A2(new_n282), .B1(\b[11] ), .B2(new_n303), .Y(new_n686));
  OAI221xp5_ASAP7_75t_L     g00430(.A1(new_n291), .A2(new_n617), .B1(new_n268), .B2(new_n685), .C(new_n686), .Y(new_n687));
  XNOR2x2_ASAP7_75t_L       g00431(.A(new_n262), .B(new_n687), .Y(new_n688));
  NAND2xp33_ASAP7_75t_L     g00432(.A(new_n688), .B(new_n676), .Y(new_n689));
  INVx1_ASAP7_75t_L         g00433(.A(new_n689), .Y(new_n690));
  INVx1_ASAP7_75t_L         g00434(.A(new_n688), .Y(new_n691));
  AND3x1_ASAP7_75t_L        g00435(.A(new_n673), .B(new_n691), .C(new_n675), .Y(new_n692));
  NOR2xp33_ASAP7_75t_L      g00436(.A(new_n692), .B(new_n690), .Y(new_n693));
  XNOR2x2_ASAP7_75t_L       g00437(.A(new_n633), .B(new_n693), .Y(\f[11] ));
  INVx1_ASAP7_75t_L         g00438(.A(\a[12] ), .Y(new_n695));
  NAND2xp33_ASAP7_75t_L     g00439(.A(\a[11] ), .B(new_n695), .Y(new_n696));
  NAND2xp33_ASAP7_75t_L     g00440(.A(\a[12] ), .B(new_n574), .Y(new_n697));
  AND2x2_ASAP7_75t_L        g00441(.A(new_n696), .B(new_n697), .Y(new_n698));
  NOR2xp33_ASAP7_75t_L      g00442(.A(new_n258), .B(new_n698), .Y(new_n699));
  OAI21xp33_ASAP7_75t_L     g00443(.A1(new_n656), .A2(new_n653), .B(new_n699), .Y(new_n700));
  OAI21xp33_ASAP7_75t_L     g00444(.A1(new_n261), .A2(new_n580), .B(new_n585), .Y(new_n701));
  A2O1A1Ixp33_ASAP7_75t_L   g00445(.A1(new_n506), .A2(new_n507), .B(new_n258), .C(\a[11] ), .Y(new_n702));
  AOI211xp5_ASAP7_75t_L     g00446(.A1(new_n578), .A2(new_n269), .B(new_n702), .C(new_n701), .Y(new_n703));
  INVx1_ASAP7_75t_L         g00447(.A(new_n699), .Y(new_n704));
  NAND4xp25_ASAP7_75t_L     g00448(.A(new_n703), .B(new_n704), .C(new_n652), .D(new_n649), .Y(new_n705));
  NAND3xp33_ASAP7_75t_L     g00449(.A(new_n508), .B(new_n576), .C(new_n583), .Y(new_n706));
  OAI22xp33_ASAP7_75t_L     g00450(.A1(new_n706), .A2(new_n261), .B1(new_n298), .B2(new_n580), .Y(new_n707));
  AOI221xp5_ASAP7_75t_L     g00451(.A1(\b[2] ), .A2(new_n584), .B1(new_n406), .B2(new_n578), .C(new_n707), .Y(new_n708));
  XNOR2x2_ASAP7_75t_L       g00452(.A(new_n574), .B(new_n708), .Y(new_n709));
  AOI21xp33_ASAP7_75t_L     g00453(.A1(new_n705), .A2(new_n700), .B(new_n709), .Y(new_n710));
  NAND2xp33_ASAP7_75t_L     g00454(.A(\a[11] ), .B(new_n708), .Y(new_n711));
  AO21x2_ASAP7_75t_L        g00455(.A1(new_n406), .A2(new_n578), .B(new_n707), .Y(new_n712));
  A2O1A1Ixp33_ASAP7_75t_L   g00456(.A1(\b[2] ), .A2(new_n584), .B(new_n712), .C(new_n574), .Y(new_n713));
  AND4x1_ASAP7_75t_L        g00457(.A(new_n700), .B(new_n713), .C(new_n705), .D(new_n711), .Y(new_n714));
  NOR2xp33_ASAP7_75t_L      g00458(.A(new_n354), .B(new_n468), .Y(new_n715));
  INVx1_ASAP7_75t_L         g00459(.A(new_n715), .Y(new_n716));
  NAND2xp33_ASAP7_75t_L     g00460(.A(new_n441), .B(new_n526), .Y(new_n717));
  AOI22xp33_ASAP7_75t_L     g00461(.A1(new_n444), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n471), .Y(new_n718));
  NAND4xp25_ASAP7_75t_L     g00462(.A(new_n717), .B(\a[8] ), .C(new_n716), .D(new_n718), .Y(new_n719));
  INVx1_ASAP7_75t_L         g00463(.A(new_n719), .Y(new_n720));
  AOI31xp33_ASAP7_75t_L     g00464(.A1(new_n717), .A2(new_n716), .A3(new_n718), .B(\a[8] ), .Y(new_n721));
  NOR4xp25_ASAP7_75t_L      g00465(.A(new_n710), .B(new_n720), .C(new_n714), .D(new_n721), .Y(new_n722));
  AO22x1_ASAP7_75t_L        g00466(.A1(new_n713), .A2(new_n711), .B1(new_n705), .B2(new_n700), .Y(new_n723));
  NAND3xp33_ASAP7_75t_L     g00467(.A(new_n709), .B(new_n705), .C(new_n700), .Y(new_n724));
  INVx1_ASAP7_75t_L         g00468(.A(new_n721), .Y(new_n725));
  AOI22xp33_ASAP7_75t_L     g00469(.A1(new_n719), .A2(new_n725), .B1(new_n723), .B2(new_n724), .Y(new_n726));
  NOR2xp33_ASAP7_75t_L      g00470(.A(new_n726), .B(new_n722), .Y(new_n727));
  NOR2xp33_ASAP7_75t_L      g00471(.A(new_n654), .B(new_n660), .Y(new_n728));
  MAJIxp5_ASAP7_75t_L       g00472(.A(new_n663), .B(new_n659), .C(new_n728), .Y(new_n729));
  XNOR2x2_ASAP7_75t_L       g00473(.A(new_n727), .B(new_n729), .Y(new_n730));
  AND2x2_ASAP7_75t_L        g00474(.A(new_n547), .B(new_n545), .Y(new_n731));
  NOR2xp33_ASAP7_75t_L      g00475(.A(new_n420), .B(new_n407), .Y(new_n732));
  AOI221xp5_ASAP7_75t_L     g00476(.A1(\b[9] ), .A2(new_n344), .B1(new_n341), .B2(new_n731), .C(new_n732), .Y(new_n733));
  OAI211xp5_ASAP7_75t_L     g00477(.A1(new_n488), .A2(new_n429), .B(new_n733), .C(\a[5] ), .Y(new_n734));
  INVx1_ASAP7_75t_L         g00478(.A(new_n734), .Y(new_n735));
  O2A1O1Ixp33_ASAP7_75t_L   g00479(.A1(new_n488), .A2(new_n429), .B(new_n733), .C(\a[5] ), .Y(new_n736));
  NOR2xp33_ASAP7_75t_L      g00480(.A(new_n736), .B(new_n735), .Y(new_n737));
  NAND2xp33_ASAP7_75t_L     g00481(.A(new_n730), .B(new_n737), .Y(new_n738));
  OR2x4_ASAP7_75t_L         g00482(.A(new_n726), .B(new_n722), .Y(new_n739));
  NAND2xp33_ASAP7_75t_L     g00483(.A(new_n659), .B(new_n728), .Y(new_n740));
  A2O1A1Ixp33_ASAP7_75t_L   g00484(.A1(new_n658), .A2(new_n661), .B(new_n641), .C(new_n740), .Y(new_n741));
  NOR2xp33_ASAP7_75t_L      g00485(.A(new_n741), .B(new_n739), .Y(new_n742));
  A2O1A1O1Ixp25_ASAP7_75t_L g00486(.A1(new_n658), .A2(new_n661), .B(new_n641), .C(new_n740), .D(new_n727), .Y(new_n743));
  NOR2xp33_ASAP7_75t_L      g00487(.A(new_n743), .B(new_n742), .Y(new_n744));
  INVx1_ASAP7_75t_L         g00488(.A(new_n736), .Y(new_n745));
  NAND2xp33_ASAP7_75t_L     g00489(.A(new_n734), .B(new_n745), .Y(new_n746));
  NAND2xp33_ASAP7_75t_L     g00490(.A(new_n746), .B(new_n744), .Y(new_n747));
  NAND2xp33_ASAP7_75t_L     g00491(.A(new_n738), .B(new_n747), .Y(new_n748));
  NOR2xp33_ASAP7_75t_L      g00492(.A(new_n637), .B(new_n639), .Y(new_n749));
  NAND2xp33_ASAP7_75t_L     g00493(.A(new_n668), .B(new_n669), .Y(new_n750));
  NOR2xp33_ASAP7_75t_L      g00494(.A(new_n749), .B(new_n750), .Y(new_n751));
  A2O1A1O1Ixp25_ASAP7_75t_L g00495(.A1(new_n611), .A2(new_n609), .B(new_n634), .C(new_n671), .D(new_n751), .Y(new_n752));
  NOR2xp33_ASAP7_75t_L      g00496(.A(new_n752), .B(new_n748), .Y(new_n753));
  NOR2xp33_ASAP7_75t_L      g00497(.A(new_n746), .B(new_n744), .Y(new_n754));
  NOR2xp33_ASAP7_75t_L      g00498(.A(new_n730), .B(new_n737), .Y(new_n755));
  NOR2xp33_ASAP7_75t_L      g00499(.A(new_n755), .B(new_n754), .Y(new_n756));
  INVx1_ASAP7_75t_L         g00500(.A(new_n752), .Y(new_n757));
  NOR2xp33_ASAP7_75t_L      g00501(.A(new_n757), .B(new_n756), .Y(new_n758));
  NOR2xp33_ASAP7_75t_L      g00502(.A(\b[11] ), .B(\b[12] ), .Y(new_n759));
  INVx1_ASAP7_75t_L         g00503(.A(\b[12] ), .Y(new_n760));
  NOR2xp33_ASAP7_75t_L      g00504(.A(new_n679), .B(new_n760), .Y(new_n761));
  NOR2xp33_ASAP7_75t_L      g00505(.A(new_n759), .B(new_n761), .Y(new_n762));
  INVx1_ASAP7_75t_L         g00506(.A(new_n762), .Y(new_n763));
  O2A1O1Ixp33_ASAP7_75t_L   g00507(.A1(new_n617), .A2(new_n679), .B(new_n682), .C(new_n763), .Y(new_n764));
  INVx1_ASAP7_75t_L         g00508(.A(new_n764), .Y(new_n765));
  A2O1A1O1Ixp25_ASAP7_75t_L g00509(.A1(new_n619), .A2(new_n677), .B(new_n618), .C(new_n681), .D(new_n680), .Y(new_n766));
  NAND2xp33_ASAP7_75t_L     g00510(.A(new_n763), .B(new_n766), .Y(new_n767));
  NAND2xp33_ASAP7_75t_L     g00511(.A(new_n767), .B(new_n765), .Y(new_n768));
  AOI22xp33_ASAP7_75t_L     g00512(.A1(\b[10] ), .A2(new_n282), .B1(\b[12] ), .B2(new_n303), .Y(new_n769));
  OAI221xp5_ASAP7_75t_L     g00513(.A1(new_n291), .A2(new_n679), .B1(new_n268), .B2(new_n768), .C(new_n769), .Y(new_n770));
  XNOR2x2_ASAP7_75t_L       g00514(.A(\a[2] ), .B(new_n770), .Y(new_n771));
  INVx1_ASAP7_75t_L         g00515(.A(new_n771), .Y(new_n772));
  NOR3xp33_ASAP7_75t_L      g00516(.A(new_n758), .B(new_n753), .C(new_n772), .Y(new_n773));
  NAND2xp33_ASAP7_75t_L     g00517(.A(new_n757), .B(new_n756), .Y(new_n774));
  NAND2xp33_ASAP7_75t_L     g00518(.A(new_n752), .B(new_n748), .Y(new_n775));
  AOI21xp33_ASAP7_75t_L     g00519(.A1(new_n774), .A2(new_n775), .B(new_n771), .Y(new_n776));
  OAI21xp33_ASAP7_75t_L     g00520(.A1(new_n692), .A2(new_n633), .B(new_n689), .Y(new_n777));
  OAI21xp33_ASAP7_75t_L     g00521(.A1(new_n773), .A2(new_n776), .B(new_n777), .Y(new_n778));
  INVx1_ASAP7_75t_L         g00522(.A(new_n778), .Y(new_n779));
  NOR3xp33_ASAP7_75t_L      g00523(.A(new_n777), .B(new_n776), .C(new_n773), .Y(new_n780));
  NOR2xp33_ASAP7_75t_L      g00524(.A(new_n780), .B(new_n779), .Y(\f[12] ));
  NOR2xp33_ASAP7_75t_L      g00525(.A(new_n753), .B(new_n758), .Y(new_n782));
  NOR2xp33_ASAP7_75t_L      g00526(.A(\b[12] ), .B(\b[13] ), .Y(new_n783));
  INVx1_ASAP7_75t_L         g00527(.A(\b[13] ), .Y(new_n784));
  NOR2xp33_ASAP7_75t_L      g00528(.A(new_n760), .B(new_n784), .Y(new_n785));
  NOR2xp33_ASAP7_75t_L      g00529(.A(new_n783), .B(new_n785), .Y(new_n786));
  A2O1A1Ixp33_ASAP7_75t_L   g00530(.A1(\b[12] ), .A2(\b[11] ), .B(new_n764), .C(new_n786), .Y(new_n787));
  INVx1_ASAP7_75t_L         g00531(.A(new_n761), .Y(new_n788));
  OAI221xp5_ASAP7_75t_L     g00532(.A1(new_n785), .A2(new_n783), .B1(new_n759), .B2(new_n766), .C(new_n788), .Y(new_n789));
  NAND2xp33_ASAP7_75t_L     g00533(.A(new_n789), .B(new_n787), .Y(new_n790));
  AOI22xp33_ASAP7_75t_L     g00534(.A1(\b[11] ), .A2(new_n282), .B1(\b[13] ), .B2(new_n303), .Y(new_n791));
  OAI221xp5_ASAP7_75t_L     g00535(.A1(new_n291), .A2(new_n760), .B1(new_n268), .B2(new_n790), .C(new_n791), .Y(new_n792));
  XNOR2x2_ASAP7_75t_L       g00536(.A(\a[2] ), .B(new_n792), .Y(new_n793));
  NOR2xp33_ASAP7_75t_L      g00537(.A(new_n656), .B(new_n653), .Y(new_n794));
  NAND2xp33_ASAP7_75t_L     g00538(.A(new_n699), .B(new_n794), .Y(new_n795));
  A2O1A1Ixp33_ASAP7_75t_L   g00539(.A1(new_n705), .A2(new_n700), .B(new_n709), .C(new_n795), .Y(new_n796));
  NAND2xp33_ASAP7_75t_L     g00540(.A(\b[3] ), .B(new_n584), .Y(new_n797));
  AOI22xp33_ASAP7_75t_L     g00541(.A1(\b[2] ), .A2(new_n651), .B1(\b[4] ), .B2(new_n581), .Y(new_n798));
  OA21x2_ASAP7_75t_L        g00542(.A1(new_n577), .A2(new_n330), .B(new_n798), .Y(new_n799));
  NAND3xp33_ASAP7_75t_L     g00543(.A(new_n799), .B(new_n797), .C(\a[11] ), .Y(new_n800));
  OAI211xp5_ASAP7_75t_L     g00544(.A1(new_n577), .A2(new_n330), .B(new_n797), .C(new_n798), .Y(new_n801));
  NAND2xp33_ASAP7_75t_L     g00545(.A(new_n574), .B(new_n801), .Y(new_n802));
  NAND2xp33_ASAP7_75t_L     g00546(.A(\a[14] ), .B(new_n699), .Y(new_n803));
  INVx1_ASAP7_75t_L         g00547(.A(\a[13] ), .Y(new_n804));
  NAND2xp33_ASAP7_75t_L     g00548(.A(\a[14] ), .B(new_n804), .Y(new_n805));
  INVx1_ASAP7_75t_L         g00549(.A(\a[14] ), .Y(new_n806));
  NAND2xp33_ASAP7_75t_L     g00550(.A(\a[13] ), .B(new_n806), .Y(new_n807));
  AOI21xp33_ASAP7_75t_L     g00551(.A1(new_n807), .A2(new_n805), .B(new_n698), .Y(new_n808));
  NAND2xp33_ASAP7_75t_L     g00552(.A(new_n269), .B(new_n808), .Y(new_n809));
  NAND2xp33_ASAP7_75t_L     g00553(.A(new_n807), .B(new_n805), .Y(new_n810));
  NOR2xp33_ASAP7_75t_L      g00554(.A(new_n810), .B(new_n698), .Y(new_n811));
  NAND2xp33_ASAP7_75t_L     g00555(.A(\b[1] ), .B(new_n811), .Y(new_n812));
  NAND2xp33_ASAP7_75t_L     g00556(.A(new_n697), .B(new_n696), .Y(new_n813));
  XNOR2x2_ASAP7_75t_L       g00557(.A(\a[13] ), .B(\a[12] ), .Y(new_n814));
  NOR2xp33_ASAP7_75t_L      g00558(.A(new_n814), .B(new_n813), .Y(new_n815));
  NAND2xp33_ASAP7_75t_L     g00559(.A(\b[0] ), .B(new_n815), .Y(new_n816));
  NAND3xp33_ASAP7_75t_L     g00560(.A(new_n809), .B(new_n812), .C(new_n816), .Y(new_n817));
  XOR2x2_ASAP7_75t_L        g00561(.A(new_n803), .B(new_n817), .Y(new_n818));
  NAND3xp33_ASAP7_75t_L     g00562(.A(new_n800), .B(new_n802), .C(new_n818), .Y(new_n819));
  NOR2xp33_ASAP7_75t_L      g00563(.A(new_n574), .B(new_n801), .Y(new_n820));
  INVx1_ASAP7_75t_L         g00564(.A(new_n584), .Y(new_n821));
  O2A1O1Ixp33_ASAP7_75t_L   g00565(.A1(new_n298), .A2(new_n821), .B(new_n799), .C(\a[11] ), .Y(new_n822));
  XNOR2x2_ASAP7_75t_L       g00566(.A(new_n803), .B(new_n817), .Y(new_n823));
  OAI21xp33_ASAP7_75t_L     g00567(.A1(new_n820), .A2(new_n822), .B(new_n823), .Y(new_n824));
  NAND3xp33_ASAP7_75t_L     g00568(.A(new_n796), .B(new_n819), .C(new_n824), .Y(new_n825));
  NAND2xp33_ASAP7_75t_L     g00569(.A(new_n711), .B(new_n713), .Y(new_n826));
  MAJIxp5_ASAP7_75t_L       g00570(.A(new_n826), .B(new_n699), .C(new_n794), .Y(new_n827));
  NOR3xp33_ASAP7_75t_L      g00571(.A(new_n822), .B(new_n823), .C(new_n820), .Y(new_n828));
  AOI21xp33_ASAP7_75t_L     g00572(.A1(new_n800), .A2(new_n802), .B(new_n818), .Y(new_n829));
  OAI21xp33_ASAP7_75t_L     g00573(.A1(new_n829), .A2(new_n828), .B(new_n827), .Y(new_n830));
  AOI22xp33_ASAP7_75t_L     g00574(.A1(new_n444), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n471), .Y(new_n831));
  OAI221xp5_ASAP7_75t_L     g00575(.A1(new_n468), .A2(new_n418), .B1(new_n469), .B2(new_n425), .C(new_n831), .Y(new_n832));
  XNOR2x2_ASAP7_75t_L       g00576(.A(\a[8] ), .B(new_n832), .Y(new_n833));
  NAND3xp33_ASAP7_75t_L     g00577(.A(new_n825), .B(new_n830), .C(new_n833), .Y(new_n834));
  NOR3xp33_ASAP7_75t_L      g00578(.A(new_n827), .B(new_n828), .C(new_n829), .Y(new_n835));
  AOI21xp33_ASAP7_75t_L     g00579(.A1(new_n824), .A2(new_n819), .B(new_n796), .Y(new_n836));
  XNOR2x2_ASAP7_75t_L       g00580(.A(new_n435), .B(new_n832), .Y(new_n837));
  OAI21xp33_ASAP7_75t_L     g00581(.A1(new_n836), .A2(new_n835), .B(new_n837), .Y(new_n838));
  AOI211xp5_ASAP7_75t_L     g00582(.A1(new_n719), .A2(new_n725), .B(new_n714), .C(new_n710), .Y(new_n839));
  O2A1O1Ixp33_ASAP7_75t_L   g00583(.A1(new_n722), .A2(new_n726), .B(new_n741), .C(new_n839), .Y(new_n840));
  NAND3xp33_ASAP7_75t_L     g00584(.A(new_n840), .B(new_n838), .C(new_n834), .Y(new_n841));
  NAND2xp33_ASAP7_75t_L     g00585(.A(new_n834), .B(new_n838), .Y(new_n842));
  A2O1A1Ixp33_ASAP7_75t_L   g00586(.A1(new_n739), .A2(new_n741), .B(new_n839), .C(new_n842), .Y(new_n843));
  AOI22xp33_ASAP7_75t_L     g00587(.A1(new_n344), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n370), .Y(new_n844));
  OAI221xp5_ASAP7_75t_L     g00588(.A1(new_n429), .A2(new_n540), .B1(new_n366), .B2(new_n624), .C(new_n844), .Y(new_n845));
  XNOR2x2_ASAP7_75t_L       g00589(.A(\a[5] ), .B(new_n845), .Y(new_n846));
  INVx1_ASAP7_75t_L         g00590(.A(new_n846), .Y(new_n847));
  AOI21xp33_ASAP7_75t_L     g00591(.A1(new_n841), .A2(new_n843), .B(new_n847), .Y(new_n848));
  INVx1_ASAP7_75t_L         g00592(.A(new_n839), .Y(new_n849));
  OAI21xp33_ASAP7_75t_L     g00593(.A1(new_n727), .A2(new_n729), .B(new_n849), .Y(new_n850));
  NOR2xp33_ASAP7_75t_L      g00594(.A(new_n842), .B(new_n850), .Y(new_n851));
  AOI21xp33_ASAP7_75t_L     g00595(.A1(new_n838), .A2(new_n834), .B(new_n840), .Y(new_n852));
  NOR3xp33_ASAP7_75t_L      g00596(.A(new_n852), .B(new_n846), .C(new_n851), .Y(new_n853));
  NOR2xp33_ASAP7_75t_L      g00597(.A(new_n853), .B(new_n848), .Y(new_n854));
  NOR3xp33_ASAP7_75t_L      g00598(.A(new_n753), .B(new_n854), .C(new_n755), .Y(new_n855));
  INVx1_ASAP7_75t_L         g00599(.A(new_n854), .Y(new_n856));
  O2A1O1Ixp33_ASAP7_75t_L   g00600(.A1(new_n754), .A2(new_n752), .B(new_n747), .C(new_n856), .Y(new_n857));
  OR3x1_ASAP7_75t_L         g00601(.A(new_n855), .B(new_n857), .C(new_n793), .Y(new_n858));
  INVx1_ASAP7_75t_L         g00602(.A(new_n858), .Y(new_n859));
  OA21x2_ASAP7_75t_L        g00603(.A1(new_n857), .A2(new_n855), .B(new_n793), .Y(new_n860));
  NOR2xp33_ASAP7_75t_L      g00604(.A(new_n860), .B(new_n859), .Y(new_n861));
  A2O1A1Ixp33_ASAP7_75t_L   g00605(.A1(new_n772), .A2(new_n782), .B(new_n779), .C(new_n861), .Y(new_n862));
  NAND2xp33_ASAP7_75t_L     g00606(.A(new_n772), .B(new_n782), .Y(new_n863));
  OAI211xp5_ASAP7_75t_L     g00607(.A1(new_n860), .A2(new_n859), .B(new_n863), .C(new_n778), .Y(new_n864));
  AND2x2_ASAP7_75t_L        g00608(.A(new_n864), .B(new_n862), .Y(\f[13] ));
  INVx1_ASAP7_75t_L         g00609(.A(new_n680), .Y(new_n866));
  A2O1A1Ixp33_ASAP7_75t_L   g00610(.A1(new_n682), .A2(new_n866), .B(new_n759), .C(new_n788), .Y(new_n867));
  NOR2xp33_ASAP7_75t_L      g00611(.A(\b[13] ), .B(\b[14] ), .Y(new_n868));
  INVx1_ASAP7_75t_L         g00612(.A(\b[14] ), .Y(new_n869));
  NOR2xp33_ASAP7_75t_L      g00613(.A(new_n784), .B(new_n869), .Y(new_n870));
  NOR2xp33_ASAP7_75t_L      g00614(.A(new_n868), .B(new_n870), .Y(new_n871));
  A2O1A1Ixp33_ASAP7_75t_L   g00615(.A1(new_n867), .A2(new_n786), .B(new_n785), .C(new_n871), .Y(new_n872));
  O2A1O1Ixp33_ASAP7_75t_L   g00616(.A1(new_n761), .A2(new_n764), .B(new_n786), .C(new_n785), .Y(new_n873));
  OAI21xp33_ASAP7_75t_L     g00617(.A1(new_n868), .A2(new_n870), .B(new_n873), .Y(new_n874));
  NAND2xp33_ASAP7_75t_L     g00618(.A(new_n872), .B(new_n874), .Y(new_n875));
  AOI22xp33_ASAP7_75t_L     g00619(.A1(\b[12] ), .A2(new_n282), .B1(\b[14] ), .B2(new_n303), .Y(new_n876));
  OAI221xp5_ASAP7_75t_L     g00620(.A1(new_n291), .A2(new_n784), .B1(new_n268), .B2(new_n875), .C(new_n876), .Y(new_n877));
  XNOR2x2_ASAP7_75t_L       g00621(.A(\a[2] ), .B(new_n877), .Y(new_n878));
  INVx1_ASAP7_75t_L         g00622(.A(new_n848), .Y(new_n879));
  AOI22xp33_ASAP7_75t_L     g00623(.A1(new_n344), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n370), .Y(new_n880));
  OAI221xp5_ASAP7_75t_L     g00624(.A1(new_n429), .A2(new_n617), .B1(new_n366), .B2(new_n685), .C(new_n880), .Y(new_n881));
  XNOR2x2_ASAP7_75t_L       g00625(.A(\a[5] ), .B(new_n881), .Y(new_n882));
  INVx1_ASAP7_75t_L         g00626(.A(new_n842), .Y(new_n883));
  NAND3xp33_ASAP7_75t_L     g00627(.A(new_n825), .B(new_n830), .C(new_n837), .Y(new_n884));
  AOI22xp33_ASAP7_75t_L     g00628(.A1(new_n444), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n471), .Y(new_n885));
  OAI221xp5_ASAP7_75t_L     g00629(.A1(new_n468), .A2(new_n420), .B1(new_n469), .B2(new_n494), .C(new_n885), .Y(new_n886));
  XNOR2x2_ASAP7_75t_L       g00630(.A(new_n435), .B(new_n886), .Y(new_n887));
  A2O1A1O1Ixp25_ASAP7_75t_L g00631(.A1(new_n794), .A2(new_n699), .B(new_n710), .C(new_n819), .D(new_n829), .Y(new_n888));
  NAND2xp33_ASAP7_75t_L     g00632(.A(\b[4] ), .B(new_n584), .Y(new_n889));
  NAND2xp33_ASAP7_75t_L     g00633(.A(new_n578), .B(new_n359), .Y(new_n890));
  AOI22xp33_ASAP7_75t_L     g00634(.A1(\b[3] ), .A2(new_n651), .B1(\b[5] ), .B2(new_n581), .Y(new_n891));
  AND3x1_ASAP7_75t_L        g00635(.A(new_n890), .B(new_n891), .C(new_n889), .Y(new_n892));
  NAND2xp33_ASAP7_75t_L     g00636(.A(\a[11] ), .B(new_n892), .Y(new_n893));
  NAND3xp33_ASAP7_75t_L     g00637(.A(new_n890), .B(new_n889), .C(new_n891), .Y(new_n894));
  NAND2xp33_ASAP7_75t_L     g00638(.A(new_n574), .B(new_n894), .Y(new_n895));
  NAND2xp33_ASAP7_75t_L     g00639(.A(new_n895), .B(new_n893), .Y(new_n896));
  NAND2xp33_ASAP7_75t_L     g00640(.A(\b[1] ), .B(new_n815), .Y(new_n897));
  NAND2xp33_ASAP7_75t_L     g00641(.A(new_n810), .B(new_n813), .Y(new_n898));
  NOR2xp33_ASAP7_75t_L      g00642(.A(new_n280), .B(new_n898), .Y(new_n899));
  AND3x1_ASAP7_75t_L        g00643(.A(new_n698), .B(new_n814), .C(new_n810), .Y(new_n900));
  AOI221xp5_ASAP7_75t_L     g00644(.A1(new_n811), .A2(\b[2] ), .B1(new_n900), .B2(\b[0] ), .C(new_n899), .Y(new_n901));
  NAND2xp33_ASAP7_75t_L     g00645(.A(new_n897), .B(new_n901), .Y(new_n902));
  O2A1O1Ixp33_ASAP7_75t_L   g00646(.A1(new_n699), .A2(new_n817), .B(\a[14] ), .C(new_n902), .Y(new_n903));
  INVx1_ASAP7_75t_L         g00647(.A(new_n815), .Y(new_n904));
  A2O1A1Ixp33_ASAP7_75t_L   g00648(.A1(\b[0] ), .A2(new_n813), .B(new_n817), .C(\a[14] ), .Y(new_n905));
  O2A1O1Ixp33_ASAP7_75t_L   g00649(.A1(new_n904), .A2(new_n261), .B(new_n901), .C(new_n905), .Y(new_n906));
  NOR2xp33_ASAP7_75t_L      g00650(.A(new_n903), .B(new_n906), .Y(new_n907));
  NOR2xp33_ASAP7_75t_L      g00651(.A(new_n907), .B(new_n896), .Y(new_n908));
  OR2x4_ASAP7_75t_L         g00652(.A(new_n903), .B(new_n906), .Y(new_n909));
  AOI21xp33_ASAP7_75t_L     g00653(.A1(new_n895), .A2(new_n893), .B(new_n909), .Y(new_n910));
  OAI21xp33_ASAP7_75t_L     g00654(.A1(new_n910), .A2(new_n908), .B(new_n888), .Y(new_n911));
  A2O1A1Ixp33_ASAP7_75t_L   g00655(.A1(new_n723), .A2(new_n795), .B(new_n828), .C(new_n824), .Y(new_n912));
  NAND3xp33_ASAP7_75t_L     g00656(.A(new_n909), .B(new_n895), .C(new_n893), .Y(new_n913));
  NAND2xp33_ASAP7_75t_L     g00657(.A(new_n907), .B(new_n896), .Y(new_n914));
  NAND3xp33_ASAP7_75t_L     g00658(.A(new_n913), .B(new_n914), .C(new_n912), .Y(new_n915));
  AO21x2_ASAP7_75t_L        g00659(.A1(new_n915), .A2(new_n911), .B(new_n887), .Y(new_n916));
  NAND3xp33_ASAP7_75t_L     g00660(.A(new_n911), .B(new_n915), .C(new_n887), .Y(new_n917));
  NAND2xp33_ASAP7_75t_L     g00661(.A(new_n917), .B(new_n916), .Y(new_n918));
  O2A1O1Ixp33_ASAP7_75t_L   g00662(.A1(new_n883), .A2(new_n840), .B(new_n884), .C(new_n918), .Y(new_n919));
  A2O1A1Ixp33_ASAP7_75t_L   g00663(.A1(new_n838), .A2(new_n834), .B(new_n840), .C(new_n884), .Y(new_n920));
  AOI21xp33_ASAP7_75t_L     g00664(.A1(new_n917), .A2(new_n916), .B(new_n920), .Y(new_n921));
  OAI21xp33_ASAP7_75t_L     g00665(.A1(new_n921), .A2(new_n919), .B(new_n882), .Y(new_n922));
  OR3x1_ASAP7_75t_L         g00666(.A(new_n919), .B(new_n921), .C(new_n882), .Y(new_n923));
  NAND3xp33_ASAP7_75t_L     g00667(.A(new_n841), .B(new_n843), .C(new_n847), .Y(new_n924));
  OAI211xp5_ASAP7_75t_L     g00668(.A1(new_n754), .A2(new_n752), .B(new_n924), .C(new_n747), .Y(new_n925));
  NAND4xp25_ASAP7_75t_L     g00669(.A(new_n923), .B(new_n879), .C(new_n922), .D(new_n925), .Y(new_n926));
  AOI22xp33_ASAP7_75t_L     g00670(.A1(new_n879), .A2(new_n925), .B1(new_n922), .B2(new_n923), .Y(new_n927));
  INVx1_ASAP7_75t_L         g00671(.A(new_n927), .Y(new_n928));
  NAND3xp33_ASAP7_75t_L     g00672(.A(new_n928), .B(new_n926), .C(new_n878), .Y(new_n929));
  INVx1_ASAP7_75t_L         g00673(.A(new_n878), .Y(new_n930));
  INVx1_ASAP7_75t_L         g00674(.A(new_n926), .Y(new_n931));
  OAI21xp33_ASAP7_75t_L     g00675(.A1(new_n927), .A2(new_n931), .B(new_n930), .Y(new_n932));
  NAND2xp33_ASAP7_75t_L     g00676(.A(new_n932), .B(new_n929), .Y(new_n933));
  INVx1_ASAP7_75t_L         g00677(.A(new_n933), .Y(new_n934));
  A2O1A1O1Ixp25_ASAP7_75t_L g00678(.A1(new_n863), .A2(new_n778), .B(new_n860), .C(new_n858), .D(new_n934), .Y(new_n935));
  A2O1A1Ixp33_ASAP7_75t_L   g00679(.A1(new_n778), .A2(new_n863), .B(new_n860), .C(new_n858), .Y(new_n936));
  NOR2xp33_ASAP7_75t_L      g00680(.A(new_n933), .B(new_n936), .Y(new_n937));
  NOR2xp33_ASAP7_75t_L      g00681(.A(new_n937), .B(new_n935), .Y(\f[14] ));
  NOR3xp33_ASAP7_75t_L      g00682(.A(new_n931), .B(new_n927), .C(new_n878), .Y(new_n939));
  AOI21xp33_ASAP7_75t_L     g00683(.A1(new_n936), .A2(new_n933), .B(new_n939), .Y(new_n940));
  NOR2xp33_ASAP7_75t_L      g00684(.A(\b[14] ), .B(\b[15] ), .Y(new_n941));
  INVx1_ASAP7_75t_L         g00685(.A(\b[15] ), .Y(new_n942));
  NOR2xp33_ASAP7_75t_L      g00686(.A(new_n869), .B(new_n942), .Y(new_n943));
  NOR2xp33_ASAP7_75t_L      g00687(.A(new_n941), .B(new_n943), .Y(new_n944));
  INVx1_ASAP7_75t_L         g00688(.A(new_n944), .Y(new_n945));
  O2A1O1Ixp33_ASAP7_75t_L   g00689(.A1(new_n784), .A2(new_n869), .B(new_n872), .C(new_n945), .Y(new_n946));
  INVx1_ASAP7_75t_L         g00690(.A(new_n946), .Y(new_n947));
  A2O1A1O1Ixp25_ASAP7_75t_L g00691(.A1(new_n786), .A2(new_n867), .B(new_n785), .C(new_n871), .D(new_n870), .Y(new_n948));
  NAND2xp33_ASAP7_75t_L     g00692(.A(new_n945), .B(new_n948), .Y(new_n949));
  NAND2xp33_ASAP7_75t_L     g00693(.A(new_n949), .B(new_n947), .Y(new_n950));
  AOI22xp33_ASAP7_75t_L     g00694(.A1(\b[13] ), .A2(new_n282), .B1(\b[15] ), .B2(new_n303), .Y(new_n951));
  OAI221xp5_ASAP7_75t_L     g00695(.A1(new_n291), .A2(new_n869), .B1(new_n268), .B2(new_n950), .C(new_n951), .Y(new_n952));
  XNOR2x2_ASAP7_75t_L       g00696(.A(\a[2] ), .B(new_n952), .Y(new_n953));
  NOR3xp33_ASAP7_75t_L      g00697(.A(new_n919), .B(new_n921), .C(new_n882), .Y(new_n954));
  AO31x2_ASAP7_75t_L        g00698(.A1(new_n925), .A2(new_n922), .A3(new_n879), .B(new_n954), .Y(new_n955));
  AOI22xp33_ASAP7_75t_L     g00699(.A1(new_n344), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n370), .Y(new_n956));
  OAI221xp5_ASAP7_75t_L     g00700(.A1(new_n429), .A2(new_n679), .B1(new_n366), .B2(new_n768), .C(new_n956), .Y(new_n957));
  XNOR2x2_ASAP7_75t_L       g00701(.A(\a[5] ), .B(new_n957), .Y(new_n958));
  AND3x1_ASAP7_75t_L        g00702(.A(new_n911), .B(new_n915), .C(new_n887), .Y(new_n959));
  AOI22xp33_ASAP7_75t_L     g00703(.A1(new_n444), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n471), .Y(new_n960));
  OAI221xp5_ASAP7_75t_L     g00704(.A1(new_n468), .A2(new_n488), .B1(new_n469), .B2(new_n548), .C(new_n960), .Y(new_n961));
  XNOR2x2_ASAP7_75t_L       g00705(.A(\a[8] ), .B(new_n961), .Y(new_n962));
  NOR2xp33_ASAP7_75t_L      g00706(.A(new_n806), .B(new_n699), .Y(new_n963));
  NAND4xp25_ASAP7_75t_L     g00707(.A(new_n963), .B(new_n809), .C(new_n812), .D(new_n816), .Y(new_n964));
  INVx1_ASAP7_75t_L         g00708(.A(\a[15] ), .Y(new_n965));
  NAND2xp33_ASAP7_75t_L     g00709(.A(\a[14] ), .B(new_n965), .Y(new_n966));
  NAND2xp33_ASAP7_75t_L     g00710(.A(\a[15] ), .B(new_n806), .Y(new_n967));
  AND2x2_ASAP7_75t_L        g00711(.A(new_n966), .B(new_n967), .Y(new_n968));
  NOR2xp33_ASAP7_75t_L      g00712(.A(new_n258), .B(new_n968), .Y(new_n969));
  OAI21xp33_ASAP7_75t_L     g00713(.A1(new_n964), .A2(new_n902), .B(new_n969), .Y(new_n970));
  AND4x1_ASAP7_75t_L        g00714(.A(new_n809), .B(new_n963), .C(new_n812), .D(new_n816), .Y(new_n971));
  INVx1_ASAP7_75t_L         g00715(.A(new_n969), .Y(new_n972));
  NAND4xp25_ASAP7_75t_L     g00716(.A(new_n971), .B(new_n972), .C(new_n901), .D(new_n897), .Y(new_n973));
  AOI22xp33_ASAP7_75t_L     g00717(.A1(new_n811), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n900), .Y(new_n974));
  OAI221xp5_ASAP7_75t_L     g00718(.A1(new_n898), .A2(new_n302), .B1(new_n276), .B2(new_n904), .C(new_n974), .Y(new_n975));
  NOR2xp33_ASAP7_75t_L      g00719(.A(new_n806), .B(new_n975), .Y(new_n976));
  NAND3xp33_ASAP7_75t_L     g00720(.A(new_n813), .B(new_n805), .C(new_n807), .Y(new_n977));
  NAND3xp33_ASAP7_75t_L     g00721(.A(new_n698), .B(new_n810), .C(new_n814), .Y(new_n978));
  OAI22xp33_ASAP7_75t_L     g00722(.A1(new_n978), .A2(new_n261), .B1(new_n298), .B2(new_n977), .Y(new_n979));
  AOI221xp5_ASAP7_75t_L     g00723(.A1(\b[2] ), .A2(new_n815), .B1(new_n406), .B2(new_n808), .C(new_n979), .Y(new_n980));
  NOR2xp33_ASAP7_75t_L      g00724(.A(\a[14] ), .B(new_n980), .Y(new_n981));
  NOR2xp33_ASAP7_75t_L      g00725(.A(new_n981), .B(new_n976), .Y(new_n982));
  AOI21xp33_ASAP7_75t_L     g00726(.A1(new_n973), .A2(new_n970), .B(new_n982), .Y(new_n983));
  AOI31xp33_ASAP7_75t_L     g00727(.A1(new_n971), .A2(new_n897), .A3(new_n901), .B(new_n972), .Y(new_n984));
  NOR3xp33_ASAP7_75t_L      g00728(.A(new_n902), .B(new_n969), .C(new_n964), .Y(new_n985));
  NOR4xp25_ASAP7_75t_L      g00729(.A(new_n985), .B(new_n981), .C(new_n984), .D(new_n976), .Y(new_n986));
  NOR2xp33_ASAP7_75t_L      g00730(.A(new_n354), .B(new_n821), .Y(new_n987));
  INVx1_ASAP7_75t_L         g00731(.A(new_n987), .Y(new_n988));
  NAND2xp33_ASAP7_75t_L     g00732(.A(new_n578), .B(new_n526), .Y(new_n989));
  AOI22xp33_ASAP7_75t_L     g00733(.A1(\b[4] ), .A2(new_n651), .B1(\b[6] ), .B2(new_n581), .Y(new_n990));
  NAND4xp25_ASAP7_75t_L     g00734(.A(new_n989), .B(\a[11] ), .C(new_n988), .D(new_n990), .Y(new_n991));
  INVx1_ASAP7_75t_L         g00735(.A(new_n991), .Y(new_n992));
  AOI31xp33_ASAP7_75t_L     g00736(.A1(new_n989), .A2(new_n988), .A3(new_n990), .B(\a[11] ), .Y(new_n993));
  NOR4xp25_ASAP7_75t_L      g00737(.A(new_n983), .B(new_n993), .C(new_n992), .D(new_n986), .Y(new_n994));
  OAI22xp33_ASAP7_75t_L     g00738(.A1(new_n985), .A2(new_n984), .B1(new_n981), .B2(new_n976), .Y(new_n995));
  NAND3xp33_ASAP7_75t_L     g00739(.A(new_n982), .B(new_n973), .C(new_n970), .Y(new_n996));
  INVx1_ASAP7_75t_L         g00740(.A(new_n993), .Y(new_n997));
  AOI22xp33_ASAP7_75t_L     g00741(.A1(new_n991), .A2(new_n997), .B1(new_n995), .B2(new_n996), .Y(new_n998));
  OAI221xp5_ASAP7_75t_L     g00742(.A1(new_n910), .A2(new_n912), .B1(new_n998), .B2(new_n994), .C(new_n913), .Y(new_n999));
  NOR2xp33_ASAP7_75t_L      g00743(.A(new_n998), .B(new_n994), .Y(new_n1000));
  A2O1A1Ixp33_ASAP7_75t_L   g00744(.A1(new_n914), .A2(new_n888), .B(new_n908), .C(new_n1000), .Y(new_n1001));
  AO21x2_ASAP7_75t_L        g00745(.A1(new_n999), .A2(new_n1001), .B(new_n962), .Y(new_n1002));
  NAND3xp33_ASAP7_75t_L     g00746(.A(new_n1001), .B(new_n999), .C(new_n962), .Y(new_n1003));
  NAND2xp33_ASAP7_75t_L     g00747(.A(new_n1003), .B(new_n1002), .Y(new_n1004));
  A2O1A1Ixp33_ASAP7_75t_L   g00748(.A1(new_n916), .A2(new_n920), .B(new_n959), .C(new_n1004), .Y(new_n1005));
  INVx1_ASAP7_75t_L         g00749(.A(new_n884), .Y(new_n1006));
  A2O1A1O1Ixp25_ASAP7_75t_L g00750(.A1(new_n842), .A2(new_n850), .B(new_n1006), .C(new_n916), .D(new_n959), .Y(new_n1007));
  AOI21xp33_ASAP7_75t_L     g00751(.A1(new_n1001), .A2(new_n999), .B(new_n962), .Y(new_n1008));
  AND3x1_ASAP7_75t_L        g00752(.A(new_n1001), .B(new_n999), .C(new_n962), .Y(new_n1009));
  NOR2xp33_ASAP7_75t_L      g00753(.A(new_n1008), .B(new_n1009), .Y(new_n1010));
  NAND2xp33_ASAP7_75t_L     g00754(.A(new_n1007), .B(new_n1010), .Y(new_n1011));
  AOI21xp33_ASAP7_75t_L     g00755(.A1(new_n1005), .A2(new_n1011), .B(new_n958), .Y(new_n1012));
  INVx1_ASAP7_75t_L         g00756(.A(new_n958), .Y(new_n1013));
  A2O1A1O1Ixp25_ASAP7_75t_L g00757(.A1(new_n884), .A2(new_n843), .B(new_n918), .C(new_n917), .D(new_n1010), .Y(new_n1014));
  NOR3xp33_ASAP7_75t_L      g00758(.A(new_n919), .B(new_n1004), .C(new_n959), .Y(new_n1015));
  NOR3xp33_ASAP7_75t_L      g00759(.A(new_n1014), .B(new_n1015), .C(new_n1013), .Y(new_n1016));
  OAI21xp33_ASAP7_75t_L     g00760(.A1(new_n1012), .A2(new_n1016), .B(new_n955), .Y(new_n1017));
  AOI31xp33_ASAP7_75t_L     g00761(.A1(new_n925), .A2(new_n922), .A3(new_n879), .B(new_n954), .Y(new_n1018));
  NOR2xp33_ASAP7_75t_L      g00762(.A(new_n1012), .B(new_n1016), .Y(new_n1019));
  NAND2xp33_ASAP7_75t_L     g00763(.A(new_n1018), .B(new_n1019), .Y(new_n1020));
  AOI21xp33_ASAP7_75t_L     g00764(.A1(new_n1020), .A2(new_n1017), .B(new_n953), .Y(new_n1021));
  INVx1_ASAP7_75t_L         g00765(.A(new_n953), .Y(new_n1022));
  INVx1_ASAP7_75t_L         g00766(.A(new_n1017), .Y(new_n1023));
  NOR3xp33_ASAP7_75t_L      g00767(.A(new_n955), .B(new_n1012), .C(new_n1016), .Y(new_n1024));
  NOR3xp33_ASAP7_75t_L      g00768(.A(new_n1023), .B(new_n1024), .C(new_n1022), .Y(new_n1025));
  NOR2xp33_ASAP7_75t_L      g00769(.A(new_n1021), .B(new_n1025), .Y(new_n1026));
  XOR2x2_ASAP7_75t_L        g00770(.A(new_n1026), .B(new_n940), .Y(\f[15] ));
  NAND3xp33_ASAP7_75t_L     g00771(.A(new_n1020), .B(new_n1017), .C(new_n1022), .Y(new_n1028));
  NOR2xp33_ASAP7_75t_L      g00772(.A(\b[15] ), .B(\b[16] ), .Y(new_n1029));
  INVx1_ASAP7_75t_L         g00773(.A(\b[16] ), .Y(new_n1030));
  NOR2xp33_ASAP7_75t_L      g00774(.A(new_n942), .B(new_n1030), .Y(new_n1031));
  NOR2xp33_ASAP7_75t_L      g00775(.A(new_n1029), .B(new_n1031), .Y(new_n1032));
  A2O1A1Ixp33_ASAP7_75t_L   g00776(.A1(\b[15] ), .A2(\b[14] ), .B(new_n946), .C(new_n1032), .Y(new_n1033));
  OR3x1_ASAP7_75t_L         g00777(.A(new_n946), .B(new_n943), .C(new_n1032), .Y(new_n1034));
  NAND2xp33_ASAP7_75t_L     g00778(.A(new_n1033), .B(new_n1034), .Y(new_n1035));
  AOI22xp33_ASAP7_75t_L     g00779(.A1(\b[14] ), .A2(new_n282), .B1(\b[16] ), .B2(new_n303), .Y(new_n1036));
  OAI221xp5_ASAP7_75t_L     g00780(.A1(new_n291), .A2(new_n942), .B1(new_n268), .B2(new_n1035), .C(new_n1036), .Y(new_n1037));
  XNOR2x2_ASAP7_75t_L       g00781(.A(\a[2] ), .B(new_n1037), .Y(new_n1038));
  NAND3xp33_ASAP7_75t_L     g00782(.A(new_n1005), .B(new_n1011), .C(new_n1013), .Y(new_n1039));
  AOI22xp33_ASAP7_75t_L     g00783(.A1(new_n344), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n370), .Y(new_n1040));
  OAI221xp5_ASAP7_75t_L     g00784(.A1(new_n429), .A2(new_n760), .B1(new_n366), .B2(new_n790), .C(new_n1040), .Y(new_n1041));
  XNOR2x2_ASAP7_75t_L       g00785(.A(\a[5] ), .B(new_n1041), .Y(new_n1042));
  NAND4xp25_ASAP7_75t_L     g00786(.A(new_n996), .B(new_n991), .C(new_n997), .D(new_n995), .Y(new_n1043));
  OAI22xp33_ASAP7_75t_L     g00787(.A1(new_n983), .A2(new_n986), .B1(new_n993), .B2(new_n992), .Y(new_n1044));
  AOI221xp5_ASAP7_75t_L     g00788(.A1(new_n1044), .A2(new_n1043), .B1(new_n914), .B2(new_n888), .C(new_n908), .Y(new_n1045));
  NAND2xp33_ASAP7_75t_L     g00789(.A(new_n1043), .B(new_n1044), .Y(new_n1046));
  O2A1O1Ixp33_ASAP7_75t_L   g00790(.A1(new_n912), .A2(new_n910), .B(new_n913), .C(new_n1046), .Y(new_n1047));
  OR3x1_ASAP7_75t_L         g00791(.A(new_n1047), .B(new_n962), .C(new_n1045), .Y(new_n1048));
  AOI22xp33_ASAP7_75t_L     g00792(.A1(new_n444), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n471), .Y(new_n1049));
  OAI221xp5_ASAP7_75t_L     g00793(.A1(new_n468), .A2(new_n540), .B1(new_n469), .B2(new_n624), .C(new_n1049), .Y(new_n1050));
  XNOR2x2_ASAP7_75t_L       g00794(.A(new_n435), .B(new_n1050), .Y(new_n1051));
  INVx1_ASAP7_75t_L         g00795(.A(new_n1051), .Y(new_n1052));
  AOI211xp5_ASAP7_75t_L     g00796(.A1(new_n991), .A2(new_n997), .B(new_n986), .C(new_n983), .Y(new_n1053));
  INVx1_ASAP7_75t_L         g00797(.A(new_n1053), .Y(new_n1054));
  AOI22xp33_ASAP7_75t_L     g00798(.A1(\b[5] ), .A2(new_n651), .B1(\b[7] ), .B2(new_n581), .Y(new_n1055));
  OAI221xp5_ASAP7_75t_L     g00799(.A1(new_n821), .A2(new_n418), .B1(new_n577), .B2(new_n425), .C(new_n1055), .Y(new_n1056));
  XNOR2x2_ASAP7_75t_L       g00800(.A(\a[11] ), .B(new_n1056), .Y(new_n1057));
  INVx1_ASAP7_75t_L         g00801(.A(new_n1057), .Y(new_n1058));
  NAND2xp33_ASAP7_75t_L     g00802(.A(new_n973), .B(new_n970), .Y(new_n1059));
  XNOR2x2_ASAP7_75t_L       g00803(.A(\a[14] ), .B(new_n980), .Y(new_n1060));
  NOR3xp33_ASAP7_75t_L      g00804(.A(new_n902), .B(new_n972), .C(new_n964), .Y(new_n1061));
  NAND2xp33_ASAP7_75t_L     g00805(.A(\b[3] ), .B(new_n815), .Y(new_n1062));
  NAND2xp33_ASAP7_75t_L     g00806(.A(new_n808), .B(new_n329), .Y(new_n1063));
  AOI22xp33_ASAP7_75t_L     g00807(.A1(new_n811), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n900), .Y(new_n1064));
  NAND4xp25_ASAP7_75t_L     g00808(.A(new_n1063), .B(\a[14] ), .C(new_n1062), .D(new_n1064), .Y(new_n1065));
  INVx1_ASAP7_75t_L         g00809(.A(new_n1065), .Y(new_n1066));
  AOI31xp33_ASAP7_75t_L     g00810(.A1(new_n1063), .A2(new_n1062), .A3(new_n1064), .B(\a[14] ), .Y(new_n1067));
  NAND2xp33_ASAP7_75t_L     g00811(.A(\a[17] ), .B(new_n969), .Y(new_n1068));
  INVx1_ASAP7_75t_L         g00812(.A(\a[16] ), .Y(new_n1069));
  NAND2xp33_ASAP7_75t_L     g00813(.A(\a[17] ), .B(new_n1069), .Y(new_n1070));
  INVx1_ASAP7_75t_L         g00814(.A(\a[17] ), .Y(new_n1071));
  NAND2xp33_ASAP7_75t_L     g00815(.A(\a[16] ), .B(new_n1071), .Y(new_n1072));
  AOI21xp33_ASAP7_75t_L     g00816(.A1(new_n1072), .A2(new_n1070), .B(new_n968), .Y(new_n1073));
  NAND2xp33_ASAP7_75t_L     g00817(.A(new_n269), .B(new_n1073), .Y(new_n1074));
  NAND2xp33_ASAP7_75t_L     g00818(.A(new_n1072), .B(new_n1070), .Y(new_n1075));
  NOR2xp33_ASAP7_75t_L      g00819(.A(new_n1075), .B(new_n968), .Y(new_n1076));
  NAND2xp33_ASAP7_75t_L     g00820(.A(\b[1] ), .B(new_n1076), .Y(new_n1077));
  NAND2xp33_ASAP7_75t_L     g00821(.A(new_n967), .B(new_n966), .Y(new_n1078));
  XNOR2x2_ASAP7_75t_L       g00822(.A(\a[16] ), .B(\a[15] ), .Y(new_n1079));
  NOR2xp33_ASAP7_75t_L      g00823(.A(new_n1079), .B(new_n1078), .Y(new_n1080));
  NAND2xp33_ASAP7_75t_L     g00824(.A(\b[0] ), .B(new_n1080), .Y(new_n1081));
  NAND3xp33_ASAP7_75t_L     g00825(.A(new_n1074), .B(new_n1077), .C(new_n1081), .Y(new_n1082));
  XNOR2x2_ASAP7_75t_L       g00826(.A(new_n1068), .B(new_n1082), .Y(new_n1083));
  NOR3xp33_ASAP7_75t_L      g00827(.A(new_n1083), .B(new_n1066), .C(new_n1067), .Y(new_n1084));
  INVx1_ASAP7_75t_L         g00828(.A(new_n1067), .Y(new_n1085));
  XOR2x2_ASAP7_75t_L        g00829(.A(new_n1068), .B(new_n1082), .Y(new_n1086));
  AOI21xp33_ASAP7_75t_L     g00830(.A1(new_n1085), .A2(new_n1065), .B(new_n1086), .Y(new_n1087));
  NOR2xp33_ASAP7_75t_L      g00831(.A(new_n1084), .B(new_n1087), .Y(new_n1088));
  A2O1A1Ixp33_ASAP7_75t_L   g00832(.A1(new_n1060), .A2(new_n1059), .B(new_n1061), .C(new_n1088), .Y(new_n1089));
  O2A1O1Ixp33_ASAP7_75t_L   g00833(.A1(new_n984), .A2(new_n985), .B(new_n1060), .C(new_n1061), .Y(new_n1090));
  OAI21xp33_ASAP7_75t_L     g00834(.A1(new_n1084), .A2(new_n1087), .B(new_n1090), .Y(new_n1091));
  AOI21xp33_ASAP7_75t_L     g00835(.A1(new_n1089), .A2(new_n1091), .B(new_n1058), .Y(new_n1092));
  NOR3xp33_ASAP7_75t_L      g00836(.A(new_n1090), .B(new_n1084), .C(new_n1087), .Y(new_n1093));
  INVx1_ASAP7_75t_L         g00837(.A(new_n1061), .Y(new_n1094));
  A2O1A1Ixp33_ASAP7_75t_L   g00838(.A1(new_n973), .A2(new_n970), .B(new_n982), .C(new_n1094), .Y(new_n1095));
  NOR2xp33_ASAP7_75t_L      g00839(.A(new_n1095), .B(new_n1088), .Y(new_n1096));
  NOR3xp33_ASAP7_75t_L      g00840(.A(new_n1096), .B(new_n1093), .C(new_n1057), .Y(new_n1097));
  AOI211xp5_ASAP7_75t_L     g00841(.A1(new_n999), .A2(new_n1054), .B(new_n1092), .C(new_n1097), .Y(new_n1098));
  OAI21xp33_ASAP7_75t_L     g00842(.A1(new_n1093), .A2(new_n1096), .B(new_n1057), .Y(new_n1099));
  NAND3xp33_ASAP7_75t_L     g00843(.A(new_n1058), .B(new_n1089), .C(new_n1091), .Y(new_n1100));
  AOI211xp5_ASAP7_75t_L     g00844(.A1(new_n1100), .A2(new_n1099), .B(new_n1045), .C(new_n1053), .Y(new_n1101));
  OAI21xp33_ASAP7_75t_L     g00845(.A1(new_n1101), .A2(new_n1098), .B(new_n1052), .Y(new_n1102));
  OAI211xp5_ASAP7_75t_L     g00846(.A1(new_n1053), .A2(new_n1045), .B(new_n1099), .C(new_n1100), .Y(new_n1103));
  OAI211xp5_ASAP7_75t_L     g00847(.A1(new_n1097), .A2(new_n1092), .B(new_n1054), .C(new_n999), .Y(new_n1104));
  NAND3xp33_ASAP7_75t_L     g00848(.A(new_n1103), .B(new_n1104), .C(new_n1051), .Y(new_n1105));
  NAND2xp33_ASAP7_75t_L     g00849(.A(new_n1105), .B(new_n1102), .Y(new_n1106));
  O2A1O1Ixp33_ASAP7_75t_L   g00850(.A1(new_n1007), .A2(new_n1010), .B(new_n1048), .C(new_n1106), .Y(new_n1107));
  A2O1A1Ixp33_ASAP7_75t_L   g00851(.A1(new_n1002), .A2(new_n1003), .B(new_n1007), .C(new_n1048), .Y(new_n1108));
  AOI21xp33_ASAP7_75t_L     g00852(.A1(new_n1105), .A2(new_n1102), .B(new_n1108), .Y(new_n1109));
  OAI21xp33_ASAP7_75t_L     g00853(.A1(new_n1109), .A2(new_n1107), .B(new_n1042), .Y(new_n1110));
  INVx1_ASAP7_75t_L         g00854(.A(new_n1042), .Y(new_n1111));
  NAND3xp33_ASAP7_75t_L     g00855(.A(new_n1108), .B(new_n1102), .C(new_n1105), .Y(new_n1112));
  OAI211xp5_ASAP7_75t_L     g00856(.A1(new_n1007), .A2(new_n1010), .B(new_n1106), .C(new_n1048), .Y(new_n1113));
  NAND3xp33_ASAP7_75t_L     g00857(.A(new_n1113), .B(new_n1112), .C(new_n1111), .Y(new_n1114));
  NAND2xp33_ASAP7_75t_L     g00858(.A(new_n1114), .B(new_n1110), .Y(new_n1115));
  O2A1O1Ixp33_ASAP7_75t_L   g00859(.A1(new_n1018), .A2(new_n1019), .B(new_n1039), .C(new_n1115), .Y(new_n1116));
  OAI21xp33_ASAP7_75t_L     g00860(.A1(new_n1015), .A2(new_n1014), .B(new_n1013), .Y(new_n1117));
  NAND3xp33_ASAP7_75t_L     g00861(.A(new_n1005), .B(new_n1011), .C(new_n958), .Y(new_n1118));
  A2O1A1Ixp33_ASAP7_75t_L   g00862(.A1(new_n1117), .A2(new_n1118), .B(new_n1018), .C(new_n1039), .Y(new_n1119));
  AOI21xp33_ASAP7_75t_L     g00863(.A1(new_n1114), .A2(new_n1110), .B(new_n1119), .Y(new_n1120));
  NOR2xp33_ASAP7_75t_L      g00864(.A(new_n1120), .B(new_n1116), .Y(new_n1121));
  NAND2xp33_ASAP7_75t_L     g00865(.A(new_n1038), .B(new_n1121), .Y(new_n1122));
  INVx1_ASAP7_75t_L         g00866(.A(new_n1038), .Y(new_n1123));
  OAI21xp33_ASAP7_75t_L     g00867(.A1(new_n1120), .A2(new_n1116), .B(new_n1123), .Y(new_n1124));
  NAND2xp33_ASAP7_75t_L     g00868(.A(new_n1124), .B(new_n1122), .Y(new_n1125));
  INVx1_ASAP7_75t_L         g00869(.A(new_n1125), .Y(new_n1126));
  O2A1O1Ixp33_ASAP7_75t_L   g00870(.A1(new_n940), .A2(new_n1026), .B(new_n1028), .C(new_n1126), .Y(new_n1127));
  OAI21xp33_ASAP7_75t_L     g00871(.A1(new_n1026), .A2(new_n940), .B(new_n1028), .Y(new_n1128));
  NOR2xp33_ASAP7_75t_L      g00872(.A(new_n1125), .B(new_n1128), .Y(new_n1129));
  NOR2xp33_ASAP7_75t_L      g00873(.A(new_n1129), .B(new_n1127), .Y(\f[16] ));
  INVx1_ASAP7_75t_L         g00874(.A(new_n1114), .Y(new_n1131));
  AOI22xp33_ASAP7_75t_L     g00875(.A1(new_n344), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n370), .Y(new_n1132));
  OAI221xp5_ASAP7_75t_L     g00876(.A1(new_n429), .A2(new_n784), .B1(new_n366), .B2(new_n875), .C(new_n1132), .Y(new_n1133));
  XNOR2x2_ASAP7_75t_L       g00877(.A(\a[5] ), .B(new_n1133), .Y(new_n1134));
  INVx1_ASAP7_75t_L         g00878(.A(new_n1134), .Y(new_n1135));
  INVx1_ASAP7_75t_L         g00879(.A(new_n1105), .Y(new_n1136));
  AOI22xp33_ASAP7_75t_L     g00880(.A1(new_n444), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n471), .Y(new_n1137));
  OAI221xp5_ASAP7_75t_L     g00881(.A1(new_n468), .A2(new_n617), .B1(new_n469), .B2(new_n685), .C(new_n1137), .Y(new_n1138));
  XNOR2x2_ASAP7_75t_L       g00882(.A(\a[8] ), .B(new_n1138), .Y(new_n1139));
  AOI21xp33_ASAP7_75t_L     g00883(.A1(new_n888), .A2(new_n914), .B(new_n908), .Y(new_n1140));
  A2O1A1O1Ixp25_ASAP7_75t_L g00884(.A1(new_n1046), .A2(new_n1140), .B(new_n1053), .C(new_n1099), .D(new_n1097), .Y(new_n1141));
  AOI22xp33_ASAP7_75t_L     g00885(.A1(\b[6] ), .A2(new_n651), .B1(\b[8] ), .B2(new_n581), .Y(new_n1142));
  OAI221xp5_ASAP7_75t_L     g00886(.A1(new_n821), .A2(new_n420), .B1(new_n577), .B2(new_n494), .C(new_n1142), .Y(new_n1143));
  XNOR2x2_ASAP7_75t_L       g00887(.A(new_n574), .B(new_n1143), .Y(new_n1144));
  NAND3xp33_ASAP7_75t_L     g00888(.A(new_n1085), .B(new_n1086), .C(new_n1065), .Y(new_n1145));
  A2O1A1O1Ixp25_ASAP7_75t_L g00889(.A1(new_n1060), .A2(new_n1059), .B(new_n1061), .C(new_n1145), .D(new_n1087), .Y(new_n1146));
  NAND2xp33_ASAP7_75t_L     g00890(.A(\b[4] ), .B(new_n815), .Y(new_n1147));
  AOI22xp33_ASAP7_75t_L     g00891(.A1(new_n811), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n900), .Y(new_n1148));
  OAI311xp33_ASAP7_75t_L    g00892(.A1(new_n357), .A2(new_n898), .A3(new_n358), .B1(new_n1147), .C1(new_n1148), .Y(new_n1149));
  NOR2xp33_ASAP7_75t_L      g00893(.A(new_n806), .B(new_n1149), .Y(new_n1150));
  NAND2xp33_ASAP7_75t_L     g00894(.A(new_n806), .B(new_n1149), .Y(new_n1151));
  INVx1_ASAP7_75t_L         g00895(.A(new_n1151), .Y(new_n1152));
  INVx1_ASAP7_75t_L         g00896(.A(new_n1082), .Y(new_n1153));
  OR2x4_ASAP7_75t_L         g00897(.A(new_n1079), .B(new_n1078), .Y(new_n1154));
  NOR2xp33_ASAP7_75t_L      g00898(.A(new_n261), .B(new_n1154), .Y(new_n1155));
  NAND2xp33_ASAP7_75t_L     g00899(.A(new_n1075), .B(new_n1078), .Y(new_n1156));
  NAND2xp33_ASAP7_75t_L     g00900(.A(\b[2] ), .B(new_n1076), .Y(new_n1157));
  NAND3xp33_ASAP7_75t_L     g00901(.A(new_n968), .B(new_n1075), .C(new_n1079), .Y(new_n1158));
  OAI221xp5_ASAP7_75t_L     g00902(.A1(new_n258), .A2(new_n1158), .B1(new_n280), .B2(new_n1156), .C(new_n1157), .Y(new_n1159));
  NOR2xp33_ASAP7_75t_L      g00903(.A(new_n1155), .B(new_n1159), .Y(new_n1160));
  A2O1A1Ixp33_ASAP7_75t_L   g00904(.A1(new_n972), .A2(new_n1153), .B(new_n1071), .C(new_n1160), .Y(new_n1161));
  A2O1A1Ixp33_ASAP7_75t_L   g00905(.A1(\b[0] ), .A2(new_n1078), .B(new_n1082), .C(\a[17] ), .Y(new_n1162));
  INVx1_ASAP7_75t_L         g00906(.A(new_n1162), .Y(new_n1163));
  A2O1A1Ixp33_ASAP7_75t_L   g00907(.A1(\b[1] ), .A2(new_n1080), .B(new_n1159), .C(new_n1163), .Y(new_n1164));
  AOI211xp5_ASAP7_75t_L     g00908(.A1(new_n1164), .A2(new_n1161), .B(new_n1150), .C(new_n1152), .Y(new_n1165));
  INVx1_ASAP7_75t_L         g00909(.A(new_n1150), .Y(new_n1166));
  XNOR2x2_ASAP7_75t_L       g00910(.A(new_n1160), .B(new_n1162), .Y(new_n1167));
  AOI21xp33_ASAP7_75t_L     g00911(.A1(new_n1151), .A2(new_n1166), .B(new_n1167), .Y(new_n1168));
  OAI21xp33_ASAP7_75t_L     g00912(.A1(new_n1168), .A2(new_n1165), .B(new_n1146), .Y(new_n1169));
  OAI21xp33_ASAP7_75t_L     g00913(.A1(new_n1067), .A2(new_n1066), .B(new_n1083), .Y(new_n1170));
  A2O1A1Ixp33_ASAP7_75t_L   g00914(.A1(new_n995), .A2(new_n1094), .B(new_n1084), .C(new_n1170), .Y(new_n1171));
  NAND3xp33_ASAP7_75t_L     g00915(.A(new_n1167), .B(new_n1151), .C(new_n1166), .Y(new_n1172));
  OAI211xp5_ASAP7_75t_L     g00916(.A1(new_n1150), .A2(new_n1152), .B(new_n1164), .C(new_n1161), .Y(new_n1173));
  NAND3xp33_ASAP7_75t_L     g00917(.A(new_n1171), .B(new_n1172), .C(new_n1173), .Y(new_n1174));
  AOI21xp33_ASAP7_75t_L     g00918(.A1(new_n1174), .A2(new_n1169), .B(new_n1144), .Y(new_n1175));
  NAND3xp33_ASAP7_75t_L     g00919(.A(new_n1174), .B(new_n1169), .C(new_n1144), .Y(new_n1176));
  INVx1_ASAP7_75t_L         g00920(.A(new_n1176), .Y(new_n1177));
  NOR3xp33_ASAP7_75t_L      g00921(.A(new_n1141), .B(new_n1175), .C(new_n1177), .Y(new_n1178));
  A2O1A1Ixp33_ASAP7_75t_L   g00922(.A1(new_n999), .A2(new_n1054), .B(new_n1092), .C(new_n1100), .Y(new_n1179));
  INVx1_ASAP7_75t_L         g00923(.A(new_n1175), .Y(new_n1180));
  AOI21xp33_ASAP7_75t_L     g00924(.A1(new_n1176), .A2(new_n1180), .B(new_n1179), .Y(new_n1181));
  OAI21xp33_ASAP7_75t_L     g00925(.A1(new_n1181), .A2(new_n1178), .B(new_n1139), .Y(new_n1182));
  NOR2xp33_ASAP7_75t_L      g00926(.A(new_n435), .B(new_n1138), .Y(new_n1183));
  AND2x2_ASAP7_75t_L        g00927(.A(new_n435), .B(new_n1138), .Y(new_n1184));
  NAND3xp33_ASAP7_75t_L     g00928(.A(new_n1179), .B(new_n1180), .C(new_n1176), .Y(new_n1185));
  OAI21xp33_ASAP7_75t_L     g00929(.A1(new_n1175), .A2(new_n1177), .B(new_n1141), .Y(new_n1186));
  OAI211xp5_ASAP7_75t_L     g00930(.A1(new_n1184), .A2(new_n1183), .B(new_n1185), .C(new_n1186), .Y(new_n1187));
  AND2x2_ASAP7_75t_L        g00931(.A(new_n1187), .B(new_n1182), .Y(new_n1188));
  OAI21xp33_ASAP7_75t_L     g00932(.A1(new_n1136), .A2(new_n1107), .B(new_n1188), .Y(new_n1189));
  AOI221xp5_ASAP7_75t_L     g00933(.A1(new_n1108), .A2(new_n1102), .B1(new_n1182), .B2(new_n1187), .C(new_n1136), .Y(new_n1190));
  INVx1_ASAP7_75t_L         g00934(.A(new_n1190), .Y(new_n1191));
  AOI21xp33_ASAP7_75t_L     g00935(.A1(new_n1189), .A2(new_n1191), .B(new_n1135), .Y(new_n1192));
  NAND2xp33_ASAP7_75t_L     g00936(.A(new_n1187), .B(new_n1182), .Y(new_n1193));
  A2O1A1O1Ixp25_ASAP7_75t_L g00937(.A1(new_n1048), .A2(new_n1005), .B(new_n1106), .C(new_n1105), .D(new_n1193), .Y(new_n1194));
  NOR3xp33_ASAP7_75t_L      g00938(.A(new_n1194), .B(new_n1190), .C(new_n1134), .Y(new_n1195));
  NOR2xp33_ASAP7_75t_L      g00939(.A(new_n1192), .B(new_n1195), .Y(new_n1196));
  A2O1A1Ixp33_ASAP7_75t_L   g00940(.A1(new_n1110), .A2(new_n1119), .B(new_n1131), .C(new_n1196), .Y(new_n1197));
  AOI21xp33_ASAP7_75t_L     g00941(.A1(new_n1119), .A2(new_n1110), .B(new_n1131), .Y(new_n1198));
  OAI21xp33_ASAP7_75t_L     g00942(.A1(new_n1192), .A2(new_n1195), .B(new_n1198), .Y(new_n1199));
  NOR2xp33_ASAP7_75t_L      g00943(.A(\b[16] ), .B(\b[17] ), .Y(new_n1200));
  INVx1_ASAP7_75t_L         g00944(.A(\b[17] ), .Y(new_n1201));
  NOR2xp33_ASAP7_75t_L      g00945(.A(new_n1030), .B(new_n1201), .Y(new_n1202));
  NOR2xp33_ASAP7_75t_L      g00946(.A(new_n1200), .B(new_n1202), .Y(new_n1203));
  INVx1_ASAP7_75t_L         g00947(.A(new_n1203), .Y(new_n1204));
  O2A1O1Ixp33_ASAP7_75t_L   g00948(.A1(new_n942), .A2(new_n1030), .B(new_n1033), .C(new_n1204), .Y(new_n1205));
  INVx1_ASAP7_75t_L         g00949(.A(new_n1205), .Y(new_n1206));
  O2A1O1Ixp33_ASAP7_75t_L   g00950(.A1(new_n943), .A2(new_n946), .B(new_n1032), .C(new_n1031), .Y(new_n1207));
  NAND2xp33_ASAP7_75t_L     g00951(.A(new_n1204), .B(new_n1207), .Y(new_n1208));
  NAND2xp33_ASAP7_75t_L     g00952(.A(new_n1208), .B(new_n1206), .Y(new_n1209));
  AOI22xp33_ASAP7_75t_L     g00953(.A1(\b[15] ), .A2(new_n282), .B1(\b[17] ), .B2(new_n303), .Y(new_n1210));
  OAI221xp5_ASAP7_75t_L     g00954(.A1(new_n291), .A2(new_n1030), .B1(new_n268), .B2(new_n1209), .C(new_n1210), .Y(new_n1211));
  XNOR2x2_ASAP7_75t_L       g00955(.A(\a[2] ), .B(new_n1211), .Y(new_n1212));
  NAND3xp33_ASAP7_75t_L     g00956(.A(new_n1197), .B(new_n1199), .C(new_n1212), .Y(new_n1213));
  NOR3xp33_ASAP7_75t_L      g00957(.A(new_n1198), .B(new_n1192), .C(new_n1195), .Y(new_n1214));
  A2O1A1Ixp33_ASAP7_75t_L   g00958(.A1(new_n1017), .A2(new_n1039), .B(new_n1115), .C(new_n1114), .Y(new_n1215));
  NOR2xp33_ASAP7_75t_L      g00959(.A(new_n1196), .B(new_n1215), .Y(new_n1216));
  INVx1_ASAP7_75t_L         g00960(.A(new_n1212), .Y(new_n1217));
  OAI21xp33_ASAP7_75t_L     g00961(.A1(new_n1214), .A2(new_n1216), .B(new_n1217), .Y(new_n1218));
  NAND2xp33_ASAP7_75t_L     g00962(.A(new_n1213), .B(new_n1218), .Y(new_n1219));
  NOR3xp33_ASAP7_75t_L      g00963(.A(new_n1116), .B(new_n1120), .C(new_n1038), .Y(new_n1220));
  A2O1A1Ixp33_ASAP7_75t_L   g00964(.A1(new_n1128), .A2(new_n1125), .B(new_n1220), .C(new_n1219), .Y(new_n1221));
  OR3x1_ASAP7_75t_L         g00965(.A(new_n1127), .B(new_n1219), .C(new_n1220), .Y(new_n1222));
  AND2x2_ASAP7_75t_L        g00966(.A(new_n1221), .B(new_n1222), .Y(\f[17] ));
  OAI21xp33_ASAP7_75t_L     g00967(.A1(new_n1190), .A2(new_n1194), .B(new_n1134), .Y(new_n1224));
  A2O1A1O1Ixp25_ASAP7_75t_L g00968(.A1(new_n1110), .A2(new_n1119), .B(new_n1131), .C(new_n1224), .D(new_n1195), .Y(new_n1225));
  AOI22xp33_ASAP7_75t_L     g00969(.A1(new_n344), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n370), .Y(new_n1226));
  OAI221xp5_ASAP7_75t_L     g00970(.A1(new_n429), .A2(new_n869), .B1(new_n366), .B2(new_n950), .C(new_n1226), .Y(new_n1227));
  XNOR2x2_ASAP7_75t_L       g00971(.A(\a[5] ), .B(new_n1227), .Y(new_n1228));
  NOR3xp33_ASAP7_75t_L      g00972(.A(new_n1178), .B(new_n1181), .C(new_n1139), .Y(new_n1229));
  A2O1A1O1Ixp25_ASAP7_75t_L g00973(.A1(new_n1102), .A2(new_n1108), .B(new_n1136), .C(new_n1182), .D(new_n1229), .Y(new_n1230));
  INVx1_ASAP7_75t_L         g00974(.A(new_n767), .Y(new_n1231));
  NOR2xp33_ASAP7_75t_L      g00975(.A(new_n764), .B(new_n1231), .Y(new_n1232));
  NOR2xp33_ASAP7_75t_L      g00976(.A(new_n679), .B(new_n468), .Y(new_n1233));
  AOI22xp33_ASAP7_75t_L     g00977(.A1(new_n444), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n471), .Y(new_n1234));
  INVx1_ASAP7_75t_L         g00978(.A(new_n1234), .Y(new_n1235));
  AOI211xp5_ASAP7_75t_L     g00979(.A1(new_n1232), .A2(new_n441), .B(new_n1233), .C(new_n1235), .Y(new_n1236));
  NAND2xp33_ASAP7_75t_L     g00980(.A(\a[8] ), .B(new_n1236), .Y(new_n1237));
  OAI21xp33_ASAP7_75t_L     g00981(.A1(new_n469), .A2(new_n768), .B(new_n1234), .Y(new_n1238));
  A2O1A1Ixp33_ASAP7_75t_L   g00982(.A1(\b[11] ), .A2(new_n447), .B(new_n1238), .C(new_n435), .Y(new_n1239));
  NAND2xp33_ASAP7_75t_L     g00983(.A(new_n1239), .B(new_n1237), .Y(new_n1240));
  OAI21xp33_ASAP7_75t_L     g00984(.A1(new_n1175), .A2(new_n1141), .B(new_n1176), .Y(new_n1241));
  NAND5xp2_ASAP7_75t_L      g00985(.A(\a[17] ), .B(new_n1074), .C(new_n1077), .D(new_n1081), .E(new_n972), .Y(new_n1242));
  INVx1_ASAP7_75t_L         g00986(.A(\a[18] ), .Y(new_n1243));
  NAND2xp33_ASAP7_75t_L     g00987(.A(\a[17] ), .B(new_n1243), .Y(new_n1244));
  NAND2xp33_ASAP7_75t_L     g00988(.A(\a[18] ), .B(new_n1071), .Y(new_n1245));
  AND2x2_ASAP7_75t_L        g00989(.A(new_n1244), .B(new_n1245), .Y(new_n1246));
  NOR2xp33_ASAP7_75t_L      g00990(.A(new_n258), .B(new_n1246), .Y(new_n1247));
  OAI31xp33_ASAP7_75t_L     g00991(.A1(new_n1242), .A2(new_n1159), .A3(new_n1155), .B(new_n1247), .Y(new_n1248));
  NOR2xp33_ASAP7_75t_L      g00992(.A(new_n1071), .B(new_n969), .Y(new_n1249));
  AND4x1_ASAP7_75t_L        g00993(.A(new_n1074), .B(new_n1249), .C(new_n1077), .D(new_n1081), .Y(new_n1250));
  INVx1_ASAP7_75t_L         g00994(.A(new_n1155), .Y(new_n1251));
  NOR2xp33_ASAP7_75t_L      g00995(.A(new_n280), .B(new_n1156), .Y(new_n1252));
  INVx1_ASAP7_75t_L         g00996(.A(new_n1158), .Y(new_n1253));
  AOI221xp5_ASAP7_75t_L     g00997(.A1(\b[2] ), .A2(new_n1076), .B1(\b[0] ), .B2(new_n1253), .C(new_n1252), .Y(new_n1254));
  NAND2xp33_ASAP7_75t_L     g00998(.A(new_n1245), .B(new_n1244), .Y(new_n1255));
  NAND2xp33_ASAP7_75t_L     g00999(.A(\b[0] ), .B(new_n1255), .Y(new_n1256));
  NAND4xp25_ASAP7_75t_L     g01000(.A(new_n1250), .B(new_n1256), .C(new_n1254), .D(new_n1251), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g01001(.A(new_n276), .B(new_n1154), .Y(new_n1258));
  NAND3xp33_ASAP7_75t_L     g01002(.A(new_n1078), .B(new_n1070), .C(new_n1072), .Y(new_n1259));
  OAI22xp33_ASAP7_75t_L     g01003(.A1(new_n1158), .A2(new_n261), .B1(new_n298), .B2(new_n1259), .Y(new_n1260));
  AOI211xp5_ASAP7_75t_L     g01004(.A1(new_n406), .A2(new_n1073), .B(new_n1258), .C(new_n1260), .Y(new_n1261));
  NAND2xp33_ASAP7_75t_L     g01005(.A(\a[17] ), .B(new_n1261), .Y(new_n1262));
  AO21x2_ASAP7_75t_L        g01006(.A1(new_n406), .A2(new_n1073), .B(new_n1260), .Y(new_n1263));
  A2O1A1Ixp33_ASAP7_75t_L   g01007(.A1(\b[2] ), .A2(new_n1080), .B(new_n1263), .C(new_n1071), .Y(new_n1264));
  AO22x1_ASAP7_75t_L        g01008(.A1(new_n1248), .A2(new_n1257), .B1(new_n1262), .B2(new_n1264), .Y(new_n1265));
  NAND4xp25_ASAP7_75t_L     g01009(.A(new_n1264), .B(new_n1248), .C(new_n1257), .D(new_n1262), .Y(new_n1266));
  NAND2xp33_ASAP7_75t_L     g01010(.A(\b[5] ), .B(new_n815), .Y(new_n1267));
  NAND2xp33_ASAP7_75t_L     g01011(.A(new_n808), .B(new_n526), .Y(new_n1268));
  AOI22xp33_ASAP7_75t_L     g01012(.A1(new_n811), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n900), .Y(new_n1269));
  NAND4xp25_ASAP7_75t_L     g01013(.A(new_n1268), .B(\a[14] ), .C(new_n1267), .D(new_n1269), .Y(new_n1270));
  NAND3xp33_ASAP7_75t_L     g01014(.A(new_n1268), .B(new_n1267), .C(new_n1269), .Y(new_n1271));
  NAND2xp33_ASAP7_75t_L     g01015(.A(new_n806), .B(new_n1271), .Y(new_n1272));
  NAND4xp25_ASAP7_75t_L     g01016(.A(new_n1272), .B(new_n1265), .C(new_n1266), .D(new_n1270), .Y(new_n1273));
  AO22x1_ASAP7_75t_L        g01017(.A1(new_n1266), .A2(new_n1265), .B1(new_n1270), .B2(new_n1272), .Y(new_n1274));
  NAND2xp33_ASAP7_75t_L     g01018(.A(new_n1273), .B(new_n1274), .Y(new_n1275));
  OAI21xp33_ASAP7_75t_L     g01019(.A1(new_n1168), .A2(new_n1171), .B(new_n1172), .Y(new_n1276));
  NOR2xp33_ASAP7_75t_L      g01020(.A(new_n1276), .B(new_n1275), .Y(new_n1277));
  AND4x1_ASAP7_75t_L        g01021(.A(new_n1265), .B(new_n1272), .C(new_n1266), .D(new_n1270), .Y(new_n1278));
  AOI22xp33_ASAP7_75t_L     g01022(.A1(new_n1265), .A2(new_n1266), .B1(new_n1270), .B2(new_n1272), .Y(new_n1279));
  NOR2xp33_ASAP7_75t_L      g01023(.A(new_n1279), .B(new_n1278), .Y(new_n1280));
  O2A1O1Ixp33_ASAP7_75t_L   g01024(.A1(new_n1171), .A2(new_n1168), .B(new_n1172), .C(new_n1280), .Y(new_n1281));
  AOI22xp33_ASAP7_75t_L     g01025(.A1(\b[7] ), .A2(new_n651), .B1(\b[9] ), .B2(new_n581), .Y(new_n1282));
  OAI221xp5_ASAP7_75t_L     g01026(.A1(new_n821), .A2(new_n488), .B1(new_n577), .B2(new_n548), .C(new_n1282), .Y(new_n1283));
  NOR2xp33_ASAP7_75t_L      g01027(.A(new_n574), .B(new_n1283), .Y(new_n1284));
  AND2x2_ASAP7_75t_L        g01028(.A(new_n574), .B(new_n1283), .Y(new_n1285));
  OAI22xp33_ASAP7_75t_L     g01029(.A1(new_n1281), .A2(new_n1277), .B1(new_n1285), .B2(new_n1284), .Y(new_n1286));
  AOI21xp33_ASAP7_75t_L     g01030(.A1(new_n1146), .A2(new_n1173), .B(new_n1165), .Y(new_n1287));
  NAND2xp33_ASAP7_75t_L     g01031(.A(new_n1287), .B(new_n1280), .Y(new_n1288));
  A2O1A1Ixp33_ASAP7_75t_L   g01032(.A1(new_n1173), .A2(new_n1146), .B(new_n1165), .C(new_n1275), .Y(new_n1289));
  OR2x4_ASAP7_75t_L         g01033(.A(new_n574), .B(new_n1283), .Y(new_n1290));
  NAND2xp33_ASAP7_75t_L     g01034(.A(new_n574), .B(new_n1283), .Y(new_n1291));
  NAND4xp25_ASAP7_75t_L     g01035(.A(new_n1289), .B(new_n1291), .C(new_n1288), .D(new_n1290), .Y(new_n1292));
  NAND3xp33_ASAP7_75t_L     g01036(.A(new_n1241), .B(new_n1286), .C(new_n1292), .Y(new_n1293));
  NAND2xp33_ASAP7_75t_L     g01037(.A(new_n1054), .B(new_n999), .Y(new_n1294));
  A2O1A1O1Ixp25_ASAP7_75t_L g01038(.A1(new_n1099), .A2(new_n1294), .B(new_n1097), .C(new_n1180), .D(new_n1177), .Y(new_n1295));
  NAND2xp33_ASAP7_75t_L     g01039(.A(new_n1292), .B(new_n1286), .Y(new_n1296));
  NAND2xp33_ASAP7_75t_L     g01040(.A(new_n1295), .B(new_n1296), .Y(new_n1297));
  AOI21xp33_ASAP7_75t_L     g01041(.A1(new_n1297), .A2(new_n1293), .B(new_n1240), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g01042(.A(new_n1295), .B(new_n1296), .Y(new_n1299));
  AOI21xp33_ASAP7_75t_L     g01043(.A1(new_n1292), .A2(new_n1286), .B(new_n1241), .Y(new_n1300));
  AOI211xp5_ASAP7_75t_L     g01044(.A1(new_n1239), .A2(new_n1237), .B(new_n1300), .C(new_n1299), .Y(new_n1301));
  NOR3xp33_ASAP7_75t_L      g01045(.A(new_n1230), .B(new_n1298), .C(new_n1301), .Y(new_n1302));
  INVx1_ASAP7_75t_L         g01046(.A(new_n1230), .Y(new_n1303));
  NOR2xp33_ASAP7_75t_L      g01047(.A(new_n1298), .B(new_n1301), .Y(new_n1304));
  NOR2xp33_ASAP7_75t_L      g01048(.A(new_n1303), .B(new_n1304), .Y(new_n1305));
  NOR3xp33_ASAP7_75t_L      g01049(.A(new_n1305), .B(new_n1302), .C(new_n1228), .Y(new_n1306));
  OA21x2_ASAP7_75t_L        g01050(.A1(new_n1302), .A2(new_n1305), .B(new_n1228), .Y(new_n1307));
  NOR3xp33_ASAP7_75t_L      g01051(.A(new_n1225), .B(new_n1307), .C(new_n1306), .Y(new_n1308));
  OAI21xp33_ASAP7_75t_L     g01052(.A1(new_n1306), .A2(new_n1307), .B(new_n1225), .Y(new_n1309));
  INVx1_ASAP7_75t_L         g01053(.A(new_n1309), .Y(new_n1310));
  INVx1_ASAP7_75t_L         g01054(.A(new_n1202), .Y(new_n1311));
  NOR2xp33_ASAP7_75t_L      g01055(.A(\b[17] ), .B(\b[18] ), .Y(new_n1312));
  INVx1_ASAP7_75t_L         g01056(.A(\b[18] ), .Y(new_n1313));
  NOR2xp33_ASAP7_75t_L      g01057(.A(new_n1201), .B(new_n1313), .Y(new_n1314));
  NOR2xp33_ASAP7_75t_L      g01058(.A(new_n1312), .B(new_n1314), .Y(new_n1315));
  INVx1_ASAP7_75t_L         g01059(.A(new_n1315), .Y(new_n1316));
  O2A1O1Ixp33_ASAP7_75t_L   g01060(.A1(new_n1204), .A2(new_n1207), .B(new_n1311), .C(new_n1316), .Y(new_n1317));
  NOR3xp33_ASAP7_75t_L      g01061(.A(new_n1205), .B(new_n1315), .C(new_n1202), .Y(new_n1318));
  NOR2xp33_ASAP7_75t_L      g01062(.A(new_n1317), .B(new_n1318), .Y(new_n1319));
  INVx1_ASAP7_75t_L         g01063(.A(new_n1319), .Y(new_n1320));
  AOI22xp33_ASAP7_75t_L     g01064(.A1(\b[16] ), .A2(new_n282), .B1(\b[18] ), .B2(new_n303), .Y(new_n1321));
  OAI221xp5_ASAP7_75t_L     g01065(.A1(new_n291), .A2(new_n1201), .B1(new_n268), .B2(new_n1320), .C(new_n1321), .Y(new_n1322));
  XNOR2x2_ASAP7_75t_L       g01066(.A(\a[2] ), .B(new_n1322), .Y(new_n1323));
  INVx1_ASAP7_75t_L         g01067(.A(new_n1323), .Y(new_n1324));
  NOR3xp33_ASAP7_75t_L      g01068(.A(new_n1310), .B(new_n1324), .C(new_n1308), .Y(new_n1325));
  INVx1_ASAP7_75t_L         g01069(.A(new_n1308), .Y(new_n1326));
  AOI21xp33_ASAP7_75t_L     g01070(.A1(new_n1326), .A2(new_n1309), .B(new_n1323), .Y(new_n1327));
  NOR2xp33_ASAP7_75t_L      g01071(.A(new_n1325), .B(new_n1327), .Y(new_n1328));
  NOR3xp33_ASAP7_75t_L      g01072(.A(new_n1216), .B(new_n1214), .C(new_n1212), .Y(new_n1329));
  A2O1A1O1Ixp25_ASAP7_75t_L g01073(.A1(new_n1125), .A2(new_n1128), .B(new_n1220), .C(new_n1219), .D(new_n1329), .Y(new_n1330));
  XOR2x2_ASAP7_75t_L        g01074(.A(new_n1328), .B(new_n1330), .Y(\f[18] ));
  OR3x1_ASAP7_75t_L         g01075(.A(new_n1305), .B(new_n1228), .C(new_n1302), .Y(new_n1332));
  NAND3xp33_ASAP7_75t_L     g01076(.A(new_n1297), .B(new_n1293), .C(new_n1240), .Y(new_n1333));
  NAND2xp33_ASAP7_75t_L     g01077(.A(new_n1270), .B(new_n1272), .Y(new_n1334));
  NAND3xp33_ASAP7_75t_L     g01078(.A(new_n1334), .B(new_n1266), .C(new_n1265), .Y(new_n1335));
  A2O1A1Ixp33_ASAP7_75t_L   g01079(.A1(new_n1274), .A2(new_n1273), .B(new_n1276), .C(new_n1335), .Y(new_n1336));
  OAI22xp33_ASAP7_75t_L     g01080(.A1(new_n978), .A2(new_n354), .B1(new_n420), .B2(new_n977), .Y(new_n1337));
  INVx1_ASAP7_75t_L         g01081(.A(new_n1337), .Y(new_n1338));
  OAI221xp5_ASAP7_75t_L     g01082(.A1(new_n904), .A2(new_n418), .B1(new_n898), .B2(new_n425), .C(new_n1338), .Y(new_n1339));
  NOR2xp33_ASAP7_75t_L      g01083(.A(new_n806), .B(new_n1339), .Y(new_n1340));
  NAND2xp33_ASAP7_75t_L     g01084(.A(new_n806), .B(new_n1339), .Y(new_n1341));
  INVx1_ASAP7_75t_L         g01085(.A(new_n1341), .Y(new_n1342));
  AOI22xp33_ASAP7_75t_L     g01086(.A1(new_n1248), .A2(new_n1257), .B1(new_n1262), .B2(new_n1264), .Y(new_n1343));
  NOR3xp33_ASAP7_75t_L      g01087(.A(new_n1242), .B(new_n1155), .C(new_n1159), .Y(new_n1344));
  NAND2xp33_ASAP7_75t_L     g01088(.A(new_n1247), .B(new_n1344), .Y(new_n1345));
  INVx1_ASAP7_75t_L         g01089(.A(new_n1345), .Y(new_n1346));
  NOR2xp33_ASAP7_75t_L      g01090(.A(new_n298), .B(new_n1154), .Y(new_n1347));
  NOR3xp33_ASAP7_75t_L      g01091(.A(new_n326), .B(new_n328), .C(new_n1156), .Y(new_n1348));
  OAI22xp33_ASAP7_75t_L     g01092(.A1(new_n1158), .A2(new_n276), .B1(new_n324), .B2(new_n1259), .Y(new_n1349));
  NOR4xp25_ASAP7_75t_L      g01093(.A(new_n1348), .B(new_n1349), .C(new_n1071), .D(new_n1347), .Y(new_n1350));
  INVx1_ASAP7_75t_L         g01094(.A(new_n1350), .Y(new_n1351));
  OAI31xp33_ASAP7_75t_L     g01095(.A1(new_n1348), .A2(new_n1349), .A3(new_n1347), .B(new_n1071), .Y(new_n1352));
  NAND2xp33_ASAP7_75t_L     g01096(.A(\a[20] ), .B(new_n1247), .Y(new_n1353));
  INVx1_ASAP7_75t_L         g01097(.A(\a[19] ), .Y(new_n1354));
  NAND2xp33_ASAP7_75t_L     g01098(.A(\a[20] ), .B(new_n1354), .Y(new_n1355));
  INVx1_ASAP7_75t_L         g01099(.A(\a[20] ), .Y(new_n1356));
  NAND2xp33_ASAP7_75t_L     g01100(.A(\a[19] ), .B(new_n1356), .Y(new_n1357));
  NAND2xp33_ASAP7_75t_L     g01101(.A(new_n1357), .B(new_n1355), .Y(new_n1358));
  NAND2xp33_ASAP7_75t_L     g01102(.A(new_n1358), .B(new_n1255), .Y(new_n1359));
  NOR2xp33_ASAP7_75t_L      g01103(.A(new_n1358), .B(new_n1246), .Y(new_n1360));
  XNOR2x2_ASAP7_75t_L       g01104(.A(\a[19] ), .B(\a[18] ), .Y(new_n1361));
  NOR2xp33_ASAP7_75t_L      g01105(.A(new_n1361), .B(new_n1255), .Y(new_n1362));
  AOI22xp33_ASAP7_75t_L     g01106(.A1(\b[0] ), .A2(new_n1362), .B1(\b[1] ), .B2(new_n1360), .Y(new_n1363));
  O2A1O1Ixp33_ASAP7_75t_L   g01107(.A1(new_n1359), .A2(new_n270), .B(new_n1363), .C(new_n1353), .Y(new_n1364));
  AOI21xp33_ASAP7_75t_L     g01108(.A1(new_n1357), .A2(new_n1355), .B(new_n1246), .Y(new_n1365));
  NAND2xp33_ASAP7_75t_L     g01109(.A(new_n269), .B(new_n1365), .Y(new_n1366));
  AND3x1_ASAP7_75t_L        g01110(.A(new_n1363), .B(new_n1366), .C(new_n1353), .Y(new_n1367));
  NOR2xp33_ASAP7_75t_L      g01111(.A(new_n1364), .B(new_n1367), .Y(new_n1368));
  NAND3xp33_ASAP7_75t_L     g01112(.A(new_n1368), .B(new_n1352), .C(new_n1351), .Y(new_n1369));
  INVx1_ASAP7_75t_L         g01113(.A(new_n1352), .Y(new_n1370));
  NOR2xp33_ASAP7_75t_L      g01114(.A(new_n1356), .B(new_n1256), .Y(new_n1371));
  NAND3xp33_ASAP7_75t_L     g01115(.A(new_n1255), .B(new_n1355), .C(new_n1357), .Y(new_n1372));
  OR2x4_ASAP7_75t_L         g01116(.A(new_n1361), .B(new_n1255), .Y(new_n1373));
  OAI22xp33_ASAP7_75t_L     g01117(.A1(new_n1373), .A2(new_n258), .B1(new_n261), .B2(new_n1372), .Y(new_n1374));
  A2O1A1Ixp33_ASAP7_75t_L   g01118(.A1(new_n269), .A2(new_n1365), .B(new_n1374), .C(new_n1371), .Y(new_n1375));
  NAND3xp33_ASAP7_75t_L     g01119(.A(new_n1363), .B(new_n1366), .C(new_n1353), .Y(new_n1376));
  NAND2xp33_ASAP7_75t_L     g01120(.A(new_n1376), .B(new_n1375), .Y(new_n1377));
  OAI21xp33_ASAP7_75t_L     g01121(.A1(new_n1350), .A2(new_n1370), .B(new_n1377), .Y(new_n1378));
  NAND2xp33_ASAP7_75t_L     g01122(.A(new_n1378), .B(new_n1369), .Y(new_n1379));
  OAI21xp33_ASAP7_75t_L     g01123(.A1(new_n1343), .A2(new_n1346), .B(new_n1379), .Y(new_n1380));
  NAND4xp25_ASAP7_75t_L     g01124(.A(new_n1265), .B(new_n1378), .C(new_n1369), .D(new_n1345), .Y(new_n1381));
  OAI211xp5_ASAP7_75t_L     g01125(.A1(new_n1342), .A2(new_n1340), .B(new_n1380), .C(new_n1381), .Y(new_n1382));
  INVx1_ASAP7_75t_L         g01126(.A(new_n1339), .Y(new_n1383));
  NAND2xp33_ASAP7_75t_L     g01127(.A(\a[14] ), .B(new_n1383), .Y(new_n1384));
  XNOR2x2_ASAP7_75t_L       g01128(.A(\a[17] ), .B(new_n1261), .Y(new_n1385));
  MAJIxp5_ASAP7_75t_L       g01129(.A(new_n1385), .B(new_n1247), .C(new_n1344), .Y(new_n1386));
  AOI21xp33_ASAP7_75t_L     g01130(.A1(new_n1378), .A2(new_n1369), .B(new_n1386), .Y(new_n1387));
  NOR3xp33_ASAP7_75t_L      g01131(.A(new_n1379), .B(new_n1346), .C(new_n1343), .Y(new_n1388));
  OAI211xp5_ASAP7_75t_L     g01132(.A1(new_n1388), .A2(new_n1387), .B(new_n1341), .C(new_n1384), .Y(new_n1389));
  NAND3xp33_ASAP7_75t_L     g01133(.A(new_n1336), .B(new_n1382), .C(new_n1389), .Y(new_n1390));
  OAI221xp5_ASAP7_75t_L     g01134(.A1(new_n1168), .A2(new_n1171), .B1(new_n1279), .B2(new_n1278), .C(new_n1172), .Y(new_n1391));
  AOI211xp5_ASAP7_75t_L     g01135(.A1(new_n1341), .A2(new_n1384), .B(new_n1388), .C(new_n1387), .Y(new_n1392));
  AOI211xp5_ASAP7_75t_L     g01136(.A1(new_n1380), .A2(new_n1381), .B(new_n1342), .C(new_n1340), .Y(new_n1393));
  OAI211xp5_ASAP7_75t_L     g01137(.A1(new_n1392), .A2(new_n1393), .B(new_n1391), .C(new_n1335), .Y(new_n1394));
  AOI22xp33_ASAP7_75t_L     g01138(.A1(\b[8] ), .A2(new_n651), .B1(\b[10] ), .B2(new_n581), .Y(new_n1395));
  OAI221xp5_ASAP7_75t_L     g01139(.A1(new_n821), .A2(new_n540), .B1(new_n577), .B2(new_n624), .C(new_n1395), .Y(new_n1396));
  XNOR2x2_ASAP7_75t_L       g01140(.A(\a[11] ), .B(new_n1396), .Y(new_n1397));
  NAND3xp33_ASAP7_75t_L     g01141(.A(new_n1390), .B(new_n1394), .C(new_n1397), .Y(new_n1398));
  AO21x2_ASAP7_75t_L        g01142(.A1(new_n1394), .A2(new_n1390), .B(new_n1397), .Y(new_n1399));
  AOI22xp33_ASAP7_75t_L     g01143(.A1(new_n1290), .A2(new_n1291), .B1(new_n1288), .B2(new_n1289), .Y(new_n1400));
  A2O1A1O1Ixp25_ASAP7_75t_L g01144(.A1(new_n1180), .A2(new_n1179), .B(new_n1177), .C(new_n1292), .D(new_n1400), .Y(new_n1401));
  AND3x1_ASAP7_75t_L        g01145(.A(new_n1401), .B(new_n1399), .C(new_n1398), .Y(new_n1402));
  AOI21xp33_ASAP7_75t_L     g01146(.A1(new_n1399), .A2(new_n1398), .B(new_n1401), .Y(new_n1403));
  AOI22xp33_ASAP7_75t_L     g01147(.A1(new_n444), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n471), .Y(new_n1404));
  OAI221xp5_ASAP7_75t_L     g01148(.A1(new_n468), .A2(new_n760), .B1(new_n469), .B2(new_n790), .C(new_n1404), .Y(new_n1405));
  NOR2xp33_ASAP7_75t_L      g01149(.A(new_n435), .B(new_n1405), .Y(new_n1406));
  AND2x2_ASAP7_75t_L        g01150(.A(new_n435), .B(new_n1405), .Y(new_n1407));
  NOR2xp33_ASAP7_75t_L      g01151(.A(new_n1406), .B(new_n1407), .Y(new_n1408));
  OAI21xp33_ASAP7_75t_L     g01152(.A1(new_n1403), .A2(new_n1402), .B(new_n1408), .Y(new_n1409));
  NAND3xp33_ASAP7_75t_L     g01153(.A(new_n1401), .B(new_n1399), .C(new_n1398), .Y(new_n1410));
  AO21x2_ASAP7_75t_L        g01154(.A1(new_n1398), .A2(new_n1399), .B(new_n1401), .Y(new_n1411));
  OAI211xp5_ASAP7_75t_L     g01155(.A1(new_n1406), .A2(new_n1407), .B(new_n1411), .C(new_n1410), .Y(new_n1412));
  NAND2xp33_ASAP7_75t_L     g01156(.A(new_n1409), .B(new_n1412), .Y(new_n1413));
  O2A1O1Ixp33_ASAP7_75t_L   g01157(.A1(new_n1230), .A2(new_n1298), .B(new_n1333), .C(new_n1413), .Y(new_n1414));
  OAI21xp33_ASAP7_75t_L     g01158(.A1(new_n1298), .A2(new_n1230), .B(new_n1333), .Y(new_n1415));
  AOI21xp33_ASAP7_75t_L     g01159(.A1(new_n1412), .A2(new_n1409), .B(new_n1415), .Y(new_n1416));
  AOI22xp33_ASAP7_75t_L     g01160(.A1(new_n344), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n370), .Y(new_n1417));
  OAI221xp5_ASAP7_75t_L     g01161(.A1(new_n429), .A2(new_n942), .B1(new_n366), .B2(new_n1035), .C(new_n1417), .Y(new_n1418));
  XNOR2x2_ASAP7_75t_L       g01162(.A(\a[5] ), .B(new_n1418), .Y(new_n1419));
  INVx1_ASAP7_75t_L         g01163(.A(new_n1419), .Y(new_n1420));
  NOR3xp33_ASAP7_75t_L      g01164(.A(new_n1414), .B(new_n1416), .C(new_n1420), .Y(new_n1421));
  NAND3xp33_ASAP7_75t_L     g01165(.A(new_n1415), .B(new_n1412), .C(new_n1409), .Y(new_n1422));
  OA21x2_ASAP7_75t_L        g01166(.A1(new_n1298), .A2(new_n1230), .B(new_n1333), .Y(new_n1423));
  NAND2xp33_ASAP7_75t_L     g01167(.A(new_n1413), .B(new_n1423), .Y(new_n1424));
  AOI21xp33_ASAP7_75t_L     g01168(.A1(new_n1424), .A2(new_n1422), .B(new_n1419), .Y(new_n1425));
  NOR2xp33_ASAP7_75t_L      g01169(.A(new_n1425), .B(new_n1421), .Y(new_n1426));
  NAND3xp33_ASAP7_75t_L     g01170(.A(new_n1326), .B(new_n1332), .C(new_n1426), .Y(new_n1427));
  INVx1_ASAP7_75t_L         g01171(.A(new_n1426), .Y(new_n1428));
  OAI21xp33_ASAP7_75t_L     g01172(.A1(new_n1307), .A2(new_n1225), .B(new_n1332), .Y(new_n1429));
  NAND2xp33_ASAP7_75t_L     g01173(.A(new_n1429), .B(new_n1428), .Y(new_n1430));
  NOR2xp33_ASAP7_75t_L      g01174(.A(\b[18] ), .B(\b[19] ), .Y(new_n1431));
  INVx1_ASAP7_75t_L         g01175(.A(\b[19] ), .Y(new_n1432));
  NOR2xp33_ASAP7_75t_L      g01176(.A(new_n1313), .B(new_n1432), .Y(new_n1433));
  NOR2xp33_ASAP7_75t_L      g01177(.A(new_n1431), .B(new_n1433), .Y(new_n1434));
  A2O1A1Ixp33_ASAP7_75t_L   g01178(.A1(\b[18] ), .A2(\b[17] ), .B(new_n1317), .C(new_n1434), .Y(new_n1435));
  NOR3xp33_ASAP7_75t_L      g01179(.A(new_n1317), .B(new_n1434), .C(new_n1314), .Y(new_n1436));
  INVx1_ASAP7_75t_L         g01180(.A(new_n1436), .Y(new_n1437));
  NAND2xp33_ASAP7_75t_L     g01181(.A(new_n1435), .B(new_n1437), .Y(new_n1438));
  AOI22xp33_ASAP7_75t_L     g01182(.A1(\b[17] ), .A2(new_n282), .B1(\b[19] ), .B2(new_n303), .Y(new_n1439));
  OAI221xp5_ASAP7_75t_L     g01183(.A1(new_n291), .A2(new_n1313), .B1(new_n268), .B2(new_n1438), .C(new_n1439), .Y(new_n1440));
  NOR2xp33_ASAP7_75t_L      g01184(.A(new_n262), .B(new_n1440), .Y(new_n1441));
  AND2x2_ASAP7_75t_L        g01185(.A(new_n262), .B(new_n1440), .Y(new_n1442));
  NOR2xp33_ASAP7_75t_L      g01186(.A(new_n1441), .B(new_n1442), .Y(new_n1443));
  NAND3xp33_ASAP7_75t_L     g01187(.A(new_n1430), .B(new_n1427), .C(new_n1443), .Y(new_n1444));
  NOR2xp33_ASAP7_75t_L      g01188(.A(new_n1429), .B(new_n1428), .Y(new_n1445));
  O2A1O1Ixp33_ASAP7_75t_L   g01189(.A1(new_n1225), .A2(new_n1307), .B(new_n1332), .C(new_n1426), .Y(new_n1446));
  OAI22xp33_ASAP7_75t_L     g01190(.A1(new_n1445), .A2(new_n1446), .B1(new_n1442), .B2(new_n1441), .Y(new_n1447));
  NAND2xp33_ASAP7_75t_L     g01191(.A(new_n1444), .B(new_n1447), .Y(new_n1448));
  INVx1_ASAP7_75t_L         g01192(.A(new_n1448), .Y(new_n1449));
  NAND3xp33_ASAP7_75t_L     g01193(.A(new_n1326), .B(new_n1309), .C(new_n1324), .Y(new_n1450));
  O2A1O1Ixp33_ASAP7_75t_L   g01194(.A1(new_n1330), .A2(new_n1328), .B(new_n1450), .C(new_n1449), .Y(new_n1451));
  OAI21xp33_ASAP7_75t_L     g01195(.A1(new_n1328), .A2(new_n1330), .B(new_n1450), .Y(new_n1452));
  NOR2xp33_ASAP7_75t_L      g01196(.A(new_n1448), .B(new_n1452), .Y(new_n1453));
  NOR2xp33_ASAP7_75t_L      g01197(.A(new_n1453), .B(new_n1451), .Y(\f[19] ));
  NOR3xp33_ASAP7_75t_L      g01198(.A(new_n1445), .B(new_n1446), .C(new_n1443), .Y(new_n1455));
  NOR2xp33_ASAP7_75t_L      g01199(.A(new_n1455), .B(new_n1451), .Y(new_n1456));
  NOR3xp33_ASAP7_75t_L      g01200(.A(new_n1414), .B(new_n1416), .C(new_n1419), .Y(new_n1457));
  AOI22xp33_ASAP7_75t_L     g01201(.A1(new_n344), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n370), .Y(new_n1458));
  OAI221xp5_ASAP7_75t_L     g01202(.A1(new_n429), .A2(new_n1030), .B1(new_n366), .B2(new_n1209), .C(new_n1458), .Y(new_n1459));
  XNOR2x2_ASAP7_75t_L       g01203(.A(new_n338), .B(new_n1459), .Y(new_n1460));
  NAND2xp33_ASAP7_75t_L     g01204(.A(new_n1394), .B(new_n1390), .Y(new_n1461));
  MAJIxp5_ASAP7_75t_L       g01205(.A(new_n1401), .B(new_n1397), .C(new_n1461), .Y(new_n1462));
  AOI22xp33_ASAP7_75t_L     g01206(.A1(\b[9] ), .A2(new_n651), .B1(\b[11] ), .B2(new_n581), .Y(new_n1463));
  OAI221xp5_ASAP7_75t_L     g01207(.A1(new_n821), .A2(new_n617), .B1(new_n577), .B2(new_n685), .C(new_n1463), .Y(new_n1464));
  XNOR2x2_ASAP7_75t_L       g01208(.A(new_n574), .B(new_n1464), .Y(new_n1465));
  A2O1A1Ixp33_ASAP7_75t_L   g01209(.A1(new_n1391), .A2(new_n1335), .B(new_n1393), .C(new_n1382), .Y(new_n1466));
  AOI22xp33_ASAP7_75t_L     g01210(.A1(new_n811), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n900), .Y(new_n1467));
  OAI221xp5_ASAP7_75t_L     g01211(.A1(new_n904), .A2(new_n420), .B1(new_n898), .B2(new_n494), .C(new_n1467), .Y(new_n1468));
  XNOR2x2_ASAP7_75t_L       g01212(.A(\a[14] ), .B(new_n1468), .Y(new_n1469));
  AOI21xp33_ASAP7_75t_L     g01213(.A1(new_n1352), .A2(new_n1351), .B(new_n1377), .Y(new_n1470));
  INVx1_ASAP7_75t_L         g01214(.A(new_n1470), .Y(new_n1471));
  A2O1A1Ixp33_ASAP7_75t_L   g01215(.A1(new_n1369), .A2(new_n1378), .B(new_n1386), .C(new_n1471), .Y(new_n1472));
  NAND2xp33_ASAP7_75t_L     g01216(.A(\b[4] ), .B(new_n1080), .Y(new_n1473));
  INVx1_ASAP7_75t_L         g01217(.A(new_n1473), .Y(new_n1474));
  NOR3xp33_ASAP7_75t_L      g01218(.A(new_n357), .B(new_n358), .C(new_n1156), .Y(new_n1475));
  OAI22xp33_ASAP7_75t_L     g01219(.A1(new_n1158), .A2(new_n298), .B1(new_n354), .B2(new_n1259), .Y(new_n1476));
  NOR4xp25_ASAP7_75t_L      g01220(.A(new_n1475), .B(new_n1071), .C(new_n1476), .D(new_n1474), .Y(new_n1477));
  NOR2xp33_ASAP7_75t_L      g01221(.A(new_n1476), .B(new_n1475), .Y(new_n1478));
  O2A1O1Ixp33_ASAP7_75t_L   g01222(.A1(new_n324), .A2(new_n1154), .B(new_n1478), .C(\a[17] ), .Y(new_n1479));
  AOI21xp33_ASAP7_75t_L     g01223(.A1(new_n1365), .A2(new_n269), .B(new_n1374), .Y(new_n1480));
  NOR2xp33_ASAP7_75t_L      g01224(.A(new_n261), .B(new_n1373), .Y(new_n1481));
  NAND2xp33_ASAP7_75t_L     g01225(.A(\b[2] ), .B(new_n1360), .Y(new_n1482));
  NAND3xp33_ASAP7_75t_L     g01226(.A(new_n1246), .B(new_n1358), .C(new_n1361), .Y(new_n1483));
  OAI221xp5_ASAP7_75t_L     g01227(.A1(new_n258), .A2(new_n1483), .B1(new_n280), .B2(new_n1359), .C(new_n1482), .Y(new_n1484));
  NOR2xp33_ASAP7_75t_L      g01228(.A(new_n1481), .B(new_n1484), .Y(new_n1485));
  A2O1A1Ixp33_ASAP7_75t_L   g01229(.A1(new_n1256), .A2(new_n1480), .B(new_n1356), .C(new_n1485), .Y(new_n1486));
  O2A1O1Ixp33_ASAP7_75t_L   g01230(.A1(new_n258), .A2(new_n1246), .B(new_n1480), .C(new_n1356), .Y(new_n1487));
  A2O1A1Ixp33_ASAP7_75t_L   g01231(.A1(\b[1] ), .A2(new_n1362), .B(new_n1484), .C(new_n1487), .Y(new_n1488));
  AOI211xp5_ASAP7_75t_L     g01232(.A1(new_n1488), .A2(new_n1486), .B(new_n1477), .C(new_n1479), .Y(new_n1489));
  INVx1_ASAP7_75t_L         g01233(.A(new_n1489), .Y(new_n1490));
  OAI211xp5_ASAP7_75t_L     g01234(.A1(new_n1477), .A2(new_n1479), .B(new_n1488), .C(new_n1486), .Y(new_n1491));
  AOI21xp33_ASAP7_75t_L     g01235(.A1(new_n1490), .A2(new_n1491), .B(new_n1472), .Y(new_n1492));
  O2A1O1Ixp33_ASAP7_75t_L   g01236(.A1(new_n1343), .A2(new_n1346), .B(new_n1379), .C(new_n1470), .Y(new_n1493));
  INVx1_ASAP7_75t_L         g01237(.A(new_n1491), .Y(new_n1494));
  NOR3xp33_ASAP7_75t_L      g01238(.A(new_n1493), .B(new_n1489), .C(new_n1494), .Y(new_n1495));
  OAI21xp33_ASAP7_75t_L     g01239(.A1(new_n1495), .A2(new_n1492), .B(new_n1469), .Y(new_n1496));
  INVx1_ASAP7_75t_L         g01240(.A(new_n1469), .Y(new_n1497));
  OAI21xp33_ASAP7_75t_L     g01241(.A1(new_n1489), .A2(new_n1494), .B(new_n1493), .Y(new_n1498));
  NAND3xp33_ASAP7_75t_L     g01242(.A(new_n1490), .B(new_n1472), .C(new_n1491), .Y(new_n1499));
  NAND3xp33_ASAP7_75t_L     g01243(.A(new_n1497), .B(new_n1498), .C(new_n1499), .Y(new_n1500));
  NAND3xp33_ASAP7_75t_L     g01244(.A(new_n1466), .B(new_n1496), .C(new_n1500), .Y(new_n1501));
  INVx1_ASAP7_75t_L         g01245(.A(new_n1335), .Y(new_n1502));
  A2O1A1O1Ixp25_ASAP7_75t_L g01246(.A1(new_n1287), .A2(new_n1275), .B(new_n1502), .C(new_n1389), .D(new_n1392), .Y(new_n1503));
  AOI21xp33_ASAP7_75t_L     g01247(.A1(new_n1499), .A2(new_n1498), .B(new_n1497), .Y(new_n1504));
  NOR3xp33_ASAP7_75t_L      g01248(.A(new_n1492), .B(new_n1495), .C(new_n1469), .Y(new_n1505));
  OAI21xp33_ASAP7_75t_L     g01249(.A1(new_n1504), .A2(new_n1505), .B(new_n1503), .Y(new_n1506));
  AOI21xp33_ASAP7_75t_L     g01250(.A1(new_n1501), .A2(new_n1506), .B(new_n1465), .Y(new_n1507));
  INVx1_ASAP7_75t_L         g01251(.A(new_n1507), .Y(new_n1508));
  NAND3xp33_ASAP7_75t_L     g01252(.A(new_n1501), .B(new_n1465), .C(new_n1506), .Y(new_n1509));
  NAND3xp33_ASAP7_75t_L     g01253(.A(new_n1462), .B(new_n1508), .C(new_n1509), .Y(new_n1510));
  AND3x1_ASAP7_75t_L        g01254(.A(new_n1390), .B(new_n1397), .C(new_n1394), .Y(new_n1511));
  AOI21xp33_ASAP7_75t_L     g01255(.A1(new_n1390), .A2(new_n1394), .B(new_n1397), .Y(new_n1512));
  NOR2xp33_ASAP7_75t_L      g01256(.A(new_n1512), .B(new_n1511), .Y(new_n1513));
  OR2x4_ASAP7_75t_L         g01257(.A(new_n1397), .B(new_n1461), .Y(new_n1514));
  AND3x1_ASAP7_75t_L        g01258(.A(new_n1501), .B(new_n1465), .C(new_n1506), .Y(new_n1515));
  OAI221xp5_ASAP7_75t_L     g01259(.A1(new_n1515), .A2(new_n1507), .B1(new_n1401), .B2(new_n1513), .C(new_n1514), .Y(new_n1516));
  AOI22xp33_ASAP7_75t_L     g01260(.A1(new_n444), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n471), .Y(new_n1517));
  OAI221xp5_ASAP7_75t_L     g01261(.A1(new_n468), .A2(new_n784), .B1(new_n469), .B2(new_n875), .C(new_n1517), .Y(new_n1518));
  XNOR2x2_ASAP7_75t_L       g01262(.A(\a[8] ), .B(new_n1518), .Y(new_n1519));
  NAND3xp33_ASAP7_75t_L     g01263(.A(new_n1510), .B(new_n1516), .C(new_n1519), .Y(new_n1520));
  AO21x2_ASAP7_75t_L        g01264(.A1(new_n1516), .A2(new_n1510), .B(new_n1519), .Y(new_n1521));
  INVx1_ASAP7_75t_L         g01265(.A(new_n1412), .Y(new_n1522));
  AOI21xp33_ASAP7_75t_L     g01266(.A1(new_n1415), .A2(new_n1409), .B(new_n1522), .Y(new_n1523));
  AOI21xp33_ASAP7_75t_L     g01267(.A1(new_n1521), .A2(new_n1520), .B(new_n1523), .Y(new_n1524));
  NAND2xp33_ASAP7_75t_L     g01268(.A(new_n1520), .B(new_n1521), .Y(new_n1525));
  OAI21xp33_ASAP7_75t_L     g01269(.A1(new_n1413), .A2(new_n1423), .B(new_n1412), .Y(new_n1526));
  NOR2xp33_ASAP7_75t_L      g01270(.A(new_n1525), .B(new_n1526), .Y(new_n1527));
  OAI21xp33_ASAP7_75t_L     g01271(.A1(new_n1524), .A2(new_n1527), .B(new_n1460), .Y(new_n1528));
  XNOR2x2_ASAP7_75t_L       g01272(.A(\a[5] ), .B(new_n1459), .Y(new_n1529));
  A2O1A1Ixp33_ASAP7_75t_L   g01273(.A1(new_n1415), .A2(new_n1409), .B(new_n1522), .C(new_n1525), .Y(new_n1530));
  NAND3xp33_ASAP7_75t_L     g01274(.A(new_n1523), .B(new_n1521), .C(new_n1520), .Y(new_n1531));
  NAND3xp33_ASAP7_75t_L     g01275(.A(new_n1530), .B(new_n1529), .C(new_n1531), .Y(new_n1532));
  NAND2xp33_ASAP7_75t_L     g01276(.A(new_n1532), .B(new_n1528), .Y(new_n1533));
  INVx1_ASAP7_75t_L         g01277(.A(new_n1533), .Y(new_n1534));
  A2O1A1Ixp33_ASAP7_75t_L   g01278(.A1(new_n1429), .A2(new_n1428), .B(new_n1457), .C(new_n1534), .Y(new_n1535));
  O2A1O1Ixp33_ASAP7_75t_L   g01279(.A1(new_n1421), .A2(new_n1425), .B(new_n1429), .C(new_n1457), .Y(new_n1536));
  NAND2xp33_ASAP7_75t_L     g01280(.A(new_n1533), .B(new_n1536), .Y(new_n1537));
  NOR2xp33_ASAP7_75t_L      g01281(.A(\b[19] ), .B(\b[20] ), .Y(new_n1538));
  INVx1_ASAP7_75t_L         g01282(.A(\b[20] ), .Y(new_n1539));
  NOR2xp33_ASAP7_75t_L      g01283(.A(new_n1432), .B(new_n1539), .Y(new_n1540));
  NOR2xp33_ASAP7_75t_L      g01284(.A(new_n1538), .B(new_n1540), .Y(new_n1541));
  INVx1_ASAP7_75t_L         g01285(.A(new_n1541), .Y(new_n1542));
  O2A1O1Ixp33_ASAP7_75t_L   g01286(.A1(new_n1313), .A2(new_n1432), .B(new_n1435), .C(new_n1542), .Y(new_n1543));
  INVx1_ASAP7_75t_L         g01287(.A(new_n1543), .Y(new_n1544));
  O2A1O1Ixp33_ASAP7_75t_L   g01288(.A1(new_n1314), .A2(new_n1317), .B(new_n1434), .C(new_n1433), .Y(new_n1545));
  NAND2xp33_ASAP7_75t_L     g01289(.A(new_n1542), .B(new_n1545), .Y(new_n1546));
  NAND2xp33_ASAP7_75t_L     g01290(.A(new_n1546), .B(new_n1544), .Y(new_n1547));
  AOI22xp33_ASAP7_75t_L     g01291(.A1(\b[18] ), .A2(new_n282), .B1(\b[20] ), .B2(new_n303), .Y(new_n1548));
  OAI221xp5_ASAP7_75t_L     g01292(.A1(new_n291), .A2(new_n1432), .B1(new_n268), .B2(new_n1547), .C(new_n1548), .Y(new_n1549));
  XNOR2x2_ASAP7_75t_L       g01293(.A(\a[2] ), .B(new_n1549), .Y(new_n1550));
  AOI21xp33_ASAP7_75t_L     g01294(.A1(new_n1535), .A2(new_n1537), .B(new_n1550), .Y(new_n1551));
  INVx1_ASAP7_75t_L         g01295(.A(new_n1551), .Y(new_n1552));
  NAND3xp33_ASAP7_75t_L     g01296(.A(new_n1535), .B(new_n1537), .C(new_n1550), .Y(new_n1553));
  NAND2xp33_ASAP7_75t_L     g01297(.A(new_n1553), .B(new_n1552), .Y(new_n1554));
  XOR2x2_ASAP7_75t_L        g01298(.A(new_n1554), .B(new_n1456), .Y(\f[20] ));
  NAND2xp33_ASAP7_75t_L     g01299(.A(new_n1516), .B(new_n1510), .Y(new_n1556));
  AOI22xp33_ASAP7_75t_L     g01300(.A1(new_n444), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n471), .Y(new_n1557));
  OAI221xp5_ASAP7_75t_L     g01301(.A1(new_n468), .A2(new_n869), .B1(new_n469), .B2(new_n950), .C(new_n1557), .Y(new_n1558));
  XNOR2x2_ASAP7_75t_L       g01302(.A(\a[8] ), .B(new_n1558), .Y(new_n1559));
  INVx1_ASAP7_75t_L         g01303(.A(new_n1559), .Y(new_n1560));
  AO21x2_ASAP7_75t_L        g01304(.A1(new_n1508), .A2(new_n1462), .B(new_n1515), .Y(new_n1561));
  NAND2xp33_ASAP7_75t_L     g01305(.A(\b[11] ), .B(new_n584), .Y(new_n1562));
  NAND3xp33_ASAP7_75t_L     g01306(.A(new_n765), .B(new_n578), .C(new_n767), .Y(new_n1563));
  AOI22xp33_ASAP7_75t_L     g01307(.A1(\b[10] ), .A2(new_n651), .B1(\b[12] ), .B2(new_n581), .Y(new_n1564));
  AND4x1_ASAP7_75t_L        g01308(.A(new_n1564), .B(new_n1563), .C(new_n1562), .D(\a[11] ), .Y(new_n1565));
  AOI31xp33_ASAP7_75t_L     g01309(.A1(new_n1563), .A2(new_n1562), .A3(new_n1564), .B(\a[11] ), .Y(new_n1566));
  NOR2xp33_ASAP7_75t_L      g01310(.A(new_n1566), .B(new_n1565), .Y(new_n1567));
  A2O1A1O1Ixp25_ASAP7_75t_L g01311(.A1(new_n1389), .A2(new_n1336), .B(new_n1392), .C(new_n1496), .D(new_n1505), .Y(new_n1568));
  NAND4xp25_ASAP7_75t_L     g01312(.A(new_n1363), .B(\a[20] ), .C(new_n1256), .D(new_n1366), .Y(new_n1569));
  INVx1_ASAP7_75t_L         g01313(.A(\a[21] ), .Y(new_n1570));
  NAND2xp33_ASAP7_75t_L     g01314(.A(\a[20] ), .B(new_n1570), .Y(new_n1571));
  NAND2xp33_ASAP7_75t_L     g01315(.A(\a[21] ), .B(new_n1356), .Y(new_n1572));
  NAND2xp33_ASAP7_75t_L     g01316(.A(new_n1572), .B(new_n1571), .Y(new_n1573));
  NAND2xp33_ASAP7_75t_L     g01317(.A(\b[0] ), .B(new_n1573), .Y(new_n1574));
  INVx1_ASAP7_75t_L         g01318(.A(new_n1574), .Y(new_n1575));
  OAI31xp33_ASAP7_75t_L     g01319(.A1(new_n1569), .A2(new_n1484), .A3(new_n1481), .B(new_n1575), .Y(new_n1576));
  A2O1A1Ixp33_ASAP7_75t_L   g01320(.A1(new_n1244), .A2(new_n1245), .B(new_n258), .C(\a[20] ), .Y(new_n1577));
  AOI211xp5_ASAP7_75t_L     g01321(.A1(new_n1365), .A2(new_n269), .B(new_n1577), .C(new_n1374), .Y(new_n1578));
  INVx1_ASAP7_75t_L         g01322(.A(new_n1481), .Y(new_n1579));
  NOR2xp33_ASAP7_75t_L      g01323(.A(new_n280), .B(new_n1359), .Y(new_n1580));
  AND3x1_ASAP7_75t_L        g01324(.A(new_n1246), .B(new_n1361), .C(new_n1358), .Y(new_n1581));
  AOI221xp5_ASAP7_75t_L     g01325(.A1(new_n1360), .A2(\b[2] ), .B1(new_n1581), .B2(\b[0] ), .C(new_n1580), .Y(new_n1582));
  NAND4xp25_ASAP7_75t_L     g01326(.A(new_n1578), .B(new_n1574), .C(new_n1582), .D(new_n1579), .Y(new_n1583));
  NOR2xp33_ASAP7_75t_L      g01327(.A(new_n276), .B(new_n1373), .Y(new_n1584));
  NOR2xp33_ASAP7_75t_L      g01328(.A(new_n1359), .B(new_n302), .Y(new_n1585));
  OAI22xp33_ASAP7_75t_L     g01329(.A1(new_n1483), .A2(new_n261), .B1(new_n298), .B2(new_n1372), .Y(new_n1586));
  OR4x2_ASAP7_75t_L         g01330(.A(new_n1586), .B(new_n1585), .C(new_n1584), .D(new_n1356), .Y(new_n1587));
  OAI31xp33_ASAP7_75t_L     g01331(.A1(new_n1585), .A2(new_n1584), .A3(new_n1586), .B(new_n1356), .Y(new_n1588));
  AOI22xp33_ASAP7_75t_L     g01332(.A1(new_n1587), .A2(new_n1588), .B1(new_n1576), .B2(new_n1583), .Y(new_n1589));
  AND4x1_ASAP7_75t_L        g01333(.A(new_n1583), .B(new_n1576), .C(new_n1588), .D(new_n1587), .Y(new_n1590));
  NAND2xp33_ASAP7_75t_L     g01334(.A(\b[5] ), .B(new_n1080), .Y(new_n1591));
  NAND2xp33_ASAP7_75t_L     g01335(.A(new_n1073), .B(new_n526), .Y(new_n1592));
  AOI22xp33_ASAP7_75t_L     g01336(.A1(new_n1076), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1253), .Y(new_n1593));
  NAND4xp25_ASAP7_75t_L     g01337(.A(new_n1592), .B(\a[17] ), .C(new_n1591), .D(new_n1593), .Y(new_n1594));
  INVx1_ASAP7_75t_L         g01338(.A(new_n1594), .Y(new_n1595));
  AOI31xp33_ASAP7_75t_L     g01339(.A1(new_n1592), .A2(new_n1591), .A3(new_n1593), .B(\a[17] ), .Y(new_n1596));
  NOR4xp25_ASAP7_75t_L      g01340(.A(new_n1595), .B(new_n1590), .C(new_n1589), .D(new_n1596), .Y(new_n1597));
  AO22x1_ASAP7_75t_L        g01341(.A1(new_n1588), .A2(new_n1587), .B1(new_n1576), .B2(new_n1583), .Y(new_n1598));
  NAND4xp25_ASAP7_75t_L     g01342(.A(new_n1583), .B(new_n1576), .C(new_n1587), .D(new_n1588), .Y(new_n1599));
  INVx1_ASAP7_75t_L         g01343(.A(new_n1596), .Y(new_n1600));
  AOI22xp33_ASAP7_75t_L     g01344(.A1(new_n1598), .A2(new_n1599), .B1(new_n1594), .B2(new_n1600), .Y(new_n1601));
  NOR2xp33_ASAP7_75t_L      g01345(.A(new_n1597), .B(new_n1601), .Y(new_n1602));
  OAI311xp33_ASAP7_75t_L    g01346(.A1(new_n1387), .A2(new_n1470), .A3(new_n1494), .B1(new_n1490), .C1(new_n1602), .Y(new_n1603));
  NAND4xp25_ASAP7_75t_L     g01347(.A(new_n1600), .B(new_n1598), .C(new_n1599), .D(new_n1594), .Y(new_n1604));
  OAI22xp33_ASAP7_75t_L     g01348(.A1(new_n1595), .A2(new_n1596), .B1(new_n1589), .B2(new_n1590), .Y(new_n1605));
  NAND2xp33_ASAP7_75t_L     g01349(.A(new_n1605), .B(new_n1604), .Y(new_n1606));
  A2O1A1Ixp33_ASAP7_75t_L   g01350(.A1(new_n1491), .A2(new_n1493), .B(new_n1489), .C(new_n1606), .Y(new_n1607));
  AOI22xp33_ASAP7_75t_L     g01351(.A1(new_n811), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n900), .Y(new_n1608));
  OAI221xp5_ASAP7_75t_L     g01352(.A1(new_n904), .A2(new_n488), .B1(new_n898), .B2(new_n548), .C(new_n1608), .Y(new_n1609));
  OR2x4_ASAP7_75t_L         g01353(.A(new_n806), .B(new_n1609), .Y(new_n1610));
  NAND2xp33_ASAP7_75t_L     g01354(.A(new_n806), .B(new_n1609), .Y(new_n1611));
  AOI22xp33_ASAP7_75t_L     g01355(.A1(new_n1610), .A2(new_n1611), .B1(new_n1607), .B2(new_n1603), .Y(new_n1612));
  NAND4xp25_ASAP7_75t_L     g01356(.A(new_n1603), .B(new_n1610), .C(new_n1607), .D(new_n1611), .Y(new_n1613));
  INVx1_ASAP7_75t_L         g01357(.A(new_n1613), .Y(new_n1614));
  NOR3xp33_ASAP7_75t_L      g01358(.A(new_n1614), .B(new_n1568), .C(new_n1612), .Y(new_n1615));
  OAI21xp33_ASAP7_75t_L     g01359(.A1(new_n1494), .A2(new_n1472), .B(new_n1490), .Y(new_n1616));
  NOR2xp33_ASAP7_75t_L      g01360(.A(new_n1606), .B(new_n1616), .Y(new_n1617));
  O2A1O1Ixp33_ASAP7_75t_L   g01361(.A1(new_n1472), .A2(new_n1494), .B(new_n1490), .C(new_n1602), .Y(new_n1618));
  XNOR2x2_ASAP7_75t_L       g01362(.A(new_n806), .B(new_n1609), .Y(new_n1619));
  OAI21xp33_ASAP7_75t_L     g01363(.A1(new_n1618), .A2(new_n1617), .B(new_n1619), .Y(new_n1620));
  AOI221xp5_ASAP7_75t_L     g01364(.A1(new_n1466), .A2(new_n1496), .B1(new_n1613), .B2(new_n1620), .C(new_n1505), .Y(new_n1621));
  OAI21xp33_ASAP7_75t_L     g01365(.A1(new_n1621), .A2(new_n1615), .B(new_n1567), .Y(new_n1622));
  NOR3xp33_ASAP7_75t_L      g01366(.A(new_n1615), .B(new_n1567), .C(new_n1621), .Y(new_n1623));
  INVx1_ASAP7_75t_L         g01367(.A(new_n1623), .Y(new_n1624));
  NAND3xp33_ASAP7_75t_L     g01368(.A(new_n1561), .B(new_n1622), .C(new_n1624), .Y(new_n1625));
  NOR2xp33_ASAP7_75t_L      g01369(.A(new_n1397), .B(new_n1461), .Y(new_n1626));
  O2A1O1Ixp33_ASAP7_75t_L   g01370(.A1(new_n1626), .A2(new_n1403), .B(new_n1508), .C(new_n1515), .Y(new_n1627));
  INVx1_ASAP7_75t_L         g01371(.A(new_n1622), .Y(new_n1628));
  OAI21xp33_ASAP7_75t_L     g01372(.A1(new_n1628), .A2(new_n1623), .B(new_n1627), .Y(new_n1629));
  NAND3xp33_ASAP7_75t_L     g01373(.A(new_n1625), .B(new_n1560), .C(new_n1629), .Y(new_n1630));
  NOR3xp33_ASAP7_75t_L      g01374(.A(new_n1627), .B(new_n1628), .C(new_n1623), .Y(new_n1631));
  AOI21xp33_ASAP7_75t_L     g01375(.A1(new_n1624), .A2(new_n1622), .B(new_n1561), .Y(new_n1632));
  OAI21xp33_ASAP7_75t_L     g01376(.A1(new_n1632), .A2(new_n1631), .B(new_n1559), .Y(new_n1633));
  NAND2xp33_ASAP7_75t_L     g01377(.A(new_n1630), .B(new_n1633), .Y(new_n1634));
  O2A1O1Ixp33_ASAP7_75t_L   g01378(.A1(new_n1556), .A2(new_n1519), .B(new_n1530), .C(new_n1634), .Y(new_n1635));
  MAJIxp5_ASAP7_75t_L       g01379(.A(new_n1523), .B(new_n1556), .C(new_n1519), .Y(new_n1636));
  AOI21xp33_ASAP7_75t_L     g01380(.A1(new_n1633), .A2(new_n1630), .B(new_n1636), .Y(new_n1637));
  AOI22xp33_ASAP7_75t_L     g01381(.A1(new_n344), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n370), .Y(new_n1638));
  OAI221xp5_ASAP7_75t_L     g01382(.A1(new_n429), .A2(new_n1201), .B1(new_n366), .B2(new_n1320), .C(new_n1638), .Y(new_n1639));
  XNOR2x2_ASAP7_75t_L       g01383(.A(new_n338), .B(new_n1639), .Y(new_n1640));
  NOR3xp33_ASAP7_75t_L      g01384(.A(new_n1635), .B(new_n1637), .C(new_n1640), .Y(new_n1641));
  NAND3xp33_ASAP7_75t_L     g01385(.A(new_n1636), .B(new_n1630), .C(new_n1633), .Y(new_n1642));
  NOR2xp33_ASAP7_75t_L      g01386(.A(new_n1519), .B(new_n1556), .Y(new_n1643));
  A2O1A1O1Ixp25_ASAP7_75t_L g01387(.A1(new_n1409), .A2(new_n1415), .B(new_n1522), .C(new_n1525), .D(new_n1643), .Y(new_n1644));
  NAND2xp33_ASAP7_75t_L     g01388(.A(new_n1634), .B(new_n1644), .Y(new_n1645));
  XNOR2x2_ASAP7_75t_L       g01389(.A(\a[5] ), .B(new_n1639), .Y(new_n1646));
  AOI21xp33_ASAP7_75t_L     g01390(.A1(new_n1645), .A2(new_n1642), .B(new_n1646), .Y(new_n1647));
  NOR2xp33_ASAP7_75t_L      g01391(.A(new_n1647), .B(new_n1641), .Y(new_n1648));
  NOR3xp33_ASAP7_75t_L      g01392(.A(new_n1527), .B(new_n1524), .C(new_n1529), .Y(new_n1649));
  INVx1_ASAP7_75t_L         g01393(.A(new_n1649), .Y(new_n1650));
  A2O1A1Ixp33_ASAP7_75t_L   g01394(.A1(new_n1528), .A2(new_n1532), .B(new_n1536), .C(new_n1650), .Y(new_n1651));
  XOR2x2_ASAP7_75t_L        g01395(.A(new_n1651), .B(new_n1648), .Y(new_n1652));
  INVx1_ASAP7_75t_L         g01396(.A(new_n1540), .Y(new_n1653));
  NOR2xp33_ASAP7_75t_L      g01397(.A(\b[20] ), .B(\b[21] ), .Y(new_n1654));
  INVx1_ASAP7_75t_L         g01398(.A(\b[21] ), .Y(new_n1655));
  NOR2xp33_ASAP7_75t_L      g01399(.A(new_n1539), .B(new_n1655), .Y(new_n1656));
  NOR2xp33_ASAP7_75t_L      g01400(.A(new_n1654), .B(new_n1656), .Y(new_n1657));
  INVx1_ASAP7_75t_L         g01401(.A(new_n1657), .Y(new_n1658));
  O2A1O1Ixp33_ASAP7_75t_L   g01402(.A1(new_n1542), .A2(new_n1545), .B(new_n1653), .C(new_n1658), .Y(new_n1659));
  NOR3xp33_ASAP7_75t_L      g01403(.A(new_n1543), .B(new_n1657), .C(new_n1540), .Y(new_n1660));
  NOR2xp33_ASAP7_75t_L      g01404(.A(new_n1659), .B(new_n1660), .Y(new_n1661));
  INVx1_ASAP7_75t_L         g01405(.A(new_n1661), .Y(new_n1662));
  AOI22xp33_ASAP7_75t_L     g01406(.A1(\b[19] ), .A2(new_n282), .B1(\b[21] ), .B2(new_n303), .Y(new_n1663));
  OAI221xp5_ASAP7_75t_L     g01407(.A1(new_n291), .A2(new_n1539), .B1(new_n268), .B2(new_n1662), .C(new_n1663), .Y(new_n1664));
  XNOR2x2_ASAP7_75t_L       g01408(.A(\a[2] ), .B(new_n1664), .Y(new_n1665));
  XOR2x2_ASAP7_75t_L        g01409(.A(new_n1665), .B(new_n1652), .Y(new_n1666));
  A2O1A1O1Ixp25_ASAP7_75t_L g01410(.A1(new_n1448), .A2(new_n1452), .B(new_n1455), .C(new_n1553), .D(new_n1551), .Y(new_n1667));
  XNOR2x2_ASAP7_75t_L       g01411(.A(new_n1667), .B(new_n1666), .Y(\f[21] ));
  MAJIxp5_ASAP7_75t_L       g01412(.A(new_n1667), .B(new_n1652), .C(new_n1665), .Y(new_n1669));
  NOR3xp33_ASAP7_75t_L      g01413(.A(new_n1631), .B(new_n1632), .C(new_n1559), .Y(new_n1670));
  AOI22xp33_ASAP7_75t_L     g01414(.A1(new_n444), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n471), .Y(new_n1671));
  OAI221xp5_ASAP7_75t_L     g01415(.A1(new_n468), .A2(new_n942), .B1(new_n469), .B2(new_n1035), .C(new_n1671), .Y(new_n1672));
  XNOR2x2_ASAP7_75t_L       g01416(.A(\a[8] ), .B(new_n1672), .Y(new_n1673));
  AOI211xp5_ASAP7_75t_L     g01417(.A1(new_n1600), .A2(new_n1594), .B(new_n1589), .C(new_n1590), .Y(new_n1674));
  AOI221xp5_ASAP7_75t_L     g01418(.A1(new_n1605), .A2(new_n1604), .B1(new_n1491), .B2(new_n1493), .C(new_n1489), .Y(new_n1675));
  NAND2xp33_ASAP7_75t_L     g01419(.A(\b[6] ), .B(new_n1080), .Y(new_n1676));
  AOI22xp33_ASAP7_75t_L     g01420(.A1(new_n1076), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1253), .Y(new_n1677));
  OAI211xp5_ASAP7_75t_L     g01421(.A1(new_n1156), .A2(new_n425), .B(new_n1676), .C(new_n1677), .Y(new_n1678));
  NOR2xp33_ASAP7_75t_L      g01422(.A(new_n1071), .B(new_n1678), .Y(new_n1679));
  INVx1_ASAP7_75t_L         g01423(.A(new_n1679), .Y(new_n1680));
  NAND2xp33_ASAP7_75t_L     g01424(.A(new_n1071), .B(new_n1678), .Y(new_n1681));
  NOR4xp25_ASAP7_75t_L      g01425(.A(new_n1569), .B(new_n1574), .C(new_n1484), .D(new_n1481), .Y(new_n1682));
  INVx1_ASAP7_75t_L         g01426(.A(new_n1682), .Y(new_n1683));
  NAND2xp33_ASAP7_75t_L     g01427(.A(\b[3] ), .B(new_n1362), .Y(new_n1684));
  NAND2xp33_ASAP7_75t_L     g01428(.A(new_n1365), .B(new_n329), .Y(new_n1685));
  AOI22xp33_ASAP7_75t_L     g01429(.A1(new_n1360), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n1581), .Y(new_n1686));
  AND4x1_ASAP7_75t_L        g01430(.A(new_n1686), .B(new_n1685), .C(new_n1684), .D(\a[20] ), .Y(new_n1687));
  AOI31xp33_ASAP7_75t_L     g01431(.A1(new_n1685), .A2(new_n1684), .A3(new_n1686), .B(\a[20] ), .Y(new_n1688));
  INVx1_ASAP7_75t_L         g01432(.A(\a[23] ), .Y(new_n1689));
  NOR2xp33_ASAP7_75t_L      g01433(.A(new_n1689), .B(new_n1574), .Y(new_n1690));
  AND2x2_ASAP7_75t_L        g01434(.A(new_n1571), .B(new_n1572), .Y(new_n1691));
  INVx1_ASAP7_75t_L         g01435(.A(\a[22] ), .Y(new_n1692));
  NAND2xp33_ASAP7_75t_L     g01436(.A(\a[23] ), .B(new_n1692), .Y(new_n1693));
  NAND2xp33_ASAP7_75t_L     g01437(.A(\a[22] ), .B(new_n1689), .Y(new_n1694));
  AOI21xp33_ASAP7_75t_L     g01438(.A1(new_n1694), .A2(new_n1693), .B(new_n1691), .Y(new_n1695));
  NAND3xp33_ASAP7_75t_L     g01439(.A(new_n1573), .B(new_n1693), .C(new_n1694), .Y(new_n1696));
  NOR2xp33_ASAP7_75t_L      g01440(.A(\a[21] ), .B(new_n1692), .Y(new_n1697));
  NOR2xp33_ASAP7_75t_L      g01441(.A(\a[22] ), .B(new_n1570), .Y(new_n1698));
  OAI21xp33_ASAP7_75t_L     g01442(.A1(new_n1697), .A2(new_n1698), .B(new_n1691), .Y(new_n1699));
  OAI22xp33_ASAP7_75t_L     g01443(.A1(new_n1699), .A2(new_n258), .B1(new_n261), .B2(new_n1696), .Y(new_n1700));
  A2O1A1Ixp33_ASAP7_75t_L   g01444(.A1(new_n269), .A2(new_n1695), .B(new_n1700), .C(new_n1690), .Y(new_n1701));
  NAND2xp33_ASAP7_75t_L     g01445(.A(new_n269), .B(new_n1695), .Y(new_n1702));
  NAND2xp33_ASAP7_75t_L     g01446(.A(new_n1694), .B(new_n1693), .Y(new_n1703));
  NOR2xp33_ASAP7_75t_L      g01447(.A(new_n1703), .B(new_n1691), .Y(new_n1704));
  NOR2xp33_ASAP7_75t_L      g01448(.A(new_n1697), .B(new_n1698), .Y(new_n1705));
  NOR2xp33_ASAP7_75t_L      g01449(.A(new_n1573), .B(new_n1705), .Y(new_n1706));
  AOI22xp33_ASAP7_75t_L     g01450(.A1(\b[0] ), .A2(new_n1706), .B1(\b[1] ), .B2(new_n1704), .Y(new_n1707));
  OAI211xp5_ASAP7_75t_L     g01451(.A1(new_n1689), .A2(new_n1574), .B(new_n1707), .C(new_n1702), .Y(new_n1708));
  NAND2xp33_ASAP7_75t_L     g01452(.A(new_n1701), .B(new_n1708), .Y(new_n1709));
  OR3x1_ASAP7_75t_L         g01453(.A(new_n1687), .B(new_n1688), .C(new_n1709), .Y(new_n1710));
  OAI21xp33_ASAP7_75t_L     g01454(.A1(new_n1688), .A2(new_n1687), .B(new_n1709), .Y(new_n1711));
  AOI22xp33_ASAP7_75t_L     g01455(.A1(new_n1710), .A2(new_n1711), .B1(new_n1683), .B2(new_n1598), .Y(new_n1712));
  NOR3xp33_ASAP7_75t_L      g01456(.A(new_n1687), .B(new_n1688), .C(new_n1709), .Y(new_n1713));
  OA21x2_ASAP7_75t_L        g01457(.A1(new_n1688), .A2(new_n1687), .B(new_n1709), .Y(new_n1714));
  NOR4xp25_ASAP7_75t_L      g01458(.A(new_n1589), .B(new_n1714), .C(new_n1713), .D(new_n1682), .Y(new_n1715));
  AOI211xp5_ASAP7_75t_L     g01459(.A1(new_n1680), .A2(new_n1681), .B(new_n1712), .C(new_n1715), .Y(new_n1716));
  INVx1_ASAP7_75t_L         g01460(.A(new_n1681), .Y(new_n1717));
  OAI22xp33_ASAP7_75t_L     g01461(.A1(new_n1682), .A2(new_n1589), .B1(new_n1713), .B2(new_n1714), .Y(new_n1718));
  NAND4xp25_ASAP7_75t_L     g01462(.A(new_n1598), .B(new_n1710), .C(new_n1711), .D(new_n1683), .Y(new_n1719));
  AOI211xp5_ASAP7_75t_L     g01463(.A1(new_n1719), .A2(new_n1718), .B(new_n1679), .C(new_n1717), .Y(new_n1720));
  NOR2xp33_ASAP7_75t_L      g01464(.A(new_n1720), .B(new_n1716), .Y(new_n1721));
  OAI21xp33_ASAP7_75t_L     g01465(.A1(new_n1674), .A2(new_n1675), .B(new_n1721), .Y(new_n1722));
  INVx1_ASAP7_75t_L         g01466(.A(new_n1674), .Y(new_n1723));
  OAI221xp5_ASAP7_75t_L     g01467(.A1(new_n1597), .A2(new_n1601), .B1(new_n1494), .B2(new_n1472), .C(new_n1490), .Y(new_n1724));
  OAI211xp5_ASAP7_75t_L     g01468(.A1(new_n1716), .A2(new_n1720), .B(new_n1724), .C(new_n1723), .Y(new_n1725));
  AOI22xp33_ASAP7_75t_L     g01469(.A1(new_n811), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n900), .Y(new_n1726));
  OAI221xp5_ASAP7_75t_L     g01470(.A1(new_n904), .A2(new_n540), .B1(new_n898), .B2(new_n624), .C(new_n1726), .Y(new_n1727));
  XNOR2x2_ASAP7_75t_L       g01471(.A(\a[14] ), .B(new_n1727), .Y(new_n1728));
  NAND3xp33_ASAP7_75t_L     g01472(.A(new_n1722), .B(new_n1725), .C(new_n1728), .Y(new_n1729));
  AO21x2_ASAP7_75t_L        g01473(.A1(new_n1725), .A2(new_n1722), .B(new_n1728), .Y(new_n1730));
  A2O1A1O1Ixp25_ASAP7_75t_L g01474(.A1(new_n1496), .A2(new_n1466), .B(new_n1505), .C(new_n1613), .D(new_n1612), .Y(new_n1731));
  AND3x1_ASAP7_75t_L        g01475(.A(new_n1731), .B(new_n1730), .C(new_n1729), .Y(new_n1732));
  AOI21xp33_ASAP7_75t_L     g01476(.A1(new_n1730), .A2(new_n1729), .B(new_n1731), .Y(new_n1733));
  AOI22xp33_ASAP7_75t_L     g01477(.A1(\b[11] ), .A2(new_n651), .B1(\b[13] ), .B2(new_n581), .Y(new_n1734));
  OAI221xp5_ASAP7_75t_L     g01478(.A1(new_n821), .A2(new_n760), .B1(new_n577), .B2(new_n790), .C(new_n1734), .Y(new_n1735));
  XNOR2x2_ASAP7_75t_L       g01479(.A(\a[11] ), .B(new_n1735), .Y(new_n1736));
  OAI21xp33_ASAP7_75t_L     g01480(.A1(new_n1733), .A2(new_n1732), .B(new_n1736), .Y(new_n1737));
  NAND3xp33_ASAP7_75t_L     g01481(.A(new_n1731), .B(new_n1730), .C(new_n1729), .Y(new_n1738));
  AO21x2_ASAP7_75t_L        g01482(.A1(new_n1729), .A2(new_n1730), .B(new_n1731), .Y(new_n1739));
  INVx1_ASAP7_75t_L         g01483(.A(new_n1736), .Y(new_n1740));
  NAND3xp33_ASAP7_75t_L     g01484(.A(new_n1740), .B(new_n1739), .C(new_n1738), .Y(new_n1741));
  NAND2xp33_ASAP7_75t_L     g01485(.A(new_n1737), .B(new_n1741), .Y(new_n1742));
  O2A1O1Ixp33_ASAP7_75t_L   g01486(.A1(new_n1627), .A2(new_n1628), .B(new_n1624), .C(new_n1742), .Y(new_n1743));
  AOI21xp33_ASAP7_75t_L     g01487(.A1(new_n1739), .A2(new_n1738), .B(new_n1740), .Y(new_n1744));
  NOR3xp33_ASAP7_75t_L      g01488(.A(new_n1732), .B(new_n1733), .C(new_n1736), .Y(new_n1745));
  NOR2xp33_ASAP7_75t_L      g01489(.A(new_n1745), .B(new_n1744), .Y(new_n1746));
  AOI211xp5_ASAP7_75t_L     g01490(.A1(new_n1561), .A2(new_n1622), .B(new_n1623), .C(new_n1746), .Y(new_n1747));
  NOR3xp33_ASAP7_75t_L      g01491(.A(new_n1747), .B(new_n1743), .C(new_n1673), .Y(new_n1748));
  INVx1_ASAP7_75t_L         g01492(.A(new_n1673), .Y(new_n1749));
  A2O1A1Ixp33_ASAP7_75t_L   g01493(.A1(new_n1622), .A2(new_n1561), .B(new_n1623), .C(new_n1746), .Y(new_n1750));
  A2O1A1O1Ixp25_ASAP7_75t_L g01494(.A1(new_n1508), .A2(new_n1462), .B(new_n1515), .C(new_n1622), .D(new_n1623), .Y(new_n1751));
  NAND2xp33_ASAP7_75t_L     g01495(.A(new_n1751), .B(new_n1742), .Y(new_n1752));
  AOI21xp33_ASAP7_75t_L     g01496(.A1(new_n1750), .A2(new_n1752), .B(new_n1749), .Y(new_n1753));
  NOR2xp33_ASAP7_75t_L      g01497(.A(new_n1753), .B(new_n1748), .Y(new_n1754));
  A2O1A1Ixp33_ASAP7_75t_L   g01498(.A1(new_n1633), .A2(new_n1636), .B(new_n1670), .C(new_n1754), .Y(new_n1755));
  A2O1A1O1Ixp25_ASAP7_75t_L g01499(.A1(new_n1525), .A2(new_n1526), .B(new_n1643), .C(new_n1633), .D(new_n1670), .Y(new_n1756));
  NAND3xp33_ASAP7_75t_L     g01500(.A(new_n1750), .B(new_n1749), .C(new_n1752), .Y(new_n1757));
  OAI21xp33_ASAP7_75t_L     g01501(.A1(new_n1743), .A2(new_n1747), .B(new_n1673), .Y(new_n1758));
  NAND2xp33_ASAP7_75t_L     g01502(.A(new_n1757), .B(new_n1758), .Y(new_n1759));
  NAND2xp33_ASAP7_75t_L     g01503(.A(new_n1756), .B(new_n1759), .Y(new_n1760));
  AOI22xp33_ASAP7_75t_L     g01504(.A1(new_n344), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n370), .Y(new_n1761));
  OAI221xp5_ASAP7_75t_L     g01505(.A1(new_n429), .A2(new_n1313), .B1(new_n366), .B2(new_n1438), .C(new_n1761), .Y(new_n1762));
  XNOR2x2_ASAP7_75t_L       g01506(.A(\a[5] ), .B(new_n1762), .Y(new_n1763));
  NAND3xp33_ASAP7_75t_L     g01507(.A(new_n1755), .B(new_n1760), .C(new_n1763), .Y(new_n1764));
  O2A1O1Ixp33_ASAP7_75t_L   g01508(.A1(new_n1644), .A2(new_n1634), .B(new_n1630), .C(new_n1759), .Y(new_n1765));
  NOR3xp33_ASAP7_75t_L      g01509(.A(new_n1635), .B(new_n1754), .C(new_n1670), .Y(new_n1766));
  INVx1_ASAP7_75t_L         g01510(.A(new_n1763), .Y(new_n1767));
  OAI21xp33_ASAP7_75t_L     g01511(.A1(new_n1765), .A2(new_n1766), .B(new_n1767), .Y(new_n1768));
  NAND2xp33_ASAP7_75t_L     g01512(.A(new_n1764), .B(new_n1768), .Y(new_n1769));
  NOR3xp33_ASAP7_75t_L      g01513(.A(new_n1635), .B(new_n1637), .C(new_n1646), .Y(new_n1770));
  O2A1O1Ixp33_ASAP7_75t_L   g01514(.A1(new_n1641), .A2(new_n1647), .B(new_n1651), .C(new_n1770), .Y(new_n1771));
  XOR2x2_ASAP7_75t_L        g01515(.A(new_n1769), .B(new_n1771), .Y(new_n1772));
  NOR2xp33_ASAP7_75t_L      g01516(.A(\b[21] ), .B(\b[22] ), .Y(new_n1773));
  INVx1_ASAP7_75t_L         g01517(.A(\b[22] ), .Y(new_n1774));
  NOR2xp33_ASAP7_75t_L      g01518(.A(new_n1655), .B(new_n1774), .Y(new_n1775));
  NOR2xp33_ASAP7_75t_L      g01519(.A(new_n1773), .B(new_n1775), .Y(new_n1776));
  A2O1A1Ixp33_ASAP7_75t_L   g01520(.A1(\b[21] ), .A2(\b[20] ), .B(new_n1659), .C(new_n1776), .Y(new_n1777));
  NOR3xp33_ASAP7_75t_L      g01521(.A(new_n1659), .B(new_n1776), .C(new_n1656), .Y(new_n1778));
  INVx1_ASAP7_75t_L         g01522(.A(new_n1778), .Y(new_n1779));
  NAND2xp33_ASAP7_75t_L     g01523(.A(new_n1777), .B(new_n1779), .Y(new_n1780));
  AOI22xp33_ASAP7_75t_L     g01524(.A1(\b[20] ), .A2(new_n282), .B1(\b[22] ), .B2(new_n303), .Y(new_n1781));
  OAI221xp5_ASAP7_75t_L     g01525(.A1(new_n291), .A2(new_n1655), .B1(new_n268), .B2(new_n1780), .C(new_n1781), .Y(new_n1782));
  XNOR2x2_ASAP7_75t_L       g01526(.A(\a[2] ), .B(new_n1782), .Y(new_n1783));
  NAND2xp33_ASAP7_75t_L     g01527(.A(new_n1783), .B(new_n1772), .Y(new_n1784));
  NOR2xp33_ASAP7_75t_L      g01528(.A(new_n1783), .B(new_n1772), .Y(new_n1785));
  INVx1_ASAP7_75t_L         g01529(.A(new_n1785), .Y(new_n1786));
  NAND2xp33_ASAP7_75t_L     g01530(.A(new_n1784), .B(new_n1786), .Y(new_n1787));
  XNOR2x2_ASAP7_75t_L       g01531(.A(new_n1669), .B(new_n1787), .Y(\f[22] ));
  NOR3xp33_ASAP7_75t_L      g01532(.A(new_n1766), .B(new_n1765), .C(new_n1767), .Y(new_n1789));
  AOI21xp33_ASAP7_75t_L     g01533(.A1(new_n1755), .A2(new_n1760), .B(new_n1763), .Y(new_n1790));
  NOR2xp33_ASAP7_75t_L      g01534(.A(new_n1790), .B(new_n1789), .Y(new_n1791));
  NOR3xp33_ASAP7_75t_L      g01535(.A(new_n1766), .B(new_n1763), .C(new_n1765), .Y(new_n1792));
  INVx1_ASAP7_75t_L         g01536(.A(new_n1792), .Y(new_n1793));
  A2O1A1O1Ixp25_ASAP7_75t_L g01537(.A1(new_n1633), .A2(new_n1636), .B(new_n1670), .C(new_n1758), .D(new_n1748), .Y(new_n1794));
  NOR2xp33_ASAP7_75t_L      g01538(.A(new_n1030), .B(new_n468), .Y(new_n1795));
  INVx1_ASAP7_75t_L         g01539(.A(new_n1208), .Y(new_n1796));
  AOI22xp33_ASAP7_75t_L     g01540(.A1(new_n444), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n471), .Y(new_n1797));
  OAI31xp33_ASAP7_75t_L     g01541(.A1(new_n1796), .A2(new_n469), .A3(new_n1205), .B(new_n1797), .Y(new_n1798));
  OR3x1_ASAP7_75t_L         g01542(.A(new_n1798), .B(new_n435), .C(new_n1795), .Y(new_n1799));
  A2O1A1Ixp33_ASAP7_75t_L   g01543(.A1(\b[16] ), .A2(new_n447), .B(new_n1798), .C(new_n435), .Y(new_n1800));
  NAND2xp33_ASAP7_75t_L     g01544(.A(new_n1800), .B(new_n1799), .Y(new_n1801));
  NAND2xp33_ASAP7_75t_L     g01545(.A(new_n1725), .B(new_n1722), .Y(new_n1802));
  MAJIxp5_ASAP7_75t_L       g01546(.A(new_n1731), .B(new_n1728), .C(new_n1802), .Y(new_n1803));
  AOI22xp33_ASAP7_75t_L     g01547(.A1(new_n811), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n900), .Y(new_n1804));
  OAI221xp5_ASAP7_75t_L     g01548(.A1(new_n904), .A2(new_n617), .B1(new_n898), .B2(new_n685), .C(new_n1804), .Y(new_n1805));
  XNOR2x2_ASAP7_75t_L       g01549(.A(\a[14] ), .B(new_n1805), .Y(new_n1806));
  INVx1_ASAP7_75t_L         g01550(.A(new_n1720), .Y(new_n1807));
  O2A1O1Ixp33_ASAP7_75t_L   g01551(.A1(new_n1674), .A2(new_n1675), .B(new_n1807), .C(new_n1716), .Y(new_n1808));
  AOI22xp33_ASAP7_75t_L     g01552(.A1(new_n1076), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1253), .Y(new_n1809));
  OAI221xp5_ASAP7_75t_L     g01553(.A1(new_n1154), .A2(new_n420), .B1(new_n1156), .B2(new_n494), .C(new_n1809), .Y(new_n1810));
  XNOR2x2_ASAP7_75t_L       g01554(.A(\a[17] ), .B(new_n1810), .Y(new_n1811));
  NOR3xp33_ASAP7_75t_L      g01555(.A(new_n1569), .B(new_n1481), .C(new_n1484), .Y(new_n1812));
  NAND2xp33_ASAP7_75t_L     g01556(.A(new_n1588), .B(new_n1587), .Y(new_n1813));
  MAJIxp5_ASAP7_75t_L       g01557(.A(new_n1813), .B(new_n1575), .C(new_n1812), .Y(new_n1814));
  NOR2xp33_ASAP7_75t_L      g01558(.A(new_n1688), .B(new_n1687), .Y(new_n1815));
  MAJIxp5_ASAP7_75t_L       g01559(.A(new_n1814), .B(new_n1815), .C(new_n1709), .Y(new_n1816));
  NAND2xp33_ASAP7_75t_L     g01560(.A(\b[4] ), .B(new_n1362), .Y(new_n1817));
  NOR3xp33_ASAP7_75t_L      g01561(.A(new_n357), .B(new_n358), .C(new_n1359), .Y(new_n1818));
  OAI22xp33_ASAP7_75t_L     g01562(.A1(new_n1483), .A2(new_n298), .B1(new_n354), .B2(new_n1372), .Y(new_n1819));
  NOR2xp33_ASAP7_75t_L      g01563(.A(new_n1819), .B(new_n1818), .Y(new_n1820));
  NAND3xp33_ASAP7_75t_L     g01564(.A(new_n1820), .B(new_n1817), .C(\a[20] ), .Y(new_n1821));
  INVx1_ASAP7_75t_L         g01565(.A(new_n1817), .Y(new_n1822));
  OAI31xp33_ASAP7_75t_L     g01566(.A1(new_n1818), .A2(new_n1822), .A3(new_n1819), .B(new_n1356), .Y(new_n1823));
  NAND4xp25_ASAP7_75t_L     g01567(.A(new_n1707), .B(\a[23] ), .C(new_n1574), .D(new_n1702), .Y(new_n1824));
  NAND2xp33_ASAP7_75t_L     g01568(.A(\a[23] ), .B(new_n1824), .Y(new_n1825));
  NOR2xp33_ASAP7_75t_L      g01569(.A(new_n261), .B(new_n1699), .Y(new_n1826));
  NAND2xp33_ASAP7_75t_L     g01570(.A(new_n1703), .B(new_n1573), .Y(new_n1827));
  NAND2xp33_ASAP7_75t_L     g01571(.A(\b[2] ), .B(new_n1704), .Y(new_n1828));
  NAND3xp33_ASAP7_75t_L     g01572(.A(new_n1691), .B(new_n1703), .C(new_n1705), .Y(new_n1829));
  OAI221xp5_ASAP7_75t_L     g01573(.A1(new_n258), .A2(new_n1829), .B1(new_n280), .B2(new_n1827), .C(new_n1828), .Y(new_n1830));
  NOR2xp33_ASAP7_75t_L      g01574(.A(new_n1826), .B(new_n1830), .Y(new_n1831));
  XNOR2x2_ASAP7_75t_L       g01575(.A(new_n1831), .B(new_n1825), .Y(new_n1832));
  NAND3xp33_ASAP7_75t_L     g01576(.A(new_n1832), .B(new_n1823), .C(new_n1821), .Y(new_n1833));
  NAND2xp33_ASAP7_75t_L     g01577(.A(new_n1823), .B(new_n1821), .Y(new_n1834));
  INVx1_ASAP7_75t_L         g01578(.A(new_n1826), .Y(new_n1835));
  NOR2xp33_ASAP7_75t_L      g01579(.A(new_n280), .B(new_n1827), .Y(new_n1836));
  AND3x1_ASAP7_75t_L        g01580(.A(new_n1691), .B(new_n1705), .C(new_n1703), .Y(new_n1837));
  AOI221xp5_ASAP7_75t_L     g01581(.A1(new_n1704), .A2(\b[2] ), .B1(new_n1837), .B2(\b[0] ), .C(new_n1836), .Y(new_n1838));
  NAND2xp33_ASAP7_75t_L     g01582(.A(new_n1835), .B(new_n1838), .Y(new_n1839));
  XNOR2x2_ASAP7_75t_L       g01583(.A(new_n1839), .B(new_n1825), .Y(new_n1840));
  NAND2xp33_ASAP7_75t_L     g01584(.A(new_n1834), .B(new_n1840), .Y(new_n1841));
  AOI21xp33_ASAP7_75t_L     g01585(.A1(new_n1841), .A2(new_n1833), .B(new_n1816), .Y(new_n1842));
  OR2x4_ASAP7_75t_L         g01586(.A(new_n1688), .B(new_n1687), .Y(new_n1843));
  INVx1_ASAP7_75t_L         g01587(.A(new_n1709), .Y(new_n1844));
  NAND2xp33_ASAP7_75t_L     g01588(.A(new_n1844), .B(new_n1843), .Y(new_n1845));
  NOR2xp33_ASAP7_75t_L      g01589(.A(new_n1834), .B(new_n1840), .Y(new_n1846));
  AOI21xp33_ASAP7_75t_L     g01590(.A1(new_n1823), .A2(new_n1821), .B(new_n1832), .Y(new_n1847));
  AOI211xp5_ASAP7_75t_L     g01591(.A1(new_n1718), .A2(new_n1845), .B(new_n1846), .C(new_n1847), .Y(new_n1848));
  OAI21xp33_ASAP7_75t_L     g01592(.A1(new_n1848), .A2(new_n1842), .B(new_n1811), .Y(new_n1849));
  INVx1_ASAP7_75t_L         g01593(.A(new_n1849), .Y(new_n1850));
  NOR3xp33_ASAP7_75t_L      g01594(.A(new_n1842), .B(new_n1848), .C(new_n1811), .Y(new_n1851));
  NOR3xp33_ASAP7_75t_L      g01595(.A(new_n1808), .B(new_n1850), .C(new_n1851), .Y(new_n1852));
  OAI211xp5_ASAP7_75t_L     g01596(.A1(new_n1679), .A2(new_n1717), .B(new_n1718), .C(new_n1719), .Y(new_n1853));
  A2O1A1Ixp33_ASAP7_75t_L   g01597(.A1(new_n1724), .A2(new_n1723), .B(new_n1720), .C(new_n1853), .Y(new_n1854));
  INVx1_ASAP7_75t_L         g01598(.A(new_n1851), .Y(new_n1855));
  AOI21xp33_ASAP7_75t_L     g01599(.A1(new_n1855), .A2(new_n1849), .B(new_n1854), .Y(new_n1856));
  OAI21xp33_ASAP7_75t_L     g01600(.A1(new_n1856), .A2(new_n1852), .B(new_n1806), .Y(new_n1857));
  OR3x1_ASAP7_75t_L         g01601(.A(new_n1852), .B(new_n1806), .C(new_n1856), .Y(new_n1858));
  NAND3xp33_ASAP7_75t_L     g01602(.A(new_n1858), .B(new_n1803), .C(new_n1857), .Y(new_n1859));
  AO21x2_ASAP7_75t_L        g01603(.A1(new_n1857), .A2(new_n1858), .B(new_n1803), .Y(new_n1860));
  AOI22xp33_ASAP7_75t_L     g01604(.A1(\b[12] ), .A2(new_n651), .B1(\b[14] ), .B2(new_n581), .Y(new_n1861));
  OAI221xp5_ASAP7_75t_L     g01605(.A1(new_n821), .A2(new_n784), .B1(new_n577), .B2(new_n875), .C(new_n1861), .Y(new_n1862));
  XNOR2x2_ASAP7_75t_L       g01606(.A(\a[11] ), .B(new_n1862), .Y(new_n1863));
  NAND3xp33_ASAP7_75t_L     g01607(.A(new_n1860), .B(new_n1859), .C(new_n1863), .Y(new_n1864));
  AOI21xp33_ASAP7_75t_L     g01608(.A1(new_n1860), .A2(new_n1859), .B(new_n1863), .Y(new_n1865));
  INVx1_ASAP7_75t_L         g01609(.A(new_n1865), .Y(new_n1866));
  A2O1A1O1Ixp25_ASAP7_75t_L g01610(.A1(new_n1622), .A2(new_n1561), .B(new_n1623), .C(new_n1737), .D(new_n1745), .Y(new_n1867));
  AOI21xp33_ASAP7_75t_L     g01611(.A1(new_n1866), .A2(new_n1864), .B(new_n1867), .Y(new_n1868));
  AND3x1_ASAP7_75t_L        g01612(.A(new_n1858), .B(new_n1803), .C(new_n1857), .Y(new_n1869));
  AOI21xp33_ASAP7_75t_L     g01613(.A1(new_n1858), .A2(new_n1857), .B(new_n1803), .Y(new_n1870));
  INVx1_ASAP7_75t_L         g01614(.A(new_n1863), .Y(new_n1871));
  NOR3xp33_ASAP7_75t_L      g01615(.A(new_n1871), .B(new_n1870), .C(new_n1869), .Y(new_n1872));
  OAI21xp33_ASAP7_75t_L     g01616(.A1(new_n1744), .A2(new_n1751), .B(new_n1741), .Y(new_n1873));
  NOR3xp33_ASAP7_75t_L      g01617(.A(new_n1873), .B(new_n1865), .C(new_n1872), .Y(new_n1874));
  OAI21xp33_ASAP7_75t_L     g01618(.A1(new_n1874), .A2(new_n1868), .B(new_n1801), .Y(new_n1875));
  AND2x2_ASAP7_75t_L        g01619(.A(new_n1800), .B(new_n1799), .Y(new_n1876));
  OAI21xp33_ASAP7_75t_L     g01620(.A1(new_n1872), .A2(new_n1865), .B(new_n1873), .Y(new_n1877));
  NAND3xp33_ASAP7_75t_L     g01621(.A(new_n1866), .B(new_n1867), .C(new_n1864), .Y(new_n1878));
  NAND3xp33_ASAP7_75t_L     g01622(.A(new_n1878), .B(new_n1877), .C(new_n1876), .Y(new_n1879));
  NAND2xp33_ASAP7_75t_L     g01623(.A(new_n1879), .B(new_n1875), .Y(new_n1880));
  NOR2xp33_ASAP7_75t_L      g01624(.A(new_n1794), .B(new_n1880), .Y(new_n1881));
  OAI21xp33_ASAP7_75t_L     g01625(.A1(new_n1753), .A2(new_n1756), .B(new_n1757), .Y(new_n1882));
  AOI21xp33_ASAP7_75t_L     g01626(.A1(new_n1879), .A2(new_n1875), .B(new_n1882), .Y(new_n1883));
  NAND2xp33_ASAP7_75t_L     g01627(.A(\b[19] ), .B(new_n347), .Y(new_n1884));
  INVx1_ASAP7_75t_L         g01628(.A(new_n1546), .Y(new_n1885));
  NOR2xp33_ASAP7_75t_L      g01629(.A(new_n1543), .B(new_n1885), .Y(new_n1886));
  NAND2xp33_ASAP7_75t_L     g01630(.A(new_n341), .B(new_n1886), .Y(new_n1887));
  AOI22xp33_ASAP7_75t_L     g01631(.A1(new_n344), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n370), .Y(new_n1888));
  NAND4xp25_ASAP7_75t_L     g01632(.A(new_n1887), .B(\a[5] ), .C(new_n1884), .D(new_n1888), .Y(new_n1889));
  OAI21xp33_ASAP7_75t_L     g01633(.A1(new_n366), .A2(new_n1547), .B(new_n1888), .Y(new_n1890));
  A2O1A1Ixp33_ASAP7_75t_L   g01634(.A1(\b[19] ), .A2(new_n347), .B(new_n1890), .C(new_n338), .Y(new_n1891));
  NAND2xp33_ASAP7_75t_L     g01635(.A(new_n1889), .B(new_n1891), .Y(new_n1892));
  OAI21xp33_ASAP7_75t_L     g01636(.A1(new_n1881), .A2(new_n1883), .B(new_n1892), .Y(new_n1893));
  NAND3xp33_ASAP7_75t_L     g01637(.A(new_n1882), .B(new_n1875), .C(new_n1879), .Y(new_n1894));
  NAND2xp33_ASAP7_75t_L     g01638(.A(new_n1794), .B(new_n1880), .Y(new_n1895));
  AND2x2_ASAP7_75t_L        g01639(.A(new_n1889), .B(new_n1891), .Y(new_n1896));
  NAND3xp33_ASAP7_75t_L     g01640(.A(new_n1894), .B(new_n1896), .C(new_n1895), .Y(new_n1897));
  NAND2xp33_ASAP7_75t_L     g01641(.A(new_n1897), .B(new_n1893), .Y(new_n1898));
  OAI211xp5_ASAP7_75t_L     g01642(.A1(new_n1791), .A2(new_n1771), .B(new_n1898), .C(new_n1793), .Y(new_n1899));
  A2O1A1Ixp33_ASAP7_75t_L   g01643(.A1(new_n1428), .A2(new_n1429), .B(new_n1457), .C(new_n1533), .Y(new_n1900));
  INVx1_ASAP7_75t_L         g01644(.A(new_n1770), .Y(new_n1901));
  A2O1A1Ixp33_ASAP7_75t_L   g01645(.A1(new_n1650), .A2(new_n1900), .B(new_n1648), .C(new_n1901), .Y(new_n1902));
  AOI21xp33_ASAP7_75t_L     g01646(.A1(new_n1894), .A2(new_n1895), .B(new_n1896), .Y(new_n1903));
  NOR3xp33_ASAP7_75t_L      g01647(.A(new_n1883), .B(new_n1881), .C(new_n1892), .Y(new_n1904));
  NOR2xp33_ASAP7_75t_L      g01648(.A(new_n1904), .B(new_n1903), .Y(new_n1905));
  A2O1A1Ixp33_ASAP7_75t_L   g01649(.A1(new_n1902), .A2(new_n1769), .B(new_n1792), .C(new_n1905), .Y(new_n1906));
  INVx1_ASAP7_75t_L         g01650(.A(new_n1777), .Y(new_n1907));
  NOR2xp33_ASAP7_75t_L      g01651(.A(\b[22] ), .B(\b[23] ), .Y(new_n1908));
  INVx1_ASAP7_75t_L         g01652(.A(\b[23] ), .Y(new_n1909));
  NOR2xp33_ASAP7_75t_L      g01653(.A(new_n1774), .B(new_n1909), .Y(new_n1910));
  NOR2xp33_ASAP7_75t_L      g01654(.A(new_n1908), .B(new_n1910), .Y(new_n1911));
  A2O1A1Ixp33_ASAP7_75t_L   g01655(.A1(\b[22] ), .A2(\b[21] ), .B(new_n1907), .C(new_n1911), .Y(new_n1912));
  O2A1O1Ixp33_ASAP7_75t_L   g01656(.A1(new_n1656), .A2(new_n1659), .B(new_n1776), .C(new_n1775), .Y(new_n1913));
  OAI21xp33_ASAP7_75t_L     g01657(.A1(new_n1908), .A2(new_n1910), .B(new_n1913), .Y(new_n1914));
  NAND2xp33_ASAP7_75t_L     g01658(.A(new_n1914), .B(new_n1912), .Y(new_n1915));
  AOI22xp33_ASAP7_75t_L     g01659(.A1(\b[21] ), .A2(new_n282), .B1(\b[23] ), .B2(new_n303), .Y(new_n1916));
  OAI221xp5_ASAP7_75t_L     g01660(.A1(new_n291), .A2(new_n1774), .B1(new_n268), .B2(new_n1915), .C(new_n1916), .Y(new_n1917));
  XNOR2x2_ASAP7_75t_L       g01661(.A(\a[2] ), .B(new_n1917), .Y(new_n1918));
  NAND3xp33_ASAP7_75t_L     g01662(.A(new_n1906), .B(new_n1899), .C(new_n1918), .Y(new_n1919));
  AOI221xp5_ASAP7_75t_L     g01663(.A1(new_n1897), .A2(new_n1893), .B1(new_n1769), .B2(new_n1902), .C(new_n1792), .Y(new_n1920));
  O2A1O1Ixp33_ASAP7_75t_L   g01664(.A1(new_n1791), .A2(new_n1771), .B(new_n1793), .C(new_n1898), .Y(new_n1921));
  INVx1_ASAP7_75t_L         g01665(.A(new_n1918), .Y(new_n1922));
  OAI21xp33_ASAP7_75t_L     g01666(.A1(new_n1920), .A2(new_n1921), .B(new_n1922), .Y(new_n1923));
  NAND2xp33_ASAP7_75t_L     g01667(.A(new_n1923), .B(new_n1919), .Y(new_n1924));
  AOI21xp33_ASAP7_75t_L     g01668(.A1(new_n1669), .A2(new_n1784), .B(new_n1785), .Y(new_n1925));
  XNOR2x2_ASAP7_75t_L       g01669(.A(new_n1924), .B(new_n1925), .Y(\f[23] ));
  INVx1_ASAP7_75t_L         g01670(.A(new_n1910), .Y(new_n1927));
  NOR2xp33_ASAP7_75t_L      g01671(.A(\b[23] ), .B(\b[24] ), .Y(new_n1928));
  INVx1_ASAP7_75t_L         g01672(.A(\b[24] ), .Y(new_n1929));
  NOR2xp33_ASAP7_75t_L      g01673(.A(new_n1909), .B(new_n1929), .Y(new_n1930));
  NOR2xp33_ASAP7_75t_L      g01674(.A(new_n1928), .B(new_n1930), .Y(new_n1931));
  INVx1_ASAP7_75t_L         g01675(.A(new_n1931), .Y(new_n1932));
  O2A1O1Ixp33_ASAP7_75t_L   g01676(.A1(new_n1908), .A2(new_n1913), .B(new_n1927), .C(new_n1932), .Y(new_n1933));
  AND3x1_ASAP7_75t_L        g01677(.A(new_n1912), .B(new_n1932), .C(new_n1927), .Y(new_n1934));
  NOR2xp33_ASAP7_75t_L      g01678(.A(new_n1933), .B(new_n1934), .Y(new_n1935));
  OAI22xp33_ASAP7_75t_L     g01679(.A1(new_n271), .A2(new_n1929), .B1(new_n1774), .B2(new_n283), .Y(new_n1936));
  AOI221xp5_ASAP7_75t_L     g01680(.A1(\b[23] ), .A2(new_n272), .B1(new_n267), .B2(new_n1935), .C(new_n1936), .Y(new_n1937));
  XNOR2x2_ASAP7_75t_L       g01681(.A(\a[2] ), .B(new_n1937), .Y(new_n1938));
  A2O1A1O1Ixp25_ASAP7_75t_L g01682(.A1(new_n1769), .A2(new_n1902), .B(new_n1792), .C(new_n1897), .D(new_n1903), .Y(new_n1939));
  AOI22xp33_ASAP7_75t_L     g01683(.A1(new_n344), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n370), .Y(new_n1940));
  OAI221xp5_ASAP7_75t_L     g01684(.A1(new_n429), .A2(new_n1539), .B1(new_n366), .B2(new_n1662), .C(new_n1940), .Y(new_n1941));
  XNOR2x2_ASAP7_75t_L       g01685(.A(\a[5] ), .B(new_n1941), .Y(new_n1942));
  NOR3xp33_ASAP7_75t_L      g01686(.A(new_n1868), .B(new_n1874), .C(new_n1876), .Y(new_n1943));
  INVx1_ASAP7_75t_L         g01687(.A(new_n1943), .Y(new_n1944));
  A2O1A1Ixp33_ASAP7_75t_L   g01688(.A1(new_n1875), .A2(new_n1879), .B(new_n1794), .C(new_n1944), .Y(new_n1945));
  NOR3xp33_ASAP7_75t_L      g01689(.A(new_n1852), .B(new_n1856), .C(new_n1806), .Y(new_n1946));
  AO21x2_ASAP7_75t_L        g01690(.A1(new_n1857), .A2(new_n1803), .B(new_n1946), .Y(new_n1947));
  NOR2xp33_ASAP7_75t_L      g01691(.A(new_n679), .B(new_n904), .Y(new_n1948));
  INVx1_ASAP7_75t_L         g01692(.A(new_n1948), .Y(new_n1949));
  NAND2xp33_ASAP7_75t_L     g01693(.A(new_n808), .B(new_n1232), .Y(new_n1950));
  AOI22xp33_ASAP7_75t_L     g01694(.A1(new_n811), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n900), .Y(new_n1951));
  AND4x1_ASAP7_75t_L        g01695(.A(new_n1951), .B(new_n1950), .C(new_n1949), .D(\a[14] ), .Y(new_n1952));
  AOI31xp33_ASAP7_75t_L     g01696(.A1(new_n1950), .A2(new_n1949), .A3(new_n1951), .B(\a[14] ), .Y(new_n1953));
  NOR2xp33_ASAP7_75t_L      g01697(.A(new_n1953), .B(new_n1952), .Y(new_n1954));
  OAI21xp33_ASAP7_75t_L     g01698(.A1(new_n1602), .A2(new_n1616), .B(new_n1723), .Y(new_n1955));
  A2O1A1O1Ixp25_ASAP7_75t_L g01699(.A1(new_n1721), .A2(new_n1955), .B(new_n1716), .C(new_n1849), .D(new_n1851), .Y(new_n1956));
  INVx1_ASAP7_75t_L         g01700(.A(\a[24] ), .Y(new_n1957));
  NAND2xp33_ASAP7_75t_L     g01701(.A(\a[23] ), .B(new_n1957), .Y(new_n1958));
  NAND2xp33_ASAP7_75t_L     g01702(.A(\a[24] ), .B(new_n1689), .Y(new_n1959));
  NAND2xp33_ASAP7_75t_L     g01703(.A(new_n1959), .B(new_n1958), .Y(new_n1960));
  NAND2xp33_ASAP7_75t_L     g01704(.A(\b[0] ), .B(new_n1960), .Y(new_n1961));
  INVx1_ASAP7_75t_L         g01705(.A(new_n1961), .Y(new_n1962));
  OAI31xp33_ASAP7_75t_L     g01706(.A1(new_n1824), .A2(new_n1830), .A3(new_n1826), .B(new_n1962), .Y(new_n1963));
  A2O1A1Ixp33_ASAP7_75t_L   g01707(.A1(new_n1571), .A2(new_n1572), .B(new_n258), .C(\a[23] ), .Y(new_n1964));
  AOI211xp5_ASAP7_75t_L     g01708(.A1(new_n1695), .A2(new_n269), .B(new_n1964), .C(new_n1700), .Y(new_n1965));
  NAND4xp25_ASAP7_75t_L     g01709(.A(new_n1965), .B(new_n1961), .C(new_n1838), .D(new_n1835), .Y(new_n1966));
  NOR2xp33_ASAP7_75t_L      g01710(.A(new_n276), .B(new_n1699), .Y(new_n1967));
  OAI22xp33_ASAP7_75t_L     g01711(.A1(new_n1829), .A2(new_n261), .B1(new_n298), .B2(new_n1696), .Y(new_n1968));
  AOI211xp5_ASAP7_75t_L     g01712(.A1(new_n406), .A2(new_n1695), .B(new_n1967), .C(new_n1968), .Y(new_n1969));
  NAND2xp33_ASAP7_75t_L     g01713(.A(\a[23] ), .B(new_n1969), .Y(new_n1970));
  NOR2xp33_ASAP7_75t_L      g01714(.A(new_n1827), .B(new_n302), .Y(new_n1971));
  OAI31xp33_ASAP7_75t_L     g01715(.A1(new_n1971), .A2(new_n1967), .A3(new_n1968), .B(new_n1689), .Y(new_n1972));
  AO22x1_ASAP7_75t_L        g01716(.A1(new_n1972), .A2(new_n1970), .B1(new_n1966), .B2(new_n1963), .Y(new_n1973));
  NAND4xp25_ASAP7_75t_L     g01717(.A(new_n1963), .B(new_n1966), .C(new_n1970), .D(new_n1972), .Y(new_n1974));
  NAND2xp33_ASAP7_75t_L     g01718(.A(\b[5] ), .B(new_n1362), .Y(new_n1975));
  NAND2xp33_ASAP7_75t_L     g01719(.A(new_n1365), .B(new_n526), .Y(new_n1976));
  AOI22xp33_ASAP7_75t_L     g01720(.A1(new_n1360), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1581), .Y(new_n1977));
  NAND4xp25_ASAP7_75t_L     g01721(.A(new_n1976), .B(\a[20] ), .C(new_n1975), .D(new_n1977), .Y(new_n1978));
  OAI21xp33_ASAP7_75t_L     g01722(.A1(new_n1359), .A2(new_n390), .B(new_n1977), .Y(new_n1979));
  A2O1A1Ixp33_ASAP7_75t_L   g01723(.A1(\b[5] ), .A2(new_n1362), .B(new_n1979), .C(new_n1356), .Y(new_n1980));
  AND4x1_ASAP7_75t_L        g01724(.A(new_n1980), .B(new_n1978), .C(new_n1974), .D(new_n1973), .Y(new_n1981));
  AOI22xp33_ASAP7_75t_L     g01725(.A1(new_n1973), .A2(new_n1974), .B1(new_n1978), .B2(new_n1980), .Y(new_n1982));
  NOR2xp33_ASAP7_75t_L      g01726(.A(new_n1982), .B(new_n1981), .Y(new_n1983));
  AOI31xp33_ASAP7_75t_L     g01727(.A1(new_n1718), .A2(new_n1841), .A3(new_n1845), .B(new_n1846), .Y(new_n1984));
  NAND2xp33_ASAP7_75t_L     g01728(.A(new_n1984), .B(new_n1983), .Y(new_n1985));
  NAND4xp25_ASAP7_75t_L     g01729(.A(new_n1980), .B(new_n1973), .C(new_n1974), .D(new_n1978), .Y(new_n1986));
  AO22x1_ASAP7_75t_L        g01730(.A1(new_n1973), .A2(new_n1974), .B1(new_n1978), .B2(new_n1980), .Y(new_n1987));
  NAND2xp33_ASAP7_75t_L     g01731(.A(new_n1986), .B(new_n1987), .Y(new_n1988));
  NOR2xp33_ASAP7_75t_L      g01732(.A(new_n1709), .B(new_n1815), .Y(new_n1989));
  OAI31xp33_ASAP7_75t_L     g01733(.A1(new_n1712), .A2(new_n1989), .A3(new_n1847), .B(new_n1833), .Y(new_n1990));
  NAND2xp33_ASAP7_75t_L     g01734(.A(new_n1988), .B(new_n1990), .Y(new_n1991));
  AOI22xp33_ASAP7_75t_L     g01735(.A1(new_n1076), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1253), .Y(new_n1992));
  OAI221xp5_ASAP7_75t_L     g01736(.A1(new_n1154), .A2(new_n488), .B1(new_n1156), .B2(new_n548), .C(new_n1992), .Y(new_n1993));
  OR2x4_ASAP7_75t_L         g01737(.A(new_n1071), .B(new_n1993), .Y(new_n1994));
  NAND2xp33_ASAP7_75t_L     g01738(.A(new_n1071), .B(new_n1993), .Y(new_n1995));
  AOI22xp33_ASAP7_75t_L     g01739(.A1(new_n1994), .A2(new_n1995), .B1(new_n1985), .B2(new_n1991), .Y(new_n1996));
  AND4x1_ASAP7_75t_L        g01740(.A(new_n1991), .B(new_n1985), .C(new_n1995), .D(new_n1994), .Y(new_n1997));
  NOR3xp33_ASAP7_75t_L      g01741(.A(new_n1956), .B(new_n1996), .C(new_n1997), .Y(new_n1998));
  AO22x1_ASAP7_75t_L        g01742(.A1(new_n1995), .A2(new_n1994), .B1(new_n1985), .B2(new_n1991), .Y(new_n1999));
  NAND4xp25_ASAP7_75t_L     g01743(.A(new_n1991), .B(new_n1985), .C(new_n1994), .D(new_n1995), .Y(new_n2000));
  AOI221xp5_ASAP7_75t_L     g01744(.A1(new_n1854), .A2(new_n1849), .B1(new_n2000), .B2(new_n1999), .C(new_n1851), .Y(new_n2001));
  OAI21xp33_ASAP7_75t_L     g01745(.A1(new_n2001), .A2(new_n1998), .B(new_n1954), .Y(new_n2002));
  OR2x4_ASAP7_75t_L         g01746(.A(new_n1953), .B(new_n1952), .Y(new_n2003));
  NOR2xp33_ASAP7_75t_L      g01747(.A(new_n1996), .B(new_n1997), .Y(new_n2004));
  A2O1A1Ixp33_ASAP7_75t_L   g01748(.A1(new_n1849), .A2(new_n1854), .B(new_n1851), .C(new_n2004), .Y(new_n2005));
  OAI21xp33_ASAP7_75t_L     g01749(.A1(new_n1996), .A2(new_n1997), .B(new_n1956), .Y(new_n2006));
  NAND3xp33_ASAP7_75t_L     g01750(.A(new_n2003), .B(new_n2005), .C(new_n2006), .Y(new_n2007));
  NAND3xp33_ASAP7_75t_L     g01751(.A(new_n1947), .B(new_n2002), .C(new_n2007), .Y(new_n2008));
  AOI21xp33_ASAP7_75t_L     g01752(.A1(new_n1803), .A2(new_n1857), .B(new_n1946), .Y(new_n2009));
  AOI21xp33_ASAP7_75t_L     g01753(.A1(new_n2005), .A2(new_n2006), .B(new_n2003), .Y(new_n2010));
  NOR3xp33_ASAP7_75t_L      g01754(.A(new_n1998), .B(new_n1954), .C(new_n2001), .Y(new_n2011));
  OAI21xp33_ASAP7_75t_L     g01755(.A1(new_n2011), .A2(new_n2010), .B(new_n2009), .Y(new_n2012));
  NAND2xp33_ASAP7_75t_L     g01756(.A(new_n2012), .B(new_n2008), .Y(new_n2013));
  AOI22xp33_ASAP7_75t_L     g01757(.A1(\b[13] ), .A2(new_n651), .B1(\b[15] ), .B2(new_n581), .Y(new_n2014));
  OAI221xp5_ASAP7_75t_L     g01758(.A1(new_n821), .A2(new_n869), .B1(new_n577), .B2(new_n950), .C(new_n2014), .Y(new_n2015));
  XNOR2x2_ASAP7_75t_L       g01759(.A(\a[11] ), .B(new_n2015), .Y(new_n2016));
  INVx1_ASAP7_75t_L         g01760(.A(new_n2016), .Y(new_n2017));
  NOR2xp33_ASAP7_75t_L      g01761(.A(new_n2017), .B(new_n2013), .Y(new_n2018));
  NOR3xp33_ASAP7_75t_L      g01762(.A(new_n2009), .B(new_n2010), .C(new_n2011), .Y(new_n2019));
  AOI21xp33_ASAP7_75t_L     g01763(.A1(new_n2007), .A2(new_n2002), .B(new_n1947), .Y(new_n2020));
  NOR2xp33_ASAP7_75t_L      g01764(.A(new_n2019), .B(new_n2020), .Y(new_n2021));
  NOR2xp33_ASAP7_75t_L      g01765(.A(new_n2016), .B(new_n2021), .Y(new_n2022));
  NAND2xp33_ASAP7_75t_L     g01766(.A(new_n1859), .B(new_n1860), .Y(new_n2023));
  MAJIxp5_ASAP7_75t_L       g01767(.A(new_n1867), .B(new_n2023), .C(new_n1863), .Y(new_n2024));
  NOR3xp33_ASAP7_75t_L      g01768(.A(new_n2024), .B(new_n2022), .C(new_n2018), .Y(new_n2025));
  NAND2xp33_ASAP7_75t_L     g01769(.A(new_n2016), .B(new_n2021), .Y(new_n2026));
  NAND2xp33_ASAP7_75t_L     g01770(.A(new_n2017), .B(new_n2013), .Y(new_n2027));
  NOR2xp33_ASAP7_75t_L      g01771(.A(new_n1870), .B(new_n1869), .Y(new_n2028));
  MAJIxp5_ASAP7_75t_L       g01772(.A(new_n1873), .B(new_n1871), .C(new_n2028), .Y(new_n2029));
  AOI21xp33_ASAP7_75t_L     g01773(.A1(new_n2026), .A2(new_n2027), .B(new_n2029), .Y(new_n2030));
  OAI22xp33_ASAP7_75t_L     g01774(.A1(new_n516), .A2(new_n1030), .B1(new_n1313), .B2(new_n515), .Y(new_n2031));
  AOI221xp5_ASAP7_75t_L     g01775(.A1(\b[17] ), .A2(new_n447), .B1(new_n441), .B2(new_n1319), .C(new_n2031), .Y(new_n2032));
  XNOR2x2_ASAP7_75t_L       g01776(.A(\a[8] ), .B(new_n2032), .Y(new_n2033));
  INVx1_ASAP7_75t_L         g01777(.A(new_n2033), .Y(new_n2034));
  OAI21xp33_ASAP7_75t_L     g01778(.A1(new_n2030), .A2(new_n2025), .B(new_n2034), .Y(new_n2035));
  NAND3xp33_ASAP7_75t_L     g01779(.A(new_n2026), .B(new_n2027), .C(new_n2029), .Y(new_n2036));
  OAI21xp33_ASAP7_75t_L     g01780(.A1(new_n2018), .A2(new_n2022), .B(new_n2024), .Y(new_n2037));
  NAND3xp33_ASAP7_75t_L     g01781(.A(new_n2037), .B(new_n2036), .C(new_n2033), .Y(new_n2038));
  NAND3xp33_ASAP7_75t_L     g01782(.A(new_n1945), .B(new_n2035), .C(new_n2038), .Y(new_n2039));
  INVx1_ASAP7_75t_L         g01783(.A(new_n1756), .Y(new_n2040));
  A2O1A1O1Ixp25_ASAP7_75t_L g01784(.A1(new_n1754), .A2(new_n2040), .B(new_n1748), .C(new_n1880), .D(new_n1943), .Y(new_n2041));
  NAND2xp33_ASAP7_75t_L     g01785(.A(new_n2038), .B(new_n2035), .Y(new_n2042));
  NAND2xp33_ASAP7_75t_L     g01786(.A(new_n2042), .B(new_n2041), .Y(new_n2043));
  AOI21xp33_ASAP7_75t_L     g01787(.A1(new_n2043), .A2(new_n2039), .B(new_n1942), .Y(new_n2044));
  XNOR2x2_ASAP7_75t_L       g01788(.A(new_n338), .B(new_n1941), .Y(new_n2045));
  NOR2xp33_ASAP7_75t_L      g01789(.A(new_n2042), .B(new_n2041), .Y(new_n2046));
  AOI21xp33_ASAP7_75t_L     g01790(.A1(new_n2038), .A2(new_n2035), .B(new_n1945), .Y(new_n2047));
  NOR3xp33_ASAP7_75t_L      g01791(.A(new_n2046), .B(new_n2047), .C(new_n2045), .Y(new_n2048));
  NOR2xp33_ASAP7_75t_L      g01792(.A(new_n2044), .B(new_n2048), .Y(new_n2049));
  NOR2xp33_ASAP7_75t_L      g01793(.A(new_n2049), .B(new_n1939), .Y(new_n2050));
  OAI21xp33_ASAP7_75t_L     g01794(.A1(new_n2047), .A2(new_n2046), .B(new_n2045), .Y(new_n2051));
  NAND3xp33_ASAP7_75t_L     g01795(.A(new_n2043), .B(new_n2039), .C(new_n1942), .Y(new_n2052));
  NAND2xp33_ASAP7_75t_L     g01796(.A(new_n2052), .B(new_n2051), .Y(new_n2053));
  NOR3xp33_ASAP7_75t_L      g01797(.A(new_n2053), .B(new_n1921), .C(new_n1903), .Y(new_n2054));
  NOR3xp33_ASAP7_75t_L      g01798(.A(new_n2054), .B(new_n2050), .C(new_n1938), .Y(new_n2055));
  XNOR2x2_ASAP7_75t_L       g01799(.A(new_n262), .B(new_n1937), .Y(new_n2056));
  NAND2xp33_ASAP7_75t_L     g01800(.A(new_n1895), .B(new_n1894), .Y(new_n2057));
  A2O1A1Ixp33_ASAP7_75t_L   g01801(.A1(new_n1892), .A2(new_n2057), .B(new_n1921), .C(new_n2053), .Y(new_n2058));
  NAND2xp33_ASAP7_75t_L     g01802(.A(new_n2049), .B(new_n1939), .Y(new_n2059));
  AOI21xp33_ASAP7_75t_L     g01803(.A1(new_n2058), .A2(new_n2059), .B(new_n2056), .Y(new_n2060));
  NOR2xp33_ASAP7_75t_L      g01804(.A(new_n2060), .B(new_n2055), .Y(new_n2061));
  NOR3xp33_ASAP7_75t_L      g01805(.A(new_n1921), .B(new_n1920), .C(new_n1918), .Y(new_n2062));
  A2O1A1O1Ixp25_ASAP7_75t_L g01806(.A1(new_n1784), .A2(new_n1669), .B(new_n1785), .C(new_n1924), .D(new_n2062), .Y(new_n2063));
  XOR2x2_ASAP7_75t_L        g01807(.A(new_n2061), .B(new_n2063), .Y(\f[24] ));
  NAND3xp33_ASAP7_75t_L     g01808(.A(new_n2058), .B(new_n2059), .C(new_n1938), .Y(new_n2065));
  NOR2xp33_ASAP7_75t_L      g01809(.A(\b[24] ), .B(\b[25] ), .Y(new_n2066));
  INVx1_ASAP7_75t_L         g01810(.A(\b[25] ), .Y(new_n2067));
  NOR2xp33_ASAP7_75t_L      g01811(.A(new_n1929), .B(new_n2067), .Y(new_n2068));
  NOR2xp33_ASAP7_75t_L      g01812(.A(new_n2066), .B(new_n2068), .Y(new_n2069));
  A2O1A1Ixp33_ASAP7_75t_L   g01813(.A1(\b[24] ), .A2(\b[23] ), .B(new_n1933), .C(new_n2069), .Y(new_n2070));
  INVx1_ASAP7_75t_L         g01814(.A(new_n2070), .Y(new_n2071));
  INVx1_ASAP7_75t_L         g01815(.A(new_n1930), .Y(new_n2072));
  A2O1A1Ixp33_ASAP7_75t_L   g01816(.A1(new_n1912), .A2(new_n1927), .B(new_n1928), .C(new_n2072), .Y(new_n2073));
  NOR2xp33_ASAP7_75t_L      g01817(.A(new_n2069), .B(new_n2073), .Y(new_n2074));
  OR2x4_ASAP7_75t_L         g01818(.A(new_n2071), .B(new_n2074), .Y(new_n2075));
  AOI22xp33_ASAP7_75t_L     g01819(.A1(\b[23] ), .A2(new_n282), .B1(\b[25] ), .B2(new_n303), .Y(new_n2076));
  OAI221xp5_ASAP7_75t_L     g01820(.A1(new_n291), .A2(new_n1929), .B1(new_n268), .B2(new_n2075), .C(new_n2076), .Y(new_n2077));
  XNOR2x2_ASAP7_75t_L       g01821(.A(\a[2] ), .B(new_n2077), .Y(new_n2078));
  NOR3xp33_ASAP7_75t_L      g01822(.A(new_n2046), .B(new_n2047), .C(new_n1942), .Y(new_n2079));
  INVx1_ASAP7_75t_L         g01823(.A(new_n2079), .Y(new_n2080));
  NAND2xp33_ASAP7_75t_L     g01824(.A(new_n1978), .B(new_n1980), .Y(new_n2081));
  AND3x1_ASAP7_75t_L        g01825(.A(new_n2081), .B(new_n1974), .C(new_n1973), .Y(new_n2082));
  NOR2xp33_ASAP7_75t_L      g01826(.A(new_n424), .B(new_n419), .Y(new_n2083));
  NOR2xp33_ASAP7_75t_L      g01827(.A(new_n492), .B(new_n2083), .Y(new_n2084));
  AOI22xp33_ASAP7_75t_L     g01828(.A1(new_n1360), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1581), .Y(new_n2085));
  INVx1_ASAP7_75t_L         g01829(.A(new_n2085), .Y(new_n2086));
  AOI221xp5_ASAP7_75t_L     g01830(.A1(new_n1362), .A2(\b[6] ), .B1(new_n1365), .B2(new_n2084), .C(new_n2086), .Y(new_n2087));
  NAND2xp33_ASAP7_75t_L     g01831(.A(\a[20] ), .B(new_n2087), .Y(new_n2088));
  OAI221xp5_ASAP7_75t_L     g01832(.A1(new_n1373), .A2(new_n418), .B1(new_n1359), .B2(new_n425), .C(new_n2085), .Y(new_n2089));
  NAND2xp33_ASAP7_75t_L     g01833(.A(new_n1356), .B(new_n2089), .Y(new_n2090));
  NOR2xp33_ASAP7_75t_L      g01834(.A(new_n1824), .B(new_n1839), .Y(new_n2091));
  NAND2xp33_ASAP7_75t_L     g01835(.A(new_n1962), .B(new_n2091), .Y(new_n2092));
  NOR2xp33_ASAP7_75t_L      g01836(.A(new_n298), .B(new_n1699), .Y(new_n2093));
  INVx1_ASAP7_75t_L         g01837(.A(new_n2093), .Y(new_n2094));
  NOR3xp33_ASAP7_75t_L      g01838(.A(new_n326), .B(new_n328), .C(new_n1827), .Y(new_n2095));
  INVx1_ASAP7_75t_L         g01839(.A(new_n2095), .Y(new_n2096));
  AOI22xp33_ASAP7_75t_L     g01840(.A1(new_n1704), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n1837), .Y(new_n2097));
  AND4x1_ASAP7_75t_L        g01841(.A(new_n2097), .B(new_n2096), .C(new_n2094), .D(\a[23] ), .Y(new_n2098));
  AOI31xp33_ASAP7_75t_L     g01842(.A1(new_n2096), .A2(new_n2094), .A3(new_n2097), .B(\a[23] ), .Y(new_n2099));
  INVx1_ASAP7_75t_L         g01843(.A(\a[26] ), .Y(new_n2100));
  NOR2xp33_ASAP7_75t_L      g01844(.A(new_n2100), .B(new_n1961), .Y(new_n2101));
  AND2x2_ASAP7_75t_L        g01845(.A(new_n1958), .B(new_n1959), .Y(new_n2102));
  INVx1_ASAP7_75t_L         g01846(.A(\a[25] ), .Y(new_n2103));
  NAND2xp33_ASAP7_75t_L     g01847(.A(\a[26] ), .B(new_n2103), .Y(new_n2104));
  NAND2xp33_ASAP7_75t_L     g01848(.A(\a[25] ), .B(new_n2100), .Y(new_n2105));
  AOI21xp33_ASAP7_75t_L     g01849(.A1(new_n2105), .A2(new_n2104), .B(new_n2102), .Y(new_n2106));
  NAND3xp33_ASAP7_75t_L     g01850(.A(new_n1960), .B(new_n2104), .C(new_n2105), .Y(new_n2107));
  XNOR2x2_ASAP7_75t_L       g01851(.A(\a[25] ), .B(\a[24] ), .Y(new_n2108));
  OR2x4_ASAP7_75t_L         g01852(.A(new_n2108), .B(new_n1960), .Y(new_n2109));
  OAI22xp33_ASAP7_75t_L     g01853(.A1(new_n2109), .A2(new_n258), .B1(new_n261), .B2(new_n2107), .Y(new_n2110));
  A2O1A1Ixp33_ASAP7_75t_L   g01854(.A1(new_n269), .A2(new_n2106), .B(new_n2110), .C(new_n2101), .Y(new_n2111));
  NAND2xp33_ASAP7_75t_L     g01855(.A(new_n269), .B(new_n2106), .Y(new_n2112));
  NAND2xp33_ASAP7_75t_L     g01856(.A(new_n2105), .B(new_n2104), .Y(new_n2113));
  NOR2xp33_ASAP7_75t_L      g01857(.A(new_n2113), .B(new_n2102), .Y(new_n2114));
  NOR2xp33_ASAP7_75t_L      g01858(.A(new_n2108), .B(new_n1960), .Y(new_n2115));
  AOI22xp33_ASAP7_75t_L     g01859(.A1(\b[0] ), .A2(new_n2115), .B1(\b[1] ), .B2(new_n2114), .Y(new_n2116));
  OAI211xp5_ASAP7_75t_L     g01860(.A1(new_n2100), .A2(new_n1961), .B(new_n2116), .C(new_n2112), .Y(new_n2117));
  NAND2xp33_ASAP7_75t_L     g01861(.A(new_n2117), .B(new_n2111), .Y(new_n2118));
  OR3x1_ASAP7_75t_L         g01862(.A(new_n2118), .B(new_n2098), .C(new_n2099), .Y(new_n2119));
  OAI21xp33_ASAP7_75t_L     g01863(.A1(new_n2099), .A2(new_n2098), .B(new_n2118), .Y(new_n2120));
  AOI22xp33_ASAP7_75t_L     g01864(.A1(new_n1973), .A2(new_n2092), .B1(new_n2119), .B2(new_n2120), .Y(new_n2121));
  AOI22xp33_ASAP7_75t_L     g01865(.A1(new_n1970), .A2(new_n1972), .B1(new_n1966), .B2(new_n1963), .Y(new_n2122));
  NAND2xp33_ASAP7_75t_L     g01866(.A(new_n1965), .B(new_n1831), .Y(new_n2123));
  NOR2xp33_ASAP7_75t_L      g01867(.A(new_n1961), .B(new_n2123), .Y(new_n2124));
  NOR3xp33_ASAP7_75t_L      g01868(.A(new_n2118), .B(new_n2098), .C(new_n2099), .Y(new_n2125));
  OA21x2_ASAP7_75t_L        g01869(.A1(new_n2099), .A2(new_n2098), .B(new_n2118), .Y(new_n2126));
  NOR4xp25_ASAP7_75t_L      g01870(.A(new_n2124), .B(new_n2126), .C(new_n2122), .D(new_n2125), .Y(new_n2127));
  AOI211xp5_ASAP7_75t_L     g01871(.A1(new_n2090), .A2(new_n2088), .B(new_n2127), .C(new_n2121), .Y(new_n2128));
  NOR2xp33_ASAP7_75t_L      g01872(.A(new_n1356), .B(new_n2089), .Y(new_n2129));
  NOR2xp33_ASAP7_75t_L      g01873(.A(\a[20] ), .B(new_n2087), .Y(new_n2130));
  OAI22xp33_ASAP7_75t_L     g01874(.A1(new_n2124), .A2(new_n2122), .B1(new_n2126), .B2(new_n2125), .Y(new_n2131));
  NAND4xp25_ASAP7_75t_L     g01875(.A(new_n2119), .B(new_n1973), .C(new_n2092), .D(new_n2120), .Y(new_n2132));
  AOI211xp5_ASAP7_75t_L     g01876(.A1(new_n2132), .A2(new_n2131), .B(new_n2129), .C(new_n2130), .Y(new_n2133));
  NOR2xp33_ASAP7_75t_L      g01877(.A(new_n2128), .B(new_n2133), .Y(new_n2134));
  A2O1A1Ixp33_ASAP7_75t_L   g01878(.A1(new_n1984), .A2(new_n1988), .B(new_n2082), .C(new_n2134), .Y(new_n2135));
  O2A1O1Ixp33_ASAP7_75t_L   g01879(.A1(new_n1981), .A2(new_n1982), .B(new_n1984), .C(new_n2082), .Y(new_n2136));
  OAI211xp5_ASAP7_75t_L     g01880(.A1(new_n2129), .A2(new_n2130), .B(new_n2132), .C(new_n2131), .Y(new_n2137));
  OAI211xp5_ASAP7_75t_L     g01881(.A1(new_n2127), .A2(new_n2121), .B(new_n2090), .C(new_n2088), .Y(new_n2138));
  NAND2xp33_ASAP7_75t_L     g01882(.A(new_n2137), .B(new_n2138), .Y(new_n2139));
  NAND2xp33_ASAP7_75t_L     g01883(.A(new_n2139), .B(new_n2136), .Y(new_n2140));
  NAND2xp33_ASAP7_75t_L     g01884(.A(\b[9] ), .B(new_n1080), .Y(new_n2141));
  INVx1_ASAP7_75t_L         g01885(.A(new_n623), .Y(new_n2142));
  NOR2xp33_ASAP7_75t_L      g01886(.A(new_n621), .B(new_n2142), .Y(new_n2143));
  NAND2xp33_ASAP7_75t_L     g01887(.A(new_n1073), .B(new_n2143), .Y(new_n2144));
  AOI22xp33_ASAP7_75t_L     g01888(.A1(new_n1076), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1253), .Y(new_n2145));
  NAND4xp25_ASAP7_75t_L     g01889(.A(new_n2144), .B(\a[17] ), .C(new_n2141), .D(new_n2145), .Y(new_n2146));
  NAND3xp33_ASAP7_75t_L     g01890(.A(new_n2144), .B(new_n2141), .C(new_n2145), .Y(new_n2147));
  NAND2xp33_ASAP7_75t_L     g01891(.A(new_n1071), .B(new_n2147), .Y(new_n2148));
  NAND4xp25_ASAP7_75t_L     g01892(.A(new_n2135), .B(new_n2148), .C(new_n2140), .D(new_n2146), .Y(new_n2149));
  NAND3xp33_ASAP7_75t_L     g01893(.A(new_n2081), .B(new_n1974), .C(new_n1973), .Y(new_n2150));
  O2A1O1Ixp33_ASAP7_75t_L   g01894(.A1(new_n1983), .A2(new_n1990), .B(new_n2150), .C(new_n2139), .Y(new_n2151));
  OAI21xp33_ASAP7_75t_L     g01895(.A1(new_n1983), .A2(new_n1990), .B(new_n2150), .Y(new_n2152));
  NOR2xp33_ASAP7_75t_L      g01896(.A(new_n2134), .B(new_n2152), .Y(new_n2153));
  NAND2xp33_ASAP7_75t_L     g01897(.A(new_n2146), .B(new_n2148), .Y(new_n2154));
  OAI21xp33_ASAP7_75t_L     g01898(.A1(new_n2151), .A2(new_n2153), .B(new_n2154), .Y(new_n2155));
  NAND2xp33_ASAP7_75t_L     g01899(.A(new_n2149), .B(new_n2155), .Y(new_n2156));
  OAI21xp33_ASAP7_75t_L     g01900(.A1(new_n1997), .A2(new_n1956), .B(new_n1999), .Y(new_n2157));
  NOR2xp33_ASAP7_75t_L      g01901(.A(new_n2157), .B(new_n2156), .Y(new_n2158));
  A2O1A1O1Ixp25_ASAP7_75t_L g01902(.A1(new_n1849), .A2(new_n1854), .B(new_n1851), .C(new_n2000), .D(new_n1996), .Y(new_n2159));
  AOI21xp33_ASAP7_75t_L     g01903(.A1(new_n2155), .A2(new_n2149), .B(new_n2159), .Y(new_n2160));
  AOI22xp33_ASAP7_75t_L     g01904(.A1(new_n811), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n900), .Y(new_n2161));
  OAI221xp5_ASAP7_75t_L     g01905(.A1(new_n904), .A2(new_n760), .B1(new_n898), .B2(new_n790), .C(new_n2161), .Y(new_n2162));
  XNOR2x2_ASAP7_75t_L       g01906(.A(\a[14] ), .B(new_n2162), .Y(new_n2163));
  OAI21xp33_ASAP7_75t_L     g01907(.A1(new_n2160), .A2(new_n2158), .B(new_n2163), .Y(new_n2164));
  NAND3xp33_ASAP7_75t_L     g01908(.A(new_n2159), .B(new_n2155), .C(new_n2149), .Y(new_n2165));
  INVx1_ASAP7_75t_L         g01909(.A(new_n2160), .Y(new_n2166));
  INVx1_ASAP7_75t_L         g01910(.A(new_n2163), .Y(new_n2167));
  NAND3xp33_ASAP7_75t_L     g01911(.A(new_n2166), .B(new_n2165), .C(new_n2167), .Y(new_n2168));
  OAI21xp33_ASAP7_75t_L     g01912(.A1(new_n2010), .A2(new_n2009), .B(new_n2007), .Y(new_n2169));
  NAND3xp33_ASAP7_75t_L     g01913(.A(new_n2169), .B(new_n2168), .C(new_n2164), .Y(new_n2170));
  AOI21xp33_ASAP7_75t_L     g01914(.A1(new_n2166), .A2(new_n2165), .B(new_n2167), .Y(new_n2171));
  NOR3xp33_ASAP7_75t_L      g01915(.A(new_n2158), .B(new_n2160), .C(new_n2163), .Y(new_n2172));
  A2O1A1O1Ixp25_ASAP7_75t_L g01916(.A1(new_n1857), .A2(new_n1803), .B(new_n1946), .C(new_n2002), .D(new_n2011), .Y(new_n2173));
  OAI21xp33_ASAP7_75t_L     g01917(.A1(new_n2172), .A2(new_n2171), .B(new_n2173), .Y(new_n2174));
  AOI22xp33_ASAP7_75t_L     g01918(.A1(\b[14] ), .A2(new_n651), .B1(\b[16] ), .B2(new_n581), .Y(new_n2175));
  OAI221xp5_ASAP7_75t_L     g01919(.A1(new_n821), .A2(new_n942), .B1(new_n577), .B2(new_n1035), .C(new_n2175), .Y(new_n2176));
  XNOR2x2_ASAP7_75t_L       g01920(.A(\a[11] ), .B(new_n2176), .Y(new_n2177));
  NAND3xp33_ASAP7_75t_L     g01921(.A(new_n2170), .B(new_n2174), .C(new_n2177), .Y(new_n2178));
  NOR3xp33_ASAP7_75t_L      g01922(.A(new_n2173), .B(new_n2172), .C(new_n2171), .Y(new_n2179));
  AOI221xp5_ASAP7_75t_L     g01923(.A1(new_n1947), .A2(new_n2002), .B1(new_n2164), .B2(new_n2168), .C(new_n2011), .Y(new_n2180));
  NOR2xp33_ASAP7_75t_L      g01924(.A(new_n574), .B(new_n2176), .Y(new_n2181));
  AND2x2_ASAP7_75t_L        g01925(.A(new_n574), .B(new_n2176), .Y(new_n2182));
  OAI22xp33_ASAP7_75t_L     g01926(.A1(new_n2180), .A2(new_n2179), .B1(new_n2182), .B2(new_n2181), .Y(new_n2183));
  NAND2xp33_ASAP7_75t_L     g01927(.A(new_n2183), .B(new_n2178), .Y(new_n2184));
  MAJIxp5_ASAP7_75t_L       g01928(.A(new_n2029), .B(new_n2013), .C(new_n2016), .Y(new_n2185));
  OR2x4_ASAP7_75t_L         g01929(.A(new_n2184), .B(new_n2185), .Y(new_n2186));
  NAND2xp33_ASAP7_75t_L     g01930(.A(new_n2184), .B(new_n2185), .Y(new_n2187));
  AOI22xp33_ASAP7_75t_L     g01931(.A1(new_n444), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n471), .Y(new_n2188));
  OAI221xp5_ASAP7_75t_L     g01932(.A1(new_n468), .A2(new_n1313), .B1(new_n469), .B2(new_n1438), .C(new_n2188), .Y(new_n2189));
  XNOR2x2_ASAP7_75t_L       g01933(.A(\a[8] ), .B(new_n2189), .Y(new_n2190));
  AND3x1_ASAP7_75t_L        g01934(.A(new_n2186), .B(new_n2190), .C(new_n2187), .Y(new_n2191));
  AOI21xp33_ASAP7_75t_L     g01935(.A1(new_n2186), .A2(new_n2187), .B(new_n2190), .Y(new_n2192));
  NOR3xp33_ASAP7_75t_L      g01936(.A(new_n2025), .B(new_n2034), .C(new_n2030), .Y(new_n2193));
  A2O1A1O1Ixp25_ASAP7_75t_L g01937(.A1(new_n1880), .A2(new_n1882), .B(new_n1943), .C(new_n2035), .D(new_n2193), .Y(new_n2194));
  OA21x2_ASAP7_75t_L        g01938(.A1(new_n2192), .A2(new_n2191), .B(new_n2194), .Y(new_n2195));
  NOR3xp33_ASAP7_75t_L      g01939(.A(new_n2191), .B(new_n2194), .C(new_n2192), .Y(new_n2196));
  AOI22xp33_ASAP7_75t_L     g01940(.A1(new_n344), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n370), .Y(new_n2197));
  OAI221xp5_ASAP7_75t_L     g01941(.A1(new_n429), .A2(new_n1655), .B1(new_n366), .B2(new_n1780), .C(new_n2197), .Y(new_n2198));
  XNOR2x2_ASAP7_75t_L       g01942(.A(\a[5] ), .B(new_n2198), .Y(new_n2199));
  INVx1_ASAP7_75t_L         g01943(.A(new_n2199), .Y(new_n2200));
  OAI21xp33_ASAP7_75t_L     g01944(.A1(new_n2196), .A2(new_n2195), .B(new_n2200), .Y(new_n2201));
  OAI21xp33_ASAP7_75t_L     g01945(.A1(new_n2192), .A2(new_n2191), .B(new_n2194), .Y(new_n2202));
  OR3x1_ASAP7_75t_L         g01946(.A(new_n2191), .B(new_n2194), .C(new_n2192), .Y(new_n2203));
  NAND3xp33_ASAP7_75t_L     g01947(.A(new_n2203), .B(new_n2202), .C(new_n2199), .Y(new_n2204));
  NAND2xp33_ASAP7_75t_L     g01948(.A(new_n2201), .B(new_n2204), .Y(new_n2205));
  O2A1O1Ixp33_ASAP7_75t_L   g01949(.A1(new_n1939), .A2(new_n2049), .B(new_n2080), .C(new_n2205), .Y(new_n2206));
  INVx1_ASAP7_75t_L         g01950(.A(new_n1939), .Y(new_n2207));
  AOI221xp5_ASAP7_75t_L     g01951(.A1(new_n2204), .A2(new_n2201), .B1(new_n2053), .B2(new_n2207), .C(new_n2079), .Y(new_n2208));
  NOR3xp33_ASAP7_75t_L      g01952(.A(new_n2208), .B(new_n2206), .C(new_n2078), .Y(new_n2209));
  XNOR2x2_ASAP7_75t_L       g01953(.A(new_n262), .B(new_n2077), .Y(new_n2210));
  A2O1A1Ixp33_ASAP7_75t_L   g01954(.A1(new_n2051), .A2(new_n2052), .B(new_n1939), .C(new_n2080), .Y(new_n2211));
  NAND3xp33_ASAP7_75t_L     g01955(.A(new_n2211), .B(new_n2201), .C(new_n2204), .Y(new_n2212));
  O2A1O1Ixp33_ASAP7_75t_L   g01956(.A1(new_n1903), .A2(new_n1921), .B(new_n2053), .C(new_n2079), .Y(new_n2213));
  NAND2xp33_ASAP7_75t_L     g01957(.A(new_n2205), .B(new_n2213), .Y(new_n2214));
  AOI21xp33_ASAP7_75t_L     g01958(.A1(new_n2212), .A2(new_n2214), .B(new_n2210), .Y(new_n2215));
  NOR2xp33_ASAP7_75t_L      g01959(.A(new_n2209), .B(new_n2215), .Y(new_n2216));
  INVx1_ASAP7_75t_L         g01960(.A(new_n2216), .Y(new_n2217));
  O2A1O1Ixp33_ASAP7_75t_L   g01961(.A1(new_n2061), .A2(new_n2063), .B(new_n2065), .C(new_n2217), .Y(new_n2218));
  OAI21xp33_ASAP7_75t_L     g01962(.A1(new_n2061), .A2(new_n2063), .B(new_n2065), .Y(new_n2219));
  NOR2xp33_ASAP7_75t_L      g01963(.A(new_n2216), .B(new_n2219), .Y(new_n2220));
  NOR2xp33_ASAP7_75t_L      g01964(.A(new_n2220), .B(new_n2218), .Y(\f[25] ));
  NOR2xp33_ASAP7_75t_L      g01965(.A(new_n2209), .B(new_n2218), .Y(new_n2222));
  AOI21xp33_ASAP7_75t_L     g01966(.A1(new_n2203), .A2(new_n2202), .B(new_n2199), .Y(new_n2223));
  NAND2xp33_ASAP7_75t_L     g01967(.A(new_n2174), .B(new_n2170), .Y(new_n2224));
  NOR2xp33_ASAP7_75t_L      g01968(.A(new_n2177), .B(new_n2224), .Y(new_n2225));
  NOR2xp33_ASAP7_75t_L      g01969(.A(new_n1030), .B(new_n821), .Y(new_n2226));
  AOI22xp33_ASAP7_75t_L     g01970(.A1(\b[15] ), .A2(new_n651), .B1(\b[17] ), .B2(new_n581), .Y(new_n2227));
  OAI31xp33_ASAP7_75t_L     g01971(.A1(new_n1796), .A2(new_n577), .A3(new_n1205), .B(new_n2227), .Y(new_n2228));
  OR3x1_ASAP7_75t_L         g01972(.A(new_n2228), .B(new_n574), .C(new_n2226), .Y(new_n2229));
  A2O1A1Ixp33_ASAP7_75t_L   g01973(.A1(\b[16] ), .A2(new_n584), .B(new_n2228), .C(new_n574), .Y(new_n2230));
  NAND2xp33_ASAP7_75t_L     g01974(.A(new_n2230), .B(new_n2229), .Y(new_n2231));
  OAI21xp33_ASAP7_75t_L     g01975(.A1(new_n2171), .A2(new_n2173), .B(new_n2168), .Y(new_n2232));
  NAND3xp33_ASAP7_75t_L     g01976(.A(new_n2154), .B(new_n2135), .C(new_n2140), .Y(new_n2233));
  AOI22xp33_ASAP7_75t_L     g01977(.A1(new_n1076), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1253), .Y(new_n2234));
  OAI221xp5_ASAP7_75t_L     g01978(.A1(new_n1154), .A2(new_n617), .B1(new_n1156), .B2(new_n685), .C(new_n2234), .Y(new_n2235));
  XNOR2x2_ASAP7_75t_L       g01979(.A(\a[17] ), .B(new_n2235), .Y(new_n2236));
  A2O1A1O1Ixp25_ASAP7_75t_L g01980(.A1(new_n1984), .A2(new_n1988), .B(new_n2082), .C(new_n2138), .D(new_n2128), .Y(new_n2237));
  AOI22xp33_ASAP7_75t_L     g01981(.A1(new_n1360), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1581), .Y(new_n2238));
  OAI221xp5_ASAP7_75t_L     g01982(.A1(new_n1373), .A2(new_n420), .B1(new_n1359), .B2(new_n494), .C(new_n2238), .Y(new_n2239));
  XNOR2x2_ASAP7_75t_L       g01983(.A(\a[20] ), .B(new_n2239), .Y(new_n2240));
  INVx1_ASAP7_75t_L         g01984(.A(new_n2240), .Y(new_n2241));
  XNOR2x2_ASAP7_75t_L       g01985(.A(new_n1689), .B(new_n1969), .Y(new_n2242));
  MAJIxp5_ASAP7_75t_L       g01986(.A(new_n2242), .B(new_n1961), .C(new_n2123), .Y(new_n2243));
  NOR2xp33_ASAP7_75t_L      g01987(.A(new_n2099), .B(new_n2098), .Y(new_n2244));
  NOR2xp33_ASAP7_75t_L      g01988(.A(new_n2118), .B(new_n2244), .Y(new_n2245));
  O2A1O1Ixp33_ASAP7_75t_L   g01989(.A1(new_n2125), .A2(new_n2126), .B(new_n2243), .C(new_n2245), .Y(new_n2246));
  NAND2xp33_ASAP7_75t_L     g01990(.A(\b[4] ), .B(new_n1706), .Y(new_n2247));
  INVx1_ASAP7_75t_L         g01991(.A(new_n2247), .Y(new_n2248));
  NOR3xp33_ASAP7_75t_L      g01992(.A(new_n357), .B(new_n358), .C(new_n1827), .Y(new_n2249));
  OAI22xp33_ASAP7_75t_L     g01993(.A1(new_n1829), .A2(new_n298), .B1(new_n354), .B2(new_n1696), .Y(new_n2250));
  NOR4xp25_ASAP7_75t_L      g01994(.A(new_n2249), .B(new_n1689), .C(new_n2250), .D(new_n2248), .Y(new_n2251));
  INVx1_ASAP7_75t_L         g01995(.A(new_n2251), .Y(new_n2252));
  OAI31xp33_ASAP7_75t_L     g01996(.A1(new_n2249), .A2(new_n2248), .A3(new_n2250), .B(new_n1689), .Y(new_n2253));
  NAND2xp33_ASAP7_75t_L     g01997(.A(new_n2112), .B(new_n2116), .Y(new_n2254));
  NOR2xp33_ASAP7_75t_L      g01998(.A(new_n261), .B(new_n2109), .Y(new_n2255));
  INVx1_ASAP7_75t_L         g01999(.A(new_n2255), .Y(new_n2256));
  NAND2xp33_ASAP7_75t_L     g02000(.A(new_n2113), .B(new_n1960), .Y(new_n2257));
  NOR2xp33_ASAP7_75t_L      g02001(.A(new_n280), .B(new_n2257), .Y(new_n2258));
  AND3x1_ASAP7_75t_L        g02002(.A(new_n2102), .B(new_n2108), .C(new_n2113), .Y(new_n2259));
  AOI221xp5_ASAP7_75t_L     g02003(.A1(new_n2114), .A2(\b[2] ), .B1(new_n2259), .B2(\b[0] ), .C(new_n2258), .Y(new_n2260));
  NAND2xp33_ASAP7_75t_L     g02004(.A(new_n2256), .B(new_n2260), .Y(new_n2261));
  O2A1O1Ixp33_ASAP7_75t_L   g02005(.A1(new_n1962), .A2(new_n2254), .B(\a[26] ), .C(new_n2261), .Y(new_n2262));
  A2O1A1Ixp33_ASAP7_75t_L   g02006(.A1(\b[0] ), .A2(new_n1960), .B(new_n2254), .C(\a[26] ), .Y(new_n2263));
  O2A1O1Ixp33_ASAP7_75t_L   g02007(.A1(new_n2109), .A2(new_n261), .B(new_n2260), .C(new_n2263), .Y(new_n2264));
  OAI211xp5_ASAP7_75t_L     g02008(.A1(new_n2262), .A2(new_n2264), .B(new_n2253), .C(new_n2252), .Y(new_n2265));
  INVx1_ASAP7_75t_L         g02009(.A(new_n2253), .Y(new_n2266));
  AOI21xp33_ASAP7_75t_L     g02010(.A1(new_n2106), .A2(new_n269), .B(new_n2110), .Y(new_n2267));
  NAND2xp33_ASAP7_75t_L     g02011(.A(\b[2] ), .B(new_n2114), .Y(new_n2268));
  NAND3xp33_ASAP7_75t_L     g02012(.A(new_n2102), .B(new_n2113), .C(new_n2108), .Y(new_n2269));
  OAI221xp5_ASAP7_75t_L     g02013(.A1(new_n258), .A2(new_n2269), .B1(new_n280), .B2(new_n2257), .C(new_n2268), .Y(new_n2270));
  NOR2xp33_ASAP7_75t_L      g02014(.A(new_n2255), .B(new_n2270), .Y(new_n2271));
  A2O1A1Ixp33_ASAP7_75t_L   g02015(.A1(new_n1961), .A2(new_n2267), .B(new_n2100), .C(new_n2271), .Y(new_n2272));
  O2A1O1Ixp33_ASAP7_75t_L   g02016(.A1(new_n258), .A2(new_n2102), .B(new_n2267), .C(new_n2100), .Y(new_n2273));
  A2O1A1Ixp33_ASAP7_75t_L   g02017(.A1(\b[1] ), .A2(new_n2115), .B(new_n2270), .C(new_n2273), .Y(new_n2274));
  OAI211xp5_ASAP7_75t_L     g02018(.A1(new_n2251), .A2(new_n2266), .B(new_n2274), .C(new_n2272), .Y(new_n2275));
  NAND2xp33_ASAP7_75t_L     g02019(.A(new_n2265), .B(new_n2275), .Y(new_n2276));
  NAND2xp33_ASAP7_75t_L     g02020(.A(new_n2276), .B(new_n2246), .Y(new_n2277));
  NAND2xp33_ASAP7_75t_L     g02021(.A(new_n1972), .B(new_n1970), .Y(new_n2278));
  MAJIxp5_ASAP7_75t_L       g02022(.A(new_n2278), .B(new_n1962), .C(new_n2091), .Y(new_n2279));
  MAJIxp5_ASAP7_75t_L       g02023(.A(new_n2279), .B(new_n2244), .C(new_n2118), .Y(new_n2280));
  NAND3xp33_ASAP7_75t_L     g02024(.A(new_n2280), .B(new_n2265), .C(new_n2275), .Y(new_n2281));
  AOI21xp33_ASAP7_75t_L     g02025(.A1(new_n2281), .A2(new_n2277), .B(new_n2241), .Y(new_n2282));
  AOI21xp33_ASAP7_75t_L     g02026(.A1(new_n2275), .A2(new_n2265), .B(new_n2280), .Y(new_n2283));
  O2A1O1Ixp33_ASAP7_75t_L   g02027(.A1(new_n2244), .A2(new_n2118), .B(new_n2131), .C(new_n2276), .Y(new_n2284));
  NOR3xp33_ASAP7_75t_L      g02028(.A(new_n2284), .B(new_n2283), .C(new_n2240), .Y(new_n2285));
  NOR3xp33_ASAP7_75t_L      g02029(.A(new_n2282), .B(new_n2237), .C(new_n2285), .Y(new_n2286));
  OAI221xp5_ASAP7_75t_L     g02030(.A1(new_n1981), .A2(new_n1982), .B1(new_n1847), .B2(new_n1816), .C(new_n1833), .Y(new_n2287));
  A2O1A1Ixp33_ASAP7_75t_L   g02031(.A1(new_n2287), .A2(new_n2150), .B(new_n2133), .C(new_n2137), .Y(new_n2288));
  OAI21xp33_ASAP7_75t_L     g02032(.A1(new_n2283), .A2(new_n2284), .B(new_n2240), .Y(new_n2289));
  NAND3xp33_ASAP7_75t_L     g02033(.A(new_n2241), .B(new_n2277), .C(new_n2281), .Y(new_n2290));
  AOI21xp33_ASAP7_75t_L     g02034(.A1(new_n2290), .A2(new_n2289), .B(new_n2288), .Y(new_n2291));
  OAI21xp33_ASAP7_75t_L     g02035(.A1(new_n2286), .A2(new_n2291), .B(new_n2236), .Y(new_n2292));
  NOR2xp33_ASAP7_75t_L      g02036(.A(new_n1071), .B(new_n2235), .Y(new_n2293));
  AND2x2_ASAP7_75t_L        g02037(.A(new_n1071), .B(new_n2235), .Y(new_n2294));
  NAND3xp33_ASAP7_75t_L     g02038(.A(new_n2288), .B(new_n2289), .C(new_n2290), .Y(new_n2295));
  OAI21xp33_ASAP7_75t_L     g02039(.A1(new_n2285), .A2(new_n2282), .B(new_n2237), .Y(new_n2296));
  OAI211xp5_ASAP7_75t_L     g02040(.A1(new_n2294), .A2(new_n2293), .B(new_n2295), .C(new_n2296), .Y(new_n2297));
  NAND2xp33_ASAP7_75t_L     g02041(.A(new_n2292), .B(new_n2297), .Y(new_n2298));
  A2O1A1O1Ixp25_ASAP7_75t_L g02042(.A1(new_n2155), .A2(new_n2149), .B(new_n2159), .C(new_n2233), .D(new_n2298), .Y(new_n2299));
  A2O1A1Ixp33_ASAP7_75t_L   g02043(.A1(new_n2155), .A2(new_n2149), .B(new_n2159), .C(new_n2233), .Y(new_n2300));
  AOI21xp33_ASAP7_75t_L     g02044(.A1(new_n2297), .A2(new_n2292), .B(new_n2300), .Y(new_n2301));
  AOI22xp33_ASAP7_75t_L     g02045(.A1(new_n811), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n900), .Y(new_n2302));
  OAI221xp5_ASAP7_75t_L     g02046(.A1(new_n904), .A2(new_n784), .B1(new_n898), .B2(new_n875), .C(new_n2302), .Y(new_n2303));
  XNOR2x2_ASAP7_75t_L       g02047(.A(\a[14] ), .B(new_n2303), .Y(new_n2304));
  INVx1_ASAP7_75t_L         g02048(.A(new_n2304), .Y(new_n2305));
  NOR3xp33_ASAP7_75t_L      g02049(.A(new_n2299), .B(new_n2305), .C(new_n2301), .Y(new_n2306));
  NAND3xp33_ASAP7_75t_L     g02050(.A(new_n2300), .B(new_n2292), .C(new_n2297), .Y(new_n2307));
  AO21x2_ASAP7_75t_L        g02051(.A1(new_n2297), .A2(new_n2292), .B(new_n2300), .Y(new_n2308));
  AOI21xp33_ASAP7_75t_L     g02052(.A1(new_n2308), .A2(new_n2307), .B(new_n2304), .Y(new_n2309));
  OAI21xp33_ASAP7_75t_L     g02053(.A1(new_n2309), .A2(new_n2306), .B(new_n2232), .Y(new_n2310));
  A2O1A1O1Ixp25_ASAP7_75t_L g02054(.A1(new_n2002), .A2(new_n1947), .B(new_n2011), .C(new_n2164), .D(new_n2172), .Y(new_n2311));
  NAND3xp33_ASAP7_75t_L     g02055(.A(new_n2308), .B(new_n2307), .C(new_n2304), .Y(new_n2312));
  OAI21xp33_ASAP7_75t_L     g02056(.A1(new_n2301), .A2(new_n2299), .B(new_n2305), .Y(new_n2313));
  NAND3xp33_ASAP7_75t_L     g02057(.A(new_n2311), .B(new_n2312), .C(new_n2313), .Y(new_n2314));
  NAND3xp33_ASAP7_75t_L     g02058(.A(new_n2314), .B(new_n2310), .C(new_n2231), .Y(new_n2315));
  AO21x2_ASAP7_75t_L        g02059(.A1(new_n2310), .A2(new_n2314), .B(new_n2231), .Y(new_n2316));
  AOI221xp5_ASAP7_75t_L     g02060(.A1(new_n2185), .A2(new_n2184), .B1(new_n2315), .B2(new_n2316), .C(new_n2225), .Y(new_n2317));
  NAND2xp33_ASAP7_75t_L     g02061(.A(new_n2315), .B(new_n2316), .Y(new_n2318));
  O2A1O1Ixp33_ASAP7_75t_L   g02062(.A1(new_n2224), .A2(new_n2177), .B(new_n2187), .C(new_n2318), .Y(new_n2319));
  AOI22xp33_ASAP7_75t_L     g02063(.A1(new_n444), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n471), .Y(new_n2320));
  INVx1_ASAP7_75t_L         g02064(.A(new_n2320), .Y(new_n2321));
  AOI221xp5_ASAP7_75t_L     g02065(.A1(\b[19] ), .A2(new_n447), .B1(new_n441), .B2(new_n1886), .C(new_n2321), .Y(new_n2322));
  XNOR2x2_ASAP7_75t_L       g02066(.A(\a[8] ), .B(new_n2322), .Y(new_n2323));
  NOR3xp33_ASAP7_75t_L      g02067(.A(new_n2319), .B(new_n2323), .C(new_n2317), .Y(new_n2324));
  OAI211xp5_ASAP7_75t_L     g02068(.A1(new_n2224), .A2(new_n2177), .B(new_n2318), .C(new_n2187), .Y(new_n2325));
  AND3x1_ASAP7_75t_L        g02069(.A(new_n2314), .B(new_n2310), .C(new_n2231), .Y(new_n2326));
  AOI21xp33_ASAP7_75t_L     g02070(.A1(new_n2314), .A2(new_n2310), .B(new_n2231), .Y(new_n2327));
  NOR2xp33_ASAP7_75t_L      g02071(.A(new_n2327), .B(new_n2326), .Y(new_n2328));
  A2O1A1Ixp33_ASAP7_75t_L   g02072(.A1(new_n2185), .A2(new_n2184), .B(new_n2225), .C(new_n2328), .Y(new_n2329));
  XNOR2x2_ASAP7_75t_L       g02073(.A(new_n435), .B(new_n2322), .Y(new_n2330));
  AOI21xp33_ASAP7_75t_L     g02074(.A1(new_n2325), .A2(new_n2329), .B(new_n2330), .Y(new_n2331));
  NOR2xp33_ASAP7_75t_L      g02075(.A(new_n2331), .B(new_n2324), .Y(new_n2332));
  XNOR2x2_ASAP7_75t_L       g02076(.A(new_n2184), .B(new_n2185), .Y(new_n2333));
  MAJx2_ASAP7_75t_L         g02077(.A(new_n2194), .B(new_n2190), .C(new_n2333), .Y(new_n2334));
  NAND2xp33_ASAP7_75t_L     g02078(.A(new_n2332), .B(new_n2334), .Y(new_n2335));
  MAJIxp5_ASAP7_75t_L       g02079(.A(new_n2194), .B(new_n2333), .C(new_n2190), .Y(new_n2336));
  OAI21xp33_ASAP7_75t_L     g02080(.A1(new_n2324), .A2(new_n2331), .B(new_n2336), .Y(new_n2337));
  AOI22xp33_ASAP7_75t_L     g02081(.A1(new_n344), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n370), .Y(new_n2338));
  OAI221xp5_ASAP7_75t_L     g02082(.A1(new_n429), .A2(new_n1774), .B1(new_n366), .B2(new_n1915), .C(new_n2338), .Y(new_n2339));
  XNOR2x2_ASAP7_75t_L       g02083(.A(\a[5] ), .B(new_n2339), .Y(new_n2340));
  NAND3xp33_ASAP7_75t_L     g02084(.A(new_n2335), .B(new_n2337), .C(new_n2340), .Y(new_n2341));
  AO21x2_ASAP7_75t_L        g02085(.A1(new_n2337), .A2(new_n2335), .B(new_n2340), .Y(new_n2342));
  OAI211xp5_ASAP7_75t_L     g02086(.A1(new_n2223), .A2(new_n2206), .B(new_n2341), .C(new_n2342), .Y(new_n2343));
  A2O1A1O1Ixp25_ASAP7_75t_L g02087(.A1(new_n2053), .A2(new_n2207), .B(new_n2079), .C(new_n2204), .D(new_n2223), .Y(new_n2344));
  NAND2xp33_ASAP7_75t_L     g02088(.A(new_n2341), .B(new_n2342), .Y(new_n2345));
  NAND2xp33_ASAP7_75t_L     g02089(.A(new_n2345), .B(new_n2344), .Y(new_n2346));
  NOR2xp33_ASAP7_75t_L      g02090(.A(\b[25] ), .B(\b[26] ), .Y(new_n2347));
  INVx1_ASAP7_75t_L         g02091(.A(\b[26] ), .Y(new_n2348));
  NOR2xp33_ASAP7_75t_L      g02092(.A(new_n2067), .B(new_n2348), .Y(new_n2349));
  NOR2xp33_ASAP7_75t_L      g02093(.A(new_n2347), .B(new_n2349), .Y(new_n2350));
  A2O1A1Ixp33_ASAP7_75t_L   g02094(.A1(new_n2073), .A2(new_n2069), .B(new_n2068), .C(new_n2350), .Y(new_n2351));
  O2A1O1Ixp33_ASAP7_75t_L   g02095(.A1(new_n1930), .A2(new_n1933), .B(new_n2069), .C(new_n2068), .Y(new_n2352));
  INVx1_ASAP7_75t_L         g02096(.A(new_n2350), .Y(new_n2353));
  NAND2xp33_ASAP7_75t_L     g02097(.A(new_n2353), .B(new_n2352), .Y(new_n2354));
  NAND2xp33_ASAP7_75t_L     g02098(.A(new_n2354), .B(new_n2351), .Y(new_n2355));
  AOI22xp33_ASAP7_75t_L     g02099(.A1(\b[24] ), .A2(new_n282), .B1(\b[26] ), .B2(new_n303), .Y(new_n2356));
  OAI221xp5_ASAP7_75t_L     g02100(.A1(new_n291), .A2(new_n2067), .B1(new_n268), .B2(new_n2355), .C(new_n2356), .Y(new_n2357));
  XNOR2x2_ASAP7_75t_L       g02101(.A(\a[2] ), .B(new_n2357), .Y(new_n2358));
  AOI21xp33_ASAP7_75t_L     g02102(.A1(new_n2343), .A2(new_n2346), .B(new_n2358), .Y(new_n2359));
  INVx1_ASAP7_75t_L         g02103(.A(new_n2359), .Y(new_n2360));
  NAND3xp33_ASAP7_75t_L     g02104(.A(new_n2343), .B(new_n2346), .C(new_n2358), .Y(new_n2361));
  NAND2xp33_ASAP7_75t_L     g02105(.A(new_n2361), .B(new_n2360), .Y(new_n2362));
  XOR2x2_ASAP7_75t_L        g02106(.A(new_n2362), .B(new_n2222), .Y(\f[26] ));
  NAND3xp33_ASAP7_75t_L     g02107(.A(new_n2325), .B(new_n2329), .C(new_n2330), .Y(new_n2364));
  OAI21xp33_ASAP7_75t_L     g02108(.A1(new_n2317), .A2(new_n2319), .B(new_n2323), .Y(new_n2365));
  NAND2xp33_ASAP7_75t_L     g02109(.A(new_n2365), .B(new_n2364), .Y(new_n2366));
  NOR3xp33_ASAP7_75t_L      g02110(.A(new_n2291), .B(new_n2236), .C(new_n2286), .Y(new_n2367));
  AO21x2_ASAP7_75t_L        g02111(.A1(new_n2292), .A2(new_n2300), .B(new_n2367), .Y(new_n2368));
  NAND2xp33_ASAP7_75t_L     g02112(.A(\b[11] ), .B(new_n1080), .Y(new_n2369));
  NAND3xp33_ASAP7_75t_L     g02113(.A(new_n765), .B(new_n767), .C(new_n1073), .Y(new_n2370));
  AOI22xp33_ASAP7_75t_L     g02114(.A1(new_n1076), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1253), .Y(new_n2371));
  NAND4xp25_ASAP7_75t_L     g02115(.A(new_n2370), .B(\a[17] ), .C(new_n2369), .D(new_n2371), .Y(new_n2372));
  OAI31xp33_ASAP7_75t_L     g02116(.A1(new_n1231), .A2(new_n764), .A3(new_n1156), .B(new_n2371), .Y(new_n2373));
  A2O1A1Ixp33_ASAP7_75t_L   g02117(.A1(\b[11] ), .A2(new_n1080), .B(new_n2373), .C(new_n1071), .Y(new_n2374));
  NAND2xp33_ASAP7_75t_L     g02118(.A(new_n2372), .B(new_n2374), .Y(new_n2375));
  OAI21xp33_ASAP7_75t_L     g02119(.A1(new_n2237), .A2(new_n2282), .B(new_n2290), .Y(new_n2376));
  AOI211xp5_ASAP7_75t_L     g02120(.A1(new_n2253), .A2(new_n2252), .B(new_n2262), .C(new_n2264), .Y(new_n2377));
  NAND4xp25_ASAP7_75t_L     g02121(.A(new_n2116), .B(\a[26] ), .C(new_n1961), .D(new_n2112), .Y(new_n2378));
  INVx1_ASAP7_75t_L         g02122(.A(\a[27] ), .Y(new_n2379));
  NAND2xp33_ASAP7_75t_L     g02123(.A(\a[26] ), .B(new_n2379), .Y(new_n2380));
  NAND2xp33_ASAP7_75t_L     g02124(.A(\a[27] ), .B(new_n2100), .Y(new_n2381));
  NAND2xp33_ASAP7_75t_L     g02125(.A(new_n2381), .B(new_n2380), .Y(new_n2382));
  NAND2xp33_ASAP7_75t_L     g02126(.A(\b[0] ), .B(new_n2382), .Y(new_n2383));
  INVx1_ASAP7_75t_L         g02127(.A(new_n2383), .Y(new_n2384));
  OAI31xp33_ASAP7_75t_L     g02128(.A1(new_n2378), .A2(new_n2270), .A3(new_n2255), .B(new_n2384), .Y(new_n2385));
  A2O1A1Ixp33_ASAP7_75t_L   g02129(.A1(new_n1958), .A2(new_n1959), .B(new_n258), .C(\a[26] ), .Y(new_n2386));
  AOI211xp5_ASAP7_75t_L     g02130(.A1(new_n2106), .A2(new_n269), .B(new_n2386), .C(new_n2110), .Y(new_n2387));
  NAND4xp25_ASAP7_75t_L     g02131(.A(new_n2387), .B(new_n2383), .C(new_n2260), .D(new_n2256), .Y(new_n2388));
  NOR2xp33_ASAP7_75t_L      g02132(.A(new_n276), .B(new_n2109), .Y(new_n2389));
  OAI22xp33_ASAP7_75t_L     g02133(.A1(new_n2269), .A2(new_n261), .B1(new_n298), .B2(new_n2107), .Y(new_n2390));
  AOI211xp5_ASAP7_75t_L     g02134(.A1(new_n406), .A2(new_n2106), .B(new_n2389), .C(new_n2390), .Y(new_n2391));
  NAND2xp33_ASAP7_75t_L     g02135(.A(\a[26] ), .B(new_n2391), .Y(new_n2392));
  NOR2xp33_ASAP7_75t_L      g02136(.A(new_n2257), .B(new_n302), .Y(new_n2393));
  OAI31xp33_ASAP7_75t_L     g02137(.A1(new_n2393), .A2(new_n2389), .A3(new_n2390), .B(new_n2100), .Y(new_n2394));
  AOI22xp33_ASAP7_75t_L     g02138(.A1(new_n2392), .A2(new_n2394), .B1(new_n2385), .B2(new_n2388), .Y(new_n2395));
  AND4x1_ASAP7_75t_L        g02139(.A(new_n2388), .B(new_n2385), .C(new_n2394), .D(new_n2392), .Y(new_n2396));
  NAND2xp33_ASAP7_75t_L     g02140(.A(\b[5] ), .B(new_n1706), .Y(new_n2397));
  NAND2xp33_ASAP7_75t_L     g02141(.A(new_n1695), .B(new_n526), .Y(new_n2398));
  AOI22xp33_ASAP7_75t_L     g02142(.A1(new_n1704), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1837), .Y(new_n2399));
  NAND4xp25_ASAP7_75t_L     g02143(.A(new_n2398), .B(\a[23] ), .C(new_n2397), .D(new_n2399), .Y(new_n2400));
  INVx1_ASAP7_75t_L         g02144(.A(new_n2400), .Y(new_n2401));
  AOI31xp33_ASAP7_75t_L     g02145(.A1(new_n2398), .A2(new_n2397), .A3(new_n2399), .B(\a[23] ), .Y(new_n2402));
  NOR4xp25_ASAP7_75t_L      g02146(.A(new_n2401), .B(new_n2396), .C(new_n2395), .D(new_n2402), .Y(new_n2403));
  AO22x1_ASAP7_75t_L        g02147(.A1(new_n2394), .A2(new_n2392), .B1(new_n2385), .B2(new_n2388), .Y(new_n2404));
  NAND4xp25_ASAP7_75t_L     g02148(.A(new_n2388), .B(new_n2385), .C(new_n2392), .D(new_n2394), .Y(new_n2405));
  INVx1_ASAP7_75t_L         g02149(.A(new_n2402), .Y(new_n2406));
  AOI22xp33_ASAP7_75t_L     g02150(.A1(new_n2404), .A2(new_n2405), .B1(new_n2400), .B2(new_n2406), .Y(new_n2407));
  NOR2xp33_ASAP7_75t_L      g02151(.A(new_n2403), .B(new_n2407), .Y(new_n2408));
  OAI211xp5_ASAP7_75t_L     g02152(.A1(new_n2280), .A2(new_n2377), .B(new_n2408), .C(new_n2265), .Y(new_n2409));
  AOI211xp5_ASAP7_75t_L     g02153(.A1(new_n2274), .A2(new_n2272), .B(new_n2251), .C(new_n2266), .Y(new_n2410));
  NAND4xp25_ASAP7_75t_L     g02154(.A(new_n2406), .B(new_n2404), .C(new_n2405), .D(new_n2400), .Y(new_n2411));
  OAI22xp33_ASAP7_75t_L     g02155(.A1(new_n2401), .A2(new_n2402), .B1(new_n2395), .B2(new_n2396), .Y(new_n2412));
  NAND2xp33_ASAP7_75t_L     g02156(.A(new_n2412), .B(new_n2411), .Y(new_n2413));
  A2O1A1Ixp33_ASAP7_75t_L   g02157(.A1(new_n2275), .A2(new_n2246), .B(new_n2410), .C(new_n2413), .Y(new_n2414));
  AOI22xp33_ASAP7_75t_L     g02158(.A1(new_n1360), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1581), .Y(new_n2415));
  OAI221xp5_ASAP7_75t_L     g02159(.A1(new_n1373), .A2(new_n488), .B1(new_n1359), .B2(new_n548), .C(new_n2415), .Y(new_n2416));
  OR2x4_ASAP7_75t_L         g02160(.A(new_n1356), .B(new_n2416), .Y(new_n2417));
  NAND2xp33_ASAP7_75t_L     g02161(.A(new_n1356), .B(new_n2416), .Y(new_n2418));
  AO22x1_ASAP7_75t_L        g02162(.A1(new_n2418), .A2(new_n2417), .B1(new_n2414), .B2(new_n2409), .Y(new_n2419));
  NAND4xp25_ASAP7_75t_L     g02163(.A(new_n2409), .B(new_n2418), .C(new_n2414), .D(new_n2417), .Y(new_n2420));
  NAND3xp33_ASAP7_75t_L     g02164(.A(new_n2376), .B(new_n2419), .C(new_n2420), .Y(new_n2421));
  A2O1A1O1Ixp25_ASAP7_75t_L g02165(.A1(new_n2134), .A2(new_n2152), .B(new_n2128), .C(new_n2289), .D(new_n2285), .Y(new_n2422));
  AOI22xp33_ASAP7_75t_L     g02166(.A1(new_n2417), .A2(new_n2418), .B1(new_n2414), .B2(new_n2409), .Y(new_n2423));
  AND4x1_ASAP7_75t_L        g02167(.A(new_n2409), .B(new_n2418), .C(new_n2414), .D(new_n2417), .Y(new_n2424));
  OAI21xp33_ASAP7_75t_L     g02168(.A1(new_n2423), .A2(new_n2424), .B(new_n2422), .Y(new_n2425));
  AOI21xp33_ASAP7_75t_L     g02169(.A1(new_n2421), .A2(new_n2425), .B(new_n2375), .Y(new_n2426));
  INVx1_ASAP7_75t_L         g02170(.A(new_n2375), .Y(new_n2427));
  NOR3xp33_ASAP7_75t_L      g02171(.A(new_n2422), .B(new_n2423), .C(new_n2424), .Y(new_n2428));
  AOI21xp33_ASAP7_75t_L     g02172(.A1(new_n2420), .A2(new_n2419), .B(new_n2376), .Y(new_n2429));
  NOR3xp33_ASAP7_75t_L      g02173(.A(new_n2428), .B(new_n2427), .C(new_n2429), .Y(new_n2430));
  NOR2xp33_ASAP7_75t_L      g02174(.A(new_n2426), .B(new_n2430), .Y(new_n2431));
  NAND2xp33_ASAP7_75t_L     g02175(.A(new_n2368), .B(new_n2431), .Y(new_n2432));
  AOI21xp33_ASAP7_75t_L     g02176(.A1(new_n2300), .A2(new_n2292), .B(new_n2367), .Y(new_n2433));
  OAI21xp33_ASAP7_75t_L     g02177(.A1(new_n2429), .A2(new_n2428), .B(new_n2427), .Y(new_n2434));
  NAND3xp33_ASAP7_75t_L     g02178(.A(new_n2421), .B(new_n2425), .C(new_n2375), .Y(new_n2435));
  NAND2xp33_ASAP7_75t_L     g02179(.A(new_n2435), .B(new_n2434), .Y(new_n2436));
  NAND2xp33_ASAP7_75t_L     g02180(.A(new_n2433), .B(new_n2436), .Y(new_n2437));
  AOI22xp33_ASAP7_75t_L     g02181(.A1(new_n811), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n900), .Y(new_n2438));
  OAI221xp5_ASAP7_75t_L     g02182(.A1(new_n904), .A2(new_n869), .B1(new_n898), .B2(new_n950), .C(new_n2438), .Y(new_n2439));
  XNOR2x2_ASAP7_75t_L       g02183(.A(\a[14] ), .B(new_n2439), .Y(new_n2440));
  NAND3xp33_ASAP7_75t_L     g02184(.A(new_n2432), .B(new_n2437), .C(new_n2440), .Y(new_n2441));
  NOR2xp33_ASAP7_75t_L      g02185(.A(new_n2433), .B(new_n2436), .Y(new_n2442));
  AOI221xp5_ASAP7_75t_L     g02186(.A1(new_n2300), .A2(new_n2292), .B1(new_n2435), .B2(new_n2434), .C(new_n2367), .Y(new_n2443));
  XNOR2x2_ASAP7_75t_L       g02187(.A(new_n806), .B(new_n2439), .Y(new_n2444));
  OAI21xp33_ASAP7_75t_L     g02188(.A1(new_n2443), .A2(new_n2442), .B(new_n2444), .Y(new_n2445));
  NOR2xp33_ASAP7_75t_L      g02189(.A(new_n2301), .B(new_n2299), .Y(new_n2446));
  MAJIxp5_ASAP7_75t_L       g02190(.A(new_n2232), .B(new_n2305), .C(new_n2446), .Y(new_n2447));
  NAND3xp33_ASAP7_75t_L     g02191(.A(new_n2447), .B(new_n2445), .C(new_n2441), .Y(new_n2448));
  NAND2xp33_ASAP7_75t_L     g02192(.A(new_n2445), .B(new_n2441), .Y(new_n2449));
  NAND2xp33_ASAP7_75t_L     g02193(.A(new_n2307), .B(new_n2308), .Y(new_n2450));
  MAJIxp5_ASAP7_75t_L       g02194(.A(new_n2311), .B(new_n2304), .C(new_n2450), .Y(new_n2451));
  NAND2xp33_ASAP7_75t_L     g02195(.A(new_n2451), .B(new_n2449), .Y(new_n2452));
  AOI22xp33_ASAP7_75t_L     g02196(.A1(\b[16] ), .A2(new_n651), .B1(\b[18] ), .B2(new_n581), .Y(new_n2453));
  OAI221xp5_ASAP7_75t_L     g02197(.A1(new_n821), .A2(new_n1201), .B1(new_n577), .B2(new_n1320), .C(new_n2453), .Y(new_n2454));
  XNOR2x2_ASAP7_75t_L       g02198(.A(\a[11] ), .B(new_n2454), .Y(new_n2455));
  NAND3xp33_ASAP7_75t_L     g02199(.A(new_n2455), .B(new_n2452), .C(new_n2448), .Y(new_n2456));
  AO21x2_ASAP7_75t_L        g02200(.A1(new_n2448), .A2(new_n2452), .B(new_n2455), .Y(new_n2457));
  A2O1A1O1Ixp25_ASAP7_75t_L g02201(.A1(new_n2184), .A2(new_n2185), .B(new_n2225), .C(new_n2316), .D(new_n2326), .Y(new_n2458));
  NAND3xp33_ASAP7_75t_L     g02202(.A(new_n2458), .B(new_n2457), .C(new_n2456), .Y(new_n2459));
  AOI21xp33_ASAP7_75t_L     g02203(.A1(new_n2457), .A2(new_n2456), .B(new_n2458), .Y(new_n2460));
  INVx1_ASAP7_75t_L         g02204(.A(new_n2460), .Y(new_n2461));
  AOI22xp33_ASAP7_75t_L     g02205(.A1(new_n444), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n471), .Y(new_n2462));
  OAI221xp5_ASAP7_75t_L     g02206(.A1(new_n468), .A2(new_n1539), .B1(new_n469), .B2(new_n1662), .C(new_n2462), .Y(new_n2463));
  XNOR2x2_ASAP7_75t_L       g02207(.A(new_n435), .B(new_n2463), .Y(new_n2464));
  AOI21xp33_ASAP7_75t_L     g02208(.A1(new_n2461), .A2(new_n2459), .B(new_n2464), .Y(new_n2465));
  INVx1_ASAP7_75t_L         g02209(.A(new_n2459), .Y(new_n2466));
  XNOR2x2_ASAP7_75t_L       g02210(.A(\a[8] ), .B(new_n2463), .Y(new_n2467));
  NOR3xp33_ASAP7_75t_L      g02211(.A(new_n2466), .B(new_n2467), .C(new_n2460), .Y(new_n2468));
  NOR2xp33_ASAP7_75t_L      g02212(.A(new_n2465), .B(new_n2468), .Y(new_n2469));
  NOR3xp33_ASAP7_75t_L      g02213(.A(new_n2319), .B(new_n2330), .C(new_n2317), .Y(new_n2470));
  A2O1A1Ixp33_ASAP7_75t_L   g02214(.A1(new_n2366), .A2(new_n2336), .B(new_n2470), .C(new_n2469), .Y(new_n2471));
  OAI21xp33_ASAP7_75t_L     g02215(.A1(new_n2460), .A2(new_n2466), .B(new_n2467), .Y(new_n2472));
  NAND3xp33_ASAP7_75t_L     g02216(.A(new_n2461), .B(new_n2464), .C(new_n2459), .Y(new_n2473));
  NAND2xp33_ASAP7_75t_L     g02217(.A(new_n2473), .B(new_n2472), .Y(new_n2474));
  O2A1O1Ixp33_ASAP7_75t_L   g02218(.A1(new_n2324), .A2(new_n2331), .B(new_n2336), .C(new_n2470), .Y(new_n2475));
  NAND2xp33_ASAP7_75t_L     g02219(.A(new_n2475), .B(new_n2474), .Y(new_n2476));
  INVx1_ASAP7_75t_L         g02220(.A(new_n1935), .Y(new_n2477));
  AOI22xp33_ASAP7_75t_L     g02221(.A1(new_n344), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n370), .Y(new_n2478));
  OAI221xp5_ASAP7_75t_L     g02222(.A1(new_n429), .A2(new_n1909), .B1(new_n366), .B2(new_n2477), .C(new_n2478), .Y(new_n2479));
  XNOR2x2_ASAP7_75t_L       g02223(.A(\a[5] ), .B(new_n2479), .Y(new_n2480));
  NAND3xp33_ASAP7_75t_L     g02224(.A(new_n2480), .B(new_n2471), .C(new_n2476), .Y(new_n2481));
  INVx1_ASAP7_75t_L         g02225(.A(new_n2470), .Y(new_n2482));
  O2A1O1Ixp33_ASAP7_75t_L   g02226(.A1(new_n2334), .A2(new_n2332), .B(new_n2482), .C(new_n2474), .Y(new_n2483));
  A2O1A1Ixp33_ASAP7_75t_L   g02227(.A1(new_n2365), .A2(new_n2364), .B(new_n2334), .C(new_n2482), .Y(new_n2484));
  NOR2xp33_ASAP7_75t_L      g02228(.A(new_n2469), .B(new_n2484), .Y(new_n2485));
  XNOR2x2_ASAP7_75t_L       g02229(.A(new_n338), .B(new_n2479), .Y(new_n2486));
  OAI21xp33_ASAP7_75t_L     g02230(.A1(new_n2485), .A2(new_n2483), .B(new_n2486), .Y(new_n2487));
  NAND2xp33_ASAP7_75t_L     g02231(.A(new_n2337), .B(new_n2335), .Y(new_n2488));
  NOR2xp33_ASAP7_75t_L      g02232(.A(new_n2340), .B(new_n2488), .Y(new_n2489));
  A2O1A1O1Ixp25_ASAP7_75t_L g02233(.A1(new_n2211), .A2(new_n2204), .B(new_n2223), .C(new_n2345), .D(new_n2489), .Y(new_n2490));
  NAND3xp33_ASAP7_75t_L     g02234(.A(new_n2490), .B(new_n2487), .C(new_n2481), .Y(new_n2491));
  INVx1_ASAP7_75t_L         g02235(.A(new_n2344), .Y(new_n2492));
  NAND2xp33_ASAP7_75t_L     g02236(.A(new_n2487), .B(new_n2481), .Y(new_n2493));
  A2O1A1Ixp33_ASAP7_75t_L   g02237(.A1(new_n2492), .A2(new_n2345), .B(new_n2489), .C(new_n2493), .Y(new_n2494));
  INVx1_ASAP7_75t_L         g02238(.A(new_n2349), .Y(new_n2495));
  NOR2xp33_ASAP7_75t_L      g02239(.A(\b[26] ), .B(\b[27] ), .Y(new_n2496));
  INVx1_ASAP7_75t_L         g02240(.A(\b[27] ), .Y(new_n2497));
  NOR2xp33_ASAP7_75t_L      g02241(.A(new_n2348), .B(new_n2497), .Y(new_n2498));
  NOR2xp33_ASAP7_75t_L      g02242(.A(new_n2496), .B(new_n2498), .Y(new_n2499));
  INVx1_ASAP7_75t_L         g02243(.A(new_n2499), .Y(new_n2500));
  O2A1O1Ixp33_ASAP7_75t_L   g02244(.A1(new_n2353), .A2(new_n2352), .B(new_n2495), .C(new_n2500), .Y(new_n2501));
  O2A1O1Ixp33_ASAP7_75t_L   g02245(.A1(new_n1929), .A2(new_n2067), .B(new_n2070), .C(new_n2353), .Y(new_n2502));
  NOR3xp33_ASAP7_75t_L      g02246(.A(new_n2502), .B(new_n2499), .C(new_n2349), .Y(new_n2503));
  NOR2xp33_ASAP7_75t_L      g02247(.A(new_n2501), .B(new_n2503), .Y(new_n2504));
  INVx1_ASAP7_75t_L         g02248(.A(new_n2504), .Y(new_n2505));
  AOI22xp33_ASAP7_75t_L     g02249(.A1(\b[25] ), .A2(new_n282), .B1(\b[27] ), .B2(new_n303), .Y(new_n2506));
  OAI221xp5_ASAP7_75t_L     g02250(.A1(new_n291), .A2(new_n2348), .B1(new_n268), .B2(new_n2505), .C(new_n2506), .Y(new_n2507));
  XNOR2x2_ASAP7_75t_L       g02251(.A(new_n262), .B(new_n2507), .Y(new_n2508));
  AOI21xp33_ASAP7_75t_L     g02252(.A1(new_n2491), .A2(new_n2494), .B(new_n2508), .Y(new_n2509));
  NAND3xp33_ASAP7_75t_L     g02253(.A(new_n2491), .B(new_n2494), .C(new_n2508), .Y(new_n2510));
  INVx1_ASAP7_75t_L         g02254(.A(new_n2510), .Y(new_n2511));
  NOR2xp33_ASAP7_75t_L      g02255(.A(new_n2509), .B(new_n2511), .Y(new_n2512));
  INVx1_ASAP7_75t_L         g02256(.A(new_n2512), .Y(new_n2513));
  O2A1O1Ixp33_ASAP7_75t_L   g02257(.A1(new_n2222), .A2(new_n2362), .B(new_n2360), .C(new_n2513), .Y(new_n2514));
  A2O1A1O1Ixp25_ASAP7_75t_L g02258(.A1(new_n2216), .A2(new_n2219), .B(new_n2209), .C(new_n2361), .D(new_n2359), .Y(new_n2515));
  INVx1_ASAP7_75t_L         g02259(.A(new_n2515), .Y(new_n2516));
  NOR2xp33_ASAP7_75t_L      g02260(.A(new_n2516), .B(new_n2512), .Y(new_n2517));
  NOR2xp33_ASAP7_75t_L      g02261(.A(new_n2517), .B(new_n2514), .Y(\f[27] ));
  NOR3xp33_ASAP7_75t_L      g02262(.A(new_n2442), .B(new_n2443), .C(new_n2440), .Y(new_n2519));
  AOI211xp5_ASAP7_75t_L     g02263(.A1(new_n2406), .A2(new_n2400), .B(new_n2395), .C(new_n2396), .Y(new_n2520));
  AOI221xp5_ASAP7_75t_L     g02264(.A1(new_n2412), .A2(new_n2411), .B1(new_n2275), .B2(new_n2246), .C(new_n2410), .Y(new_n2521));
  AOI22xp33_ASAP7_75t_L     g02265(.A1(new_n1704), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1837), .Y(new_n2522));
  INVx1_ASAP7_75t_L         g02266(.A(new_n2522), .Y(new_n2523));
  AOI221xp5_ASAP7_75t_L     g02267(.A1(new_n1706), .A2(\b[6] ), .B1(new_n1695), .B2(new_n2084), .C(new_n2523), .Y(new_n2524));
  NAND2xp33_ASAP7_75t_L     g02268(.A(\a[23] ), .B(new_n2524), .Y(new_n2525));
  OAI21xp33_ASAP7_75t_L     g02269(.A1(new_n1827), .A2(new_n425), .B(new_n2522), .Y(new_n2526));
  A2O1A1Ixp33_ASAP7_75t_L   g02270(.A1(\b[6] ), .A2(new_n1706), .B(new_n2526), .C(new_n1689), .Y(new_n2527));
  NOR3xp33_ASAP7_75t_L      g02271(.A(new_n2261), .B(new_n2383), .C(new_n2378), .Y(new_n2528));
  INVx1_ASAP7_75t_L         g02272(.A(new_n2528), .Y(new_n2529));
  NOR2xp33_ASAP7_75t_L      g02273(.A(new_n298), .B(new_n2109), .Y(new_n2530));
  INVx1_ASAP7_75t_L         g02274(.A(new_n2530), .Y(new_n2531));
  NOR3xp33_ASAP7_75t_L      g02275(.A(new_n326), .B(new_n328), .C(new_n2257), .Y(new_n2532));
  INVx1_ASAP7_75t_L         g02276(.A(new_n2532), .Y(new_n2533));
  OAI22xp33_ASAP7_75t_L     g02277(.A1(new_n2269), .A2(new_n276), .B1(new_n324), .B2(new_n2107), .Y(new_n2534));
  INVx1_ASAP7_75t_L         g02278(.A(new_n2534), .Y(new_n2535));
  NAND4xp25_ASAP7_75t_L     g02279(.A(new_n2533), .B(new_n2535), .C(\a[26] ), .D(new_n2531), .Y(new_n2536));
  OAI31xp33_ASAP7_75t_L     g02280(.A1(new_n2532), .A2(new_n2534), .A3(new_n2530), .B(new_n2100), .Y(new_n2537));
  INVx1_ASAP7_75t_L         g02281(.A(\a[29] ), .Y(new_n2538));
  NOR2xp33_ASAP7_75t_L      g02282(.A(new_n2538), .B(new_n2383), .Y(new_n2539));
  AND2x2_ASAP7_75t_L        g02283(.A(new_n2380), .B(new_n2381), .Y(new_n2540));
  INVx1_ASAP7_75t_L         g02284(.A(\a[28] ), .Y(new_n2541));
  NAND2xp33_ASAP7_75t_L     g02285(.A(\a[29] ), .B(new_n2541), .Y(new_n2542));
  NAND2xp33_ASAP7_75t_L     g02286(.A(\a[28] ), .B(new_n2538), .Y(new_n2543));
  AOI21xp33_ASAP7_75t_L     g02287(.A1(new_n2543), .A2(new_n2542), .B(new_n2540), .Y(new_n2544));
  NAND3xp33_ASAP7_75t_L     g02288(.A(new_n2382), .B(new_n2542), .C(new_n2543), .Y(new_n2545));
  XNOR2x2_ASAP7_75t_L       g02289(.A(\a[28] ), .B(\a[27] ), .Y(new_n2546));
  OR2x4_ASAP7_75t_L         g02290(.A(new_n2546), .B(new_n2382), .Y(new_n2547));
  OAI22xp33_ASAP7_75t_L     g02291(.A1(new_n2547), .A2(new_n258), .B1(new_n261), .B2(new_n2545), .Y(new_n2548));
  A2O1A1Ixp33_ASAP7_75t_L   g02292(.A1(new_n269), .A2(new_n2544), .B(new_n2548), .C(new_n2539), .Y(new_n2549));
  NAND2xp33_ASAP7_75t_L     g02293(.A(new_n269), .B(new_n2544), .Y(new_n2550));
  NAND2xp33_ASAP7_75t_L     g02294(.A(new_n2543), .B(new_n2542), .Y(new_n2551));
  NOR2xp33_ASAP7_75t_L      g02295(.A(new_n2551), .B(new_n2540), .Y(new_n2552));
  NOR2xp33_ASAP7_75t_L      g02296(.A(new_n2546), .B(new_n2382), .Y(new_n2553));
  AOI22xp33_ASAP7_75t_L     g02297(.A1(\b[0] ), .A2(new_n2553), .B1(\b[1] ), .B2(new_n2552), .Y(new_n2554));
  OAI211xp5_ASAP7_75t_L     g02298(.A1(new_n2538), .A2(new_n2383), .B(new_n2554), .C(new_n2550), .Y(new_n2555));
  AND2x2_ASAP7_75t_L        g02299(.A(new_n2555), .B(new_n2549), .Y(new_n2556));
  NAND3xp33_ASAP7_75t_L     g02300(.A(new_n2556), .B(new_n2537), .C(new_n2536), .Y(new_n2557));
  NAND2xp33_ASAP7_75t_L     g02301(.A(new_n2537), .B(new_n2536), .Y(new_n2558));
  NAND2xp33_ASAP7_75t_L     g02302(.A(new_n2555), .B(new_n2549), .Y(new_n2559));
  NAND2xp33_ASAP7_75t_L     g02303(.A(new_n2559), .B(new_n2558), .Y(new_n2560));
  AOI22xp33_ASAP7_75t_L     g02304(.A1(new_n2557), .A2(new_n2560), .B1(new_n2529), .B2(new_n2404), .Y(new_n2561));
  AND4x1_ASAP7_75t_L        g02305(.A(new_n2536), .B(new_n2555), .C(new_n2537), .D(new_n2549), .Y(new_n2562));
  AOI21xp33_ASAP7_75t_L     g02306(.A1(new_n2537), .A2(new_n2536), .B(new_n2556), .Y(new_n2563));
  NOR4xp25_ASAP7_75t_L      g02307(.A(new_n2395), .B(new_n2563), .C(new_n2562), .D(new_n2528), .Y(new_n2564));
  AOI211xp5_ASAP7_75t_L     g02308(.A1(new_n2527), .A2(new_n2525), .B(new_n2564), .C(new_n2561), .Y(new_n2565));
  INVx1_ASAP7_75t_L         g02309(.A(new_n2525), .Y(new_n2566));
  INVx1_ASAP7_75t_L         g02310(.A(new_n2527), .Y(new_n2567));
  OAI22xp33_ASAP7_75t_L     g02311(.A1(new_n2395), .A2(new_n2528), .B1(new_n2562), .B2(new_n2563), .Y(new_n2568));
  NAND4xp25_ASAP7_75t_L     g02312(.A(new_n2404), .B(new_n2529), .C(new_n2560), .D(new_n2557), .Y(new_n2569));
  AOI211xp5_ASAP7_75t_L     g02313(.A1(new_n2568), .A2(new_n2569), .B(new_n2567), .C(new_n2566), .Y(new_n2570));
  NOR2xp33_ASAP7_75t_L      g02314(.A(new_n2565), .B(new_n2570), .Y(new_n2571));
  OAI21xp33_ASAP7_75t_L     g02315(.A1(new_n2520), .A2(new_n2521), .B(new_n2571), .Y(new_n2572));
  INVx1_ASAP7_75t_L         g02316(.A(new_n2520), .Y(new_n2573));
  OAI221xp5_ASAP7_75t_L     g02317(.A1(new_n2403), .A2(new_n2407), .B1(new_n2377), .B2(new_n2280), .C(new_n2265), .Y(new_n2574));
  OAI211xp5_ASAP7_75t_L     g02318(.A1(new_n2565), .A2(new_n2570), .B(new_n2574), .C(new_n2573), .Y(new_n2575));
  NAND2xp33_ASAP7_75t_L     g02319(.A(\b[9] ), .B(new_n1362), .Y(new_n2576));
  NAND2xp33_ASAP7_75t_L     g02320(.A(new_n1365), .B(new_n2143), .Y(new_n2577));
  AOI22xp33_ASAP7_75t_L     g02321(.A1(new_n1360), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1581), .Y(new_n2578));
  NAND4xp25_ASAP7_75t_L     g02322(.A(new_n2577), .B(\a[20] ), .C(new_n2576), .D(new_n2578), .Y(new_n2579));
  OAI211xp5_ASAP7_75t_L     g02323(.A1(new_n1359), .A2(new_n624), .B(new_n2576), .C(new_n2578), .Y(new_n2580));
  NAND2xp33_ASAP7_75t_L     g02324(.A(new_n1356), .B(new_n2580), .Y(new_n2581));
  AND2x2_ASAP7_75t_L        g02325(.A(new_n2579), .B(new_n2581), .Y(new_n2582));
  NAND3xp33_ASAP7_75t_L     g02326(.A(new_n2572), .B(new_n2582), .C(new_n2575), .Y(new_n2583));
  AOI211xp5_ASAP7_75t_L     g02327(.A1(new_n2574), .A2(new_n2573), .B(new_n2565), .C(new_n2570), .Y(new_n2584));
  OAI211xp5_ASAP7_75t_L     g02328(.A1(new_n2567), .A2(new_n2566), .B(new_n2569), .C(new_n2568), .Y(new_n2585));
  OAI211xp5_ASAP7_75t_L     g02329(.A1(new_n2564), .A2(new_n2561), .B(new_n2527), .C(new_n2525), .Y(new_n2586));
  AOI211xp5_ASAP7_75t_L     g02330(.A1(new_n2586), .A2(new_n2585), .B(new_n2520), .C(new_n2521), .Y(new_n2587));
  NAND2xp33_ASAP7_75t_L     g02331(.A(new_n2579), .B(new_n2581), .Y(new_n2588));
  OAI21xp33_ASAP7_75t_L     g02332(.A1(new_n2584), .A2(new_n2587), .B(new_n2588), .Y(new_n2589));
  NAND2xp33_ASAP7_75t_L     g02333(.A(new_n2589), .B(new_n2583), .Y(new_n2590));
  OAI21xp33_ASAP7_75t_L     g02334(.A1(new_n2424), .A2(new_n2422), .B(new_n2419), .Y(new_n2591));
  NOR2xp33_ASAP7_75t_L      g02335(.A(new_n2591), .B(new_n2590), .Y(new_n2592));
  A2O1A1O1Ixp25_ASAP7_75t_L g02336(.A1(new_n2289), .A2(new_n2288), .B(new_n2285), .C(new_n2420), .D(new_n2423), .Y(new_n2593));
  AOI21xp33_ASAP7_75t_L     g02337(.A1(new_n2589), .A2(new_n2583), .B(new_n2593), .Y(new_n2594));
  AOI22xp33_ASAP7_75t_L     g02338(.A1(new_n1076), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1253), .Y(new_n2595));
  OAI221xp5_ASAP7_75t_L     g02339(.A1(new_n1154), .A2(new_n760), .B1(new_n1156), .B2(new_n790), .C(new_n2595), .Y(new_n2596));
  XNOR2x2_ASAP7_75t_L       g02340(.A(\a[17] ), .B(new_n2596), .Y(new_n2597));
  INVx1_ASAP7_75t_L         g02341(.A(new_n2597), .Y(new_n2598));
  NOR3xp33_ASAP7_75t_L      g02342(.A(new_n2598), .B(new_n2592), .C(new_n2594), .Y(new_n2599));
  OA21x2_ASAP7_75t_L        g02343(.A1(new_n2594), .A2(new_n2592), .B(new_n2598), .Y(new_n2600));
  A2O1A1O1Ixp25_ASAP7_75t_L g02344(.A1(new_n2292), .A2(new_n2300), .B(new_n2367), .C(new_n2434), .D(new_n2430), .Y(new_n2601));
  OA21x2_ASAP7_75t_L        g02345(.A1(new_n2599), .A2(new_n2600), .B(new_n2601), .Y(new_n2602));
  NOR3xp33_ASAP7_75t_L      g02346(.A(new_n2600), .B(new_n2601), .C(new_n2599), .Y(new_n2603));
  AOI22xp33_ASAP7_75t_L     g02347(.A1(new_n811), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n900), .Y(new_n2604));
  OAI221xp5_ASAP7_75t_L     g02348(.A1(new_n904), .A2(new_n942), .B1(new_n898), .B2(new_n1035), .C(new_n2604), .Y(new_n2605));
  XNOR2x2_ASAP7_75t_L       g02349(.A(new_n806), .B(new_n2605), .Y(new_n2606));
  OAI21xp33_ASAP7_75t_L     g02350(.A1(new_n2603), .A2(new_n2602), .B(new_n2606), .Y(new_n2607));
  OAI21xp33_ASAP7_75t_L     g02351(.A1(new_n2599), .A2(new_n2600), .B(new_n2601), .Y(new_n2608));
  OR3x1_ASAP7_75t_L         g02352(.A(new_n2600), .B(new_n2601), .C(new_n2599), .Y(new_n2609));
  XNOR2x2_ASAP7_75t_L       g02353(.A(\a[14] ), .B(new_n2605), .Y(new_n2610));
  NAND3xp33_ASAP7_75t_L     g02354(.A(new_n2609), .B(new_n2608), .C(new_n2610), .Y(new_n2611));
  AOI221xp5_ASAP7_75t_L     g02355(.A1(new_n2449), .A2(new_n2451), .B1(new_n2607), .B2(new_n2611), .C(new_n2519), .Y(new_n2612));
  NOR2xp33_ASAP7_75t_L      g02356(.A(new_n2443), .B(new_n2442), .Y(new_n2613));
  MAJIxp5_ASAP7_75t_L       g02357(.A(new_n2451), .B(new_n2613), .C(new_n2444), .Y(new_n2614));
  NAND2xp33_ASAP7_75t_L     g02358(.A(new_n2607), .B(new_n2611), .Y(new_n2615));
  NOR2xp33_ASAP7_75t_L      g02359(.A(new_n2614), .B(new_n2615), .Y(new_n2616));
  AOI22xp33_ASAP7_75t_L     g02360(.A1(\b[17] ), .A2(new_n651), .B1(\b[19] ), .B2(new_n581), .Y(new_n2617));
  OAI221xp5_ASAP7_75t_L     g02361(.A1(new_n821), .A2(new_n1313), .B1(new_n577), .B2(new_n1438), .C(new_n2617), .Y(new_n2618));
  XNOR2x2_ASAP7_75t_L       g02362(.A(new_n574), .B(new_n2618), .Y(new_n2619));
  NOR3xp33_ASAP7_75t_L      g02363(.A(new_n2616), .B(new_n2619), .C(new_n2612), .Y(new_n2620));
  NAND2xp33_ASAP7_75t_L     g02364(.A(new_n2614), .B(new_n2615), .Y(new_n2621));
  INVx1_ASAP7_75t_L         g02365(.A(new_n2519), .Y(new_n2622));
  A2O1A1Ixp33_ASAP7_75t_L   g02366(.A1(new_n2445), .A2(new_n2441), .B(new_n2447), .C(new_n2622), .Y(new_n2623));
  AOI21xp33_ASAP7_75t_L     g02367(.A1(new_n2609), .A2(new_n2608), .B(new_n2610), .Y(new_n2624));
  NOR3xp33_ASAP7_75t_L      g02368(.A(new_n2602), .B(new_n2603), .C(new_n2606), .Y(new_n2625));
  NOR2xp33_ASAP7_75t_L      g02369(.A(new_n2625), .B(new_n2624), .Y(new_n2626));
  NAND2xp33_ASAP7_75t_L     g02370(.A(new_n2626), .B(new_n2623), .Y(new_n2627));
  INVx1_ASAP7_75t_L         g02371(.A(new_n2619), .Y(new_n2628));
  AOI21xp33_ASAP7_75t_L     g02372(.A1(new_n2627), .A2(new_n2621), .B(new_n2628), .Y(new_n2629));
  NAND2xp33_ASAP7_75t_L     g02373(.A(new_n2452), .B(new_n2448), .Y(new_n2630));
  MAJIxp5_ASAP7_75t_L       g02374(.A(new_n2458), .B(new_n2630), .C(new_n2455), .Y(new_n2631));
  NOR3xp33_ASAP7_75t_L      g02375(.A(new_n2631), .B(new_n2629), .C(new_n2620), .Y(new_n2632));
  OAI21xp33_ASAP7_75t_L     g02376(.A1(new_n2620), .A2(new_n2629), .B(new_n2631), .Y(new_n2633));
  INVx1_ASAP7_75t_L         g02377(.A(new_n2633), .Y(new_n2634));
  AOI22xp33_ASAP7_75t_L     g02378(.A1(new_n444), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n471), .Y(new_n2635));
  OAI221xp5_ASAP7_75t_L     g02379(.A1(new_n468), .A2(new_n1655), .B1(new_n469), .B2(new_n1780), .C(new_n2635), .Y(new_n2636));
  XNOR2x2_ASAP7_75t_L       g02380(.A(\a[8] ), .B(new_n2636), .Y(new_n2637));
  OAI21xp33_ASAP7_75t_L     g02381(.A1(new_n2632), .A2(new_n2634), .B(new_n2637), .Y(new_n2638));
  INVx1_ASAP7_75t_L         g02382(.A(new_n2632), .Y(new_n2639));
  INVx1_ASAP7_75t_L         g02383(.A(new_n2637), .Y(new_n2640));
  NAND3xp33_ASAP7_75t_L     g02384(.A(new_n2639), .B(new_n2633), .C(new_n2640), .Y(new_n2641));
  A2O1A1Ixp33_ASAP7_75t_L   g02385(.A1(new_n2337), .A2(new_n2482), .B(new_n2465), .C(new_n2473), .Y(new_n2642));
  NAND3xp33_ASAP7_75t_L     g02386(.A(new_n2642), .B(new_n2641), .C(new_n2638), .Y(new_n2643));
  AOI21xp33_ASAP7_75t_L     g02387(.A1(new_n2639), .A2(new_n2633), .B(new_n2640), .Y(new_n2644));
  NOR3xp33_ASAP7_75t_L      g02388(.A(new_n2634), .B(new_n2637), .C(new_n2632), .Y(new_n2645));
  A2O1A1O1Ixp25_ASAP7_75t_L g02389(.A1(new_n2336), .A2(new_n2366), .B(new_n2470), .C(new_n2472), .D(new_n2468), .Y(new_n2646));
  OAI21xp33_ASAP7_75t_L     g02390(.A1(new_n2645), .A2(new_n2644), .B(new_n2646), .Y(new_n2647));
  NOR2xp33_ASAP7_75t_L      g02391(.A(new_n2071), .B(new_n2074), .Y(new_n2648));
  OAI22xp33_ASAP7_75t_L     g02392(.A1(new_n407), .A2(new_n1909), .B1(new_n2067), .B2(new_n343), .Y(new_n2649));
  AOI221xp5_ASAP7_75t_L     g02393(.A1(\b[24] ), .A2(new_n347), .B1(new_n341), .B2(new_n2648), .C(new_n2649), .Y(new_n2650));
  XNOR2x2_ASAP7_75t_L       g02394(.A(new_n338), .B(new_n2650), .Y(new_n2651));
  NAND3xp33_ASAP7_75t_L     g02395(.A(new_n2643), .B(new_n2651), .C(new_n2647), .Y(new_n2652));
  NOR3xp33_ASAP7_75t_L      g02396(.A(new_n2646), .B(new_n2644), .C(new_n2645), .Y(new_n2653));
  AOI21xp33_ASAP7_75t_L     g02397(.A1(new_n2641), .A2(new_n2638), .B(new_n2642), .Y(new_n2654));
  XNOR2x2_ASAP7_75t_L       g02398(.A(\a[5] ), .B(new_n2650), .Y(new_n2655));
  OAI21xp33_ASAP7_75t_L     g02399(.A1(new_n2653), .A2(new_n2654), .B(new_n2655), .Y(new_n2656));
  NAND2xp33_ASAP7_75t_L     g02400(.A(new_n2652), .B(new_n2656), .Y(new_n2657));
  NOR3xp33_ASAP7_75t_L      g02401(.A(new_n2485), .B(new_n2480), .C(new_n2483), .Y(new_n2658));
  INVx1_ASAP7_75t_L         g02402(.A(new_n2658), .Y(new_n2659));
  A2O1A1Ixp33_ASAP7_75t_L   g02403(.A1(new_n2487), .A2(new_n2481), .B(new_n2490), .C(new_n2659), .Y(new_n2660));
  NOR2xp33_ASAP7_75t_L      g02404(.A(new_n2657), .B(new_n2660), .Y(new_n2661));
  MAJIxp5_ASAP7_75t_L       g02405(.A(new_n2344), .B(new_n2488), .C(new_n2340), .Y(new_n2662));
  A2O1A1Ixp33_ASAP7_75t_L   g02406(.A1(new_n2662), .A2(new_n2493), .B(new_n2658), .C(new_n2657), .Y(new_n2663));
  INVx1_ASAP7_75t_L         g02407(.A(new_n2663), .Y(new_n2664));
  NOR2xp33_ASAP7_75t_L      g02408(.A(\b[27] ), .B(\b[28] ), .Y(new_n2665));
  INVx1_ASAP7_75t_L         g02409(.A(\b[28] ), .Y(new_n2666));
  NOR2xp33_ASAP7_75t_L      g02410(.A(new_n2497), .B(new_n2666), .Y(new_n2667));
  NOR2xp33_ASAP7_75t_L      g02411(.A(new_n2665), .B(new_n2667), .Y(new_n2668));
  A2O1A1Ixp33_ASAP7_75t_L   g02412(.A1(\b[27] ), .A2(\b[26] ), .B(new_n2501), .C(new_n2668), .Y(new_n2669));
  O2A1O1Ixp33_ASAP7_75t_L   g02413(.A1(new_n2349), .A2(new_n2502), .B(new_n2499), .C(new_n2498), .Y(new_n2670));
  OAI21xp33_ASAP7_75t_L     g02414(.A1(new_n2665), .A2(new_n2667), .B(new_n2670), .Y(new_n2671));
  NAND2xp33_ASAP7_75t_L     g02415(.A(new_n2669), .B(new_n2671), .Y(new_n2672));
  AOI22xp33_ASAP7_75t_L     g02416(.A1(\b[26] ), .A2(new_n282), .B1(\b[28] ), .B2(new_n303), .Y(new_n2673));
  OAI221xp5_ASAP7_75t_L     g02417(.A1(new_n291), .A2(new_n2497), .B1(new_n268), .B2(new_n2672), .C(new_n2673), .Y(new_n2674));
  XNOR2x2_ASAP7_75t_L       g02418(.A(\a[2] ), .B(new_n2674), .Y(new_n2675));
  OAI21xp33_ASAP7_75t_L     g02419(.A1(new_n2661), .A2(new_n2664), .B(new_n2675), .Y(new_n2676));
  NOR3xp33_ASAP7_75t_L      g02420(.A(new_n2664), .B(new_n2661), .C(new_n2675), .Y(new_n2677));
  INVx1_ASAP7_75t_L         g02421(.A(new_n2677), .Y(new_n2678));
  NAND2xp33_ASAP7_75t_L     g02422(.A(new_n2676), .B(new_n2678), .Y(new_n2679));
  O2A1O1Ixp33_ASAP7_75t_L   g02423(.A1(new_n2515), .A2(new_n2509), .B(new_n2510), .C(new_n2679), .Y(new_n2680));
  OAI21xp33_ASAP7_75t_L     g02424(.A1(new_n2509), .A2(new_n2515), .B(new_n2510), .Y(new_n2681));
  AOI21xp33_ASAP7_75t_L     g02425(.A1(new_n2678), .A2(new_n2676), .B(new_n2681), .Y(new_n2682));
  NOR2xp33_ASAP7_75t_L      g02426(.A(new_n2682), .B(new_n2680), .Y(\f[28] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02427(.A1(new_n2516), .A2(new_n2512), .B(new_n2511), .C(new_n2676), .D(new_n2677), .Y(new_n2684));
  INVx1_ASAP7_75t_L         g02428(.A(new_n2498), .Y(new_n2685));
  A2O1A1Ixp33_ASAP7_75t_L   g02429(.A1(new_n2351), .A2(new_n2495), .B(new_n2496), .C(new_n2685), .Y(new_n2686));
  NOR2xp33_ASAP7_75t_L      g02430(.A(\b[28] ), .B(\b[29] ), .Y(new_n2687));
  INVx1_ASAP7_75t_L         g02431(.A(\b[29] ), .Y(new_n2688));
  NOR2xp33_ASAP7_75t_L      g02432(.A(new_n2666), .B(new_n2688), .Y(new_n2689));
  NOR2xp33_ASAP7_75t_L      g02433(.A(new_n2687), .B(new_n2689), .Y(new_n2690));
  A2O1A1Ixp33_ASAP7_75t_L   g02434(.A1(new_n2686), .A2(new_n2668), .B(new_n2667), .C(new_n2690), .Y(new_n2691));
  O2A1O1Ixp33_ASAP7_75t_L   g02435(.A1(new_n2498), .A2(new_n2501), .B(new_n2668), .C(new_n2667), .Y(new_n2692));
  INVx1_ASAP7_75t_L         g02436(.A(new_n2690), .Y(new_n2693));
  NAND2xp33_ASAP7_75t_L     g02437(.A(new_n2693), .B(new_n2692), .Y(new_n2694));
  NAND2xp33_ASAP7_75t_L     g02438(.A(new_n2694), .B(new_n2691), .Y(new_n2695));
  AOI22xp33_ASAP7_75t_L     g02439(.A1(\b[27] ), .A2(new_n282), .B1(\b[29] ), .B2(new_n303), .Y(new_n2696));
  OAI221xp5_ASAP7_75t_L     g02440(.A1(new_n291), .A2(new_n2666), .B1(new_n268), .B2(new_n2695), .C(new_n2696), .Y(new_n2697));
  XNOR2x2_ASAP7_75t_L       g02441(.A(\a[2] ), .B(new_n2697), .Y(new_n2698));
  INVx1_ASAP7_75t_L         g02442(.A(new_n2657), .Y(new_n2699));
  A2O1A1O1Ixp25_ASAP7_75t_L g02443(.A1(new_n2345), .A2(new_n2492), .B(new_n2489), .C(new_n2493), .D(new_n2658), .Y(new_n2700));
  NOR3xp33_ASAP7_75t_L      g02444(.A(new_n2654), .B(new_n2651), .C(new_n2653), .Y(new_n2701));
  INVx1_ASAP7_75t_L         g02445(.A(new_n2701), .Y(new_n2702));
  AOI22xp33_ASAP7_75t_L     g02446(.A1(new_n344), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n370), .Y(new_n2703));
  OAI221xp5_ASAP7_75t_L     g02447(.A1(new_n429), .A2(new_n2067), .B1(new_n366), .B2(new_n2355), .C(new_n2703), .Y(new_n2704));
  XNOR2x2_ASAP7_75t_L       g02448(.A(\a[5] ), .B(new_n2704), .Y(new_n2705));
  OAI21xp33_ASAP7_75t_L     g02449(.A1(new_n2644), .A2(new_n2646), .B(new_n2641), .Y(new_n2706));
  AOI22xp33_ASAP7_75t_L     g02450(.A1(new_n444), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n471), .Y(new_n2707));
  OAI221xp5_ASAP7_75t_L     g02451(.A1(new_n468), .A2(new_n1774), .B1(new_n469), .B2(new_n1915), .C(new_n2707), .Y(new_n2708));
  XNOR2x2_ASAP7_75t_L       g02452(.A(\a[8] ), .B(new_n2708), .Y(new_n2709));
  INVx1_ASAP7_75t_L         g02453(.A(new_n2709), .Y(new_n2710));
  NOR3xp33_ASAP7_75t_L      g02454(.A(new_n2628), .B(new_n2616), .C(new_n2612), .Y(new_n2711));
  O2A1O1Ixp33_ASAP7_75t_L   g02455(.A1(new_n2620), .A2(new_n2629), .B(new_n2631), .C(new_n2711), .Y(new_n2712));
  NAND3xp33_ASAP7_75t_L     g02456(.A(new_n2572), .B(new_n2575), .C(new_n2588), .Y(new_n2713));
  A2O1A1Ixp33_ASAP7_75t_L   g02457(.A1(new_n2589), .A2(new_n2583), .B(new_n2593), .C(new_n2713), .Y(new_n2714));
  AOI22xp33_ASAP7_75t_L     g02458(.A1(new_n1360), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1581), .Y(new_n2715));
  OAI221xp5_ASAP7_75t_L     g02459(.A1(new_n1373), .A2(new_n617), .B1(new_n1359), .B2(new_n685), .C(new_n2715), .Y(new_n2716));
  XNOR2x2_ASAP7_75t_L       g02460(.A(new_n1356), .B(new_n2716), .Y(new_n2717));
  A2O1A1Ixp33_ASAP7_75t_L   g02461(.A1(new_n2574), .A2(new_n2573), .B(new_n2570), .C(new_n2585), .Y(new_n2718));
  AOI22xp33_ASAP7_75t_L     g02462(.A1(new_n1704), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1837), .Y(new_n2719));
  OAI221xp5_ASAP7_75t_L     g02463(.A1(new_n1699), .A2(new_n420), .B1(new_n1827), .B2(new_n494), .C(new_n2719), .Y(new_n2720));
  XNOR2x2_ASAP7_75t_L       g02464(.A(\a[23] ), .B(new_n2720), .Y(new_n2721));
  NOR2xp33_ASAP7_75t_L      g02465(.A(new_n2378), .B(new_n2261), .Y(new_n2722));
  NAND2xp33_ASAP7_75t_L     g02466(.A(new_n2394), .B(new_n2392), .Y(new_n2723));
  MAJIxp5_ASAP7_75t_L       g02467(.A(new_n2723), .B(new_n2384), .C(new_n2722), .Y(new_n2724));
  NAND2xp33_ASAP7_75t_L     g02468(.A(new_n2556), .B(new_n2558), .Y(new_n2725));
  A2O1A1Ixp33_ASAP7_75t_L   g02469(.A1(new_n2557), .A2(new_n2560), .B(new_n2724), .C(new_n2725), .Y(new_n2726));
  OAI22xp33_ASAP7_75t_L     g02470(.A1(new_n2269), .A2(new_n298), .B1(new_n354), .B2(new_n2107), .Y(new_n2727));
  AOI221xp5_ASAP7_75t_L     g02471(.A1(new_n2115), .A2(\b[4] ), .B1(new_n2106), .B2(new_n359), .C(new_n2727), .Y(new_n2728));
  NAND2xp33_ASAP7_75t_L     g02472(.A(\a[26] ), .B(new_n2728), .Y(new_n2729));
  OR2x4_ASAP7_75t_L         g02473(.A(\a[26] ), .B(new_n2728), .Y(new_n2730));
  NAND2xp33_ASAP7_75t_L     g02474(.A(new_n2550), .B(new_n2554), .Y(new_n2731));
  NOR2xp33_ASAP7_75t_L      g02475(.A(new_n261), .B(new_n2547), .Y(new_n2732));
  INVx1_ASAP7_75t_L         g02476(.A(new_n2732), .Y(new_n2733));
  NAND2xp33_ASAP7_75t_L     g02477(.A(new_n2551), .B(new_n2382), .Y(new_n2734));
  NOR2xp33_ASAP7_75t_L      g02478(.A(new_n280), .B(new_n2734), .Y(new_n2735));
  AND3x1_ASAP7_75t_L        g02479(.A(new_n2540), .B(new_n2546), .C(new_n2551), .Y(new_n2736));
  AOI221xp5_ASAP7_75t_L     g02480(.A1(new_n2552), .A2(\b[2] ), .B1(new_n2736), .B2(\b[0] ), .C(new_n2735), .Y(new_n2737));
  NAND2xp33_ASAP7_75t_L     g02481(.A(new_n2733), .B(new_n2737), .Y(new_n2738));
  O2A1O1Ixp33_ASAP7_75t_L   g02482(.A1(new_n2384), .A2(new_n2731), .B(\a[29] ), .C(new_n2738), .Y(new_n2739));
  A2O1A1Ixp33_ASAP7_75t_L   g02483(.A1(\b[0] ), .A2(new_n2382), .B(new_n2731), .C(\a[29] ), .Y(new_n2740));
  O2A1O1Ixp33_ASAP7_75t_L   g02484(.A1(new_n2547), .A2(new_n261), .B(new_n2737), .C(new_n2740), .Y(new_n2741));
  OAI211xp5_ASAP7_75t_L     g02485(.A1(new_n2739), .A2(new_n2741), .B(new_n2730), .C(new_n2729), .Y(new_n2742));
  AND2x2_ASAP7_75t_L        g02486(.A(\a[26] ), .B(new_n2728), .Y(new_n2743));
  NOR2xp33_ASAP7_75t_L      g02487(.A(\a[26] ), .B(new_n2728), .Y(new_n2744));
  AOI21xp33_ASAP7_75t_L     g02488(.A1(new_n2544), .A2(new_n269), .B(new_n2548), .Y(new_n2745));
  NAND2xp33_ASAP7_75t_L     g02489(.A(\b[2] ), .B(new_n2552), .Y(new_n2746));
  NAND3xp33_ASAP7_75t_L     g02490(.A(new_n2540), .B(new_n2551), .C(new_n2546), .Y(new_n2747));
  OAI221xp5_ASAP7_75t_L     g02491(.A1(new_n258), .A2(new_n2747), .B1(new_n280), .B2(new_n2734), .C(new_n2746), .Y(new_n2748));
  NOR2xp33_ASAP7_75t_L      g02492(.A(new_n2732), .B(new_n2748), .Y(new_n2749));
  A2O1A1Ixp33_ASAP7_75t_L   g02493(.A1(new_n2383), .A2(new_n2745), .B(new_n2538), .C(new_n2749), .Y(new_n2750));
  O2A1O1Ixp33_ASAP7_75t_L   g02494(.A1(new_n258), .A2(new_n2540), .B(new_n2745), .C(new_n2538), .Y(new_n2751));
  A2O1A1Ixp33_ASAP7_75t_L   g02495(.A1(\b[1] ), .A2(new_n2553), .B(new_n2748), .C(new_n2751), .Y(new_n2752));
  OAI211xp5_ASAP7_75t_L     g02496(.A1(new_n2744), .A2(new_n2743), .B(new_n2752), .C(new_n2750), .Y(new_n2753));
  AOI21xp33_ASAP7_75t_L     g02497(.A1(new_n2753), .A2(new_n2742), .B(new_n2726), .Y(new_n2754));
  NAND2xp33_ASAP7_75t_L     g02498(.A(new_n2753), .B(new_n2742), .Y(new_n2755));
  A2O1A1O1Ixp25_ASAP7_75t_L g02499(.A1(new_n2537), .A2(new_n2536), .B(new_n2559), .C(new_n2568), .D(new_n2755), .Y(new_n2756));
  OAI21xp33_ASAP7_75t_L     g02500(.A1(new_n2754), .A2(new_n2756), .B(new_n2721), .Y(new_n2757));
  INVx1_ASAP7_75t_L         g02501(.A(new_n2721), .Y(new_n2758));
  NAND3xp33_ASAP7_75t_L     g02502(.A(new_n2755), .B(new_n2725), .C(new_n2568), .Y(new_n2759));
  AOI211xp5_ASAP7_75t_L     g02503(.A1(new_n2752), .A2(new_n2750), .B(new_n2743), .C(new_n2744), .Y(new_n2760));
  AOI211xp5_ASAP7_75t_L     g02504(.A1(new_n2730), .A2(new_n2729), .B(new_n2739), .C(new_n2741), .Y(new_n2761));
  NOR2xp33_ASAP7_75t_L      g02505(.A(new_n2760), .B(new_n2761), .Y(new_n2762));
  A2O1A1Ixp33_ASAP7_75t_L   g02506(.A1(new_n2556), .A2(new_n2558), .B(new_n2561), .C(new_n2762), .Y(new_n2763));
  NAND3xp33_ASAP7_75t_L     g02507(.A(new_n2758), .B(new_n2763), .C(new_n2759), .Y(new_n2764));
  NAND3xp33_ASAP7_75t_L     g02508(.A(new_n2718), .B(new_n2764), .C(new_n2757), .Y(new_n2765));
  AOI21xp33_ASAP7_75t_L     g02509(.A1(new_n2246), .A2(new_n2275), .B(new_n2410), .Y(new_n2766));
  A2O1A1O1Ixp25_ASAP7_75t_L g02510(.A1(new_n2413), .A2(new_n2766), .B(new_n2520), .C(new_n2586), .D(new_n2565), .Y(new_n2767));
  AOI21xp33_ASAP7_75t_L     g02511(.A1(new_n2763), .A2(new_n2759), .B(new_n2758), .Y(new_n2768));
  NOR3xp33_ASAP7_75t_L      g02512(.A(new_n2756), .B(new_n2754), .C(new_n2721), .Y(new_n2769));
  OAI21xp33_ASAP7_75t_L     g02513(.A1(new_n2768), .A2(new_n2769), .B(new_n2767), .Y(new_n2770));
  AO21x2_ASAP7_75t_L        g02514(.A1(new_n2765), .A2(new_n2770), .B(new_n2717), .Y(new_n2771));
  NAND3xp33_ASAP7_75t_L     g02515(.A(new_n2770), .B(new_n2765), .C(new_n2717), .Y(new_n2772));
  NAND3xp33_ASAP7_75t_L     g02516(.A(new_n2714), .B(new_n2771), .C(new_n2772), .Y(new_n2773));
  AO21x2_ASAP7_75t_L        g02517(.A1(new_n2772), .A2(new_n2771), .B(new_n2714), .Y(new_n2774));
  AOI22xp33_ASAP7_75t_L     g02518(.A1(new_n1076), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1253), .Y(new_n2775));
  OAI221xp5_ASAP7_75t_L     g02519(.A1(new_n1154), .A2(new_n784), .B1(new_n1156), .B2(new_n875), .C(new_n2775), .Y(new_n2776));
  XNOR2x2_ASAP7_75t_L       g02520(.A(\a[17] ), .B(new_n2776), .Y(new_n2777));
  NAND3xp33_ASAP7_75t_L     g02521(.A(new_n2774), .B(new_n2773), .C(new_n2777), .Y(new_n2778));
  AO21x2_ASAP7_75t_L        g02522(.A1(new_n2773), .A2(new_n2774), .B(new_n2777), .Y(new_n2779));
  OR3x1_ASAP7_75t_L         g02523(.A(new_n2592), .B(new_n2594), .C(new_n2597), .Y(new_n2780));
  OAI21xp33_ASAP7_75t_L     g02524(.A1(new_n2426), .A2(new_n2433), .B(new_n2435), .Y(new_n2781));
  OAI21xp33_ASAP7_75t_L     g02525(.A1(new_n2599), .A2(new_n2600), .B(new_n2781), .Y(new_n2782));
  NAND4xp25_ASAP7_75t_L     g02526(.A(new_n2782), .B(new_n2778), .C(new_n2779), .D(new_n2780), .Y(new_n2783));
  AND3x1_ASAP7_75t_L        g02527(.A(new_n2774), .B(new_n2777), .C(new_n2773), .Y(new_n2784));
  AOI21xp33_ASAP7_75t_L     g02528(.A1(new_n2774), .A2(new_n2773), .B(new_n2777), .Y(new_n2785));
  XNOR2x2_ASAP7_75t_L       g02529(.A(new_n2591), .B(new_n2590), .Y(new_n2786));
  MAJIxp5_ASAP7_75t_L       g02530(.A(new_n2601), .B(new_n2597), .C(new_n2786), .Y(new_n2787));
  OAI21xp33_ASAP7_75t_L     g02531(.A1(new_n2785), .A2(new_n2784), .B(new_n2787), .Y(new_n2788));
  AOI22xp33_ASAP7_75t_L     g02532(.A1(new_n811), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n900), .Y(new_n2789));
  OAI221xp5_ASAP7_75t_L     g02533(.A1(new_n904), .A2(new_n1030), .B1(new_n898), .B2(new_n1209), .C(new_n2789), .Y(new_n2790));
  XNOR2x2_ASAP7_75t_L       g02534(.A(\a[14] ), .B(new_n2790), .Y(new_n2791));
  NAND3xp33_ASAP7_75t_L     g02535(.A(new_n2791), .B(new_n2783), .C(new_n2788), .Y(new_n2792));
  AO21x2_ASAP7_75t_L        g02536(.A1(new_n2788), .A2(new_n2783), .B(new_n2791), .Y(new_n2793));
  A2O1A1O1Ixp25_ASAP7_75t_L g02537(.A1(new_n2451), .A2(new_n2449), .B(new_n2519), .C(new_n2611), .D(new_n2624), .Y(new_n2794));
  NAND3xp33_ASAP7_75t_L     g02538(.A(new_n2794), .B(new_n2793), .C(new_n2792), .Y(new_n2795));
  NAND2xp33_ASAP7_75t_L     g02539(.A(new_n2792), .B(new_n2793), .Y(new_n2796));
  A2O1A1Ixp33_ASAP7_75t_L   g02540(.A1(new_n2611), .A2(new_n2623), .B(new_n2624), .C(new_n2796), .Y(new_n2797));
  AOI22xp33_ASAP7_75t_L     g02541(.A1(\b[18] ), .A2(new_n651), .B1(\b[20] ), .B2(new_n581), .Y(new_n2798));
  OAI221xp5_ASAP7_75t_L     g02542(.A1(new_n821), .A2(new_n1432), .B1(new_n577), .B2(new_n1547), .C(new_n2798), .Y(new_n2799));
  XNOR2x2_ASAP7_75t_L       g02543(.A(new_n574), .B(new_n2799), .Y(new_n2800));
  AOI21xp33_ASAP7_75t_L     g02544(.A1(new_n2797), .A2(new_n2795), .B(new_n2800), .Y(new_n2801));
  AND3x1_ASAP7_75t_L        g02545(.A(new_n2797), .B(new_n2800), .C(new_n2795), .Y(new_n2802));
  OAI21xp33_ASAP7_75t_L     g02546(.A1(new_n2801), .A2(new_n2802), .B(new_n2712), .Y(new_n2803));
  NOR3xp33_ASAP7_75t_L      g02547(.A(new_n2712), .B(new_n2801), .C(new_n2802), .Y(new_n2804));
  INVx1_ASAP7_75t_L         g02548(.A(new_n2804), .Y(new_n2805));
  NAND3xp33_ASAP7_75t_L     g02549(.A(new_n2805), .B(new_n2803), .C(new_n2710), .Y(new_n2806));
  OA21x2_ASAP7_75t_L        g02550(.A1(new_n2801), .A2(new_n2802), .B(new_n2712), .Y(new_n2807));
  OAI21xp33_ASAP7_75t_L     g02551(.A1(new_n2804), .A2(new_n2807), .B(new_n2709), .Y(new_n2808));
  NAND3xp33_ASAP7_75t_L     g02552(.A(new_n2706), .B(new_n2806), .C(new_n2808), .Y(new_n2809));
  A2O1A1O1Ixp25_ASAP7_75t_L g02553(.A1(new_n2472), .A2(new_n2484), .B(new_n2468), .C(new_n2638), .D(new_n2645), .Y(new_n2810));
  NOR3xp33_ASAP7_75t_L      g02554(.A(new_n2807), .B(new_n2709), .C(new_n2804), .Y(new_n2811));
  AOI21xp33_ASAP7_75t_L     g02555(.A1(new_n2805), .A2(new_n2803), .B(new_n2710), .Y(new_n2812));
  OAI21xp33_ASAP7_75t_L     g02556(.A1(new_n2811), .A2(new_n2812), .B(new_n2810), .Y(new_n2813));
  AOI21xp33_ASAP7_75t_L     g02557(.A1(new_n2813), .A2(new_n2809), .B(new_n2705), .Y(new_n2814));
  AND3x1_ASAP7_75t_L        g02558(.A(new_n2813), .B(new_n2809), .C(new_n2705), .Y(new_n2815));
  NOR2xp33_ASAP7_75t_L      g02559(.A(new_n2814), .B(new_n2815), .Y(new_n2816));
  O2A1O1Ixp33_ASAP7_75t_L   g02560(.A1(new_n2699), .A2(new_n2700), .B(new_n2702), .C(new_n2816), .Y(new_n2817));
  AO21x2_ASAP7_75t_L        g02561(.A1(new_n2809), .A2(new_n2813), .B(new_n2705), .Y(new_n2818));
  NAND3xp33_ASAP7_75t_L     g02562(.A(new_n2813), .B(new_n2809), .C(new_n2705), .Y(new_n2819));
  NAND2xp33_ASAP7_75t_L     g02563(.A(new_n2819), .B(new_n2818), .Y(new_n2820));
  AOI211xp5_ASAP7_75t_L     g02564(.A1(new_n2657), .A2(new_n2660), .B(new_n2701), .C(new_n2820), .Y(new_n2821));
  NOR3xp33_ASAP7_75t_L      g02565(.A(new_n2821), .B(new_n2817), .C(new_n2698), .Y(new_n2822));
  INVx1_ASAP7_75t_L         g02566(.A(new_n2822), .Y(new_n2823));
  OAI21xp33_ASAP7_75t_L     g02567(.A1(new_n2817), .A2(new_n2821), .B(new_n2698), .Y(new_n2824));
  NAND2xp33_ASAP7_75t_L     g02568(.A(new_n2824), .B(new_n2823), .Y(new_n2825));
  XOR2x2_ASAP7_75t_L        g02569(.A(new_n2684), .B(new_n2825), .Y(\f[29] ));
  AND3x1_ASAP7_75t_L        g02570(.A(new_n2770), .B(new_n2765), .C(new_n2717), .Y(new_n2827));
  AO21x2_ASAP7_75t_L        g02571(.A1(new_n2771), .A2(new_n2714), .B(new_n2827), .Y(new_n2828));
  AOI22xp33_ASAP7_75t_L     g02572(.A1(new_n1360), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1581), .Y(new_n2829));
  OAI21xp33_ASAP7_75t_L     g02573(.A1(new_n1359), .A2(new_n768), .B(new_n2829), .Y(new_n2830));
  AOI211xp5_ASAP7_75t_L     g02574(.A1(\b[11] ), .A2(new_n1362), .B(new_n1356), .C(new_n2830), .Y(new_n2831));
  NAND2xp33_ASAP7_75t_L     g02575(.A(\b[11] ), .B(new_n1362), .Y(new_n2832));
  NAND2xp33_ASAP7_75t_L     g02576(.A(new_n1365), .B(new_n1232), .Y(new_n2833));
  AOI31xp33_ASAP7_75t_L     g02577(.A1(new_n2833), .A2(new_n2832), .A3(new_n2829), .B(\a[20] ), .Y(new_n2834));
  NOR2xp33_ASAP7_75t_L      g02578(.A(new_n2834), .B(new_n2831), .Y(new_n2835));
  AOI21xp33_ASAP7_75t_L     g02579(.A1(new_n2718), .A2(new_n2757), .B(new_n2769), .Y(new_n2836));
  NAND4xp25_ASAP7_75t_L     g02580(.A(new_n2554), .B(\a[29] ), .C(new_n2383), .D(new_n2550), .Y(new_n2837));
  INVx1_ASAP7_75t_L         g02581(.A(\a[30] ), .Y(new_n2838));
  NAND2xp33_ASAP7_75t_L     g02582(.A(\a[29] ), .B(new_n2838), .Y(new_n2839));
  NAND2xp33_ASAP7_75t_L     g02583(.A(\a[30] ), .B(new_n2538), .Y(new_n2840));
  NAND2xp33_ASAP7_75t_L     g02584(.A(new_n2840), .B(new_n2839), .Y(new_n2841));
  NAND2xp33_ASAP7_75t_L     g02585(.A(\b[0] ), .B(new_n2841), .Y(new_n2842));
  INVx1_ASAP7_75t_L         g02586(.A(new_n2842), .Y(new_n2843));
  OAI31xp33_ASAP7_75t_L     g02587(.A1(new_n2837), .A2(new_n2748), .A3(new_n2732), .B(new_n2843), .Y(new_n2844));
  A2O1A1Ixp33_ASAP7_75t_L   g02588(.A1(new_n2380), .A2(new_n2381), .B(new_n258), .C(\a[29] ), .Y(new_n2845));
  AOI211xp5_ASAP7_75t_L     g02589(.A1(new_n2544), .A2(new_n269), .B(new_n2845), .C(new_n2548), .Y(new_n2846));
  NAND4xp25_ASAP7_75t_L     g02590(.A(new_n2846), .B(new_n2842), .C(new_n2737), .D(new_n2733), .Y(new_n2847));
  NOR2xp33_ASAP7_75t_L      g02591(.A(new_n276), .B(new_n2547), .Y(new_n2848));
  OAI22xp33_ASAP7_75t_L     g02592(.A1(new_n2747), .A2(new_n261), .B1(new_n298), .B2(new_n2545), .Y(new_n2849));
  AOI211xp5_ASAP7_75t_L     g02593(.A1(new_n406), .A2(new_n2544), .B(new_n2848), .C(new_n2849), .Y(new_n2850));
  NAND2xp33_ASAP7_75t_L     g02594(.A(\a[29] ), .B(new_n2850), .Y(new_n2851));
  NOR2xp33_ASAP7_75t_L      g02595(.A(new_n2734), .B(new_n302), .Y(new_n2852));
  OAI31xp33_ASAP7_75t_L     g02596(.A1(new_n2852), .A2(new_n2848), .A3(new_n2849), .B(new_n2538), .Y(new_n2853));
  AO22x1_ASAP7_75t_L        g02597(.A1(new_n2853), .A2(new_n2851), .B1(new_n2844), .B2(new_n2847), .Y(new_n2854));
  NAND4xp25_ASAP7_75t_L     g02598(.A(new_n2847), .B(new_n2844), .C(new_n2851), .D(new_n2853), .Y(new_n2855));
  NAND2xp33_ASAP7_75t_L     g02599(.A(\b[5] ), .B(new_n2115), .Y(new_n2856));
  NAND2xp33_ASAP7_75t_L     g02600(.A(new_n2106), .B(new_n526), .Y(new_n2857));
  AOI22xp33_ASAP7_75t_L     g02601(.A1(new_n2114), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n2259), .Y(new_n2858));
  NAND4xp25_ASAP7_75t_L     g02602(.A(new_n2857), .B(\a[26] ), .C(new_n2856), .D(new_n2858), .Y(new_n2859));
  OAI21xp33_ASAP7_75t_L     g02603(.A1(new_n2257), .A2(new_n390), .B(new_n2858), .Y(new_n2860));
  A2O1A1Ixp33_ASAP7_75t_L   g02604(.A1(\b[5] ), .A2(new_n2115), .B(new_n2860), .C(new_n2100), .Y(new_n2861));
  NAND4xp25_ASAP7_75t_L     g02605(.A(new_n2861), .B(new_n2854), .C(new_n2855), .D(new_n2859), .Y(new_n2862));
  AO22x1_ASAP7_75t_L        g02606(.A1(new_n2855), .A2(new_n2854), .B1(new_n2861), .B2(new_n2859), .Y(new_n2863));
  AOI31xp33_ASAP7_75t_L     g02607(.A1(new_n2568), .A2(new_n2753), .A3(new_n2725), .B(new_n2760), .Y(new_n2864));
  NAND3xp33_ASAP7_75t_L     g02608(.A(new_n2864), .B(new_n2863), .C(new_n2862), .Y(new_n2865));
  NAND2xp33_ASAP7_75t_L     g02609(.A(new_n2862), .B(new_n2863), .Y(new_n2866));
  AO31x2_ASAP7_75t_L        g02610(.A1(new_n2568), .A2(new_n2753), .A3(new_n2725), .B(new_n2760), .Y(new_n2867));
  NAND2xp33_ASAP7_75t_L     g02611(.A(new_n2867), .B(new_n2866), .Y(new_n2868));
  AOI22xp33_ASAP7_75t_L     g02612(.A1(new_n1704), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1837), .Y(new_n2869));
  OAI221xp5_ASAP7_75t_L     g02613(.A1(new_n1699), .A2(new_n488), .B1(new_n1827), .B2(new_n548), .C(new_n2869), .Y(new_n2870));
  OR2x4_ASAP7_75t_L         g02614(.A(new_n1689), .B(new_n2870), .Y(new_n2871));
  NAND2xp33_ASAP7_75t_L     g02615(.A(new_n1689), .B(new_n2870), .Y(new_n2872));
  AOI22xp33_ASAP7_75t_L     g02616(.A1(new_n2871), .A2(new_n2872), .B1(new_n2865), .B2(new_n2868), .Y(new_n2873));
  NAND4xp25_ASAP7_75t_L     g02617(.A(new_n2868), .B(new_n2865), .C(new_n2871), .D(new_n2872), .Y(new_n2874));
  INVx1_ASAP7_75t_L         g02618(.A(new_n2874), .Y(new_n2875));
  NOR3xp33_ASAP7_75t_L      g02619(.A(new_n2836), .B(new_n2873), .C(new_n2875), .Y(new_n2876));
  AO22x1_ASAP7_75t_L        g02620(.A1(new_n2872), .A2(new_n2871), .B1(new_n2865), .B2(new_n2868), .Y(new_n2877));
  AOI221xp5_ASAP7_75t_L     g02621(.A1(new_n2718), .A2(new_n2757), .B1(new_n2874), .B2(new_n2877), .C(new_n2769), .Y(new_n2878));
  OAI21xp33_ASAP7_75t_L     g02622(.A1(new_n2878), .A2(new_n2876), .B(new_n2835), .Y(new_n2879));
  NAND4xp25_ASAP7_75t_L     g02623(.A(new_n2833), .B(\a[20] ), .C(new_n2832), .D(new_n2829), .Y(new_n2880));
  A2O1A1Ixp33_ASAP7_75t_L   g02624(.A1(\b[11] ), .A2(new_n1362), .B(new_n2830), .C(new_n1356), .Y(new_n2881));
  NAND2xp33_ASAP7_75t_L     g02625(.A(new_n2880), .B(new_n2881), .Y(new_n2882));
  OAI21xp33_ASAP7_75t_L     g02626(.A1(new_n2768), .A2(new_n2767), .B(new_n2764), .Y(new_n2883));
  NAND3xp33_ASAP7_75t_L     g02627(.A(new_n2883), .B(new_n2877), .C(new_n2874), .Y(new_n2884));
  OAI21xp33_ASAP7_75t_L     g02628(.A1(new_n2873), .A2(new_n2875), .B(new_n2836), .Y(new_n2885));
  NAND3xp33_ASAP7_75t_L     g02629(.A(new_n2884), .B(new_n2882), .C(new_n2885), .Y(new_n2886));
  NAND3xp33_ASAP7_75t_L     g02630(.A(new_n2828), .B(new_n2879), .C(new_n2886), .Y(new_n2887));
  NAND2xp33_ASAP7_75t_L     g02631(.A(new_n2575), .B(new_n2572), .Y(new_n2888));
  NOR2xp33_ASAP7_75t_L      g02632(.A(new_n2582), .B(new_n2888), .Y(new_n2889));
  A2O1A1O1Ixp25_ASAP7_75t_L g02633(.A1(new_n2591), .A2(new_n2590), .B(new_n2889), .C(new_n2771), .D(new_n2827), .Y(new_n2890));
  NAND2xp33_ASAP7_75t_L     g02634(.A(new_n2879), .B(new_n2886), .Y(new_n2891));
  NAND2xp33_ASAP7_75t_L     g02635(.A(new_n2890), .B(new_n2891), .Y(new_n2892));
  AOI22xp33_ASAP7_75t_L     g02636(.A1(new_n1076), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1253), .Y(new_n2893));
  OAI221xp5_ASAP7_75t_L     g02637(.A1(new_n1154), .A2(new_n869), .B1(new_n1156), .B2(new_n950), .C(new_n2893), .Y(new_n2894));
  XNOR2x2_ASAP7_75t_L       g02638(.A(\a[17] ), .B(new_n2894), .Y(new_n2895));
  NAND3xp33_ASAP7_75t_L     g02639(.A(new_n2887), .B(new_n2892), .C(new_n2895), .Y(new_n2896));
  NOR2xp33_ASAP7_75t_L      g02640(.A(new_n2890), .B(new_n2891), .Y(new_n2897));
  AOI21xp33_ASAP7_75t_L     g02641(.A1(new_n2886), .A2(new_n2879), .B(new_n2828), .Y(new_n2898));
  INVx1_ASAP7_75t_L         g02642(.A(new_n2895), .Y(new_n2899));
  OAI21xp33_ASAP7_75t_L     g02643(.A1(new_n2898), .A2(new_n2897), .B(new_n2899), .Y(new_n2900));
  INVx1_ASAP7_75t_L         g02644(.A(new_n2777), .Y(new_n2901));
  AND3x1_ASAP7_75t_L        g02645(.A(new_n2901), .B(new_n2774), .C(new_n2773), .Y(new_n2902));
  O2A1O1Ixp33_ASAP7_75t_L   g02646(.A1(new_n2785), .A2(new_n2784), .B(new_n2787), .C(new_n2902), .Y(new_n2903));
  NAND3xp33_ASAP7_75t_L     g02647(.A(new_n2903), .B(new_n2900), .C(new_n2896), .Y(new_n2904));
  INVx1_ASAP7_75t_L         g02648(.A(new_n2902), .Y(new_n2905));
  AO22x1_ASAP7_75t_L        g02649(.A1(new_n2896), .A2(new_n2900), .B1(new_n2905), .B2(new_n2788), .Y(new_n2906));
  OAI22xp33_ASAP7_75t_L     g02650(.A1(new_n978), .A2(new_n1030), .B1(new_n1313), .B2(new_n977), .Y(new_n2907));
  AOI221xp5_ASAP7_75t_L     g02651(.A1(\b[17] ), .A2(new_n815), .B1(new_n808), .B2(new_n1319), .C(new_n2907), .Y(new_n2908));
  XNOR2x2_ASAP7_75t_L       g02652(.A(new_n806), .B(new_n2908), .Y(new_n2909));
  NAND3xp33_ASAP7_75t_L     g02653(.A(new_n2906), .B(new_n2904), .C(new_n2909), .Y(new_n2910));
  AND4x1_ASAP7_75t_L        g02654(.A(new_n2788), .B(new_n2905), .C(new_n2896), .D(new_n2900), .Y(new_n2911));
  AOI21xp33_ASAP7_75t_L     g02655(.A1(new_n2900), .A2(new_n2896), .B(new_n2903), .Y(new_n2912));
  XNOR2x2_ASAP7_75t_L       g02656(.A(\a[14] ), .B(new_n2908), .Y(new_n2913));
  OAI21xp33_ASAP7_75t_L     g02657(.A1(new_n2912), .A2(new_n2911), .B(new_n2913), .Y(new_n2914));
  NAND2xp33_ASAP7_75t_L     g02658(.A(new_n2914), .B(new_n2910), .Y(new_n2915));
  NAND2xp33_ASAP7_75t_L     g02659(.A(new_n2788), .B(new_n2783), .Y(new_n2916));
  MAJIxp5_ASAP7_75t_L       g02660(.A(new_n2794), .B(new_n2916), .C(new_n2791), .Y(new_n2917));
  NOR2xp33_ASAP7_75t_L      g02661(.A(new_n2917), .B(new_n2915), .Y(new_n2918));
  NOR3xp33_ASAP7_75t_L      g02662(.A(new_n2911), .B(new_n2912), .C(new_n2913), .Y(new_n2919));
  AOI21xp33_ASAP7_75t_L     g02663(.A1(new_n2906), .A2(new_n2904), .B(new_n2909), .Y(new_n2920));
  OA21x2_ASAP7_75t_L        g02664(.A1(new_n2919), .A2(new_n2920), .B(new_n2917), .Y(new_n2921));
  AOI22xp33_ASAP7_75t_L     g02665(.A1(\b[19] ), .A2(new_n651), .B1(\b[21] ), .B2(new_n581), .Y(new_n2922));
  OAI221xp5_ASAP7_75t_L     g02666(.A1(new_n821), .A2(new_n1539), .B1(new_n577), .B2(new_n1662), .C(new_n2922), .Y(new_n2923));
  XNOR2x2_ASAP7_75t_L       g02667(.A(new_n574), .B(new_n2923), .Y(new_n2924));
  NOR3xp33_ASAP7_75t_L      g02668(.A(new_n2921), .B(new_n2918), .C(new_n2924), .Y(new_n2925));
  NOR2xp33_ASAP7_75t_L      g02669(.A(new_n2919), .B(new_n2920), .Y(new_n2926));
  MAJx2_ASAP7_75t_L         g02670(.A(new_n2794), .B(new_n2791), .C(new_n2916), .Y(new_n2927));
  NAND2xp33_ASAP7_75t_L     g02671(.A(new_n2926), .B(new_n2927), .Y(new_n2928));
  NAND2xp33_ASAP7_75t_L     g02672(.A(new_n2917), .B(new_n2915), .Y(new_n2929));
  XNOR2x2_ASAP7_75t_L       g02673(.A(\a[11] ), .B(new_n2923), .Y(new_n2930));
  AOI21xp33_ASAP7_75t_L     g02674(.A1(new_n2928), .A2(new_n2929), .B(new_n2930), .Y(new_n2931));
  INVx1_ASAP7_75t_L         g02675(.A(new_n2711), .Y(new_n2932));
  NAND3xp33_ASAP7_75t_L     g02676(.A(new_n2797), .B(new_n2795), .C(new_n2800), .Y(new_n2933));
  AO31x2_ASAP7_75t_L        g02677(.A1(new_n2633), .A2(new_n2933), .A3(new_n2932), .B(new_n2801), .Y(new_n2934));
  NOR3xp33_ASAP7_75t_L      g02678(.A(new_n2934), .B(new_n2931), .C(new_n2925), .Y(new_n2935));
  NAND3xp33_ASAP7_75t_L     g02679(.A(new_n2928), .B(new_n2929), .C(new_n2930), .Y(new_n2936));
  OAI21xp33_ASAP7_75t_L     g02680(.A1(new_n2918), .A2(new_n2921), .B(new_n2924), .Y(new_n2937));
  AOI31xp33_ASAP7_75t_L     g02681(.A1(new_n2633), .A2(new_n2932), .A3(new_n2933), .B(new_n2801), .Y(new_n2938));
  AOI21xp33_ASAP7_75t_L     g02682(.A1(new_n2937), .A2(new_n2936), .B(new_n2938), .Y(new_n2939));
  AOI22xp33_ASAP7_75t_L     g02683(.A1(new_n444), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n471), .Y(new_n2940));
  OAI31xp33_ASAP7_75t_L     g02684(.A1(new_n1934), .A2(new_n469), .A3(new_n1933), .B(new_n2940), .Y(new_n2941));
  AOI21xp33_ASAP7_75t_L     g02685(.A1(new_n447), .A2(\b[23] ), .B(new_n2941), .Y(new_n2942));
  NAND2xp33_ASAP7_75t_L     g02686(.A(\a[8] ), .B(new_n2942), .Y(new_n2943));
  A2O1A1Ixp33_ASAP7_75t_L   g02687(.A1(\b[23] ), .A2(new_n447), .B(new_n2941), .C(new_n435), .Y(new_n2944));
  NAND2xp33_ASAP7_75t_L     g02688(.A(new_n2944), .B(new_n2943), .Y(new_n2945));
  OAI21xp33_ASAP7_75t_L     g02689(.A1(new_n2939), .A2(new_n2935), .B(new_n2945), .Y(new_n2946));
  NAND3xp33_ASAP7_75t_L     g02690(.A(new_n2938), .B(new_n2937), .C(new_n2936), .Y(new_n2947));
  OAI21xp33_ASAP7_75t_L     g02691(.A1(new_n2925), .A2(new_n2931), .B(new_n2934), .Y(new_n2948));
  XNOR2x2_ASAP7_75t_L       g02692(.A(new_n435), .B(new_n2942), .Y(new_n2949));
  NAND3xp33_ASAP7_75t_L     g02693(.A(new_n2948), .B(new_n2947), .C(new_n2949), .Y(new_n2950));
  AOI221xp5_ASAP7_75t_L     g02694(.A1(new_n2808), .A2(new_n2706), .B1(new_n2950), .B2(new_n2946), .C(new_n2811), .Y(new_n2951));
  A2O1A1O1Ixp25_ASAP7_75t_L g02695(.A1(new_n2638), .A2(new_n2642), .B(new_n2645), .C(new_n2808), .D(new_n2811), .Y(new_n2952));
  AOI21xp33_ASAP7_75t_L     g02696(.A1(new_n2948), .A2(new_n2947), .B(new_n2949), .Y(new_n2953));
  NOR3xp33_ASAP7_75t_L      g02697(.A(new_n2935), .B(new_n2939), .C(new_n2945), .Y(new_n2954));
  NOR3xp33_ASAP7_75t_L      g02698(.A(new_n2952), .B(new_n2953), .C(new_n2954), .Y(new_n2955));
  NAND2xp33_ASAP7_75t_L     g02699(.A(\b[26] ), .B(new_n347), .Y(new_n2956));
  NAND2xp33_ASAP7_75t_L     g02700(.A(new_n341), .B(new_n2504), .Y(new_n2957));
  AOI22xp33_ASAP7_75t_L     g02701(.A1(new_n344), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n370), .Y(new_n2958));
  AND4x1_ASAP7_75t_L        g02702(.A(new_n2958), .B(new_n2957), .C(new_n2956), .D(\a[5] ), .Y(new_n2959));
  AOI31xp33_ASAP7_75t_L     g02703(.A1(new_n2957), .A2(new_n2956), .A3(new_n2958), .B(\a[5] ), .Y(new_n2960));
  NOR2xp33_ASAP7_75t_L      g02704(.A(new_n2960), .B(new_n2959), .Y(new_n2961));
  INVx1_ASAP7_75t_L         g02705(.A(new_n2961), .Y(new_n2962));
  NOR3xp33_ASAP7_75t_L      g02706(.A(new_n2955), .B(new_n2951), .C(new_n2962), .Y(new_n2963));
  OA21x2_ASAP7_75t_L        g02707(.A1(new_n2951), .A2(new_n2955), .B(new_n2962), .Y(new_n2964));
  NOR2xp33_ASAP7_75t_L      g02708(.A(new_n2963), .B(new_n2964), .Y(new_n2965));
  INVx1_ASAP7_75t_L         g02709(.A(new_n2705), .Y(new_n2966));
  NAND3xp33_ASAP7_75t_L     g02710(.A(new_n2813), .B(new_n2809), .C(new_n2966), .Y(new_n2967));
  INVx1_ASAP7_75t_L         g02711(.A(new_n2967), .Y(new_n2968));
  A2O1A1O1Ixp25_ASAP7_75t_L g02712(.A1(new_n2657), .A2(new_n2660), .B(new_n2701), .C(new_n2820), .D(new_n2968), .Y(new_n2969));
  NAND2xp33_ASAP7_75t_L     g02713(.A(new_n2965), .B(new_n2969), .Y(new_n2970));
  A2O1A1Ixp33_ASAP7_75t_L   g02714(.A1(new_n2494), .A2(new_n2659), .B(new_n2699), .C(new_n2702), .Y(new_n2971));
  OAI21xp33_ASAP7_75t_L     g02715(.A1(new_n2953), .A2(new_n2954), .B(new_n2952), .Y(new_n2972));
  NOR2xp33_ASAP7_75t_L      g02716(.A(new_n2953), .B(new_n2954), .Y(new_n2973));
  A2O1A1Ixp33_ASAP7_75t_L   g02717(.A1(new_n2808), .A2(new_n2706), .B(new_n2811), .C(new_n2973), .Y(new_n2974));
  NAND3xp33_ASAP7_75t_L     g02718(.A(new_n2974), .B(new_n2972), .C(new_n2961), .Y(new_n2975));
  OAI21xp33_ASAP7_75t_L     g02719(.A1(new_n2951), .A2(new_n2955), .B(new_n2962), .Y(new_n2976));
  NAND2xp33_ASAP7_75t_L     g02720(.A(new_n2976), .B(new_n2975), .Y(new_n2977));
  A2O1A1Ixp33_ASAP7_75t_L   g02721(.A1(new_n2971), .A2(new_n2820), .B(new_n2968), .C(new_n2977), .Y(new_n2978));
  NAND2xp33_ASAP7_75t_L     g02722(.A(new_n2978), .B(new_n2970), .Y(new_n2979));
  INVx1_ASAP7_75t_L         g02723(.A(new_n2689), .Y(new_n2980));
  NOR2xp33_ASAP7_75t_L      g02724(.A(\b[29] ), .B(\b[30] ), .Y(new_n2981));
  INVx1_ASAP7_75t_L         g02725(.A(\b[30] ), .Y(new_n2982));
  NOR2xp33_ASAP7_75t_L      g02726(.A(new_n2688), .B(new_n2982), .Y(new_n2983));
  NOR2xp33_ASAP7_75t_L      g02727(.A(new_n2981), .B(new_n2983), .Y(new_n2984));
  INVx1_ASAP7_75t_L         g02728(.A(new_n2984), .Y(new_n2985));
  O2A1O1Ixp33_ASAP7_75t_L   g02729(.A1(new_n2693), .A2(new_n2692), .B(new_n2980), .C(new_n2985), .Y(new_n2986));
  O2A1O1Ixp33_ASAP7_75t_L   g02730(.A1(new_n2497), .A2(new_n2666), .B(new_n2669), .C(new_n2693), .Y(new_n2987));
  NOR3xp33_ASAP7_75t_L      g02731(.A(new_n2987), .B(new_n2984), .C(new_n2689), .Y(new_n2988));
  NOR2xp33_ASAP7_75t_L      g02732(.A(new_n2986), .B(new_n2988), .Y(new_n2989));
  INVx1_ASAP7_75t_L         g02733(.A(new_n2989), .Y(new_n2990));
  AOI22xp33_ASAP7_75t_L     g02734(.A1(\b[28] ), .A2(new_n282), .B1(\b[30] ), .B2(new_n303), .Y(new_n2991));
  OAI221xp5_ASAP7_75t_L     g02735(.A1(new_n291), .A2(new_n2688), .B1(new_n268), .B2(new_n2990), .C(new_n2991), .Y(new_n2992));
  XNOR2x2_ASAP7_75t_L       g02736(.A(\a[2] ), .B(new_n2992), .Y(new_n2993));
  XNOR2x2_ASAP7_75t_L       g02737(.A(new_n2993), .B(new_n2979), .Y(new_n2994));
  O2A1O1Ixp33_ASAP7_75t_L   g02738(.A1(new_n2684), .A2(new_n2825), .B(new_n2823), .C(new_n2994), .Y(new_n2995));
  A2O1A1O1Ixp25_ASAP7_75t_L g02739(.A1(new_n2676), .A2(new_n2681), .B(new_n2677), .C(new_n2824), .D(new_n2822), .Y(new_n2996));
  AND2x2_ASAP7_75t_L        g02740(.A(new_n2996), .B(new_n2994), .Y(new_n2997));
  NOR2xp33_ASAP7_75t_L      g02741(.A(new_n2995), .B(new_n2997), .Y(\f[30] ));
  NAND2xp33_ASAP7_75t_L     g02742(.A(new_n2859), .B(new_n2861), .Y(new_n2999));
  AND3x1_ASAP7_75t_L        g02743(.A(new_n2999), .B(new_n2855), .C(new_n2854), .Y(new_n3000));
  AOI22xp33_ASAP7_75t_L     g02744(.A1(new_n2114), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n2259), .Y(new_n3001));
  INVx1_ASAP7_75t_L         g02745(.A(new_n3001), .Y(new_n3002));
  AOI221xp5_ASAP7_75t_L     g02746(.A1(new_n2115), .A2(\b[6] ), .B1(new_n2106), .B2(new_n2084), .C(new_n3002), .Y(new_n3003));
  NAND2xp33_ASAP7_75t_L     g02747(.A(\a[26] ), .B(new_n3003), .Y(new_n3004));
  OAI21xp33_ASAP7_75t_L     g02748(.A1(new_n2257), .A2(new_n425), .B(new_n3001), .Y(new_n3005));
  A2O1A1Ixp33_ASAP7_75t_L   g02749(.A1(\b[6] ), .A2(new_n2115), .B(new_n3005), .C(new_n2100), .Y(new_n3006));
  NOR3xp33_ASAP7_75t_L      g02750(.A(new_n2738), .B(new_n2842), .C(new_n2837), .Y(new_n3007));
  INVx1_ASAP7_75t_L         g02751(.A(new_n3007), .Y(new_n3008));
  NOR2xp33_ASAP7_75t_L      g02752(.A(new_n298), .B(new_n2547), .Y(new_n3009));
  NOR3xp33_ASAP7_75t_L      g02753(.A(new_n326), .B(new_n328), .C(new_n2734), .Y(new_n3010));
  OAI22xp33_ASAP7_75t_L     g02754(.A1(new_n2747), .A2(new_n276), .B1(new_n324), .B2(new_n2545), .Y(new_n3011));
  NOR4xp25_ASAP7_75t_L      g02755(.A(new_n3010), .B(new_n3011), .C(new_n2538), .D(new_n3009), .Y(new_n3012));
  OA31x2_ASAP7_75t_L        g02756(.A1(new_n3009), .A2(new_n3011), .A3(new_n3010), .B1(new_n2538), .Y(new_n3013));
  NOR2xp33_ASAP7_75t_L      g02757(.A(new_n3012), .B(new_n3013), .Y(new_n3014));
  INVx1_ASAP7_75t_L         g02758(.A(\a[32] ), .Y(new_n3015));
  NOR2xp33_ASAP7_75t_L      g02759(.A(new_n3015), .B(new_n2842), .Y(new_n3016));
  AND2x2_ASAP7_75t_L        g02760(.A(new_n2839), .B(new_n2840), .Y(new_n3017));
  INVx1_ASAP7_75t_L         g02761(.A(\a[31] ), .Y(new_n3018));
  NAND2xp33_ASAP7_75t_L     g02762(.A(\a[32] ), .B(new_n3018), .Y(new_n3019));
  NAND2xp33_ASAP7_75t_L     g02763(.A(\a[31] ), .B(new_n3015), .Y(new_n3020));
  AOI21xp33_ASAP7_75t_L     g02764(.A1(new_n3020), .A2(new_n3019), .B(new_n3017), .Y(new_n3021));
  NAND3xp33_ASAP7_75t_L     g02765(.A(new_n2841), .B(new_n3019), .C(new_n3020), .Y(new_n3022));
  XNOR2x2_ASAP7_75t_L       g02766(.A(\a[31] ), .B(\a[30] ), .Y(new_n3023));
  OR2x4_ASAP7_75t_L         g02767(.A(new_n3023), .B(new_n2841), .Y(new_n3024));
  OAI22xp33_ASAP7_75t_L     g02768(.A1(new_n3024), .A2(new_n258), .B1(new_n261), .B2(new_n3022), .Y(new_n3025));
  A2O1A1Ixp33_ASAP7_75t_L   g02769(.A1(new_n269), .A2(new_n3021), .B(new_n3025), .C(new_n3016), .Y(new_n3026));
  NAND2xp33_ASAP7_75t_L     g02770(.A(new_n269), .B(new_n3021), .Y(new_n3027));
  NAND2xp33_ASAP7_75t_L     g02771(.A(new_n3020), .B(new_n3019), .Y(new_n3028));
  NOR2xp33_ASAP7_75t_L      g02772(.A(new_n3028), .B(new_n3017), .Y(new_n3029));
  NOR2xp33_ASAP7_75t_L      g02773(.A(new_n3023), .B(new_n2841), .Y(new_n3030));
  AOI22xp33_ASAP7_75t_L     g02774(.A1(\b[0] ), .A2(new_n3030), .B1(\b[1] ), .B2(new_n3029), .Y(new_n3031));
  OAI211xp5_ASAP7_75t_L     g02775(.A1(new_n3015), .A2(new_n2842), .B(new_n3031), .C(new_n3027), .Y(new_n3032));
  AND2x2_ASAP7_75t_L        g02776(.A(new_n3032), .B(new_n3026), .Y(new_n3033));
  NAND2xp33_ASAP7_75t_L     g02777(.A(new_n3033), .B(new_n3014), .Y(new_n3034));
  NAND2xp33_ASAP7_75t_L     g02778(.A(new_n3032), .B(new_n3026), .Y(new_n3035));
  OAI21xp33_ASAP7_75t_L     g02779(.A1(new_n3012), .A2(new_n3013), .B(new_n3035), .Y(new_n3036));
  AOI22xp33_ASAP7_75t_L     g02780(.A1(new_n3034), .A2(new_n3036), .B1(new_n3008), .B2(new_n2854), .Y(new_n3037));
  AOI22xp33_ASAP7_75t_L     g02781(.A1(new_n2851), .A2(new_n2853), .B1(new_n2844), .B2(new_n2847), .Y(new_n3038));
  NOR3xp33_ASAP7_75t_L      g02782(.A(new_n3035), .B(new_n3013), .C(new_n3012), .Y(new_n3039));
  OA21x2_ASAP7_75t_L        g02783(.A1(new_n3013), .A2(new_n3012), .B(new_n3035), .Y(new_n3040));
  NOR4xp25_ASAP7_75t_L      g02784(.A(new_n3038), .B(new_n3040), .C(new_n3039), .D(new_n3007), .Y(new_n3041));
  AOI211xp5_ASAP7_75t_L     g02785(.A1(new_n3006), .A2(new_n3004), .B(new_n3041), .C(new_n3037), .Y(new_n3042));
  INVx1_ASAP7_75t_L         g02786(.A(new_n3004), .Y(new_n3043));
  INVx1_ASAP7_75t_L         g02787(.A(new_n3006), .Y(new_n3044));
  OAI22xp33_ASAP7_75t_L     g02788(.A1(new_n3038), .A2(new_n3007), .B1(new_n3039), .B2(new_n3040), .Y(new_n3045));
  NAND4xp25_ASAP7_75t_L     g02789(.A(new_n2854), .B(new_n3034), .C(new_n3036), .D(new_n3008), .Y(new_n3046));
  AOI211xp5_ASAP7_75t_L     g02790(.A1(new_n3045), .A2(new_n3046), .B(new_n3044), .C(new_n3043), .Y(new_n3047));
  NOR2xp33_ASAP7_75t_L      g02791(.A(new_n3042), .B(new_n3047), .Y(new_n3048));
  A2O1A1Ixp33_ASAP7_75t_L   g02792(.A1(new_n2864), .A2(new_n2866), .B(new_n3000), .C(new_n3048), .Y(new_n3049));
  AND4x1_ASAP7_75t_L        g02793(.A(new_n2854), .B(new_n2861), .C(new_n2855), .D(new_n2859), .Y(new_n3050));
  AOI22xp33_ASAP7_75t_L     g02794(.A1(new_n2854), .A2(new_n2855), .B1(new_n2859), .B2(new_n2861), .Y(new_n3051));
  O2A1O1Ixp33_ASAP7_75t_L   g02795(.A1(new_n3050), .A2(new_n3051), .B(new_n2864), .C(new_n3000), .Y(new_n3052));
  OAI21xp33_ASAP7_75t_L     g02796(.A1(new_n3042), .A2(new_n3047), .B(new_n3052), .Y(new_n3053));
  NOR2xp33_ASAP7_75t_L      g02797(.A(new_n540), .B(new_n1699), .Y(new_n3054));
  INVx1_ASAP7_75t_L         g02798(.A(new_n3054), .Y(new_n3055));
  NAND2xp33_ASAP7_75t_L     g02799(.A(new_n1695), .B(new_n2143), .Y(new_n3056));
  AOI22xp33_ASAP7_75t_L     g02800(.A1(new_n1704), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1837), .Y(new_n3057));
  NAND4xp25_ASAP7_75t_L     g02801(.A(new_n3056), .B(\a[23] ), .C(new_n3055), .D(new_n3057), .Y(new_n3058));
  OAI21xp33_ASAP7_75t_L     g02802(.A1(new_n1827), .A2(new_n624), .B(new_n3057), .Y(new_n3059));
  A2O1A1Ixp33_ASAP7_75t_L   g02803(.A1(\b[9] ), .A2(new_n1706), .B(new_n3059), .C(new_n1689), .Y(new_n3060));
  AND2x2_ASAP7_75t_L        g02804(.A(new_n3058), .B(new_n3060), .Y(new_n3061));
  NAND3xp33_ASAP7_75t_L     g02805(.A(new_n3049), .B(new_n3061), .C(new_n3053), .Y(new_n3062));
  NAND3xp33_ASAP7_75t_L     g02806(.A(new_n2999), .B(new_n2855), .C(new_n2854), .Y(new_n3063));
  OAI221xp5_ASAP7_75t_L     g02807(.A1(new_n3050), .A2(new_n3051), .B1(new_n2761), .B2(new_n2726), .C(new_n2742), .Y(new_n3064));
  AOI211xp5_ASAP7_75t_L     g02808(.A1(new_n3064), .A2(new_n3063), .B(new_n3042), .C(new_n3047), .Y(new_n3065));
  OAI211xp5_ASAP7_75t_L     g02809(.A1(new_n3044), .A2(new_n3043), .B(new_n3046), .C(new_n3045), .Y(new_n3066));
  OAI211xp5_ASAP7_75t_L     g02810(.A1(new_n3041), .A2(new_n3037), .B(new_n3006), .C(new_n3004), .Y(new_n3067));
  AOI221xp5_ASAP7_75t_L     g02811(.A1(new_n2866), .A2(new_n2864), .B1(new_n3067), .B2(new_n3066), .C(new_n3000), .Y(new_n3068));
  NAND2xp33_ASAP7_75t_L     g02812(.A(new_n3058), .B(new_n3060), .Y(new_n3069));
  OAI21xp33_ASAP7_75t_L     g02813(.A1(new_n3068), .A2(new_n3065), .B(new_n3069), .Y(new_n3070));
  NAND2xp33_ASAP7_75t_L     g02814(.A(new_n3070), .B(new_n3062), .Y(new_n3071));
  A2O1A1O1Ixp25_ASAP7_75t_L g02815(.A1(new_n2757), .A2(new_n2718), .B(new_n2769), .C(new_n2874), .D(new_n2873), .Y(new_n3072));
  INVx1_ASAP7_75t_L         g02816(.A(new_n3072), .Y(new_n3073));
  NOR2xp33_ASAP7_75t_L      g02817(.A(new_n3071), .B(new_n3073), .Y(new_n3074));
  NOR3xp33_ASAP7_75t_L      g02818(.A(new_n3065), .B(new_n3068), .C(new_n3069), .Y(new_n3075));
  AOI21xp33_ASAP7_75t_L     g02819(.A1(new_n3049), .A2(new_n3053), .B(new_n3061), .Y(new_n3076));
  NOR2xp33_ASAP7_75t_L      g02820(.A(new_n3075), .B(new_n3076), .Y(new_n3077));
  NOR2xp33_ASAP7_75t_L      g02821(.A(new_n3072), .B(new_n3077), .Y(new_n3078));
  AOI22xp33_ASAP7_75t_L     g02822(.A1(new_n1360), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1581), .Y(new_n3079));
  OAI221xp5_ASAP7_75t_L     g02823(.A1(new_n1373), .A2(new_n760), .B1(new_n1359), .B2(new_n790), .C(new_n3079), .Y(new_n3080));
  XNOR2x2_ASAP7_75t_L       g02824(.A(\a[20] ), .B(new_n3080), .Y(new_n3081));
  OAI21xp33_ASAP7_75t_L     g02825(.A1(new_n3074), .A2(new_n3078), .B(new_n3081), .Y(new_n3082));
  NAND2xp33_ASAP7_75t_L     g02826(.A(new_n3072), .B(new_n3077), .Y(new_n3083));
  A2O1A1Ixp33_ASAP7_75t_L   g02827(.A1(new_n2874), .A2(new_n2883), .B(new_n2873), .C(new_n3071), .Y(new_n3084));
  INVx1_ASAP7_75t_L         g02828(.A(new_n3081), .Y(new_n3085));
  NAND3xp33_ASAP7_75t_L     g02829(.A(new_n3084), .B(new_n3083), .C(new_n3085), .Y(new_n3086));
  AOI21xp33_ASAP7_75t_L     g02830(.A1(new_n2884), .A2(new_n2885), .B(new_n2882), .Y(new_n3087));
  OAI21xp33_ASAP7_75t_L     g02831(.A1(new_n3087), .A2(new_n2890), .B(new_n2886), .Y(new_n3088));
  NAND3xp33_ASAP7_75t_L     g02832(.A(new_n3088), .B(new_n3086), .C(new_n3082), .Y(new_n3089));
  AOI21xp33_ASAP7_75t_L     g02833(.A1(new_n3084), .A2(new_n3083), .B(new_n3085), .Y(new_n3090));
  NOR3xp33_ASAP7_75t_L      g02834(.A(new_n3078), .B(new_n3074), .C(new_n3081), .Y(new_n3091));
  NOR3xp33_ASAP7_75t_L      g02835(.A(new_n2876), .B(new_n2835), .C(new_n2878), .Y(new_n3092));
  A2O1A1O1Ixp25_ASAP7_75t_L g02836(.A1(new_n2771), .A2(new_n2714), .B(new_n2827), .C(new_n2879), .D(new_n3092), .Y(new_n3093));
  OAI21xp33_ASAP7_75t_L     g02837(.A1(new_n3090), .A2(new_n3091), .B(new_n3093), .Y(new_n3094));
  AOI22xp33_ASAP7_75t_L     g02838(.A1(new_n1076), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1253), .Y(new_n3095));
  OAI221xp5_ASAP7_75t_L     g02839(.A1(new_n1154), .A2(new_n942), .B1(new_n1156), .B2(new_n1035), .C(new_n3095), .Y(new_n3096));
  XNOR2x2_ASAP7_75t_L       g02840(.A(\a[17] ), .B(new_n3096), .Y(new_n3097));
  NAND3xp33_ASAP7_75t_L     g02841(.A(new_n3089), .B(new_n3094), .C(new_n3097), .Y(new_n3098));
  NOR3xp33_ASAP7_75t_L      g02842(.A(new_n3093), .B(new_n3091), .C(new_n3090), .Y(new_n3099));
  AOI21xp33_ASAP7_75t_L     g02843(.A1(new_n3086), .A2(new_n3082), .B(new_n3088), .Y(new_n3100));
  NOR2xp33_ASAP7_75t_L      g02844(.A(new_n1071), .B(new_n3096), .Y(new_n3101));
  AND2x2_ASAP7_75t_L        g02845(.A(new_n1071), .B(new_n3096), .Y(new_n3102));
  OAI22xp33_ASAP7_75t_L     g02846(.A1(new_n3100), .A2(new_n3099), .B1(new_n3102), .B2(new_n3101), .Y(new_n3103));
  NAND3xp33_ASAP7_75t_L     g02847(.A(new_n2899), .B(new_n2892), .C(new_n2887), .Y(new_n3104));
  NAND4xp25_ASAP7_75t_L     g02848(.A(new_n2906), .B(new_n3104), .C(new_n3103), .D(new_n3098), .Y(new_n3105));
  NOR2xp33_ASAP7_75t_L      g02849(.A(new_n2898), .B(new_n2897), .Y(new_n3106));
  NAND2xp33_ASAP7_75t_L     g02850(.A(new_n3098), .B(new_n3103), .Y(new_n3107));
  A2O1A1Ixp33_ASAP7_75t_L   g02851(.A1(new_n2899), .A2(new_n3106), .B(new_n2912), .C(new_n3107), .Y(new_n3108));
  AOI22xp33_ASAP7_75t_L     g02852(.A1(new_n811), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n900), .Y(new_n3109));
  OAI221xp5_ASAP7_75t_L     g02853(.A1(new_n904), .A2(new_n1313), .B1(new_n898), .B2(new_n1438), .C(new_n3109), .Y(new_n3110));
  XNOR2x2_ASAP7_75t_L       g02854(.A(\a[14] ), .B(new_n3110), .Y(new_n3111));
  NAND3xp33_ASAP7_75t_L     g02855(.A(new_n3105), .B(new_n3108), .C(new_n3111), .Y(new_n3112));
  A2O1A1Ixp33_ASAP7_75t_L   g02856(.A1(new_n2900), .A2(new_n2896), .B(new_n2903), .C(new_n3104), .Y(new_n3113));
  NOR2xp33_ASAP7_75t_L      g02857(.A(new_n3107), .B(new_n3113), .Y(new_n3114));
  AOI22xp33_ASAP7_75t_L     g02858(.A1(new_n3098), .A2(new_n3103), .B1(new_n3104), .B2(new_n2906), .Y(new_n3115));
  INVx1_ASAP7_75t_L         g02859(.A(new_n3111), .Y(new_n3116));
  OAI21xp33_ASAP7_75t_L     g02860(.A1(new_n3114), .A2(new_n3115), .B(new_n3116), .Y(new_n3117));
  NOR3xp33_ASAP7_75t_L      g02861(.A(new_n2911), .B(new_n2912), .C(new_n2909), .Y(new_n3118));
  O2A1O1Ixp33_ASAP7_75t_L   g02862(.A1(new_n2919), .A2(new_n2920), .B(new_n2917), .C(new_n3118), .Y(new_n3119));
  NAND3xp33_ASAP7_75t_L     g02863(.A(new_n3119), .B(new_n3117), .C(new_n3112), .Y(new_n3120));
  NAND2xp33_ASAP7_75t_L     g02864(.A(new_n3112), .B(new_n3117), .Y(new_n3121));
  A2O1A1Ixp33_ASAP7_75t_L   g02865(.A1(new_n2915), .A2(new_n2917), .B(new_n3118), .C(new_n3121), .Y(new_n3122));
  AOI22xp33_ASAP7_75t_L     g02866(.A1(\b[20] ), .A2(new_n651), .B1(\b[22] ), .B2(new_n581), .Y(new_n3123));
  OAI221xp5_ASAP7_75t_L     g02867(.A1(new_n821), .A2(new_n1655), .B1(new_n577), .B2(new_n1780), .C(new_n3123), .Y(new_n3124));
  XNOR2x2_ASAP7_75t_L       g02868(.A(\a[11] ), .B(new_n3124), .Y(new_n3125));
  NAND3xp33_ASAP7_75t_L     g02869(.A(new_n3122), .B(new_n3125), .C(new_n3120), .Y(new_n3126));
  INVx1_ASAP7_75t_L         g02870(.A(new_n3118), .Y(new_n3127));
  A2O1A1Ixp33_ASAP7_75t_L   g02871(.A1(new_n2914), .A2(new_n2910), .B(new_n2927), .C(new_n3127), .Y(new_n3128));
  NOR2xp33_ASAP7_75t_L      g02872(.A(new_n3121), .B(new_n3128), .Y(new_n3129));
  AOI21xp33_ASAP7_75t_L     g02873(.A1(new_n3117), .A2(new_n3112), .B(new_n3119), .Y(new_n3130));
  INVx1_ASAP7_75t_L         g02874(.A(new_n3125), .Y(new_n3131));
  OAI21xp33_ASAP7_75t_L     g02875(.A1(new_n3130), .A2(new_n3129), .B(new_n3131), .Y(new_n3132));
  NOR3xp33_ASAP7_75t_L      g02876(.A(new_n2921), .B(new_n2930), .C(new_n2918), .Y(new_n3133));
  INVx1_ASAP7_75t_L         g02877(.A(new_n3133), .Y(new_n3134));
  INVx1_ASAP7_75t_L         g02878(.A(new_n2801), .Y(new_n3135));
  NOR2xp33_ASAP7_75t_L      g02879(.A(new_n2620), .B(new_n2629), .Y(new_n3136));
  MAJx2_ASAP7_75t_L         g02880(.A(new_n2458), .B(new_n2455), .C(new_n2630), .Y(new_n3137));
  OAI211xp5_ASAP7_75t_L     g02881(.A1(new_n3137), .A2(new_n3136), .B(new_n2933), .C(new_n2932), .Y(new_n3138));
  OAI211xp5_ASAP7_75t_L     g02882(.A1(new_n2925), .A2(new_n2931), .B(new_n3138), .C(new_n3135), .Y(new_n3139));
  NAND4xp25_ASAP7_75t_L     g02883(.A(new_n3139), .B(new_n3126), .C(new_n3132), .D(new_n3134), .Y(new_n3140));
  NOR3xp33_ASAP7_75t_L      g02884(.A(new_n3129), .B(new_n3131), .C(new_n3130), .Y(new_n3141));
  AOI21xp33_ASAP7_75t_L     g02885(.A1(new_n3122), .A2(new_n3120), .B(new_n3125), .Y(new_n3142));
  AOI221xp5_ASAP7_75t_L     g02886(.A1(new_n2933), .A2(new_n2712), .B1(new_n2937), .B2(new_n2936), .C(new_n2801), .Y(new_n3143));
  OAI22xp33_ASAP7_75t_L     g02887(.A1(new_n3143), .A2(new_n3133), .B1(new_n3142), .B2(new_n3141), .Y(new_n3144));
  AOI22xp33_ASAP7_75t_L     g02888(.A1(new_n444), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n471), .Y(new_n3145));
  INVx1_ASAP7_75t_L         g02889(.A(new_n3145), .Y(new_n3146));
  AOI221xp5_ASAP7_75t_L     g02890(.A1(\b[24] ), .A2(new_n447), .B1(new_n441), .B2(new_n2648), .C(new_n3146), .Y(new_n3147));
  XNOR2x2_ASAP7_75t_L       g02891(.A(new_n435), .B(new_n3147), .Y(new_n3148));
  NAND3xp33_ASAP7_75t_L     g02892(.A(new_n3148), .B(new_n3144), .C(new_n3140), .Y(new_n3149));
  NAND2xp33_ASAP7_75t_L     g02893(.A(new_n3126), .B(new_n3132), .Y(new_n3150));
  A2O1A1Ixp33_ASAP7_75t_L   g02894(.A1(new_n2937), .A2(new_n2936), .B(new_n2934), .C(new_n3134), .Y(new_n3151));
  NOR2xp33_ASAP7_75t_L      g02895(.A(new_n3151), .B(new_n3150), .Y(new_n3152));
  AOI22xp33_ASAP7_75t_L     g02896(.A1(new_n3126), .A2(new_n3132), .B1(new_n3134), .B2(new_n3139), .Y(new_n3153));
  INVx1_ASAP7_75t_L         g02897(.A(new_n3148), .Y(new_n3154));
  OAI21xp33_ASAP7_75t_L     g02898(.A1(new_n3153), .A2(new_n3152), .B(new_n3154), .Y(new_n3155));
  A2O1A1O1Ixp25_ASAP7_75t_L g02899(.A1(new_n2808), .A2(new_n2706), .B(new_n2811), .C(new_n2950), .D(new_n2953), .Y(new_n3156));
  AND3x1_ASAP7_75t_L        g02900(.A(new_n3155), .B(new_n3156), .C(new_n3149), .Y(new_n3157));
  AOI21xp33_ASAP7_75t_L     g02901(.A1(new_n3155), .A2(new_n3149), .B(new_n3156), .Y(new_n3158));
  NOR2xp33_ASAP7_75t_L      g02902(.A(new_n2497), .B(new_n429), .Y(new_n3159));
  AOI22xp33_ASAP7_75t_L     g02903(.A1(new_n344), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n370), .Y(new_n3160));
  OAI21xp33_ASAP7_75t_L     g02904(.A1(new_n366), .A2(new_n2672), .B(new_n3160), .Y(new_n3161));
  OR3x1_ASAP7_75t_L         g02905(.A(new_n3161), .B(new_n338), .C(new_n3159), .Y(new_n3162));
  A2O1A1Ixp33_ASAP7_75t_L   g02906(.A1(\b[27] ), .A2(new_n347), .B(new_n3161), .C(new_n338), .Y(new_n3163));
  NAND2xp33_ASAP7_75t_L     g02907(.A(new_n3163), .B(new_n3162), .Y(new_n3164));
  NOR3xp33_ASAP7_75t_L      g02908(.A(new_n3157), .B(new_n3158), .C(new_n3164), .Y(new_n3165));
  NAND3xp33_ASAP7_75t_L     g02909(.A(new_n3155), .B(new_n3156), .C(new_n3149), .Y(new_n3166));
  AO21x2_ASAP7_75t_L        g02910(.A1(new_n3149), .A2(new_n3155), .B(new_n3156), .Y(new_n3167));
  AND2x2_ASAP7_75t_L        g02911(.A(new_n3163), .B(new_n3162), .Y(new_n3168));
  AOI21xp33_ASAP7_75t_L     g02912(.A1(new_n3167), .A2(new_n3166), .B(new_n3168), .Y(new_n3169));
  NOR2xp33_ASAP7_75t_L      g02913(.A(new_n3169), .B(new_n3165), .Y(new_n3170));
  NOR3xp33_ASAP7_75t_L      g02914(.A(new_n2955), .B(new_n2951), .C(new_n2961), .Y(new_n3171));
  INVx1_ASAP7_75t_L         g02915(.A(new_n3171), .Y(new_n3172));
  OAI211xp5_ASAP7_75t_L     g02916(.A1(new_n2969), .A2(new_n2965), .B(new_n3170), .C(new_n3172), .Y(new_n3173));
  A2O1A1Ixp33_ASAP7_75t_L   g02917(.A1(new_n2663), .A2(new_n2702), .B(new_n2816), .C(new_n2967), .Y(new_n3174));
  NAND3xp33_ASAP7_75t_L     g02918(.A(new_n3167), .B(new_n3166), .C(new_n3168), .Y(new_n3175));
  OAI21xp33_ASAP7_75t_L     g02919(.A1(new_n3158), .A2(new_n3157), .B(new_n3164), .Y(new_n3176));
  NAND2xp33_ASAP7_75t_L     g02920(.A(new_n3175), .B(new_n3176), .Y(new_n3177));
  A2O1A1Ixp33_ASAP7_75t_L   g02921(.A1(new_n2977), .A2(new_n3174), .B(new_n3171), .C(new_n3177), .Y(new_n3178));
  NOR2xp33_ASAP7_75t_L      g02922(.A(\b[30] ), .B(\b[31] ), .Y(new_n3179));
  INVx1_ASAP7_75t_L         g02923(.A(\b[31] ), .Y(new_n3180));
  NOR2xp33_ASAP7_75t_L      g02924(.A(new_n2982), .B(new_n3180), .Y(new_n3181));
  NOR2xp33_ASAP7_75t_L      g02925(.A(new_n3179), .B(new_n3181), .Y(new_n3182));
  A2O1A1Ixp33_ASAP7_75t_L   g02926(.A1(\b[30] ), .A2(\b[29] ), .B(new_n2986), .C(new_n3182), .Y(new_n3183));
  O2A1O1Ixp33_ASAP7_75t_L   g02927(.A1(new_n2689), .A2(new_n2987), .B(new_n2984), .C(new_n2983), .Y(new_n3184));
  INVx1_ASAP7_75t_L         g02928(.A(new_n3182), .Y(new_n3185));
  NAND2xp33_ASAP7_75t_L     g02929(.A(new_n3185), .B(new_n3184), .Y(new_n3186));
  NAND2xp33_ASAP7_75t_L     g02930(.A(new_n3183), .B(new_n3186), .Y(new_n3187));
  AOI22xp33_ASAP7_75t_L     g02931(.A1(\b[29] ), .A2(new_n282), .B1(\b[31] ), .B2(new_n303), .Y(new_n3188));
  OAI221xp5_ASAP7_75t_L     g02932(.A1(new_n291), .A2(new_n2982), .B1(new_n268), .B2(new_n3187), .C(new_n3188), .Y(new_n3189));
  XNOR2x2_ASAP7_75t_L       g02933(.A(\a[2] ), .B(new_n3189), .Y(new_n3190));
  NAND3xp33_ASAP7_75t_L     g02934(.A(new_n3173), .B(new_n3178), .C(new_n3190), .Y(new_n3191));
  AOI211xp5_ASAP7_75t_L     g02935(.A1(new_n3174), .A2(new_n2977), .B(new_n3171), .C(new_n3177), .Y(new_n3192));
  O2A1O1Ixp33_ASAP7_75t_L   g02936(.A1(new_n2969), .A2(new_n2965), .B(new_n3172), .C(new_n3170), .Y(new_n3193));
  INVx1_ASAP7_75t_L         g02937(.A(new_n3190), .Y(new_n3194));
  OAI21xp33_ASAP7_75t_L     g02938(.A1(new_n3193), .A2(new_n3192), .B(new_n3194), .Y(new_n3195));
  NAND2xp33_ASAP7_75t_L     g02939(.A(new_n3191), .B(new_n3195), .Y(new_n3196));
  MAJIxp5_ASAP7_75t_L       g02940(.A(new_n2996), .B(new_n2993), .C(new_n2979), .Y(new_n3197));
  XOR2x2_ASAP7_75t_L        g02941(.A(new_n3196), .B(new_n3197), .Y(\f[31] ));
  INVx1_ASAP7_75t_L         g02942(.A(new_n3197), .Y(new_n3199));
  NOR3xp33_ASAP7_75t_L      g02943(.A(new_n3192), .B(new_n3193), .C(new_n3190), .Y(new_n3200));
  INVx1_ASAP7_75t_L         g02944(.A(new_n3200), .Y(new_n3201));
  NOR2xp33_ASAP7_75t_L      g02945(.A(new_n3180), .B(new_n291), .Y(new_n3202));
  INVx1_ASAP7_75t_L         g02946(.A(new_n3202), .Y(new_n3203));
  INVx1_ASAP7_75t_L         g02947(.A(new_n2983), .Y(new_n3204));
  A2O1A1Ixp33_ASAP7_75t_L   g02948(.A1(new_n2691), .A2(new_n2980), .B(new_n2981), .C(new_n3204), .Y(new_n3205));
  NOR2xp33_ASAP7_75t_L      g02949(.A(\b[31] ), .B(\b[32] ), .Y(new_n3206));
  INVx1_ASAP7_75t_L         g02950(.A(\b[32] ), .Y(new_n3207));
  NOR2xp33_ASAP7_75t_L      g02951(.A(new_n3180), .B(new_n3207), .Y(new_n3208));
  NOR2xp33_ASAP7_75t_L      g02952(.A(new_n3206), .B(new_n3208), .Y(new_n3209));
  A2O1A1Ixp33_ASAP7_75t_L   g02953(.A1(new_n3205), .A2(new_n3182), .B(new_n3181), .C(new_n3209), .Y(new_n3210));
  O2A1O1Ixp33_ASAP7_75t_L   g02954(.A1(new_n2983), .A2(new_n2986), .B(new_n3182), .C(new_n3181), .Y(new_n3211));
  INVx1_ASAP7_75t_L         g02955(.A(new_n3209), .Y(new_n3212));
  NAND2xp33_ASAP7_75t_L     g02956(.A(new_n3212), .B(new_n3211), .Y(new_n3213));
  NAND3xp33_ASAP7_75t_L     g02957(.A(new_n3210), .B(new_n267), .C(new_n3213), .Y(new_n3214));
  AOI22xp33_ASAP7_75t_L     g02958(.A1(\b[30] ), .A2(new_n282), .B1(\b[32] ), .B2(new_n303), .Y(new_n3215));
  NAND4xp25_ASAP7_75t_L     g02959(.A(new_n3214), .B(\a[2] ), .C(new_n3203), .D(new_n3215), .Y(new_n3216));
  NAND2xp33_ASAP7_75t_L     g02960(.A(new_n3215), .B(new_n3214), .Y(new_n3217));
  A2O1A1Ixp33_ASAP7_75t_L   g02961(.A1(\b[31] ), .A2(new_n272), .B(new_n3217), .C(new_n262), .Y(new_n3218));
  AND2x2_ASAP7_75t_L        g02962(.A(new_n3216), .B(new_n3218), .Y(new_n3219));
  A2O1A1Ixp33_ASAP7_75t_L   g02963(.A1(new_n2660), .A2(new_n2657), .B(new_n2701), .C(new_n2820), .Y(new_n3220));
  A2O1A1Ixp33_ASAP7_75t_L   g02964(.A1(new_n3220), .A2(new_n2967), .B(new_n2965), .C(new_n3172), .Y(new_n3221));
  NAND2xp33_ASAP7_75t_L     g02965(.A(new_n3166), .B(new_n3167), .Y(new_n3222));
  NOR2xp33_ASAP7_75t_L      g02966(.A(new_n3168), .B(new_n3222), .Y(new_n3223));
  NAND3xp33_ASAP7_75t_L     g02967(.A(new_n3122), .B(new_n3120), .C(new_n3131), .Y(new_n3224));
  AOI22xp33_ASAP7_75t_L     g02968(.A1(\b[21] ), .A2(new_n651), .B1(\b[23] ), .B2(new_n581), .Y(new_n3225));
  OAI221xp5_ASAP7_75t_L     g02969(.A1(new_n821), .A2(new_n1774), .B1(new_n577), .B2(new_n1915), .C(new_n3225), .Y(new_n3226));
  XNOR2x2_ASAP7_75t_L       g02970(.A(\a[11] ), .B(new_n3226), .Y(new_n3227));
  INVx1_ASAP7_75t_L         g02971(.A(new_n3227), .Y(new_n3228));
  NAND2xp33_ASAP7_75t_L     g02972(.A(new_n3108), .B(new_n3105), .Y(new_n3229));
  NOR2xp33_ASAP7_75t_L      g02973(.A(new_n3111), .B(new_n3229), .Y(new_n3230));
  O2A1O1Ixp33_ASAP7_75t_L   g02974(.A1(new_n3118), .A2(new_n2921), .B(new_n3121), .C(new_n3230), .Y(new_n3231));
  AOI22xp33_ASAP7_75t_L     g02975(.A1(new_n1360), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1581), .Y(new_n3232));
  OAI221xp5_ASAP7_75t_L     g02976(.A1(new_n1373), .A2(new_n784), .B1(new_n1359), .B2(new_n875), .C(new_n3232), .Y(new_n3233));
  XNOR2x2_ASAP7_75t_L       g02977(.A(new_n1356), .B(new_n3233), .Y(new_n3234));
  NAND3xp33_ASAP7_75t_L     g02978(.A(new_n3049), .B(new_n3053), .C(new_n3069), .Y(new_n3235));
  A2O1A1O1Ixp25_ASAP7_75t_L g02979(.A1(new_n2864), .A2(new_n2866), .B(new_n3000), .C(new_n3067), .D(new_n3042), .Y(new_n3236));
  AOI22xp33_ASAP7_75t_L     g02980(.A1(new_n2114), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n2259), .Y(new_n3237));
  OAI221xp5_ASAP7_75t_L     g02981(.A1(new_n2109), .A2(new_n420), .B1(new_n2257), .B2(new_n494), .C(new_n3237), .Y(new_n3238));
  XNOR2x2_ASAP7_75t_L       g02982(.A(\a[26] ), .B(new_n3238), .Y(new_n3239));
  NOR2xp33_ASAP7_75t_L      g02983(.A(new_n2837), .B(new_n2738), .Y(new_n3240));
  NAND2xp33_ASAP7_75t_L     g02984(.A(new_n2853), .B(new_n2851), .Y(new_n3241));
  MAJIxp5_ASAP7_75t_L       g02985(.A(new_n3241), .B(new_n2843), .C(new_n3240), .Y(new_n3242));
  NOR2xp33_ASAP7_75t_L      g02986(.A(new_n3035), .B(new_n3014), .Y(new_n3243));
  INVx1_ASAP7_75t_L         g02987(.A(new_n3243), .Y(new_n3244));
  A2O1A1Ixp33_ASAP7_75t_L   g02988(.A1(new_n3034), .A2(new_n3036), .B(new_n3242), .C(new_n3244), .Y(new_n3245));
  NAND2xp33_ASAP7_75t_L     g02989(.A(\b[4] ), .B(new_n2553), .Y(new_n3246));
  INVx1_ASAP7_75t_L         g02990(.A(new_n3246), .Y(new_n3247));
  NOR3xp33_ASAP7_75t_L      g02991(.A(new_n357), .B(new_n358), .C(new_n2734), .Y(new_n3248));
  OAI22xp33_ASAP7_75t_L     g02992(.A1(new_n2747), .A2(new_n298), .B1(new_n354), .B2(new_n2545), .Y(new_n3249));
  NOR4xp25_ASAP7_75t_L      g02993(.A(new_n3248), .B(new_n2538), .C(new_n3249), .D(new_n3247), .Y(new_n3250));
  INVx1_ASAP7_75t_L         g02994(.A(new_n3250), .Y(new_n3251));
  OAI31xp33_ASAP7_75t_L     g02995(.A1(new_n3248), .A2(new_n3247), .A3(new_n3249), .B(new_n2538), .Y(new_n3252));
  NAND2xp33_ASAP7_75t_L     g02996(.A(new_n3027), .B(new_n3031), .Y(new_n3253));
  NOR2xp33_ASAP7_75t_L      g02997(.A(new_n261), .B(new_n3024), .Y(new_n3254));
  INVx1_ASAP7_75t_L         g02998(.A(new_n3254), .Y(new_n3255));
  NAND2xp33_ASAP7_75t_L     g02999(.A(new_n3028), .B(new_n2841), .Y(new_n3256));
  NOR2xp33_ASAP7_75t_L      g03000(.A(new_n280), .B(new_n3256), .Y(new_n3257));
  AND3x1_ASAP7_75t_L        g03001(.A(new_n3017), .B(new_n3023), .C(new_n3028), .Y(new_n3258));
  AOI221xp5_ASAP7_75t_L     g03002(.A1(new_n3029), .A2(\b[2] ), .B1(new_n3258), .B2(\b[0] ), .C(new_n3257), .Y(new_n3259));
  NAND2xp33_ASAP7_75t_L     g03003(.A(new_n3255), .B(new_n3259), .Y(new_n3260));
  O2A1O1Ixp33_ASAP7_75t_L   g03004(.A1(new_n2843), .A2(new_n3253), .B(\a[32] ), .C(new_n3260), .Y(new_n3261));
  A2O1A1Ixp33_ASAP7_75t_L   g03005(.A1(\b[0] ), .A2(new_n2841), .B(new_n3253), .C(\a[32] ), .Y(new_n3262));
  O2A1O1Ixp33_ASAP7_75t_L   g03006(.A1(new_n3024), .A2(new_n261), .B(new_n3259), .C(new_n3262), .Y(new_n3263));
  OAI211xp5_ASAP7_75t_L     g03007(.A1(new_n3261), .A2(new_n3263), .B(new_n3252), .C(new_n3251), .Y(new_n3264));
  AO211x2_ASAP7_75t_L       g03008(.A1(new_n3252), .A2(new_n3251), .B(new_n3261), .C(new_n3263), .Y(new_n3265));
  AOI21xp33_ASAP7_75t_L     g03009(.A1(new_n3265), .A2(new_n3264), .B(new_n3245), .Y(new_n3266));
  NAND2xp33_ASAP7_75t_L     g03010(.A(new_n3264), .B(new_n3265), .Y(new_n3267));
  O2A1O1Ixp33_ASAP7_75t_L   g03011(.A1(new_n3014), .A2(new_n3035), .B(new_n3045), .C(new_n3267), .Y(new_n3268));
  NOR3xp33_ASAP7_75t_L      g03012(.A(new_n3268), .B(new_n3266), .C(new_n3239), .Y(new_n3269));
  XNOR2x2_ASAP7_75t_L       g03013(.A(new_n2100), .B(new_n3238), .Y(new_n3270));
  NAND2xp33_ASAP7_75t_L     g03014(.A(new_n3036), .B(new_n3034), .Y(new_n3271));
  O2A1O1Ixp33_ASAP7_75t_L   g03015(.A1(new_n3038), .A2(new_n3007), .B(new_n3271), .C(new_n3243), .Y(new_n3272));
  NAND2xp33_ASAP7_75t_L     g03016(.A(new_n3267), .B(new_n3272), .Y(new_n3273));
  NAND3xp33_ASAP7_75t_L     g03017(.A(new_n3245), .B(new_n3264), .C(new_n3265), .Y(new_n3274));
  AOI21xp33_ASAP7_75t_L     g03018(.A1(new_n3273), .A2(new_n3274), .B(new_n3270), .Y(new_n3275));
  OAI21xp33_ASAP7_75t_L     g03019(.A1(new_n3275), .A2(new_n3269), .B(new_n3236), .Y(new_n3276));
  A2O1A1Ixp33_ASAP7_75t_L   g03020(.A1(new_n3064), .A2(new_n3063), .B(new_n3047), .C(new_n3066), .Y(new_n3277));
  NAND3xp33_ASAP7_75t_L     g03021(.A(new_n3273), .B(new_n3274), .C(new_n3270), .Y(new_n3278));
  OAI21xp33_ASAP7_75t_L     g03022(.A1(new_n3266), .A2(new_n3268), .B(new_n3239), .Y(new_n3279));
  NAND3xp33_ASAP7_75t_L     g03023(.A(new_n3277), .B(new_n3278), .C(new_n3279), .Y(new_n3280));
  AOI22xp33_ASAP7_75t_L     g03024(.A1(new_n1704), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1837), .Y(new_n3281));
  OAI221xp5_ASAP7_75t_L     g03025(.A1(new_n1699), .A2(new_n617), .B1(new_n1827), .B2(new_n685), .C(new_n3281), .Y(new_n3282));
  XNOR2x2_ASAP7_75t_L       g03026(.A(new_n1689), .B(new_n3282), .Y(new_n3283));
  AOI21xp33_ASAP7_75t_L     g03027(.A1(new_n3280), .A2(new_n3276), .B(new_n3283), .Y(new_n3284));
  AOI21xp33_ASAP7_75t_L     g03028(.A1(new_n3279), .A2(new_n3278), .B(new_n3277), .Y(new_n3285));
  NOR3xp33_ASAP7_75t_L      g03029(.A(new_n3236), .B(new_n3269), .C(new_n3275), .Y(new_n3286));
  XNOR2x2_ASAP7_75t_L       g03030(.A(\a[23] ), .B(new_n3282), .Y(new_n3287));
  NOR3xp33_ASAP7_75t_L      g03031(.A(new_n3285), .B(new_n3287), .C(new_n3286), .Y(new_n3288));
  OAI221xp5_ASAP7_75t_L     g03032(.A1(new_n3288), .A2(new_n3284), .B1(new_n3072), .B2(new_n3077), .C(new_n3235), .Y(new_n3289));
  A2O1A1Ixp33_ASAP7_75t_L   g03033(.A1(new_n3070), .A2(new_n3062), .B(new_n3072), .C(new_n3235), .Y(new_n3290));
  OAI21xp33_ASAP7_75t_L     g03034(.A1(new_n3286), .A2(new_n3285), .B(new_n3287), .Y(new_n3291));
  NAND3xp33_ASAP7_75t_L     g03035(.A(new_n3280), .B(new_n3283), .C(new_n3276), .Y(new_n3292));
  NAND3xp33_ASAP7_75t_L     g03036(.A(new_n3290), .B(new_n3291), .C(new_n3292), .Y(new_n3293));
  AOI21xp33_ASAP7_75t_L     g03037(.A1(new_n3293), .A2(new_n3289), .B(new_n3234), .Y(new_n3294));
  AND3x1_ASAP7_75t_L        g03038(.A(new_n3293), .B(new_n3289), .C(new_n3234), .Y(new_n3295));
  NOR2xp33_ASAP7_75t_L      g03039(.A(new_n3294), .B(new_n3295), .Y(new_n3296));
  A2O1A1Ixp33_ASAP7_75t_L   g03040(.A1(new_n3088), .A2(new_n3082), .B(new_n3091), .C(new_n3296), .Y(new_n3297));
  A2O1A1O1Ixp25_ASAP7_75t_L g03041(.A1(new_n2879), .A2(new_n2828), .B(new_n3092), .C(new_n3082), .D(new_n3091), .Y(new_n3298));
  AO21x2_ASAP7_75t_L        g03042(.A1(new_n3289), .A2(new_n3293), .B(new_n3234), .Y(new_n3299));
  NAND3xp33_ASAP7_75t_L     g03043(.A(new_n3293), .B(new_n3289), .C(new_n3234), .Y(new_n3300));
  NAND2xp33_ASAP7_75t_L     g03044(.A(new_n3300), .B(new_n3299), .Y(new_n3301));
  NAND2xp33_ASAP7_75t_L     g03045(.A(new_n3298), .B(new_n3301), .Y(new_n3302));
  NOR2xp33_ASAP7_75t_L      g03046(.A(new_n1030), .B(new_n1154), .Y(new_n3303));
  INVx1_ASAP7_75t_L         g03047(.A(new_n3303), .Y(new_n3304));
  NOR2xp33_ASAP7_75t_L      g03048(.A(new_n1205), .B(new_n1796), .Y(new_n3305));
  NAND2xp33_ASAP7_75t_L     g03049(.A(new_n1073), .B(new_n3305), .Y(new_n3306));
  AOI22xp33_ASAP7_75t_L     g03050(.A1(new_n1076), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1253), .Y(new_n3307));
  NAND4xp25_ASAP7_75t_L     g03051(.A(new_n3306), .B(\a[17] ), .C(new_n3304), .D(new_n3307), .Y(new_n3308));
  OAI21xp33_ASAP7_75t_L     g03052(.A1(new_n1156), .A2(new_n1209), .B(new_n3307), .Y(new_n3309));
  A2O1A1Ixp33_ASAP7_75t_L   g03053(.A1(\b[16] ), .A2(new_n1080), .B(new_n3309), .C(new_n1071), .Y(new_n3310));
  AND2x2_ASAP7_75t_L        g03054(.A(new_n3308), .B(new_n3310), .Y(new_n3311));
  NAND3xp33_ASAP7_75t_L     g03055(.A(new_n3311), .B(new_n3297), .C(new_n3302), .Y(new_n3312));
  O2A1O1Ixp33_ASAP7_75t_L   g03056(.A1(new_n3090), .A2(new_n3093), .B(new_n3086), .C(new_n3301), .Y(new_n3313));
  AOI211xp5_ASAP7_75t_L     g03057(.A1(new_n3300), .A2(new_n3299), .B(new_n3091), .C(new_n3099), .Y(new_n3314));
  NAND2xp33_ASAP7_75t_L     g03058(.A(new_n3308), .B(new_n3310), .Y(new_n3315));
  OAI21xp33_ASAP7_75t_L     g03059(.A1(new_n3314), .A2(new_n3313), .B(new_n3315), .Y(new_n3316));
  NAND2xp33_ASAP7_75t_L     g03060(.A(new_n3316), .B(new_n3312), .Y(new_n3317));
  NOR3xp33_ASAP7_75t_L      g03061(.A(new_n3100), .B(new_n3097), .C(new_n3099), .Y(new_n3318));
  AO21x2_ASAP7_75t_L        g03062(.A1(new_n3107), .A2(new_n3113), .B(new_n3318), .Y(new_n3319));
  NOR2xp33_ASAP7_75t_L      g03063(.A(new_n3317), .B(new_n3319), .Y(new_n3320));
  NOR3xp33_ASAP7_75t_L      g03064(.A(new_n3313), .B(new_n3315), .C(new_n3314), .Y(new_n3321));
  AOI21xp33_ASAP7_75t_L     g03065(.A1(new_n3297), .A2(new_n3302), .B(new_n3311), .Y(new_n3322));
  NOR2xp33_ASAP7_75t_L      g03066(.A(new_n3321), .B(new_n3322), .Y(new_n3323));
  A2O1A1O1Ixp25_ASAP7_75t_L g03067(.A1(new_n2899), .A2(new_n3106), .B(new_n2912), .C(new_n3107), .D(new_n3318), .Y(new_n3324));
  NOR2xp33_ASAP7_75t_L      g03068(.A(new_n3323), .B(new_n3324), .Y(new_n3325));
  AOI22xp33_ASAP7_75t_L     g03069(.A1(new_n811), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n900), .Y(new_n3326));
  OAI221xp5_ASAP7_75t_L     g03070(.A1(new_n904), .A2(new_n1432), .B1(new_n898), .B2(new_n1547), .C(new_n3326), .Y(new_n3327));
  XNOR2x2_ASAP7_75t_L       g03071(.A(\a[14] ), .B(new_n3327), .Y(new_n3328));
  OAI21xp33_ASAP7_75t_L     g03072(.A1(new_n3325), .A2(new_n3320), .B(new_n3328), .Y(new_n3329));
  NAND2xp33_ASAP7_75t_L     g03073(.A(new_n3323), .B(new_n3324), .Y(new_n3330));
  A2O1A1Ixp33_ASAP7_75t_L   g03074(.A1(new_n3107), .A2(new_n3113), .B(new_n3318), .C(new_n3317), .Y(new_n3331));
  XNOR2x2_ASAP7_75t_L       g03075(.A(new_n806), .B(new_n3327), .Y(new_n3332));
  NAND3xp33_ASAP7_75t_L     g03076(.A(new_n3331), .B(new_n3330), .C(new_n3332), .Y(new_n3333));
  NAND2xp33_ASAP7_75t_L     g03077(.A(new_n3333), .B(new_n3329), .Y(new_n3334));
  NAND2xp33_ASAP7_75t_L     g03078(.A(new_n3334), .B(new_n3231), .Y(new_n3335));
  AOI21xp33_ASAP7_75t_L     g03079(.A1(new_n3331), .A2(new_n3330), .B(new_n3332), .Y(new_n3336));
  NOR3xp33_ASAP7_75t_L      g03080(.A(new_n3320), .B(new_n3325), .C(new_n3328), .Y(new_n3337));
  NOR2xp33_ASAP7_75t_L      g03081(.A(new_n3336), .B(new_n3337), .Y(new_n3338));
  A2O1A1Ixp33_ASAP7_75t_L   g03082(.A1(new_n3128), .A2(new_n3121), .B(new_n3230), .C(new_n3338), .Y(new_n3339));
  AOI21xp33_ASAP7_75t_L     g03083(.A1(new_n3339), .A2(new_n3335), .B(new_n3228), .Y(new_n3340));
  MAJIxp5_ASAP7_75t_L       g03084(.A(new_n3119), .B(new_n3229), .C(new_n3111), .Y(new_n3341));
  NOR2xp33_ASAP7_75t_L      g03085(.A(new_n3341), .B(new_n3338), .Y(new_n3342));
  AND2x2_ASAP7_75t_L        g03086(.A(new_n3112), .B(new_n3117), .Y(new_n3343));
  INVx1_ASAP7_75t_L         g03087(.A(new_n3230), .Y(new_n3344));
  O2A1O1Ixp33_ASAP7_75t_L   g03088(.A1(new_n3343), .A2(new_n3119), .B(new_n3344), .C(new_n3334), .Y(new_n3345));
  NOR3xp33_ASAP7_75t_L      g03089(.A(new_n3345), .B(new_n3342), .C(new_n3227), .Y(new_n3346));
  AOI211xp5_ASAP7_75t_L     g03090(.A1(new_n3144), .A2(new_n3224), .B(new_n3340), .C(new_n3346), .Y(new_n3347));
  INVx1_ASAP7_75t_L         g03091(.A(new_n3224), .Y(new_n3348));
  OAI21xp33_ASAP7_75t_L     g03092(.A1(new_n3342), .A2(new_n3345), .B(new_n3227), .Y(new_n3349));
  NAND3xp33_ASAP7_75t_L     g03093(.A(new_n3339), .B(new_n3335), .C(new_n3228), .Y(new_n3350));
  AOI211xp5_ASAP7_75t_L     g03094(.A1(new_n3349), .A2(new_n3350), .B(new_n3348), .C(new_n3153), .Y(new_n3351));
  AOI22xp33_ASAP7_75t_L     g03095(.A1(new_n444), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n471), .Y(new_n3352));
  OAI221xp5_ASAP7_75t_L     g03096(.A1(new_n468), .A2(new_n2067), .B1(new_n469), .B2(new_n2355), .C(new_n3352), .Y(new_n3353));
  XNOR2x2_ASAP7_75t_L       g03097(.A(\a[8] ), .B(new_n3353), .Y(new_n3354));
  INVx1_ASAP7_75t_L         g03098(.A(new_n3354), .Y(new_n3355));
  NOR3xp33_ASAP7_75t_L      g03099(.A(new_n3347), .B(new_n3351), .C(new_n3355), .Y(new_n3356));
  OAI211xp5_ASAP7_75t_L     g03100(.A1(new_n3348), .A2(new_n3153), .B(new_n3349), .C(new_n3350), .Y(new_n3357));
  OAI211xp5_ASAP7_75t_L     g03101(.A1(new_n3346), .A2(new_n3340), .B(new_n3144), .C(new_n3224), .Y(new_n3358));
  AOI21xp33_ASAP7_75t_L     g03102(.A1(new_n3357), .A2(new_n3358), .B(new_n3354), .Y(new_n3359));
  NAND2xp33_ASAP7_75t_L     g03103(.A(new_n3140), .B(new_n3144), .Y(new_n3360));
  MAJIxp5_ASAP7_75t_L       g03104(.A(new_n3156), .B(new_n3360), .C(new_n3148), .Y(new_n3361));
  NOR3xp33_ASAP7_75t_L      g03105(.A(new_n3361), .B(new_n3359), .C(new_n3356), .Y(new_n3362));
  OA21x2_ASAP7_75t_L        g03106(.A1(new_n3356), .A2(new_n3359), .B(new_n3361), .Y(new_n3363));
  AOI22xp33_ASAP7_75t_L     g03107(.A1(new_n344), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n370), .Y(new_n3364));
  OAI221xp5_ASAP7_75t_L     g03108(.A1(new_n429), .A2(new_n2666), .B1(new_n366), .B2(new_n2695), .C(new_n3364), .Y(new_n3365));
  XNOR2x2_ASAP7_75t_L       g03109(.A(\a[5] ), .B(new_n3365), .Y(new_n3366));
  OAI21xp33_ASAP7_75t_L     g03110(.A1(new_n3362), .A2(new_n3363), .B(new_n3366), .Y(new_n3367));
  OR3x1_ASAP7_75t_L         g03111(.A(new_n3361), .B(new_n3356), .C(new_n3359), .Y(new_n3368));
  OAI21xp33_ASAP7_75t_L     g03112(.A1(new_n3359), .A2(new_n3356), .B(new_n3361), .Y(new_n3369));
  INVx1_ASAP7_75t_L         g03113(.A(new_n3366), .Y(new_n3370));
  NAND3xp33_ASAP7_75t_L     g03114(.A(new_n3368), .B(new_n3369), .C(new_n3370), .Y(new_n3371));
  AOI221xp5_ASAP7_75t_L     g03115(.A1(new_n3371), .A2(new_n3367), .B1(new_n3177), .B2(new_n3221), .C(new_n3223), .Y(new_n3372));
  NAND2xp33_ASAP7_75t_L     g03116(.A(new_n3367), .B(new_n3371), .Y(new_n3373));
  O2A1O1Ixp33_ASAP7_75t_L   g03117(.A1(new_n3222), .A2(new_n3168), .B(new_n3178), .C(new_n3373), .Y(new_n3374));
  NOR3xp33_ASAP7_75t_L      g03118(.A(new_n3374), .B(new_n3372), .C(new_n3219), .Y(new_n3375));
  INVx1_ASAP7_75t_L         g03119(.A(new_n3375), .Y(new_n3376));
  OAI21xp33_ASAP7_75t_L     g03120(.A1(new_n3372), .A2(new_n3374), .B(new_n3219), .Y(new_n3377));
  NAND2xp33_ASAP7_75t_L     g03121(.A(new_n3377), .B(new_n3376), .Y(new_n3378));
  A2O1A1O1Ixp25_ASAP7_75t_L g03122(.A1(new_n3195), .A2(new_n3191), .B(new_n3199), .C(new_n3201), .D(new_n3378), .Y(new_n3379));
  A2O1A1Ixp33_ASAP7_75t_L   g03123(.A1(new_n3195), .A2(new_n3191), .B(new_n3199), .C(new_n3201), .Y(new_n3380));
  AOI21xp33_ASAP7_75t_L     g03124(.A1(new_n3377), .A2(new_n3376), .B(new_n3380), .Y(new_n3381));
  NOR2xp33_ASAP7_75t_L      g03125(.A(new_n3381), .B(new_n3379), .Y(\f[32] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03126(.A1(new_n3196), .A2(new_n3197), .B(new_n3200), .C(new_n3377), .D(new_n3375), .Y(new_n3383));
  NAND2xp33_ASAP7_75t_L     g03127(.A(new_n3120), .B(new_n3122), .Y(new_n3384));
  NOR2xp33_ASAP7_75t_L      g03128(.A(new_n2918), .B(new_n2921), .Y(new_n3385));
  MAJIxp5_ASAP7_75t_L       g03129(.A(new_n2938), .B(new_n3385), .C(new_n2924), .Y(new_n3386));
  MAJIxp5_ASAP7_75t_L       g03130(.A(new_n3386), .B(new_n3384), .C(new_n3125), .Y(new_n3387));
  AOI22xp33_ASAP7_75t_L     g03131(.A1(\b[22] ), .A2(new_n651), .B1(\b[24] ), .B2(new_n581), .Y(new_n3388));
  OAI31xp33_ASAP7_75t_L     g03132(.A1(new_n1934), .A2(new_n577), .A3(new_n1933), .B(new_n3388), .Y(new_n3389));
  AOI21xp33_ASAP7_75t_L     g03133(.A1(new_n584), .A2(\b[23] ), .B(new_n3389), .Y(new_n3390));
  NAND2xp33_ASAP7_75t_L     g03134(.A(\a[11] ), .B(new_n3390), .Y(new_n3391));
  A2O1A1Ixp33_ASAP7_75t_L   g03135(.A1(\b[23] ), .A2(new_n584), .B(new_n3389), .C(new_n574), .Y(new_n3392));
  NAND2xp33_ASAP7_75t_L     g03136(.A(new_n3392), .B(new_n3391), .Y(new_n3393));
  NOR3xp33_ASAP7_75t_L      g03137(.A(new_n3311), .B(new_n3313), .C(new_n3314), .Y(new_n3394));
  OAI22xp33_ASAP7_75t_L     g03138(.A1(new_n1158), .A2(new_n1030), .B1(new_n1313), .B2(new_n1259), .Y(new_n3395));
  AOI221xp5_ASAP7_75t_L     g03139(.A1(\b[17] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n1319), .C(new_n3395), .Y(new_n3396));
  XNOR2x2_ASAP7_75t_L       g03140(.A(\a[17] ), .B(new_n3396), .Y(new_n3397));
  OAI21xp33_ASAP7_75t_L     g03141(.A1(new_n3294), .A2(new_n3298), .B(new_n3300), .Y(new_n3398));
  OAI21xp33_ASAP7_75t_L     g03142(.A1(new_n3275), .A2(new_n3236), .B(new_n3278), .Y(new_n3399));
  NAND4xp25_ASAP7_75t_L     g03143(.A(new_n3031), .B(\a[32] ), .C(new_n2842), .D(new_n3027), .Y(new_n3400));
  NAND2xp33_ASAP7_75t_L     g03144(.A(\b[2] ), .B(new_n3029), .Y(new_n3401));
  NAND3xp33_ASAP7_75t_L     g03145(.A(new_n3017), .B(new_n3028), .C(new_n3023), .Y(new_n3402));
  OAI221xp5_ASAP7_75t_L     g03146(.A1(new_n258), .A2(new_n3402), .B1(new_n280), .B2(new_n3256), .C(new_n3401), .Y(new_n3403));
  INVx1_ASAP7_75t_L         g03147(.A(\a[33] ), .Y(new_n3404));
  NAND2xp33_ASAP7_75t_L     g03148(.A(\a[32] ), .B(new_n3404), .Y(new_n3405));
  NAND2xp33_ASAP7_75t_L     g03149(.A(\a[33] ), .B(new_n3015), .Y(new_n3406));
  AND2x2_ASAP7_75t_L        g03150(.A(new_n3405), .B(new_n3406), .Y(new_n3407));
  NOR2xp33_ASAP7_75t_L      g03151(.A(new_n258), .B(new_n3407), .Y(new_n3408));
  OAI31xp33_ASAP7_75t_L     g03152(.A1(new_n3400), .A2(new_n3403), .A3(new_n3254), .B(new_n3408), .Y(new_n3409));
  A2O1A1Ixp33_ASAP7_75t_L   g03153(.A1(new_n2839), .A2(new_n2840), .B(new_n258), .C(\a[32] ), .Y(new_n3410));
  AOI211xp5_ASAP7_75t_L     g03154(.A1(new_n3021), .A2(new_n269), .B(new_n3410), .C(new_n3025), .Y(new_n3411));
  INVx1_ASAP7_75t_L         g03155(.A(new_n3408), .Y(new_n3412));
  NAND4xp25_ASAP7_75t_L     g03156(.A(new_n3411), .B(new_n3412), .C(new_n3259), .D(new_n3255), .Y(new_n3413));
  OAI22xp33_ASAP7_75t_L     g03157(.A1(new_n3402), .A2(new_n261), .B1(new_n298), .B2(new_n3022), .Y(new_n3414));
  AOI221xp5_ASAP7_75t_L     g03158(.A1(\b[2] ), .A2(new_n3030), .B1(new_n406), .B2(new_n3021), .C(new_n3414), .Y(new_n3415));
  NAND2xp33_ASAP7_75t_L     g03159(.A(\a[32] ), .B(new_n3415), .Y(new_n3416));
  NAND2xp33_ASAP7_75t_L     g03160(.A(\b[3] ), .B(new_n3029), .Y(new_n3417));
  OAI221xp5_ASAP7_75t_L     g03161(.A1(new_n3402), .A2(new_n261), .B1(new_n3256), .B2(new_n302), .C(new_n3417), .Y(new_n3418));
  A2O1A1Ixp33_ASAP7_75t_L   g03162(.A1(\b[2] ), .A2(new_n3030), .B(new_n3418), .C(new_n3015), .Y(new_n3419));
  AO22x1_ASAP7_75t_L        g03163(.A1(new_n3419), .A2(new_n3416), .B1(new_n3409), .B2(new_n3413), .Y(new_n3420));
  NAND4xp25_ASAP7_75t_L     g03164(.A(new_n3413), .B(new_n3409), .C(new_n3416), .D(new_n3419), .Y(new_n3421));
  NAND2xp33_ASAP7_75t_L     g03165(.A(\b[5] ), .B(new_n2553), .Y(new_n3422));
  NAND2xp33_ASAP7_75t_L     g03166(.A(new_n2544), .B(new_n526), .Y(new_n3423));
  AOI22xp33_ASAP7_75t_L     g03167(.A1(new_n2552), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n2736), .Y(new_n3424));
  NAND4xp25_ASAP7_75t_L     g03168(.A(new_n3423), .B(\a[29] ), .C(new_n3422), .D(new_n3424), .Y(new_n3425));
  OAI21xp33_ASAP7_75t_L     g03169(.A1(new_n2734), .A2(new_n390), .B(new_n3424), .Y(new_n3426));
  A2O1A1Ixp33_ASAP7_75t_L   g03170(.A1(\b[5] ), .A2(new_n2553), .B(new_n3426), .C(new_n2538), .Y(new_n3427));
  NAND4xp25_ASAP7_75t_L     g03171(.A(new_n3427), .B(new_n3420), .C(new_n3421), .D(new_n3425), .Y(new_n3428));
  AO22x1_ASAP7_75t_L        g03172(.A1(new_n3421), .A2(new_n3420), .B1(new_n3427), .B2(new_n3425), .Y(new_n3429));
  INVx1_ASAP7_75t_L         g03173(.A(new_n3264), .Y(new_n3430));
  AOI31xp33_ASAP7_75t_L     g03174(.A1(new_n3045), .A2(new_n3265), .A3(new_n3244), .B(new_n3430), .Y(new_n3431));
  NAND3xp33_ASAP7_75t_L     g03175(.A(new_n3431), .B(new_n3429), .C(new_n3428), .Y(new_n3432));
  NAND2xp33_ASAP7_75t_L     g03176(.A(new_n3428), .B(new_n3429), .Y(new_n3433));
  A2O1A1Ixp33_ASAP7_75t_L   g03177(.A1(new_n3265), .A2(new_n3272), .B(new_n3430), .C(new_n3433), .Y(new_n3434));
  AOI22xp33_ASAP7_75t_L     g03178(.A1(new_n2114), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n2259), .Y(new_n3435));
  OAI221xp5_ASAP7_75t_L     g03179(.A1(new_n2109), .A2(new_n488), .B1(new_n2257), .B2(new_n548), .C(new_n3435), .Y(new_n3436));
  XNOR2x2_ASAP7_75t_L       g03180(.A(\a[26] ), .B(new_n3436), .Y(new_n3437));
  AO21x2_ASAP7_75t_L        g03181(.A1(new_n3432), .A2(new_n3434), .B(new_n3437), .Y(new_n3438));
  OR2x4_ASAP7_75t_L         g03182(.A(new_n2100), .B(new_n3436), .Y(new_n3439));
  NAND2xp33_ASAP7_75t_L     g03183(.A(new_n2100), .B(new_n3436), .Y(new_n3440));
  NAND4xp25_ASAP7_75t_L     g03184(.A(new_n3434), .B(new_n3432), .C(new_n3439), .D(new_n3440), .Y(new_n3441));
  AOI21xp33_ASAP7_75t_L     g03185(.A1(new_n3441), .A2(new_n3438), .B(new_n3399), .Y(new_n3442));
  A2O1A1Ixp33_ASAP7_75t_L   g03186(.A1(new_n2863), .A2(new_n2862), .B(new_n2867), .C(new_n3063), .Y(new_n3443));
  A2O1A1O1Ixp25_ASAP7_75t_L g03187(.A1(new_n3048), .A2(new_n3443), .B(new_n3042), .C(new_n3279), .D(new_n3269), .Y(new_n3444));
  AOI21xp33_ASAP7_75t_L     g03188(.A1(new_n3434), .A2(new_n3432), .B(new_n3437), .Y(new_n3445));
  AND3x1_ASAP7_75t_L        g03189(.A(new_n3437), .B(new_n3434), .C(new_n3432), .Y(new_n3446));
  NOR3xp33_ASAP7_75t_L      g03190(.A(new_n3444), .B(new_n3445), .C(new_n3446), .Y(new_n3447));
  NAND2xp33_ASAP7_75t_L     g03191(.A(\b[11] ), .B(new_n1706), .Y(new_n3448));
  NAND2xp33_ASAP7_75t_L     g03192(.A(new_n1695), .B(new_n1232), .Y(new_n3449));
  AOI22xp33_ASAP7_75t_L     g03193(.A1(new_n1704), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1837), .Y(new_n3450));
  NAND4xp25_ASAP7_75t_L     g03194(.A(new_n3449), .B(\a[23] ), .C(new_n3448), .D(new_n3450), .Y(new_n3451));
  OAI21xp33_ASAP7_75t_L     g03195(.A1(new_n1827), .A2(new_n768), .B(new_n3450), .Y(new_n3452));
  A2O1A1Ixp33_ASAP7_75t_L   g03196(.A1(\b[11] ), .A2(new_n1706), .B(new_n3452), .C(new_n1689), .Y(new_n3453));
  AND2x2_ASAP7_75t_L        g03197(.A(new_n3451), .B(new_n3453), .Y(new_n3454));
  OAI21xp33_ASAP7_75t_L     g03198(.A1(new_n3442), .A2(new_n3447), .B(new_n3454), .Y(new_n3455));
  OAI21xp33_ASAP7_75t_L     g03199(.A1(new_n3445), .A2(new_n3446), .B(new_n3444), .Y(new_n3456));
  NAND3xp33_ASAP7_75t_L     g03200(.A(new_n3399), .B(new_n3438), .C(new_n3441), .Y(new_n3457));
  NAND2xp33_ASAP7_75t_L     g03201(.A(new_n3451), .B(new_n3453), .Y(new_n3458));
  NAND3xp33_ASAP7_75t_L     g03202(.A(new_n3458), .B(new_n3457), .C(new_n3456), .Y(new_n3459));
  OAI211xp5_ASAP7_75t_L     g03203(.A1(new_n3072), .A2(new_n3077), .B(new_n3235), .C(new_n3292), .Y(new_n3460));
  NAND4xp25_ASAP7_75t_L     g03204(.A(new_n3460), .B(new_n3291), .C(new_n3455), .D(new_n3459), .Y(new_n3461));
  AOI21xp33_ASAP7_75t_L     g03205(.A1(new_n3457), .A2(new_n3456), .B(new_n3458), .Y(new_n3462));
  NOR3xp33_ASAP7_75t_L      g03206(.A(new_n3454), .B(new_n3447), .C(new_n3442), .Y(new_n3463));
  OAI21xp33_ASAP7_75t_L     g03207(.A1(new_n3288), .A2(new_n3290), .B(new_n3291), .Y(new_n3464));
  OAI21xp33_ASAP7_75t_L     g03208(.A1(new_n3462), .A2(new_n3463), .B(new_n3464), .Y(new_n3465));
  NOR2xp33_ASAP7_75t_L      g03209(.A(new_n869), .B(new_n1373), .Y(new_n3466));
  INVx1_ASAP7_75t_L         g03210(.A(new_n3466), .Y(new_n3467));
  NAND3xp33_ASAP7_75t_L     g03211(.A(new_n947), .B(new_n949), .C(new_n1365), .Y(new_n3468));
  AOI22xp33_ASAP7_75t_L     g03212(.A1(new_n1360), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1581), .Y(new_n3469));
  NAND4xp25_ASAP7_75t_L     g03213(.A(new_n3468), .B(\a[20] ), .C(new_n3467), .D(new_n3469), .Y(new_n3470));
  AOI31xp33_ASAP7_75t_L     g03214(.A1(new_n3468), .A2(new_n3467), .A3(new_n3469), .B(\a[20] ), .Y(new_n3471));
  INVx1_ASAP7_75t_L         g03215(.A(new_n3471), .Y(new_n3472));
  AND2x2_ASAP7_75t_L        g03216(.A(new_n3470), .B(new_n3472), .Y(new_n3473));
  NAND3xp33_ASAP7_75t_L     g03217(.A(new_n3465), .B(new_n3461), .C(new_n3473), .Y(new_n3474));
  NOR3xp33_ASAP7_75t_L      g03218(.A(new_n3464), .B(new_n3463), .C(new_n3462), .Y(new_n3475));
  AOI22xp33_ASAP7_75t_L     g03219(.A1(new_n3459), .A2(new_n3455), .B1(new_n3291), .B2(new_n3460), .Y(new_n3476));
  NAND2xp33_ASAP7_75t_L     g03220(.A(new_n3470), .B(new_n3472), .Y(new_n3477));
  OAI21xp33_ASAP7_75t_L     g03221(.A1(new_n3476), .A2(new_n3475), .B(new_n3477), .Y(new_n3478));
  NAND2xp33_ASAP7_75t_L     g03222(.A(new_n3474), .B(new_n3478), .Y(new_n3479));
  NAND2xp33_ASAP7_75t_L     g03223(.A(new_n3398), .B(new_n3479), .Y(new_n3480));
  A2O1A1O1Ixp25_ASAP7_75t_L g03224(.A1(new_n3082), .A2(new_n3088), .B(new_n3091), .C(new_n3299), .D(new_n3295), .Y(new_n3481));
  NAND3xp33_ASAP7_75t_L     g03225(.A(new_n3481), .B(new_n3474), .C(new_n3478), .Y(new_n3482));
  NAND3xp33_ASAP7_75t_L     g03226(.A(new_n3480), .B(new_n3397), .C(new_n3482), .Y(new_n3483));
  XNOR2x2_ASAP7_75t_L       g03227(.A(new_n1071), .B(new_n3396), .Y(new_n3484));
  AOI21xp33_ASAP7_75t_L     g03228(.A1(new_n3478), .A2(new_n3474), .B(new_n3481), .Y(new_n3485));
  NOR2xp33_ASAP7_75t_L      g03229(.A(new_n3398), .B(new_n3479), .Y(new_n3486));
  OAI21xp33_ASAP7_75t_L     g03230(.A1(new_n3485), .A2(new_n3486), .B(new_n3484), .Y(new_n3487));
  AOI221xp5_ASAP7_75t_L     g03231(.A1(new_n3487), .A2(new_n3483), .B1(new_n3317), .B2(new_n3319), .C(new_n3394), .Y(new_n3488));
  INVx1_ASAP7_75t_L         g03232(.A(new_n3394), .Y(new_n3489));
  NAND2xp33_ASAP7_75t_L     g03233(.A(new_n3483), .B(new_n3487), .Y(new_n3490));
  O2A1O1Ixp33_ASAP7_75t_L   g03234(.A1(new_n3323), .A2(new_n3324), .B(new_n3489), .C(new_n3490), .Y(new_n3491));
  NOR2xp33_ASAP7_75t_L      g03235(.A(new_n1539), .B(new_n904), .Y(new_n3492));
  INVx1_ASAP7_75t_L         g03236(.A(new_n3492), .Y(new_n3493));
  NAND2xp33_ASAP7_75t_L     g03237(.A(new_n808), .B(new_n1661), .Y(new_n3494));
  AOI22xp33_ASAP7_75t_L     g03238(.A1(new_n811), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n900), .Y(new_n3495));
  NAND4xp25_ASAP7_75t_L     g03239(.A(new_n3494), .B(\a[14] ), .C(new_n3493), .D(new_n3495), .Y(new_n3496));
  AOI31xp33_ASAP7_75t_L     g03240(.A1(new_n3494), .A2(new_n3493), .A3(new_n3495), .B(\a[14] ), .Y(new_n3497));
  INVx1_ASAP7_75t_L         g03241(.A(new_n3497), .Y(new_n3498));
  NAND2xp33_ASAP7_75t_L     g03242(.A(new_n3496), .B(new_n3498), .Y(new_n3499));
  NOR3xp33_ASAP7_75t_L      g03243(.A(new_n3491), .B(new_n3499), .C(new_n3488), .Y(new_n3500));
  OAI211xp5_ASAP7_75t_L     g03244(.A1(new_n3323), .A2(new_n3324), .B(new_n3490), .C(new_n3489), .Y(new_n3501));
  NOR3xp33_ASAP7_75t_L      g03245(.A(new_n3486), .B(new_n3485), .C(new_n3484), .Y(new_n3502));
  AOI21xp33_ASAP7_75t_L     g03246(.A1(new_n3480), .A2(new_n3482), .B(new_n3397), .Y(new_n3503));
  NOR2xp33_ASAP7_75t_L      g03247(.A(new_n3503), .B(new_n3502), .Y(new_n3504));
  A2O1A1Ixp33_ASAP7_75t_L   g03248(.A1(new_n3319), .A2(new_n3317), .B(new_n3394), .C(new_n3504), .Y(new_n3505));
  AND2x2_ASAP7_75t_L        g03249(.A(new_n3496), .B(new_n3498), .Y(new_n3506));
  AOI21xp33_ASAP7_75t_L     g03250(.A1(new_n3505), .A2(new_n3501), .B(new_n3506), .Y(new_n3507));
  OAI221xp5_ASAP7_75t_L     g03251(.A1(new_n3341), .A2(new_n3337), .B1(new_n3500), .B2(new_n3507), .C(new_n3329), .Y(new_n3508));
  NOR2xp33_ASAP7_75t_L      g03252(.A(new_n3500), .B(new_n3507), .Y(new_n3509));
  OAI21xp33_ASAP7_75t_L     g03253(.A1(new_n3337), .A2(new_n3341), .B(new_n3329), .Y(new_n3510));
  NAND2xp33_ASAP7_75t_L     g03254(.A(new_n3509), .B(new_n3510), .Y(new_n3511));
  AOI21xp33_ASAP7_75t_L     g03255(.A1(new_n3511), .A2(new_n3508), .B(new_n3393), .Y(new_n3512));
  AND2x2_ASAP7_75t_L        g03256(.A(new_n3392), .B(new_n3391), .Y(new_n3513));
  NAND3xp33_ASAP7_75t_L     g03257(.A(new_n3506), .B(new_n3505), .C(new_n3501), .Y(new_n3514));
  OAI21xp33_ASAP7_75t_L     g03258(.A1(new_n3488), .A2(new_n3491), .B(new_n3499), .Y(new_n3515));
  AOI221xp5_ASAP7_75t_L     g03259(.A1(new_n3515), .A2(new_n3514), .B1(new_n3333), .B2(new_n3231), .C(new_n3336), .Y(new_n3516));
  NAND2xp33_ASAP7_75t_L     g03260(.A(new_n3515), .B(new_n3514), .Y(new_n3517));
  OAI211xp5_ASAP7_75t_L     g03261(.A1(new_n3119), .A2(new_n3343), .B(new_n3344), .C(new_n3333), .Y(new_n3518));
  AOI21xp33_ASAP7_75t_L     g03262(.A1(new_n3329), .A2(new_n3518), .B(new_n3517), .Y(new_n3519));
  NOR3xp33_ASAP7_75t_L      g03263(.A(new_n3519), .B(new_n3513), .C(new_n3516), .Y(new_n3520));
  NOR2xp33_ASAP7_75t_L      g03264(.A(new_n3512), .B(new_n3520), .Y(new_n3521));
  A2O1A1Ixp33_ASAP7_75t_L   g03265(.A1(new_n3349), .A2(new_n3387), .B(new_n3346), .C(new_n3521), .Y(new_n3522));
  A2O1A1O1Ixp25_ASAP7_75t_L g03266(.A1(new_n3151), .A2(new_n3150), .B(new_n3348), .C(new_n3349), .D(new_n3346), .Y(new_n3523));
  OAI21xp33_ASAP7_75t_L     g03267(.A1(new_n3516), .A2(new_n3519), .B(new_n3513), .Y(new_n3524));
  NAND3xp33_ASAP7_75t_L     g03268(.A(new_n3511), .B(new_n3508), .C(new_n3393), .Y(new_n3525));
  NAND2xp33_ASAP7_75t_L     g03269(.A(new_n3525), .B(new_n3524), .Y(new_n3526));
  NAND2xp33_ASAP7_75t_L     g03270(.A(new_n3523), .B(new_n3526), .Y(new_n3527));
  AOI22xp33_ASAP7_75t_L     g03271(.A1(new_n444), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n471), .Y(new_n3528));
  OAI221xp5_ASAP7_75t_L     g03272(.A1(new_n468), .A2(new_n2348), .B1(new_n469), .B2(new_n2505), .C(new_n3528), .Y(new_n3529));
  XNOR2x2_ASAP7_75t_L       g03273(.A(\a[8] ), .B(new_n3529), .Y(new_n3530));
  NAND3xp33_ASAP7_75t_L     g03274(.A(new_n3522), .B(new_n3527), .C(new_n3530), .Y(new_n3531));
  A2O1A1O1Ixp25_ASAP7_75t_L g03275(.A1(new_n3224), .A2(new_n3144), .B(new_n3340), .C(new_n3350), .D(new_n3526), .Y(new_n3532));
  A2O1A1Ixp33_ASAP7_75t_L   g03276(.A1(new_n3144), .A2(new_n3224), .B(new_n3340), .C(new_n3350), .Y(new_n3533));
  NOR2xp33_ASAP7_75t_L      g03277(.A(new_n3533), .B(new_n3521), .Y(new_n3534));
  INVx1_ASAP7_75t_L         g03278(.A(new_n3530), .Y(new_n3535));
  OAI21xp33_ASAP7_75t_L     g03279(.A1(new_n3534), .A2(new_n3532), .B(new_n3535), .Y(new_n3536));
  NOR3xp33_ASAP7_75t_L      g03280(.A(new_n3347), .B(new_n3351), .C(new_n3354), .Y(new_n3537));
  O2A1O1Ixp33_ASAP7_75t_L   g03281(.A1(new_n3359), .A2(new_n3356), .B(new_n3361), .C(new_n3537), .Y(new_n3538));
  NAND3xp33_ASAP7_75t_L     g03282(.A(new_n3538), .B(new_n3536), .C(new_n3531), .Y(new_n3539));
  NOR3xp33_ASAP7_75t_L      g03283(.A(new_n3532), .B(new_n3534), .C(new_n3535), .Y(new_n3540));
  AOI21xp33_ASAP7_75t_L     g03284(.A1(new_n3522), .A2(new_n3527), .B(new_n3530), .Y(new_n3541));
  NAND2xp33_ASAP7_75t_L     g03285(.A(new_n3358), .B(new_n3357), .Y(new_n3542));
  MAJx2_ASAP7_75t_L         g03286(.A(new_n3156), .B(new_n3148), .C(new_n3360), .Y(new_n3543));
  MAJIxp5_ASAP7_75t_L       g03287(.A(new_n3543), .B(new_n3542), .C(new_n3354), .Y(new_n3544));
  OAI21xp33_ASAP7_75t_L     g03288(.A1(new_n3540), .A2(new_n3541), .B(new_n3544), .Y(new_n3545));
  AOI22xp33_ASAP7_75t_L     g03289(.A1(new_n344), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n370), .Y(new_n3546));
  OAI221xp5_ASAP7_75t_L     g03290(.A1(new_n429), .A2(new_n2688), .B1(new_n366), .B2(new_n2990), .C(new_n3546), .Y(new_n3547));
  XNOR2x2_ASAP7_75t_L       g03291(.A(\a[5] ), .B(new_n3547), .Y(new_n3548));
  NAND3xp33_ASAP7_75t_L     g03292(.A(new_n3545), .B(new_n3539), .C(new_n3548), .Y(new_n3549));
  NOR4xp25_ASAP7_75t_L      g03293(.A(new_n3363), .B(new_n3537), .C(new_n3541), .D(new_n3540), .Y(new_n3550));
  AOI21xp33_ASAP7_75t_L     g03294(.A1(new_n3536), .A2(new_n3531), .B(new_n3538), .Y(new_n3551));
  INVx1_ASAP7_75t_L         g03295(.A(new_n3548), .Y(new_n3552));
  OAI21xp33_ASAP7_75t_L     g03296(.A1(new_n3551), .A2(new_n3550), .B(new_n3552), .Y(new_n3553));
  NAND2xp33_ASAP7_75t_L     g03297(.A(new_n3549), .B(new_n3553), .Y(new_n3554));
  A2O1A1O1Ixp25_ASAP7_75t_L g03298(.A1(new_n2977), .A2(new_n3174), .B(new_n3171), .C(new_n3177), .D(new_n3223), .Y(new_n3555));
  INVx1_ASAP7_75t_L         g03299(.A(new_n3367), .Y(new_n3556));
  AO21x2_ASAP7_75t_L        g03300(.A1(new_n3371), .A2(new_n3555), .B(new_n3556), .Y(new_n3557));
  NOR2xp33_ASAP7_75t_L      g03301(.A(new_n3554), .B(new_n3557), .Y(new_n3558));
  AND2x2_ASAP7_75t_L        g03302(.A(new_n3549), .B(new_n3553), .Y(new_n3559));
  INVx1_ASAP7_75t_L         g03303(.A(new_n3223), .Y(new_n3560));
  AOI31xp33_ASAP7_75t_L     g03304(.A1(new_n3178), .A2(new_n3560), .A3(new_n3371), .B(new_n3556), .Y(new_n3561));
  NOR2xp33_ASAP7_75t_L      g03305(.A(new_n3561), .B(new_n3559), .Y(new_n3562));
  INVx1_ASAP7_75t_L         g03306(.A(new_n3211), .Y(new_n3563));
  NOR2xp33_ASAP7_75t_L      g03307(.A(\b[32] ), .B(\b[33] ), .Y(new_n3564));
  INVx1_ASAP7_75t_L         g03308(.A(\b[33] ), .Y(new_n3565));
  NOR2xp33_ASAP7_75t_L      g03309(.A(new_n3207), .B(new_n3565), .Y(new_n3566));
  NOR2xp33_ASAP7_75t_L      g03310(.A(new_n3564), .B(new_n3566), .Y(new_n3567));
  A2O1A1Ixp33_ASAP7_75t_L   g03311(.A1(new_n3563), .A2(new_n3209), .B(new_n3208), .C(new_n3567), .Y(new_n3568));
  O2A1O1Ixp33_ASAP7_75t_L   g03312(.A1(new_n2982), .A2(new_n3180), .B(new_n3183), .C(new_n3212), .Y(new_n3569));
  NOR3xp33_ASAP7_75t_L      g03313(.A(new_n3569), .B(new_n3567), .C(new_n3208), .Y(new_n3570));
  INVx1_ASAP7_75t_L         g03314(.A(new_n3570), .Y(new_n3571));
  NAND2xp33_ASAP7_75t_L     g03315(.A(new_n3568), .B(new_n3571), .Y(new_n3572));
  AOI22xp33_ASAP7_75t_L     g03316(.A1(\b[31] ), .A2(new_n282), .B1(\b[33] ), .B2(new_n303), .Y(new_n3573));
  OAI221xp5_ASAP7_75t_L     g03317(.A1(new_n291), .A2(new_n3207), .B1(new_n268), .B2(new_n3572), .C(new_n3573), .Y(new_n3574));
  XNOR2x2_ASAP7_75t_L       g03318(.A(new_n262), .B(new_n3574), .Y(new_n3575));
  OAI21xp33_ASAP7_75t_L     g03319(.A1(new_n3558), .A2(new_n3562), .B(new_n3575), .Y(new_n3576));
  INVx1_ASAP7_75t_L         g03320(.A(new_n3576), .Y(new_n3577));
  NOR3xp33_ASAP7_75t_L      g03321(.A(new_n3562), .B(new_n3558), .C(new_n3575), .Y(new_n3578));
  NOR2xp33_ASAP7_75t_L      g03322(.A(new_n3578), .B(new_n3577), .Y(new_n3579));
  XNOR2x2_ASAP7_75t_L       g03323(.A(new_n3383), .B(new_n3579), .Y(\f[33] ));
  INVx1_ASAP7_75t_L         g03324(.A(new_n3567), .Y(new_n3581));
  O2A1O1Ixp33_ASAP7_75t_L   g03325(.A1(new_n3180), .A2(new_n3207), .B(new_n3210), .C(new_n3581), .Y(new_n3582));
  NOR2xp33_ASAP7_75t_L      g03326(.A(\b[33] ), .B(\b[34] ), .Y(new_n3583));
  INVx1_ASAP7_75t_L         g03327(.A(\b[34] ), .Y(new_n3584));
  NOR2xp33_ASAP7_75t_L      g03328(.A(new_n3565), .B(new_n3584), .Y(new_n3585));
  NOR2xp33_ASAP7_75t_L      g03329(.A(new_n3583), .B(new_n3585), .Y(new_n3586));
  A2O1A1Ixp33_ASAP7_75t_L   g03330(.A1(\b[33] ), .A2(\b[32] ), .B(new_n3582), .C(new_n3586), .Y(new_n3587));
  A2O1A1O1Ixp25_ASAP7_75t_L g03331(.A1(new_n3209), .A2(new_n3563), .B(new_n3208), .C(new_n3567), .D(new_n3566), .Y(new_n3588));
  INVx1_ASAP7_75t_L         g03332(.A(new_n3586), .Y(new_n3589));
  NAND2xp33_ASAP7_75t_L     g03333(.A(new_n3589), .B(new_n3588), .Y(new_n3590));
  NAND2xp33_ASAP7_75t_L     g03334(.A(new_n3590), .B(new_n3587), .Y(new_n3591));
  AOI22xp33_ASAP7_75t_L     g03335(.A1(\b[32] ), .A2(new_n282), .B1(\b[34] ), .B2(new_n303), .Y(new_n3592));
  OAI221xp5_ASAP7_75t_L     g03336(.A1(new_n291), .A2(new_n3565), .B1(new_n268), .B2(new_n3591), .C(new_n3592), .Y(new_n3593));
  XNOR2x2_ASAP7_75t_L       g03337(.A(\a[2] ), .B(new_n3593), .Y(new_n3594));
  NOR3xp33_ASAP7_75t_L      g03338(.A(new_n3550), .B(new_n3551), .C(new_n3548), .Y(new_n3595));
  AOI21xp33_ASAP7_75t_L     g03339(.A1(new_n3561), .A2(new_n3554), .B(new_n3595), .Y(new_n3596));
  AOI22xp33_ASAP7_75t_L     g03340(.A1(new_n444), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n471), .Y(new_n3597));
  OAI221xp5_ASAP7_75t_L     g03341(.A1(new_n468), .A2(new_n2497), .B1(new_n469), .B2(new_n2672), .C(new_n3597), .Y(new_n3598));
  XNOR2x2_ASAP7_75t_L       g03342(.A(\a[8] ), .B(new_n3598), .Y(new_n3599));
  A2O1A1O1Ixp25_ASAP7_75t_L g03343(.A1(new_n3349), .A2(new_n3387), .B(new_n3346), .C(new_n3524), .D(new_n3520), .Y(new_n3600));
  NOR3xp33_ASAP7_75t_L      g03344(.A(new_n3475), .B(new_n3476), .C(new_n3477), .Y(new_n3601));
  AOI21xp33_ASAP7_75t_L     g03345(.A1(new_n3461), .A2(new_n3465), .B(new_n3473), .Y(new_n3602));
  NOR2xp33_ASAP7_75t_L      g03346(.A(new_n3602), .B(new_n3601), .Y(new_n3603));
  NAND3xp33_ASAP7_75t_L     g03347(.A(new_n3461), .B(new_n3465), .C(new_n3477), .Y(new_n3604));
  AOI22xp33_ASAP7_75t_L     g03348(.A1(new_n1360), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1581), .Y(new_n3605));
  OAI221xp5_ASAP7_75t_L     g03349(.A1(new_n1373), .A2(new_n942), .B1(new_n1359), .B2(new_n1035), .C(new_n3605), .Y(new_n3606));
  XNOR2x2_ASAP7_75t_L       g03350(.A(\a[20] ), .B(new_n3606), .Y(new_n3607));
  OAI21xp33_ASAP7_75t_L     g03351(.A1(new_n3462), .A2(new_n3464), .B(new_n3459), .Y(new_n3608));
  NAND2xp33_ASAP7_75t_L     g03352(.A(new_n3425), .B(new_n3427), .Y(new_n3609));
  AND3x1_ASAP7_75t_L        g03353(.A(new_n3609), .B(new_n3421), .C(new_n3420), .Y(new_n3610));
  AOI221xp5_ASAP7_75t_L     g03354(.A1(new_n3429), .A2(new_n3428), .B1(new_n3265), .B2(new_n3272), .C(new_n3430), .Y(new_n3611));
  AOI22xp33_ASAP7_75t_L     g03355(.A1(new_n2552), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n2736), .Y(new_n3612));
  OAI221xp5_ASAP7_75t_L     g03356(.A1(new_n2547), .A2(new_n418), .B1(new_n2734), .B2(new_n425), .C(new_n3612), .Y(new_n3613));
  OR2x4_ASAP7_75t_L         g03357(.A(new_n2538), .B(new_n3613), .Y(new_n3614));
  NAND2xp33_ASAP7_75t_L     g03358(.A(new_n2538), .B(new_n3613), .Y(new_n3615));
  NOR2xp33_ASAP7_75t_L      g03359(.A(new_n3400), .B(new_n3260), .Y(new_n3616));
  NAND2xp33_ASAP7_75t_L     g03360(.A(new_n3419), .B(new_n3416), .Y(new_n3617));
  MAJIxp5_ASAP7_75t_L       g03361(.A(new_n3617), .B(new_n3408), .C(new_n3616), .Y(new_n3618));
  NOR2xp33_ASAP7_75t_L      g03362(.A(new_n298), .B(new_n3024), .Y(new_n3619));
  NOR3xp33_ASAP7_75t_L      g03363(.A(new_n326), .B(new_n328), .C(new_n3256), .Y(new_n3620));
  OAI22xp33_ASAP7_75t_L     g03364(.A1(new_n3402), .A2(new_n276), .B1(new_n324), .B2(new_n3022), .Y(new_n3621));
  NOR4xp25_ASAP7_75t_L      g03365(.A(new_n3620), .B(new_n3621), .C(new_n3015), .D(new_n3619), .Y(new_n3622));
  OAI31xp33_ASAP7_75t_L     g03366(.A1(new_n3620), .A2(new_n3621), .A3(new_n3619), .B(new_n3015), .Y(new_n3623));
  INVx1_ASAP7_75t_L         g03367(.A(new_n3623), .Y(new_n3624));
  NAND2xp33_ASAP7_75t_L     g03368(.A(\a[35] ), .B(new_n3408), .Y(new_n3625));
  INVx1_ASAP7_75t_L         g03369(.A(\a[34] ), .Y(new_n3626));
  NAND2xp33_ASAP7_75t_L     g03370(.A(\a[35] ), .B(new_n3626), .Y(new_n3627));
  INVx1_ASAP7_75t_L         g03371(.A(\a[35] ), .Y(new_n3628));
  NAND2xp33_ASAP7_75t_L     g03372(.A(\a[34] ), .B(new_n3628), .Y(new_n3629));
  AOI21xp33_ASAP7_75t_L     g03373(.A1(new_n3629), .A2(new_n3627), .B(new_n3407), .Y(new_n3630));
  NAND2xp33_ASAP7_75t_L     g03374(.A(new_n269), .B(new_n3630), .Y(new_n3631));
  NAND2xp33_ASAP7_75t_L     g03375(.A(new_n3629), .B(new_n3627), .Y(new_n3632));
  NOR2xp33_ASAP7_75t_L      g03376(.A(new_n3632), .B(new_n3407), .Y(new_n3633));
  NAND2xp33_ASAP7_75t_L     g03377(.A(\b[1] ), .B(new_n3633), .Y(new_n3634));
  NAND2xp33_ASAP7_75t_L     g03378(.A(new_n3406), .B(new_n3405), .Y(new_n3635));
  NOR2xp33_ASAP7_75t_L      g03379(.A(\a[33] ), .B(new_n3626), .Y(new_n3636));
  NOR2xp33_ASAP7_75t_L      g03380(.A(\a[34] ), .B(new_n3404), .Y(new_n3637));
  NOR2xp33_ASAP7_75t_L      g03381(.A(new_n3636), .B(new_n3637), .Y(new_n3638));
  NOR2xp33_ASAP7_75t_L      g03382(.A(new_n3635), .B(new_n3638), .Y(new_n3639));
  NAND2xp33_ASAP7_75t_L     g03383(.A(\b[0] ), .B(new_n3639), .Y(new_n3640));
  NAND3xp33_ASAP7_75t_L     g03384(.A(new_n3631), .B(new_n3634), .C(new_n3640), .Y(new_n3641));
  XNOR2x2_ASAP7_75t_L       g03385(.A(new_n3625), .B(new_n3641), .Y(new_n3642));
  NOR3xp33_ASAP7_75t_L      g03386(.A(new_n3642), .B(new_n3624), .C(new_n3622), .Y(new_n3643));
  INVx1_ASAP7_75t_L         g03387(.A(new_n3622), .Y(new_n3644));
  XOR2x2_ASAP7_75t_L        g03388(.A(new_n3625), .B(new_n3641), .Y(new_n3645));
  AOI21xp33_ASAP7_75t_L     g03389(.A1(new_n3623), .A2(new_n3644), .B(new_n3645), .Y(new_n3646));
  NOR3xp33_ASAP7_75t_L      g03390(.A(new_n3618), .B(new_n3643), .C(new_n3646), .Y(new_n3647));
  AOI22xp33_ASAP7_75t_L     g03391(.A1(new_n3419), .A2(new_n3416), .B1(new_n3409), .B2(new_n3413), .Y(new_n3648));
  NAND3xp33_ASAP7_75t_L     g03392(.A(new_n3645), .B(new_n3623), .C(new_n3644), .Y(new_n3649));
  OAI21xp33_ASAP7_75t_L     g03393(.A1(new_n3622), .A2(new_n3624), .B(new_n3642), .Y(new_n3650));
  AOI221xp5_ASAP7_75t_L     g03394(.A1(new_n3408), .A2(new_n3616), .B1(new_n3650), .B2(new_n3649), .C(new_n3648), .Y(new_n3651));
  OAI211xp5_ASAP7_75t_L     g03395(.A1(new_n3651), .A2(new_n3647), .B(new_n3615), .C(new_n3614), .Y(new_n3652));
  NAND2xp33_ASAP7_75t_L     g03396(.A(new_n3615), .B(new_n3614), .Y(new_n3653));
  NOR2xp33_ASAP7_75t_L      g03397(.A(new_n3646), .B(new_n3643), .Y(new_n3654));
  A2O1A1Ixp33_ASAP7_75t_L   g03398(.A1(new_n3616), .A2(new_n3408), .B(new_n3648), .C(new_n3654), .Y(new_n3655));
  INVx1_ASAP7_75t_L         g03399(.A(new_n3651), .Y(new_n3656));
  NAND3xp33_ASAP7_75t_L     g03400(.A(new_n3656), .B(new_n3655), .C(new_n3653), .Y(new_n3657));
  OAI211xp5_ASAP7_75t_L     g03401(.A1(new_n3610), .A2(new_n3611), .B(new_n3652), .C(new_n3657), .Y(new_n3658));
  AND4x1_ASAP7_75t_L        g03402(.A(new_n3420), .B(new_n3427), .C(new_n3421), .D(new_n3425), .Y(new_n3659));
  AOI22xp33_ASAP7_75t_L     g03403(.A1(new_n3420), .A2(new_n3421), .B1(new_n3425), .B2(new_n3427), .Y(new_n3660));
  O2A1O1Ixp33_ASAP7_75t_L   g03404(.A1(new_n3659), .A2(new_n3660), .B(new_n3431), .C(new_n3610), .Y(new_n3661));
  AOI21xp33_ASAP7_75t_L     g03405(.A1(new_n3656), .A2(new_n3655), .B(new_n3653), .Y(new_n3662));
  AOI211xp5_ASAP7_75t_L     g03406(.A1(new_n3615), .A2(new_n3614), .B(new_n3651), .C(new_n3647), .Y(new_n3663));
  OAI21xp33_ASAP7_75t_L     g03407(.A1(new_n3662), .A2(new_n3663), .B(new_n3661), .Y(new_n3664));
  AOI22xp33_ASAP7_75t_L     g03408(.A1(new_n2114), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n2259), .Y(new_n3665));
  OAI221xp5_ASAP7_75t_L     g03409(.A1(new_n2109), .A2(new_n540), .B1(new_n2257), .B2(new_n624), .C(new_n3665), .Y(new_n3666));
  XNOR2x2_ASAP7_75t_L       g03410(.A(\a[26] ), .B(new_n3666), .Y(new_n3667));
  NAND3xp33_ASAP7_75t_L     g03411(.A(new_n3664), .B(new_n3658), .C(new_n3667), .Y(new_n3668));
  NOR3xp33_ASAP7_75t_L      g03412(.A(new_n3661), .B(new_n3662), .C(new_n3663), .Y(new_n3669));
  AOI211xp5_ASAP7_75t_L     g03413(.A1(new_n3252), .A2(new_n3251), .B(new_n3261), .C(new_n3263), .Y(new_n3670));
  OAI21xp33_ASAP7_75t_L     g03414(.A1(new_n3670), .A2(new_n3245), .B(new_n3264), .Y(new_n3671));
  NAND3xp33_ASAP7_75t_L     g03415(.A(new_n3609), .B(new_n3421), .C(new_n3420), .Y(new_n3672));
  A2O1A1Ixp33_ASAP7_75t_L   g03416(.A1(new_n3429), .A2(new_n3428), .B(new_n3671), .C(new_n3672), .Y(new_n3673));
  AOI21xp33_ASAP7_75t_L     g03417(.A1(new_n3657), .A2(new_n3652), .B(new_n3673), .Y(new_n3674));
  INVx1_ASAP7_75t_L         g03418(.A(new_n3667), .Y(new_n3675));
  OAI21xp33_ASAP7_75t_L     g03419(.A1(new_n3669), .A2(new_n3674), .B(new_n3675), .Y(new_n3676));
  A2O1A1O1Ixp25_ASAP7_75t_L g03420(.A1(new_n3279), .A2(new_n3277), .B(new_n3269), .C(new_n3441), .D(new_n3445), .Y(new_n3677));
  AND3x1_ASAP7_75t_L        g03421(.A(new_n3677), .B(new_n3676), .C(new_n3668), .Y(new_n3678));
  AOI21xp33_ASAP7_75t_L     g03422(.A1(new_n3676), .A2(new_n3668), .B(new_n3677), .Y(new_n3679));
  NOR2xp33_ASAP7_75t_L      g03423(.A(new_n760), .B(new_n1699), .Y(new_n3680));
  INVx1_ASAP7_75t_L         g03424(.A(new_n3680), .Y(new_n3681));
  NAND3xp33_ASAP7_75t_L     g03425(.A(new_n787), .B(new_n789), .C(new_n1695), .Y(new_n3682));
  AOI22xp33_ASAP7_75t_L     g03426(.A1(new_n1704), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1837), .Y(new_n3683));
  NAND4xp25_ASAP7_75t_L     g03427(.A(new_n3682), .B(\a[23] ), .C(new_n3681), .D(new_n3683), .Y(new_n3684));
  NAND2xp33_ASAP7_75t_L     g03428(.A(new_n3683), .B(new_n3682), .Y(new_n3685));
  A2O1A1Ixp33_ASAP7_75t_L   g03429(.A1(\b[12] ), .A2(new_n1706), .B(new_n3685), .C(new_n1689), .Y(new_n3686));
  AND2x2_ASAP7_75t_L        g03430(.A(new_n3684), .B(new_n3686), .Y(new_n3687));
  OAI21xp33_ASAP7_75t_L     g03431(.A1(new_n3679), .A2(new_n3678), .B(new_n3687), .Y(new_n3688));
  NAND3xp33_ASAP7_75t_L     g03432(.A(new_n3677), .B(new_n3676), .C(new_n3668), .Y(new_n3689));
  AO21x2_ASAP7_75t_L        g03433(.A1(new_n3668), .A2(new_n3676), .B(new_n3677), .Y(new_n3690));
  NAND2xp33_ASAP7_75t_L     g03434(.A(new_n3684), .B(new_n3686), .Y(new_n3691));
  NAND3xp33_ASAP7_75t_L     g03435(.A(new_n3690), .B(new_n3691), .C(new_n3689), .Y(new_n3692));
  AOI21xp33_ASAP7_75t_L     g03436(.A1(new_n3692), .A2(new_n3688), .B(new_n3608), .Y(new_n3693));
  AOI31xp33_ASAP7_75t_L     g03437(.A1(new_n3460), .A2(new_n3455), .A3(new_n3291), .B(new_n3463), .Y(new_n3694));
  NAND2xp33_ASAP7_75t_L     g03438(.A(new_n3692), .B(new_n3688), .Y(new_n3695));
  NOR2xp33_ASAP7_75t_L      g03439(.A(new_n3694), .B(new_n3695), .Y(new_n3696));
  NOR3xp33_ASAP7_75t_L      g03440(.A(new_n3696), .B(new_n3693), .C(new_n3607), .Y(new_n3697));
  INVx1_ASAP7_75t_L         g03441(.A(new_n3607), .Y(new_n3698));
  NAND2xp33_ASAP7_75t_L     g03442(.A(new_n3694), .B(new_n3695), .Y(new_n3699));
  NAND3xp33_ASAP7_75t_L     g03443(.A(new_n3608), .B(new_n3688), .C(new_n3692), .Y(new_n3700));
  AOI21xp33_ASAP7_75t_L     g03444(.A1(new_n3699), .A2(new_n3700), .B(new_n3698), .Y(new_n3701));
  OAI221xp5_ASAP7_75t_L     g03445(.A1(new_n3603), .A2(new_n3481), .B1(new_n3697), .B2(new_n3701), .C(new_n3604), .Y(new_n3702));
  A2O1A1Ixp33_ASAP7_75t_L   g03446(.A1(new_n3474), .A2(new_n3478), .B(new_n3481), .C(new_n3604), .Y(new_n3703));
  NAND3xp33_ASAP7_75t_L     g03447(.A(new_n3698), .B(new_n3699), .C(new_n3700), .Y(new_n3704));
  OAI21xp33_ASAP7_75t_L     g03448(.A1(new_n3693), .A2(new_n3696), .B(new_n3607), .Y(new_n3705));
  NAND3xp33_ASAP7_75t_L     g03449(.A(new_n3703), .B(new_n3704), .C(new_n3705), .Y(new_n3706));
  NOR2xp33_ASAP7_75t_L      g03450(.A(new_n1313), .B(new_n1154), .Y(new_n3707));
  AOI22xp33_ASAP7_75t_L     g03451(.A1(new_n1076), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1253), .Y(new_n3708));
  OAI21xp33_ASAP7_75t_L     g03452(.A1(new_n1156), .A2(new_n1438), .B(new_n3708), .Y(new_n3709));
  NOR3xp33_ASAP7_75t_L      g03453(.A(new_n3709), .B(new_n3707), .C(new_n1071), .Y(new_n3710));
  INVx1_ASAP7_75t_L         g03454(.A(new_n3707), .Y(new_n3711));
  INVx1_ASAP7_75t_L         g03455(.A(new_n1435), .Y(new_n3712));
  NOR2xp33_ASAP7_75t_L      g03456(.A(new_n1436), .B(new_n3712), .Y(new_n3713));
  NAND2xp33_ASAP7_75t_L     g03457(.A(new_n1073), .B(new_n3713), .Y(new_n3714));
  AOI31xp33_ASAP7_75t_L     g03458(.A1(new_n3714), .A2(new_n3711), .A3(new_n3708), .B(\a[17] ), .Y(new_n3715));
  NOR2xp33_ASAP7_75t_L      g03459(.A(new_n3710), .B(new_n3715), .Y(new_n3716));
  NAND3xp33_ASAP7_75t_L     g03460(.A(new_n3706), .B(new_n3702), .C(new_n3716), .Y(new_n3717));
  AO21x2_ASAP7_75t_L        g03461(.A1(new_n3702), .A2(new_n3706), .B(new_n3716), .Y(new_n3718));
  NAND2xp33_ASAP7_75t_L     g03462(.A(new_n3717), .B(new_n3718), .Y(new_n3719));
  NOR3xp33_ASAP7_75t_L      g03463(.A(new_n3491), .B(new_n3719), .C(new_n3502), .Y(new_n3720));
  A2O1A1O1Ixp25_ASAP7_75t_L g03464(.A1(new_n3113), .A2(new_n3107), .B(new_n3318), .C(new_n3317), .D(new_n3394), .Y(new_n3721));
  AND3x1_ASAP7_75t_L        g03465(.A(new_n3706), .B(new_n3702), .C(new_n3716), .Y(new_n3722));
  AOI21xp33_ASAP7_75t_L     g03466(.A1(new_n3706), .A2(new_n3702), .B(new_n3716), .Y(new_n3723));
  NOR2xp33_ASAP7_75t_L      g03467(.A(new_n3723), .B(new_n3722), .Y(new_n3724));
  O2A1O1Ixp33_ASAP7_75t_L   g03468(.A1(new_n3721), .A2(new_n3503), .B(new_n3483), .C(new_n3724), .Y(new_n3725));
  NOR2xp33_ASAP7_75t_L      g03469(.A(new_n1655), .B(new_n904), .Y(new_n3726));
  INVx1_ASAP7_75t_L         g03470(.A(new_n3726), .Y(new_n3727));
  NOR2xp33_ASAP7_75t_L      g03471(.A(new_n1778), .B(new_n1907), .Y(new_n3728));
  NAND2xp33_ASAP7_75t_L     g03472(.A(new_n808), .B(new_n3728), .Y(new_n3729));
  AOI22xp33_ASAP7_75t_L     g03473(.A1(new_n811), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n900), .Y(new_n3730));
  NAND4xp25_ASAP7_75t_L     g03474(.A(new_n3729), .B(\a[14] ), .C(new_n3727), .D(new_n3730), .Y(new_n3731));
  AOI31xp33_ASAP7_75t_L     g03475(.A1(new_n3729), .A2(new_n3727), .A3(new_n3730), .B(\a[14] ), .Y(new_n3732));
  INVx1_ASAP7_75t_L         g03476(.A(new_n3732), .Y(new_n3733));
  NAND2xp33_ASAP7_75t_L     g03477(.A(new_n3731), .B(new_n3733), .Y(new_n3734));
  NOR3xp33_ASAP7_75t_L      g03478(.A(new_n3720), .B(new_n3725), .C(new_n3734), .Y(new_n3735));
  A2O1A1O1Ixp25_ASAP7_75t_L g03479(.A1(new_n3317), .A2(new_n3319), .B(new_n3394), .C(new_n3487), .D(new_n3502), .Y(new_n3736));
  NAND2xp33_ASAP7_75t_L     g03480(.A(new_n3724), .B(new_n3736), .Y(new_n3737));
  A2O1A1Ixp33_ASAP7_75t_L   g03481(.A1(new_n3316), .A2(new_n3312), .B(new_n3324), .C(new_n3489), .Y(new_n3738));
  A2O1A1Ixp33_ASAP7_75t_L   g03482(.A1(new_n3487), .A2(new_n3738), .B(new_n3502), .C(new_n3719), .Y(new_n3739));
  INVx1_ASAP7_75t_L         g03483(.A(new_n3731), .Y(new_n3740));
  NOR2xp33_ASAP7_75t_L      g03484(.A(new_n3732), .B(new_n3740), .Y(new_n3741));
  AOI21xp33_ASAP7_75t_L     g03485(.A1(new_n3739), .A2(new_n3737), .B(new_n3741), .Y(new_n3742));
  NOR2xp33_ASAP7_75t_L      g03486(.A(new_n3742), .B(new_n3735), .Y(new_n3743));
  NOR3xp33_ASAP7_75t_L      g03487(.A(new_n3506), .B(new_n3491), .C(new_n3488), .Y(new_n3744));
  INVx1_ASAP7_75t_L         g03488(.A(new_n3744), .Y(new_n3745));
  NAND3xp33_ASAP7_75t_L     g03489(.A(new_n3743), .B(new_n3508), .C(new_n3745), .Y(new_n3746));
  NAND3xp33_ASAP7_75t_L     g03490(.A(new_n3739), .B(new_n3737), .C(new_n3741), .Y(new_n3747));
  OAI21xp33_ASAP7_75t_L     g03491(.A1(new_n3725), .A2(new_n3720), .B(new_n3734), .Y(new_n3748));
  NAND2xp33_ASAP7_75t_L     g03492(.A(new_n3747), .B(new_n3748), .Y(new_n3749));
  OAI21xp33_ASAP7_75t_L     g03493(.A1(new_n3744), .A2(new_n3516), .B(new_n3749), .Y(new_n3750));
  OAI22xp33_ASAP7_75t_L     g03494(.A1(new_n706), .A2(new_n1909), .B1(new_n2067), .B2(new_n580), .Y(new_n3751));
  AOI221xp5_ASAP7_75t_L     g03495(.A1(\b[24] ), .A2(new_n584), .B1(new_n578), .B2(new_n2648), .C(new_n3751), .Y(new_n3752));
  AND2x2_ASAP7_75t_L        g03496(.A(\a[11] ), .B(new_n3752), .Y(new_n3753));
  NOR2xp33_ASAP7_75t_L      g03497(.A(\a[11] ), .B(new_n3752), .Y(new_n3754));
  OAI211xp5_ASAP7_75t_L     g03498(.A1(new_n3753), .A2(new_n3754), .B(new_n3746), .C(new_n3750), .Y(new_n3755));
  OAI21xp33_ASAP7_75t_L     g03499(.A1(new_n3509), .A2(new_n3510), .B(new_n3745), .Y(new_n3756));
  NOR2xp33_ASAP7_75t_L      g03500(.A(new_n3749), .B(new_n3756), .Y(new_n3757));
  AOI22xp33_ASAP7_75t_L     g03501(.A1(new_n3747), .A2(new_n3748), .B1(new_n3745), .B2(new_n3508), .Y(new_n3758));
  NOR2xp33_ASAP7_75t_L      g03502(.A(new_n3754), .B(new_n3753), .Y(new_n3759));
  OAI21xp33_ASAP7_75t_L     g03503(.A1(new_n3758), .A2(new_n3757), .B(new_n3759), .Y(new_n3760));
  NAND2xp33_ASAP7_75t_L     g03504(.A(new_n3760), .B(new_n3755), .Y(new_n3761));
  NAND2xp33_ASAP7_75t_L     g03505(.A(new_n3600), .B(new_n3761), .Y(new_n3762));
  OAI21xp33_ASAP7_75t_L     g03506(.A1(new_n3512), .A2(new_n3523), .B(new_n3525), .Y(new_n3763));
  NAND3xp33_ASAP7_75t_L     g03507(.A(new_n3763), .B(new_n3755), .C(new_n3760), .Y(new_n3764));
  NAND3xp33_ASAP7_75t_L     g03508(.A(new_n3762), .B(new_n3599), .C(new_n3764), .Y(new_n3765));
  INVx1_ASAP7_75t_L         g03509(.A(new_n3599), .Y(new_n3766));
  AOI21xp33_ASAP7_75t_L     g03510(.A1(new_n3760), .A2(new_n3755), .B(new_n3763), .Y(new_n3767));
  NOR2xp33_ASAP7_75t_L      g03511(.A(new_n3600), .B(new_n3761), .Y(new_n3768));
  OAI21xp33_ASAP7_75t_L     g03512(.A1(new_n3767), .A2(new_n3768), .B(new_n3766), .Y(new_n3769));
  NAND2xp33_ASAP7_75t_L     g03513(.A(new_n3765), .B(new_n3769), .Y(new_n3770));
  XNOR2x2_ASAP7_75t_L       g03514(.A(new_n3523), .B(new_n3526), .Y(new_n3771));
  MAJIxp5_ASAP7_75t_L       g03515(.A(new_n3538), .B(new_n3771), .C(new_n3530), .Y(new_n3772));
  NOR2xp33_ASAP7_75t_L      g03516(.A(new_n3772), .B(new_n3770), .Y(new_n3773));
  NOR2xp33_ASAP7_75t_L      g03517(.A(new_n3534), .B(new_n3532), .Y(new_n3774));
  NAND2xp33_ASAP7_75t_L     g03518(.A(new_n3535), .B(new_n3774), .Y(new_n3775));
  AOI22xp33_ASAP7_75t_L     g03519(.A1(new_n3765), .A2(new_n3769), .B1(new_n3775), .B2(new_n3545), .Y(new_n3776));
  AOI22xp33_ASAP7_75t_L     g03520(.A1(new_n344), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n370), .Y(new_n3777));
  OAI221xp5_ASAP7_75t_L     g03521(.A1(new_n429), .A2(new_n2982), .B1(new_n366), .B2(new_n3187), .C(new_n3777), .Y(new_n3778));
  XNOR2x2_ASAP7_75t_L       g03522(.A(\a[5] ), .B(new_n3778), .Y(new_n3779));
  OAI21xp33_ASAP7_75t_L     g03523(.A1(new_n3773), .A2(new_n3776), .B(new_n3779), .Y(new_n3780));
  NOR2xp33_ASAP7_75t_L      g03524(.A(new_n3530), .B(new_n3771), .Y(new_n3781));
  O2A1O1Ixp33_ASAP7_75t_L   g03525(.A1(new_n3540), .A2(new_n3541), .B(new_n3544), .C(new_n3781), .Y(new_n3782));
  NAND3xp33_ASAP7_75t_L     g03526(.A(new_n3782), .B(new_n3769), .C(new_n3765), .Y(new_n3783));
  A2O1A1Ixp33_ASAP7_75t_L   g03527(.A1(new_n3535), .A2(new_n3774), .B(new_n3551), .C(new_n3770), .Y(new_n3784));
  INVx1_ASAP7_75t_L         g03528(.A(new_n3779), .Y(new_n3785));
  NAND3xp33_ASAP7_75t_L     g03529(.A(new_n3783), .B(new_n3784), .C(new_n3785), .Y(new_n3786));
  NAND2xp33_ASAP7_75t_L     g03530(.A(new_n3780), .B(new_n3786), .Y(new_n3787));
  AND2x2_ASAP7_75t_L        g03531(.A(new_n3596), .B(new_n3787), .Y(new_n3788));
  INVx1_ASAP7_75t_L         g03532(.A(new_n3595), .Y(new_n3789));
  O2A1O1Ixp33_ASAP7_75t_L   g03533(.A1(new_n3559), .A2(new_n3557), .B(new_n3789), .C(new_n3787), .Y(new_n3790));
  NOR3xp33_ASAP7_75t_L      g03534(.A(new_n3788), .B(new_n3790), .C(new_n3594), .Y(new_n3791));
  INVx1_ASAP7_75t_L         g03535(.A(new_n3791), .Y(new_n3792));
  OAI21xp33_ASAP7_75t_L     g03536(.A1(new_n3790), .A2(new_n3788), .B(new_n3594), .Y(new_n3793));
  NAND2xp33_ASAP7_75t_L     g03537(.A(new_n3793), .B(new_n3792), .Y(new_n3794));
  O2A1O1Ixp33_ASAP7_75t_L   g03538(.A1(new_n3383), .A2(new_n3578), .B(new_n3576), .C(new_n3794), .Y(new_n3795));
  OAI21xp33_ASAP7_75t_L     g03539(.A1(new_n3578), .A2(new_n3383), .B(new_n3576), .Y(new_n3796));
  AOI21xp33_ASAP7_75t_L     g03540(.A1(new_n3792), .A2(new_n3793), .B(new_n3796), .Y(new_n3797));
  NOR2xp33_ASAP7_75t_L      g03541(.A(new_n3797), .B(new_n3795), .Y(\f[34] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03542(.A1(new_n3377), .A2(new_n3380), .B(new_n3375), .C(new_n3579), .Y(new_n3799));
  NOR2xp33_ASAP7_75t_L      g03543(.A(new_n3584), .B(new_n291), .Y(new_n3800));
  INVx1_ASAP7_75t_L         g03544(.A(new_n3800), .Y(new_n3801));
  INVx1_ASAP7_75t_L         g03545(.A(new_n3585), .Y(new_n3802));
  NOR2xp33_ASAP7_75t_L      g03546(.A(\b[34] ), .B(\b[35] ), .Y(new_n3803));
  INVx1_ASAP7_75t_L         g03547(.A(\b[35] ), .Y(new_n3804));
  NOR2xp33_ASAP7_75t_L      g03548(.A(new_n3584), .B(new_n3804), .Y(new_n3805));
  NOR2xp33_ASAP7_75t_L      g03549(.A(new_n3803), .B(new_n3805), .Y(new_n3806));
  INVx1_ASAP7_75t_L         g03550(.A(new_n3806), .Y(new_n3807));
  O2A1O1Ixp33_ASAP7_75t_L   g03551(.A1(new_n3589), .A2(new_n3588), .B(new_n3802), .C(new_n3807), .Y(new_n3808));
  O2A1O1Ixp33_ASAP7_75t_L   g03552(.A1(new_n3207), .A2(new_n3565), .B(new_n3568), .C(new_n3589), .Y(new_n3809));
  NOR3xp33_ASAP7_75t_L      g03553(.A(new_n3809), .B(new_n3806), .C(new_n3585), .Y(new_n3810));
  NOR2xp33_ASAP7_75t_L      g03554(.A(new_n3808), .B(new_n3810), .Y(new_n3811));
  NAND2xp33_ASAP7_75t_L     g03555(.A(new_n267), .B(new_n3811), .Y(new_n3812));
  AOI22xp33_ASAP7_75t_L     g03556(.A1(\b[33] ), .A2(new_n282), .B1(\b[35] ), .B2(new_n303), .Y(new_n3813));
  NAND4xp25_ASAP7_75t_L     g03557(.A(new_n3812), .B(\a[2] ), .C(new_n3801), .D(new_n3813), .Y(new_n3814));
  NAND2xp33_ASAP7_75t_L     g03558(.A(new_n3813), .B(new_n3812), .Y(new_n3815));
  A2O1A1Ixp33_ASAP7_75t_L   g03559(.A1(\b[34] ), .A2(new_n272), .B(new_n3815), .C(new_n262), .Y(new_n3816));
  AND2x2_ASAP7_75t_L        g03560(.A(new_n3814), .B(new_n3816), .Y(new_n3817));
  INVx1_ASAP7_75t_L         g03561(.A(new_n3780), .Y(new_n3818));
  AOI22xp33_ASAP7_75t_L     g03562(.A1(\b[24] ), .A2(new_n651), .B1(\b[26] ), .B2(new_n581), .Y(new_n3819));
  OAI221xp5_ASAP7_75t_L     g03563(.A1(new_n821), .A2(new_n2067), .B1(new_n577), .B2(new_n2355), .C(new_n3819), .Y(new_n3820));
  XNOR2x2_ASAP7_75t_L       g03564(.A(\a[11] ), .B(new_n3820), .Y(new_n3821));
  NOR3xp33_ASAP7_75t_L      g03565(.A(new_n3720), .B(new_n3725), .C(new_n3741), .Y(new_n3822));
  INVx1_ASAP7_75t_L         g03566(.A(new_n3822), .Y(new_n3823));
  AOI22xp33_ASAP7_75t_L     g03567(.A1(new_n811), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n900), .Y(new_n3824));
  OAI221xp5_ASAP7_75t_L     g03568(.A1(new_n904), .A2(new_n1774), .B1(new_n898), .B2(new_n1915), .C(new_n3824), .Y(new_n3825));
  XNOR2x2_ASAP7_75t_L       g03569(.A(new_n806), .B(new_n3825), .Y(new_n3826));
  INVx1_ASAP7_75t_L         g03570(.A(new_n3826), .Y(new_n3827));
  INVx1_ASAP7_75t_L         g03571(.A(new_n3716), .Y(new_n3828));
  NAND3xp33_ASAP7_75t_L     g03572(.A(new_n3828), .B(new_n3706), .C(new_n3702), .Y(new_n3829));
  A2O1A1Ixp33_ASAP7_75t_L   g03573(.A1(new_n3718), .A2(new_n3717), .B(new_n3736), .C(new_n3829), .Y(new_n3830));
  AOI22xp33_ASAP7_75t_L     g03574(.A1(new_n1704), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1837), .Y(new_n3831));
  OAI221xp5_ASAP7_75t_L     g03575(.A1(new_n1699), .A2(new_n784), .B1(new_n1827), .B2(new_n875), .C(new_n3831), .Y(new_n3832));
  XNOR2x2_ASAP7_75t_L       g03576(.A(\a[23] ), .B(new_n3832), .Y(new_n3833));
  NOR2xp33_ASAP7_75t_L      g03577(.A(new_n3669), .B(new_n3674), .Y(new_n3834));
  OAI21xp33_ASAP7_75t_L     g03578(.A1(new_n3446), .A2(new_n3444), .B(new_n3438), .Y(new_n3835));
  MAJIxp5_ASAP7_75t_L       g03579(.A(new_n3835), .B(new_n3675), .C(new_n3834), .Y(new_n3836));
  AOI22xp33_ASAP7_75t_L     g03580(.A1(new_n2114), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n2259), .Y(new_n3837));
  OAI221xp5_ASAP7_75t_L     g03581(.A1(new_n2109), .A2(new_n617), .B1(new_n2257), .B2(new_n685), .C(new_n3837), .Y(new_n3838));
  XNOR2x2_ASAP7_75t_L       g03582(.A(new_n2100), .B(new_n3838), .Y(new_n3839));
  A2O1A1O1Ixp25_ASAP7_75t_L g03583(.A1(new_n3431), .A2(new_n3433), .B(new_n3610), .C(new_n3652), .D(new_n3663), .Y(new_n3840));
  AOI22xp33_ASAP7_75t_L     g03584(.A1(new_n2552), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n2736), .Y(new_n3841));
  OAI221xp5_ASAP7_75t_L     g03585(.A1(new_n2547), .A2(new_n420), .B1(new_n2734), .B2(new_n494), .C(new_n3841), .Y(new_n3842));
  XNOR2x2_ASAP7_75t_L       g03586(.A(\a[29] ), .B(new_n3842), .Y(new_n3843));
  NAND2xp33_ASAP7_75t_L     g03587(.A(new_n3408), .B(new_n3616), .Y(new_n3844));
  A2O1A1Ixp33_ASAP7_75t_L   g03588(.A1(new_n3420), .A2(new_n3844), .B(new_n3643), .C(new_n3650), .Y(new_n3845));
  NOR2xp33_ASAP7_75t_L      g03589(.A(new_n324), .B(new_n3024), .Y(new_n3846));
  NOR3xp33_ASAP7_75t_L      g03590(.A(new_n357), .B(new_n358), .C(new_n3256), .Y(new_n3847));
  AOI22xp33_ASAP7_75t_L     g03591(.A1(new_n3029), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n3258), .Y(new_n3848));
  INVx1_ASAP7_75t_L         g03592(.A(new_n3848), .Y(new_n3849));
  NOR4xp25_ASAP7_75t_L      g03593(.A(new_n3849), .B(new_n3015), .C(new_n3846), .D(new_n3847), .Y(new_n3850));
  INVx1_ASAP7_75t_L         g03594(.A(new_n3850), .Y(new_n3851));
  OAI31xp33_ASAP7_75t_L     g03595(.A1(new_n3849), .A2(new_n3847), .A3(new_n3846), .B(new_n3015), .Y(new_n3852));
  OAI21xp33_ASAP7_75t_L     g03596(.A1(new_n3636), .A2(new_n3637), .B(new_n3407), .Y(new_n3853));
  NOR2xp33_ASAP7_75t_L      g03597(.A(new_n261), .B(new_n3853), .Y(new_n3854));
  INVx1_ASAP7_75t_L         g03598(.A(new_n3854), .Y(new_n3855));
  NAND2xp33_ASAP7_75t_L     g03599(.A(new_n3632), .B(new_n3635), .Y(new_n3856));
  NOR2xp33_ASAP7_75t_L      g03600(.A(new_n280), .B(new_n3856), .Y(new_n3857));
  AND3x1_ASAP7_75t_L        g03601(.A(new_n3407), .B(new_n3638), .C(new_n3632), .Y(new_n3858));
  AOI221xp5_ASAP7_75t_L     g03602(.A1(new_n3633), .A2(\b[2] ), .B1(new_n3858), .B2(\b[0] ), .C(new_n3857), .Y(new_n3859));
  NAND2xp33_ASAP7_75t_L     g03603(.A(new_n3855), .B(new_n3859), .Y(new_n3860));
  O2A1O1Ixp33_ASAP7_75t_L   g03604(.A1(new_n3408), .A2(new_n3641), .B(\a[35] ), .C(new_n3860), .Y(new_n3861));
  NAND5xp2_ASAP7_75t_L      g03605(.A(\a[35] ), .B(new_n3631), .C(new_n3634), .D(new_n3640), .E(new_n3412), .Y(new_n3862));
  NAND3xp33_ASAP7_75t_L     g03606(.A(new_n3860), .B(new_n3862), .C(\a[35] ), .Y(new_n3863));
  INVx1_ASAP7_75t_L         g03607(.A(new_n3863), .Y(new_n3864));
  OAI211xp5_ASAP7_75t_L     g03608(.A1(new_n3861), .A2(new_n3864), .B(new_n3852), .C(new_n3851), .Y(new_n3865));
  INVx1_ASAP7_75t_L         g03609(.A(new_n3852), .Y(new_n3866));
  INVx1_ASAP7_75t_L         g03610(.A(new_n3861), .Y(new_n3867));
  OAI211xp5_ASAP7_75t_L     g03611(.A1(new_n3866), .A2(new_n3850), .B(new_n3867), .C(new_n3863), .Y(new_n3868));
  AOI21xp33_ASAP7_75t_L     g03612(.A1(new_n3868), .A2(new_n3865), .B(new_n3845), .Y(new_n3869));
  NAND2xp33_ASAP7_75t_L     g03613(.A(new_n3868), .B(new_n3865), .Y(new_n3870));
  O2A1O1Ixp33_ASAP7_75t_L   g03614(.A1(new_n3618), .A2(new_n3643), .B(new_n3650), .C(new_n3870), .Y(new_n3871));
  NOR3xp33_ASAP7_75t_L      g03615(.A(new_n3871), .B(new_n3869), .C(new_n3843), .Y(new_n3872));
  INVx1_ASAP7_75t_L         g03616(.A(new_n3843), .Y(new_n3873));
  A2O1A1O1Ixp25_ASAP7_75t_L g03617(.A1(new_n3616), .A2(new_n3408), .B(new_n3648), .C(new_n3649), .D(new_n3646), .Y(new_n3874));
  NAND2xp33_ASAP7_75t_L     g03618(.A(new_n3874), .B(new_n3870), .Y(new_n3875));
  NAND3xp33_ASAP7_75t_L     g03619(.A(new_n3845), .B(new_n3865), .C(new_n3868), .Y(new_n3876));
  AOI21xp33_ASAP7_75t_L     g03620(.A1(new_n3876), .A2(new_n3875), .B(new_n3873), .Y(new_n3877));
  NOR3xp33_ASAP7_75t_L      g03621(.A(new_n3840), .B(new_n3872), .C(new_n3877), .Y(new_n3878));
  OAI221xp5_ASAP7_75t_L     g03622(.A1(new_n3659), .A2(new_n3660), .B1(new_n3670), .B2(new_n3245), .C(new_n3264), .Y(new_n3879));
  A2O1A1Ixp33_ASAP7_75t_L   g03623(.A1(new_n3879), .A2(new_n3672), .B(new_n3662), .C(new_n3657), .Y(new_n3880));
  NAND3xp33_ASAP7_75t_L     g03624(.A(new_n3873), .B(new_n3875), .C(new_n3876), .Y(new_n3881));
  OAI21xp33_ASAP7_75t_L     g03625(.A1(new_n3869), .A2(new_n3871), .B(new_n3843), .Y(new_n3882));
  AOI21xp33_ASAP7_75t_L     g03626(.A1(new_n3882), .A2(new_n3881), .B(new_n3880), .Y(new_n3883));
  OAI21xp33_ASAP7_75t_L     g03627(.A1(new_n3878), .A2(new_n3883), .B(new_n3839), .Y(new_n3884));
  XNOR2x2_ASAP7_75t_L       g03628(.A(\a[26] ), .B(new_n3838), .Y(new_n3885));
  NAND3xp33_ASAP7_75t_L     g03629(.A(new_n3880), .B(new_n3881), .C(new_n3882), .Y(new_n3886));
  OAI21xp33_ASAP7_75t_L     g03630(.A1(new_n3872), .A2(new_n3877), .B(new_n3840), .Y(new_n3887));
  NAND3xp33_ASAP7_75t_L     g03631(.A(new_n3886), .B(new_n3885), .C(new_n3887), .Y(new_n3888));
  AOI21xp33_ASAP7_75t_L     g03632(.A1(new_n3888), .A2(new_n3884), .B(new_n3836), .Y(new_n3889));
  NAND2xp33_ASAP7_75t_L     g03633(.A(new_n3658), .B(new_n3664), .Y(new_n3890));
  MAJIxp5_ASAP7_75t_L       g03634(.A(new_n3677), .B(new_n3667), .C(new_n3890), .Y(new_n3891));
  NAND2xp33_ASAP7_75t_L     g03635(.A(new_n3888), .B(new_n3884), .Y(new_n3892));
  NOR2xp33_ASAP7_75t_L      g03636(.A(new_n3891), .B(new_n3892), .Y(new_n3893));
  OAI21xp33_ASAP7_75t_L     g03637(.A1(new_n3893), .A2(new_n3889), .B(new_n3833), .Y(new_n3894));
  XNOR2x2_ASAP7_75t_L       g03638(.A(new_n1689), .B(new_n3832), .Y(new_n3895));
  NAND2xp33_ASAP7_75t_L     g03639(.A(new_n3891), .B(new_n3892), .Y(new_n3896));
  NAND2xp33_ASAP7_75t_L     g03640(.A(new_n3675), .B(new_n3834), .Y(new_n3897));
  NAND4xp25_ASAP7_75t_L     g03641(.A(new_n3690), .B(new_n3888), .C(new_n3884), .D(new_n3897), .Y(new_n3898));
  NAND3xp33_ASAP7_75t_L     g03642(.A(new_n3898), .B(new_n3896), .C(new_n3895), .Y(new_n3899));
  NOR2xp33_ASAP7_75t_L      g03643(.A(new_n3288), .B(new_n3290), .Y(new_n3900));
  OAI311xp33_ASAP7_75t_L    g03644(.A1(new_n3900), .A2(new_n3284), .A3(new_n3462), .B1(new_n3459), .C1(new_n3692), .Y(new_n3901));
  NAND4xp25_ASAP7_75t_L     g03645(.A(new_n3894), .B(new_n3901), .C(new_n3899), .D(new_n3688), .Y(new_n3902));
  INVx1_ASAP7_75t_L         g03646(.A(new_n3688), .Y(new_n3903));
  AOI21xp33_ASAP7_75t_L     g03647(.A1(new_n3898), .A2(new_n3896), .B(new_n3895), .Y(new_n3904));
  NOR3xp33_ASAP7_75t_L      g03648(.A(new_n3889), .B(new_n3893), .C(new_n3833), .Y(new_n3905));
  NOR3xp33_ASAP7_75t_L      g03649(.A(new_n3678), .B(new_n3687), .C(new_n3679), .Y(new_n3906));
  AOI311xp33_ASAP7_75t_L    g03650(.A1(new_n3291), .A2(new_n3460), .A3(new_n3455), .B(new_n3463), .C(new_n3906), .Y(new_n3907));
  OAI22xp33_ASAP7_75t_L     g03651(.A1(new_n3907), .A2(new_n3903), .B1(new_n3904), .B2(new_n3905), .Y(new_n3908));
  NAND2xp33_ASAP7_75t_L     g03652(.A(\b[16] ), .B(new_n1362), .Y(new_n3909));
  NAND3xp33_ASAP7_75t_L     g03653(.A(new_n1206), .B(new_n1208), .C(new_n1365), .Y(new_n3910));
  AOI22xp33_ASAP7_75t_L     g03654(.A1(new_n1360), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1581), .Y(new_n3911));
  NAND4xp25_ASAP7_75t_L     g03655(.A(new_n3910), .B(\a[20] ), .C(new_n3909), .D(new_n3911), .Y(new_n3912));
  INVx1_ASAP7_75t_L         g03656(.A(new_n3912), .Y(new_n3913));
  AOI31xp33_ASAP7_75t_L     g03657(.A1(new_n3910), .A2(new_n3909), .A3(new_n3911), .B(\a[20] ), .Y(new_n3914));
  NOR2xp33_ASAP7_75t_L      g03658(.A(new_n3914), .B(new_n3913), .Y(new_n3915));
  NAND3xp33_ASAP7_75t_L     g03659(.A(new_n3908), .B(new_n3915), .C(new_n3902), .Y(new_n3916));
  NOR4xp25_ASAP7_75t_L      g03660(.A(new_n3907), .B(new_n3905), .C(new_n3904), .D(new_n3903), .Y(new_n3917));
  AOI22xp33_ASAP7_75t_L     g03661(.A1(new_n3901), .A2(new_n3688), .B1(new_n3899), .B2(new_n3894), .Y(new_n3918));
  INVx1_ASAP7_75t_L         g03662(.A(new_n3914), .Y(new_n3919));
  NAND2xp33_ASAP7_75t_L     g03663(.A(new_n3912), .B(new_n3919), .Y(new_n3920));
  OAI21xp33_ASAP7_75t_L     g03664(.A1(new_n3918), .A2(new_n3917), .B(new_n3920), .Y(new_n3921));
  INVx1_ASAP7_75t_L         g03665(.A(new_n3604), .Y(new_n3922));
  A2O1A1O1Ixp25_ASAP7_75t_L g03666(.A1(new_n3398), .A2(new_n3479), .B(new_n3922), .C(new_n3705), .D(new_n3697), .Y(new_n3923));
  NAND3xp33_ASAP7_75t_L     g03667(.A(new_n3923), .B(new_n3921), .C(new_n3916), .Y(new_n3924));
  NAND2xp33_ASAP7_75t_L     g03668(.A(new_n3916), .B(new_n3921), .Y(new_n3925));
  A2O1A1Ixp33_ASAP7_75t_L   g03669(.A1(new_n3705), .A2(new_n3703), .B(new_n3697), .C(new_n3925), .Y(new_n3926));
  NOR2xp33_ASAP7_75t_L      g03670(.A(new_n1432), .B(new_n1154), .Y(new_n3927));
  AOI22xp33_ASAP7_75t_L     g03671(.A1(new_n1076), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1253), .Y(new_n3928));
  OAI31xp33_ASAP7_75t_L     g03672(.A1(new_n1885), .A2(new_n1156), .A3(new_n1543), .B(new_n3928), .Y(new_n3929));
  OR3x1_ASAP7_75t_L         g03673(.A(new_n3929), .B(new_n1071), .C(new_n3927), .Y(new_n3930));
  A2O1A1Ixp33_ASAP7_75t_L   g03674(.A1(\b[19] ), .A2(new_n1080), .B(new_n3929), .C(new_n1071), .Y(new_n3931));
  NAND2xp33_ASAP7_75t_L     g03675(.A(new_n3931), .B(new_n3930), .Y(new_n3932));
  AOI21xp33_ASAP7_75t_L     g03676(.A1(new_n3926), .A2(new_n3924), .B(new_n3932), .Y(new_n3933));
  AO21x2_ASAP7_75t_L        g03677(.A1(new_n3705), .A2(new_n3703), .B(new_n3697), .Y(new_n3934));
  NOR2xp33_ASAP7_75t_L      g03678(.A(new_n3925), .B(new_n3934), .Y(new_n3935));
  AND2x2_ASAP7_75t_L        g03679(.A(new_n3916), .B(new_n3921), .Y(new_n3936));
  NOR2xp33_ASAP7_75t_L      g03680(.A(new_n3923), .B(new_n3936), .Y(new_n3937));
  AND2x2_ASAP7_75t_L        g03681(.A(new_n3931), .B(new_n3930), .Y(new_n3938));
  NOR3xp33_ASAP7_75t_L      g03682(.A(new_n3937), .B(new_n3935), .C(new_n3938), .Y(new_n3939));
  NOR2xp33_ASAP7_75t_L      g03683(.A(new_n3933), .B(new_n3939), .Y(new_n3940));
  NOR2xp33_ASAP7_75t_L      g03684(.A(new_n3940), .B(new_n3830), .Y(new_n3941));
  OAI21xp33_ASAP7_75t_L     g03685(.A1(new_n3935), .A2(new_n3937), .B(new_n3938), .Y(new_n3942));
  NAND3xp33_ASAP7_75t_L     g03686(.A(new_n3926), .B(new_n3924), .C(new_n3932), .Y(new_n3943));
  NAND2xp33_ASAP7_75t_L     g03687(.A(new_n3943), .B(new_n3942), .Y(new_n3944));
  O2A1O1Ixp33_ASAP7_75t_L   g03688(.A1(new_n3724), .A2(new_n3736), .B(new_n3829), .C(new_n3944), .Y(new_n3945));
  OAI21xp33_ASAP7_75t_L     g03689(.A1(new_n3941), .A2(new_n3945), .B(new_n3827), .Y(new_n3946));
  INVx1_ASAP7_75t_L         g03690(.A(new_n3829), .Y(new_n3947));
  A2O1A1O1Ixp25_ASAP7_75t_L g03691(.A1(new_n3738), .A2(new_n3504), .B(new_n3502), .C(new_n3719), .D(new_n3947), .Y(new_n3948));
  NAND2xp33_ASAP7_75t_L     g03692(.A(new_n3944), .B(new_n3948), .Y(new_n3949));
  NAND2xp33_ASAP7_75t_L     g03693(.A(new_n3940), .B(new_n3830), .Y(new_n3950));
  NAND3xp33_ASAP7_75t_L     g03694(.A(new_n3949), .B(new_n3950), .C(new_n3826), .Y(new_n3951));
  NAND2xp33_ASAP7_75t_L     g03695(.A(new_n3951), .B(new_n3946), .Y(new_n3952));
  AOI21xp33_ASAP7_75t_L     g03696(.A1(new_n3750), .A2(new_n3823), .B(new_n3952), .Y(new_n3953));
  AOI211xp5_ASAP7_75t_L     g03697(.A1(new_n3946), .A2(new_n3951), .B(new_n3822), .C(new_n3758), .Y(new_n3954));
  OAI21xp33_ASAP7_75t_L     g03698(.A1(new_n3954), .A2(new_n3953), .B(new_n3821), .Y(new_n3955));
  INVx1_ASAP7_75t_L         g03699(.A(new_n3821), .Y(new_n3956));
  A2O1A1Ixp33_ASAP7_75t_L   g03700(.A1(new_n3745), .A2(new_n3508), .B(new_n3743), .C(new_n3823), .Y(new_n3957));
  AOI21xp33_ASAP7_75t_L     g03701(.A1(new_n3949), .A2(new_n3950), .B(new_n3826), .Y(new_n3958));
  NOR3xp33_ASAP7_75t_L      g03702(.A(new_n3827), .B(new_n3945), .C(new_n3941), .Y(new_n3959));
  NOR2xp33_ASAP7_75t_L      g03703(.A(new_n3958), .B(new_n3959), .Y(new_n3960));
  NAND2xp33_ASAP7_75t_L     g03704(.A(new_n3960), .B(new_n3957), .Y(new_n3961));
  NAND3xp33_ASAP7_75t_L     g03705(.A(new_n3952), .B(new_n3750), .C(new_n3823), .Y(new_n3962));
  NAND3xp33_ASAP7_75t_L     g03706(.A(new_n3961), .B(new_n3962), .C(new_n3956), .Y(new_n3963));
  AOI211xp5_ASAP7_75t_L     g03707(.A1(new_n3746), .A2(new_n3750), .B(new_n3753), .C(new_n3754), .Y(new_n3964));
  OAI21xp33_ASAP7_75t_L     g03708(.A1(new_n3964), .A2(new_n3600), .B(new_n3755), .Y(new_n3965));
  NAND3xp33_ASAP7_75t_L     g03709(.A(new_n3965), .B(new_n3963), .C(new_n3955), .Y(new_n3966));
  AOI21xp33_ASAP7_75t_L     g03710(.A1(new_n3961), .A2(new_n3962), .B(new_n3956), .Y(new_n3967));
  NOR3xp33_ASAP7_75t_L      g03711(.A(new_n3953), .B(new_n3954), .C(new_n3821), .Y(new_n3968));
  NOR3xp33_ASAP7_75t_L      g03712(.A(new_n3757), .B(new_n3759), .C(new_n3758), .Y(new_n3969));
  A2O1A1O1Ixp25_ASAP7_75t_L g03713(.A1(new_n3524), .A2(new_n3533), .B(new_n3520), .C(new_n3760), .D(new_n3969), .Y(new_n3970));
  OAI21xp33_ASAP7_75t_L     g03714(.A1(new_n3967), .A2(new_n3968), .B(new_n3970), .Y(new_n3971));
  AOI22xp33_ASAP7_75t_L     g03715(.A1(new_n444), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n471), .Y(new_n3972));
  OAI221xp5_ASAP7_75t_L     g03716(.A1(new_n468), .A2(new_n2666), .B1(new_n469), .B2(new_n2695), .C(new_n3972), .Y(new_n3973));
  XNOR2x2_ASAP7_75t_L       g03717(.A(\a[8] ), .B(new_n3973), .Y(new_n3974));
  NAND3xp33_ASAP7_75t_L     g03718(.A(new_n3966), .B(new_n3971), .C(new_n3974), .Y(new_n3975));
  NOR3xp33_ASAP7_75t_L      g03719(.A(new_n3970), .B(new_n3968), .C(new_n3967), .Y(new_n3976));
  AOI221xp5_ASAP7_75t_L     g03720(.A1(new_n3763), .A2(new_n3760), .B1(new_n3955), .B2(new_n3963), .C(new_n3969), .Y(new_n3977));
  INVx1_ASAP7_75t_L         g03721(.A(new_n3974), .Y(new_n3978));
  OAI21xp33_ASAP7_75t_L     g03722(.A1(new_n3977), .A2(new_n3976), .B(new_n3978), .Y(new_n3979));
  NAND2xp33_ASAP7_75t_L     g03723(.A(new_n3979), .B(new_n3975), .Y(new_n3980));
  NOR2xp33_ASAP7_75t_L      g03724(.A(new_n3767), .B(new_n3768), .Y(new_n3981));
  NAND2xp33_ASAP7_75t_L     g03725(.A(new_n3766), .B(new_n3981), .Y(new_n3982));
  A2O1A1Ixp33_ASAP7_75t_L   g03726(.A1(new_n3769), .A2(new_n3765), .B(new_n3782), .C(new_n3982), .Y(new_n3983));
  NOR2xp33_ASAP7_75t_L      g03727(.A(new_n3980), .B(new_n3983), .Y(new_n3984));
  NOR3xp33_ASAP7_75t_L      g03728(.A(new_n3976), .B(new_n3977), .C(new_n3978), .Y(new_n3985));
  AOI21xp33_ASAP7_75t_L     g03729(.A1(new_n3966), .A2(new_n3971), .B(new_n3974), .Y(new_n3986));
  NOR2xp33_ASAP7_75t_L      g03730(.A(new_n3985), .B(new_n3986), .Y(new_n3987));
  A2O1A1O1Ixp25_ASAP7_75t_L g03731(.A1(new_n3769), .A2(new_n3765), .B(new_n3782), .C(new_n3982), .D(new_n3987), .Y(new_n3988));
  NOR2xp33_ASAP7_75t_L      g03732(.A(new_n3180), .B(new_n429), .Y(new_n3989));
  INVx1_ASAP7_75t_L         g03733(.A(new_n3989), .Y(new_n3990));
  NAND3xp33_ASAP7_75t_L     g03734(.A(new_n3210), .B(new_n341), .C(new_n3213), .Y(new_n3991));
  AOI22xp33_ASAP7_75t_L     g03735(.A1(new_n344), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n370), .Y(new_n3992));
  AND4x1_ASAP7_75t_L        g03736(.A(new_n3992), .B(new_n3991), .C(new_n3990), .D(\a[5] ), .Y(new_n3993));
  AOI31xp33_ASAP7_75t_L     g03737(.A1(new_n3991), .A2(new_n3990), .A3(new_n3992), .B(\a[5] ), .Y(new_n3994));
  NOR2xp33_ASAP7_75t_L      g03738(.A(new_n3994), .B(new_n3993), .Y(new_n3995));
  OAI21xp33_ASAP7_75t_L     g03739(.A1(new_n3988), .A2(new_n3984), .B(new_n3995), .Y(new_n3996));
  MAJIxp5_ASAP7_75t_L       g03740(.A(new_n3772), .B(new_n3766), .C(new_n3981), .Y(new_n3997));
  NAND2xp33_ASAP7_75t_L     g03741(.A(new_n3987), .B(new_n3997), .Y(new_n3998));
  INVx1_ASAP7_75t_L         g03742(.A(new_n3981), .Y(new_n3999));
  NOR2xp33_ASAP7_75t_L      g03743(.A(new_n3599), .B(new_n3999), .Y(new_n4000));
  A2O1A1Ixp33_ASAP7_75t_L   g03744(.A1(new_n3770), .A2(new_n3772), .B(new_n4000), .C(new_n3980), .Y(new_n4001));
  INVx1_ASAP7_75t_L         g03745(.A(new_n3995), .Y(new_n4002));
  NAND3xp33_ASAP7_75t_L     g03746(.A(new_n4001), .B(new_n3998), .C(new_n4002), .Y(new_n4003));
  NOR2xp33_ASAP7_75t_L      g03747(.A(new_n3773), .B(new_n3776), .Y(new_n4004));
  AOI221xp5_ASAP7_75t_L     g03748(.A1(new_n3561), .A2(new_n3554), .B1(new_n3785), .B2(new_n4004), .C(new_n3595), .Y(new_n4005));
  OAI211xp5_ASAP7_75t_L     g03749(.A1(new_n3818), .A2(new_n4005), .B(new_n3996), .C(new_n4003), .Y(new_n4006));
  AOI21xp33_ASAP7_75t_L     g03750(.A1(new_n4001), .A2(new_n3998), .B(new_n4002), .Y(new_n4007));
  NOR3xp33_ASAP7_75t_L      g03751(.A(new_n3984), .B(new_n3988), .C(new_n3995), .Y(new_n4008));
  OAI211xp5_ASAP7_75t_L     g03752(.A1(new_n3557), .A2(new_n3559), .B(new_n3789), .C(new_n3786), .Y(new_n4009));
  OAI211xp5_ASAP7_75t_L     g03753(.A1(new_n4007), .A2(new_n4008), .B(new_n4009), .C(new_n3780), .Y(new_n4010));
  AOI21xp33_ASAP7_75t_L     g03754(.A1(new_n4006), .A2(new_n4010), .B(new_n3817), .Y(new_n4011));
  INVx1_ASAP7_75t_L         g03755(.A(new_n4011), .Y(new_n4012));
  NAND3xp33_ASAP7_75t_L     g03756(.A(new_n4006), .B(new_n4010), .C(new_n3817), .Y(new_n4013));
  NAND2xp33_ASAP7_75t_L     g03757(.A(new_n4013), .B(new_n4012), .Y(new_n4014));
  A2O1A1O1Ixp25_ASAP7_75t_L g03758(.A1(new_n3799), .A2(new_n3576), .B(new_n3794), .C(new_n3792), .D(new_n4014), .Y(new_n4015));
  A2O1A1Ixp33_ASAP7_75t_L   g03759(.A1(new_n3799), .A2(new_n3576), .B(new_n3794), .C(new_n3792), .Y(new_n4016));
  AOI21xp33_ASAP7_75t_L     g03760(.A1(new_n4013), .A2(new_n4012), .B(new_n4016), .Y(new_n4017));
  NOR2xp33_ASAP7_75t_L      g03761(.A(new_n4015), .B(new_n4017), .Y(\f[35] ));
  AOI22xp33_ASAP7_75t_L     g03762(.A1(new_n344), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n370), .Y(new_n4019));
  OAI221xp5_ASAP7_75t_L     g03763(.A1(new_n429), .A2(new_n3207), .B1(new_n366), .B2(new_n3572), .C(new_n4019), .Y(new_n4020));
  XNOR2x2_ASAP7_75t_L       g03764(.A(\a[5] ), .B(new_n4020), .Y(new_n4021));
  INVx1_ASAP7_75t_L         g03765(.A(new_n4021), .Y(new_n4022));
  NOR3xp33_ASAP7_75t_L      g03766(.A(new_n3976), .B(new_n3977), .C(new_n3974), .Y(new_n4023));
  NOR2xp33_ASAP7_75t_L      g03767(.A(new_n2688), .B(new_n468), .Y(new_n4024));
  INVx1_ASAP7_75t_L         g03768(.A(new_n4024), .Y(new_n4025));
  NAND2xp33_ASAP7_75t_L     g03769(.A(new_n441), .B(new_n2989), .Y(new_n4026));
  AOI22xp33_ASAP7_75t_L     g03770(.A1(new_n444), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n471), .Y(new_n4027));
  AND4x1_ASAP7_75t_L        g03771(.A(new_n4027), .B(new_n4026), .C(new_n4025), .D(\a[8] ), .Y(new_n4028));
  AOI31xp33_ASAP7_75t_L     g03772(.A1(new_n4026), .A2(new_n4025), .A3(new_n4027), .B(\a[8] ), .Y(new_n4029));
  NOR2xp33_ASAP7_75t_L      g03773(.A(new_n4029), .B(new_n4028), .Y(new_n4030));
  INVx1_ASAP7_75t_L         g03774(.A(new_n4030), .Y(new_n4031));
  OAI21xp33_ASAP7_75t_L     g03775(.A1(new_n3967), .A2(new_n3970), .B(new_n3963), .Y(new_n4032));
  NAND2xp33_ASAP7_75t_L     g03776(.A(\b[23] ), .B(new_n815), .Y(new_n4033));
  OR3x1_ASAP7_75t_L         g03777(.A(new_n1934), .B(new_n898), .C(new_n1933), .Y(new_n4034));
  AOI22xp33_ASAP7_75t_L     g03778(.A1(new_n811), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n900), .Y(new_n4035));
  NAND4xp25_ASAP7_75t_L     g03779(.A(new_n4034), .B(\a[14] ), .C(new_n4033), .D(new_n4035), .Y(new_n4036));
  OAI31xp33_ASAP7_75t_L     g03780(.A1(new_n1934), .A2(new_n898), .A3(new_n1933), .B(new_n4035), .Y(new_n4037));
  A2O1A1Ixp33_ASAP7_75t_L   g03781(.A1(\b[23] ), .A2(new_n815), .B(new_n4037), .C(new_n806), .Y(new_n4038));
  NAND2xp33_ASAP7_75t_L     g03782(.A(new_n4038), .B(new_n4036), .Y(new_n4039));
  NOR3xp33_ASAP7_75t_L      g03783(.A(new_n3917), .B(new_n3918), .C(new_n3915), .Y(new_n4040));
  INVx1_ASAP7_75t_L         g03784(.A(new_n4040), .Y(new_n4041));
  A2O1A1Ixp33_ASAP7_75t_L   g03785(.A1(new_n3921), .A2(new_n3916), .B(new_n3923), .C(new_n4041), .Y(new_n4042));
  AOI22xp33_ASAP7_75t_L     g03786(.A1(new_n1360), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n1581), .Y(new_n4043));
  OAI31xp33_ASAP7_75t_L     g03787(.A1(new_n1318), .A2(new_n1317), .A3(new_n1359), .B(new_n4043), .Y(new_n4044));
  AOI21xp33_ASAP7_75t_L     g03788(.A1(new_n1362), .A2(\b[17] ), .B(new_n4044), .Y(new_n4045));
  NAND2xp33_ASAP7_75t_L     g03789(.A(\a[20] ), .B(new_n4045), .Y(new_n4046));
  A2O1A1Ixp33_ASAP7_75t_L   g03790(.A1(\b[17] ), .A2(new_n1362), .B(new_n4044), .C(new_n1356), .Y(new_n4047));
  NAND2xp33_ASAP7_75t_L     g03791(.A(new_n4047), .B(new_n4046), .Y(new_n4048));
  OAI31xp33_ASAP7_75t_L     g03792(.A1(new_n3907), .A2(new_n3904), .A3(new_n3903), .B(new_n3899), .Y(new_n4049));
  OAI21xp33_ASAP7_75t_L     g03793(.A1(new_n3877), .A2(new_n3840), .B(new_n3881), .Y(new_n4050));
  NAND2xp33_ASAP7_75t_L     g03794(.A(\b[2] ), .B(new_n3633), .Y(new_n4051));
  NAND3xp33_ASAP7_75t_L     g03795(.A(new_n3407), .B(new_n3632), .C(new_n3638), .Y(new_n4052));
  OAI221xp5_ASAP7_75t_L     g03796(.A1(new_n258), .A2(new_n4052), .B1(new_n280), .B2(new_n3856), .C(new_n4051), .Y(new_n4053));
  INVx1_ASAP7_75t_L         g03797(.A(\a[36] ), .Y(new_n4054));
  NAND2xp33_ASAP7_75t_L     g03798(.A(\a[35] ), .B(new_n4054), .Y(new_n4055));
  NAND2xp33_ASAP7_75t_L     g03799(.A(\a[36] ), .B(new_n3628), .Y(new_n4056));
  NAND2xp33_ASAP7_75t_L     g03800(.A(new_n4056), .B(new_n4055), .Y(new_n4057));
  NAND2xp33_ASAP7_75t_L     g03801(.A(\b[0] ), .B(new_n4057), .Y(new_n4058));
  INVx1_ASAP7_75t_L         g03802(.A(new_n4058), .Y(new_n4059));
  OAI31xp33_ASAP7_75t_L     g03803(.A1(new_n3862), .A2(new_n4053), .A3(new_n3854), .B(new_n4059), .Y(new_n4060));
  NAND3xp33_ASAP7_75t_L     g03804(.A(new_n3635), .B(new_n3627), .C(new_n3629), .Y(new_n4061));
  OAI22xp33_ASAP7_75t_L     g03805(.A1(new_n3853), .A2(new_n258), .B1(new_n261), .B2(new_n4061), .Y(new_n4062));
  A2O1A1Ixp33_ASAP7_75t_L   g03806(.A1(new_n3405), .A2(new_n3406), .B(new_n258), .C(\a[35] ), .Y(new_n4063));
  AOI211xp5_ASAP7_75t_L     g03807(.A1(new_n3630), .A2(new_n269), .B(new_n4063), .C(new_n4062), .Y(new_n4064));
  NAND4xp25_ASAP7_75t_L     g03808(.A(new_n4064), .B(new_n4058), .C(new_n3859), .D(new_n3855), .Y(new_n4065));
  NAND2xp33_ASAP7_75t_L     g03809(.A(\b[2] ), .B(new_n3639), .Y(new_n4066));
  NAND2xp33_ASAP7_75t_L     g03810(.A(new_n3630), .B(new_n406), .Y(new_n4067));
  AOI22xp33_ASAP7_75t_L     g03811(.A1(new_n3633), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n3858), .Y(new_n4068));
  NAND4xp25_ASAP7_75t_L     g03812(.A(new_n4067), .B(\a[35] ), .C(new_n4068), .D(new_n4066), .Y(new_n4069));
  OAI21xp33_ASAP7_75t_L     g03813(.A1(new_n302), .A2(new_n3856), .B(new_n4068), .Y(new_n4070));
  A2O1A1Ixp33_ASAP7_75t_L   g03814(.A1(\b[2] ), .A2(new_n3639), .B(new_n4070), .C(new_n3628), .Y(new_n4071));
  AO22x1_ASAP7_75t_L        g03815(.A1(new_n4065), .A2(new_n4060), .B1(new_n4069), .B2(new_n4071), .Y(new_n4072));
  NAND4xp25_ASAP7_75t_L     g03816(.A(new_n4071), .B(new_n4060), .C(new_n4065), .D(new_n4069), .Y(new_n4073));
  NAND2xp33_ASAP7_75t_L     g03817(.A(\b[5] ), .B(new_n3030), .Y(new_n4074));
  NAND2xp33_ASAP7_75t_L     g03818(.A(new_n3021), .B(new_n526), .Y(new_n4075));
  AOI22xp33_ASAP7_75t_L     g03819(.A1(new_n3029), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n3258), .Y(new_n4076));
  NAND4xp25_ASAP7_75t_L     g03820(.A(new_n4075), .B(\a[32] ), .C(new_n4074), .D(new_n4076), .Y(new_n4077));
  OAI21xp33_ASAP7_75t_L     g03821(.A1(new_n3256), .A2(new_n390), .B(new_n4076), .Y(new_n4078));
  A2O1A1Ixp33_ASAP7_75t_L   g03822(.A1(\b[5] ), .A2(new_n3030), .B(new_n4078), .C(new_n3015), .Y(new_n4079));
  NAND4xp25_ASAP7_75t_L     g03823(.A(new_n4079), .B(new_n4072), .C(new_n4073), .D(new_n4077), .Y(new_n4080));
  AO22x1_ASAP7_75t_L        g03824(.A1(new_n4073), .A2(new_n4072), .B1(new_n4079), .B2(new_n4077), .Y(new_n4081));
  OAI211xp5_ASAP7_75t_L     g03825(.A1(new_n3618), .A2(new_n3643), .B(new_n3868), .C(new_n3650), .Y(new_n4082));
  AND4x1_ASAP7_75t_L        g03826(.A(new_n4082), .B(new_n4081), .C(new_n4080), .D(new_n3865), .Y(new_n4083));
  AOI211xp5_ASAP7_75t_L     g03827(.A1(new_n3867), .A2(new_n3863), .B(new_n3866), .C(new_n3850), .Y(new_n4084));
  AOI21xp33_ASAP7_75t_L     g03828(.A1(new_n3874), .A2(new_n3868), .B(new_n4084), .Y(new_n4085));
  AOI21xp33_ASAP7_75t_L     g03829(.A1(new_n4081), .A2(new_n4080), .B(new_n4085), .Y(new_n4086));
  AOI22xp33_ASAP7_75t_L     g03830(.A1(new_n2552), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n2736), .Y(new_n4087));
  OAI221xp5_ASAP7_75t_L     g03831(.A1(new_n2547), .A2(new_n488), .B1(new_n2734), .B2(new_n548), .C(new_n4087), .Y(new_n4088));
  NOR2xp33_ASAP7_75t_L      g03832(.A(new_n2538), .B(new_n4088), .Y(new_n4089));
  INVx1_ASAP7_75t_L         g03833(.A(new_n4087), .Y(new_n4090));
  AOI221xp5_ASAP7_75t_L     g03834(.A1(new_n2553), .A2(\b[8] ), .B1(new_n2544), .B2(new_n731), .C(new_n4090), .Y(new_n4091));
  NOR2xp33_ASAP7_75t_L      g03835(.A(\a[29] ), .B(new_n4091), .Y(new_n4092));
  OAI22xp33_ASAP7_75t_L     g03836(.A1(new_n4086), .A2(new_n4083), .B1(new_n4092), .B2(new_n4089), .Y(new_n4093));
  NAND4xp25_ASAP7_75t_L     g03837(.A(new_n4082), .B(new_n3865), .C(new_n4080), .D(new_n4081), .Y(new_n4094));
  NAND2xp33_ASAP7_75t_L     g03838(.A(new_n4080), .B(new_n4081), .Y(new_n4095));
  AOI211xp5_ASAP7_75t_L     g03839(.A1(new_n3851), .A2(new_n3852), .B(new_n3861), .C(new_n3864), .Y(new_n4096));
  OAI21xp33_ASAP7_75t_L     g03840(.A1(new_n4096), .A2(new_n3845), .B(new_n3865), .Y(new_n4097));
  NAND2xp33_ASAP7_75t_L     g03841(.A(new_n4097), .B(new_n4095), .Y(new_n4098));
  NAND2xp33_ASAP7_75t_L     g03842(.A(\a[29] ), .B(new_n4091), .Y(new_n4099));
  NAND2xp33_ASAP7_75t_L     g03843(.A(new_n2538), .B(new_n4088), .Y(new_n4100));
  NAND4xp25_ASAP7_75t_L     g03844(.A(new_n4098), .B(new_n4099), .C(new_n4100), .D(new_n4094), .Y(new_n4101));
  AOI21xp33_ASAP7_75t_L     g03845(.A1(new_n4101), .A2(new_n4093), .B(new_n4050), .Y(new_n4102));
  A2O1A1O1Ixp25_ASAP7_75t_L g03846(.A1(new_n3652), .A2(new_n3673), .B(new_n3663), .C(new_n3882), .D(new_n3872), .Y(new_n4103));
  NAND2xp33_ASAP7_75t_L     g03847(.A(new_n4101), .B(new_n4093), .Y(new_n4104));
  NOR2xp33_ASAP7_75t_L      g03848(.A(new_n4103), .B(new_n4104), .Y(new_n4105));
  NOR2xp33_ASAP7_75t_L      g03849(.A(new_n679), .B(new_n2109), .Y(new_n4106));
  AOI22xp33_ASAP7_75t_L     g03850(.A1(new_n2114), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n2259), .Y(new_n4107));
  OAI31xp33_ASAP7_75t_L     g03851(.A1(new_n1231), .A2(new_n764), .A3(new_n2257), .B(new_n4107), .Y(new_n4108));
  OR3x1_ASAP7_75t_L         g03852(.A(new_n4108), .B(new_n2100), .C(new_n4106), .Y(new_n4109));
  A2O1A1Ixp33_ASAP7_75t_L   g03853(.A1(\b[11] ), .A2(new_n2115), .B(new_n4108), .C(new_n2100), .Y(new_n4110));
  AND2x2_ASAP7_75t_L        g03854(.A(new_n4110), .B(new_n4109), .Y(new_n4111));
  OAI21xp33_ASAP7_75t_L     g03855(.A1(new_n4102), .A2(new_n4105), .B(new_n4111), .Y(new_n4112));
  NAND2xp33_ASAP7_75t_L     g03856(.A(new_n4103), .B(new_n4104), .Y(new_n4113));
  NAND3xp33_ASAP7_75t_L     g03857(.A(new_n4050), .B(new_n4093), .C(new_n4101), .Y(new_n4114));
  NAND2xp33_ASAP7_75t_L     g03858(.A(new_n4110), .B(new_n4109), .Y(new_n4115));
  NAND3xp33_ASAP7_75t_L     g03859(.A(new_n4113), .B(new_n4114), .C(new_n4115), .Y(new_n4116));
  NAND2xp33_ASAP7_75t_L     g03860(.A(new_n4116), .B(new_n4112), .Y(new_n4117));
  NOR2xp33_ASAP7_75t_L      g03861(.A(new_n3878), .B(new_n3883), .Y(new_n4118));
  MAJIxp5_ASAP7_75t_L       g03862(.A(new_n3891), .B(new_n3839), .C(new_n4118), .Y(new_n4119));
  NOR2xp33_ASAP7_75t_L      g03863(.A(new_n4119), .B(new_n4117), .Y(new_n4120));
  NOR3xp33_ASAP7_75t_L      g03864(.A(new_n3883), .B(new_n3885), .C(new_n3878), .Y(new_n4121));
  AOI221xp5_ASAP7_75t_L     g03865(.A1(new_n3892), .A2(new_n3891), .B1(new_n4116), .B2(new_n4112), .C(new_n4121), .Y(new_n4122));
  AOI22xp33_ASAP7_75t_L     g03866(.A1(new_n1704), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1837), .Y(new_n4123));
  OAI221xp5_ASAP7_75t_L     g03867(.A1(new_n1699), .A2(new_n869), .B1(new_n1827), .B2(new_n950), .C(new_n4123), .Y(new_n4124));
  XNOR2x2_ASAP7_75t_L       g03868(.A(new_n1689), .B(new_n4124), .Y(new_n4125));
  NOR3xp33_ASAP7_75t_L      g03869(.A(new_n4120), .B(new_n4122), .C(new_n4125), .Y(new_n4126));
  AOI21xp33_ASAP7_75t_L     g03870(.A1(new_n4113), .A2(new_n4114), .B(new_n4115), .Y(new_n4127));
  NOR3xp33_ASAP7_75t_L      g03871(.A(new_n4105), .B(new_n4102), .C(new_n4111), .Y(new_n4128));
  NOR2xp33_ASAP7_75t_L      g03872(.A(new_n4127), .B(new_n4128), .Y(new_n4129));
  INVx1_ASAP7_75t_L         g03873(.A(new_n4121), .Y(new_n4130));
  A2O1A1Ixp33_ASAP7_75t_L   g03874(.A1(new_n3884), .A2(new_n3888), .B(new_n3836), .C(new_n4130), .Y(new_n4131));
  NAND2xp33_ASAP7_75t_L     g03875(.A(new_n4129), .B(new_n4131), .Y(new_n4132));
  NAND2xp33_ASAP7_75t_L     g03876(.A(new_n4119), .B(new_n4117), .Y(new_n4133));
  XNOR2x2_ASAP7_75t_L       g03877(.A(\a[23] ), .B(new_n4124), .Y(new_n4134));
  AOI21xp33_ASAP7_75t_L     g03878(.A1(new_n4132), .A2(new_n4133), .B(new_n4134), .Y(new_n4135));
  OAI21xp33_ASAP7_75t_L     g03879(.A1(new_n4135), .A2(new_n4126), .B(new_n4049), .Y(new_n4136));
  AOI31xp33_ASAP7_75t_L     g03880(.A1(new_n3894), .A2(new_n3901), .A3(new_n3688), .B(new_n3905), .Y(new_n4137));
  NAND3xp33_ASAP7_75t_L     g03881(.A(new_n4132), .B(new_n4133), .C(new_n4134), .Y(new_n4138));
  OAI21xp33_ASAP7_75t_L     g03882(.A1(new_n4122), .A2(new_n4120), .B(new_n4125), .Y(new_n4139));
  NAND3xp33_ASAP7_75t_L     g03883(.A(new_n4137), .B(new_n4138), .C(new_n4139), .Y(new_n4140));
  NAND3xp33_ASAP7_75t_L     g03884(.A(new_n4136), .B(new_n4140), .C(new_n4048), .Y(new_n4141));
  AND2x2_ASAP7_75t_L        g03885(.A(new_n4047), .B(new_n4046), .Y(new_n4142));
  AOI21xp33_ASAP7_75t_L     g03886(.A1(new_n4139), .A2(new_n4138), .B(new_n4137), .Y(new_n4143));
  AND4x1_ASAP7_75t_L        g03887(.A(new_n3902), .B(new_n4138), .C(new_n3899), .D(new_n4139), .Y(new_n4144));
  OAI21xp33_ASAP7_75t_L     g03888(.A1(new_n4143), .A2(new_n4144), .B(new_n4142), .Y(new_n4145));
  AOI21xp33_ASAP7_75t_L     g03889(.A1(new_n4145), .A2(new_n4141), .B(new_n4042), .Y(new_n4146));
  NAND2xp33_ASAP7_75t_L     g03890(.A(new_n4141), .B(new_n4145), .Y(new_n4147));
  O2A1O1Ixp33_ASAP7_75t_L   g03891(.A1(new_n3936), .A2(new_n3923), .B(new_n4041), .C(new_n4147), .Y(new_n4148));
  AOI22xp33_ASAP7_75t_L     g03892(.A1(new_n1076), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1253), .Y(new_n4149));
  OAI31xp33_ASAP7_75t_L     g03893(.A1(new_n1660), .A2(new_n1156), .A3(new_n1659), .B(new_n4149), .Y(new_n4150));
  AOI21xp33_ASAP7_75t_L     g03894(.A1(new_n1080), .A2(\b[20] ), .B(new_n4150), .Y(new_n4151));
  NAND2xp33_ASAP7_75t_L     g03895(.A(\a[17] ), .B(new_n4151), .Y(new_n4152));
  A2O1A1Ixp33_ASAP7_75t_L   g03896(.A1(\b[20] ), .A2(new_n1080), .B(new_n4150), .C(new_n1071), .Y(new_n4153));
  NAND2xp33_ASAP7_75t_L     g03897(.A(new_n4153), .B(new_n4152), .Y(new_n4154));
  NOR3xp33_ASAP7_75t_L      g03898(.A(new_n4148), .B(new_n4146), .C(new_n4154), .Y(new_n4155));
  AO221x2_ASAP7_75t_L       g03899(.A1(new_n4145), .A2(new_n4141), .B1(new_n3925), .B2(new_n3934), .C(new_n4040), .Y(new_n4156));
  NAND3xp33_ASAP7_75t_L     g03900(.A(new_n4042), .B(new_n4141), .C(new_n4145), .Y(new_n4157));
  AND2x2_ASAP7_75t_L        g03901(.A(new_n4153), .B(new_n4152), .Y(new_n4158));
  AOI21xp33_ASAP7_75t_L     g03902(.A1(new_n4157), .A2(new_n4156), .B(new_n4158), .Y(new_n4159));
  OAI211xp5_ASAP7_75t_L     g03903(.A1(new_n3724), .A2(new_n3736), .B(new_n3829), .C(new_n3943), .Y(new_n4160));
  OAI211xp5_ASAP7_75t_L     g03904(.A1(new_n4155), .A2(new_n4159), .B(new_n4160), .C(new_n3942), .Y(new_n4161));
  NOR2xp33_ASAP7_75t_L      g03905(.A(new_n4159), .B(new_n4155), .Y(new_n4162));
  OA211x2_ASAP7_75t_L       g03906(.A1(new_n3736), .A2(new_n3724), .B(new_n3943), .C(new_n3829), .Y(new_n4163));
  OAI21xp33_ASAP7_75t_L     g03907(.A1(new_n4163), .A2(new_n3933), .B(new_n4162), .Y(new_n4164));
  AOI21xp33_ASAP7_75t_L     g03908(.A1(new_n4164), .A2(new_n4161), .B(new_n4039), .Y(new_n4165));
  AND2x2_ASAP7_75t_L        g03909(.A(new_n4038), .B(new_n4036), .Y(new_n4166));
  NAND3xp33_ASAP7_75t_L     g03910(.A(new_n4157), .B(new_n4156), .C(new_n4158), .Y(new_n4167));
  OAI21xp33_ASAP7_75t_L     g03911(.A1(new_n4146), .A2(new_n4148), .B(new_n4154), .Y(new_n4168));
  AOI221xp5_ASAP7_75t_L     g03912(.A1(new_n4168), .A2(new_n4167), .B1(new_n3943), .B2(new_n3948), .C(new_n3933), .Y(new_n4169));
  AOI211xp5_ASAP7_75t_L     g03913(.A1(new_n4160), .A2(new_n3942), .B(new_n4155), .C(new_n4159), .Y(new_n4170));
  NOR3xp33_ASAP7_75t_L      g03914(.A(new_n4170), .B(new_n4169), .C(new_n4166), .Y(new_n4171));
  NOR2xp33_ASAP7_75t_L      g03915(.A(new_n4171), .B(new_n4165), .Y(new_n4172));
  A2O1A1Ixp33_ASAP7_75t_L   g03916(.A1(new_n3960), .A2(new_n3957), .B(new_n3959), .C(new_n4172), .Y(new_n4173));
  A2O1A1O1Ixp25_ASAP7_75t_L g03917(.A1(new_n3749), .A2(new_n3756), .B(new_n3822), .C(new_n3946), .D(new_n3959), .Y(new_n4174));
  OAI21xp33_ASAP7_75t_L     g03918(.A1(new_n4169), .A2(new_n4170), .B(new_n4166), .Y(new_n4175));
  NAND3xp33_ASAP7_75t_L     g03919(.A(new_n4164), .B(new_n4161), .C(new_n4039), .Y(new_n4176));
  NAND2xp33_ASAP7_75t_L     g03920(.A(new_n4175), .B(new_n4176), .Y(new_n4177));
  NAND2xp33_ASAP7_75t_L     g03921(.A(new_n4177), .B(new_n4174), .Y(new_n4178));
  NAND2xp33_ASAP7_75t_L     g03922(.A(\b[26] ), .B(new_n584), .Y(new_n4179));
  NAND2xp33_ASAP7_75t_L     g03923(.A(new_n578), .B(new_n2504), .Y(new_n4180));
  AOI22xp33_ASAP7_75t_L     g03924(.A1(\b[25] ), .A2(new_n651), .B1(\b[27] ), .B2(new_n581), .Y(new_n4181));
  AND4x1_ASAP7_75t_L        g03925(.A(new_n4181), .B(new_n4180), .C(new_n4179), .D(\a[11] ), .Y(new_n4182));
  AOI31xp33_ASAP7_75t_L     g03926(.A1(new_n4180), .A2(new_n4179), .A3(new_n4181), .B(\a[11] ), .Y(new_n4183));
  NOR2xp33_ASAP7_75t_L      g03927(.A(new_n4183), .B(new_n4182), .Y(new_n4184));
  NAND3xp33_ASAP7_75t_L     g03928(.A(new_n4173), .B(new_n4178), .C(new_n4184), .Y(new_n4185));
  NOR2xp33_ASAP7_75t_L      g03929(.A(new_n4177), .B(new_n4174), .Y(new_n4186));
  AOI221xp5_ASAP7_75t_L     g03930(.A1(new_n4176), .A2(new_n4175), .B1(new_n3960), .B2(new_n3957), .C(new_n3959), .Y(new_n4187));
  INVx1_ASAP7_75t_L         g03931(.A(new_n4184), .Y(new_n4188));
  OAI21xp33_ASAP7_75t_L     g03932(.A1(new_n4187), .A2(new_n4186), .B(new_n4188), .Y(new_n4189));
  NAND2xp33_ASAP7_75t_L     g03933(.A(new_n4189), .B(new_n4185), .Y(new_n4190));
  NAND2xp33_ASAP7_75t_L     g03934(.A(new_n4032), .B(new_n4190), .Y(new_n4191));
  A2O1A1O1Ixp25_ASAP7_75t_L g03935(.A1(new_n3760), .A2(new_n3763), .B(new_n3969), .C(new_n3955), .D(new_n3968), .Y(new_n4192));
  NAND3xp33_ASAP7_75t_L     g03936(.A(new_n4192), .B(new_n4185), .C(new_n4189), .Y(new_n4193));
  AOI21xp33_ASAP7_75t_L     g03937(.A1(new_n4191), .A2(new_n4193), .B(new_n4031), .Y(new_n4194));
  AOI21xp33_ASAP7_75t_L     g03938(.A1(new_n4189), .A2(new_n4185), .B(new_n4192), .Y(new_n4195));
  NOR2xp33_ASAP7_75t_L      g03939(.A(new_n4032), .B(new_n4190), .Y(new_n4196));
  NOR3xp33_ASAP7_75t_L      g03940(.A(new_n4196), .B(new_n4195), .C(new_n4030), .Y(new_n4197));
  NOR2xp33_ASAP7_75t_L      g03941(.A(new_n4194), .B(new_n4197), .Y(new_n4198));
  A2O1A1Ixp33_ASAP7_75t_L   g03942(.A1(new_n3983), .A2(new_n3980), .B(new_n4023), .C(new_n4198), .Y(new_n4199));
  A2O1A1O1Ixp25_ASAP7_75t_L g03943(.A1(new_n3772), .A2(new_n3770), .B(new_n4000), .C(new_n3980), .D(new_n4023), .Y(new_n4200));
  OAI21xp33_ASAP7_75t_L     g03944(.A1(new_n4195), .A2(new_n4196), .B(new_n4030), .Y(new_n4201));
  NAND3xp33_ASAP7_75t_L     g03945(.A(new_n4191), .B(new_n4031), .C(new_n4193), .Y(new_n4202));
  NAND2xp33_ASAP7_75t_L     g03946(.A(new_n4202), .B(new_n4201), .Y(new_n4203));
  NAND2xp33_ASAP7_75t_L     g03947(.A(new_n4203), .B(new_n4200), .Y(new_n4204));
  NAND3xp33_ASAP7_75t_L     g03948(.A(new_n4204), .B(new_n4199), .C(new_n4022), .Y(new_n4205));
  INVx1_ASAP7_75t_L         g03949(.A(new_n4023), .Y(new_n4206));
  O2A1O1Ixp33_ASAP7_75t_L   g03950(.A1(new_n3987), .A2(new_n3997), .B(new_n4206), .C(new_n4203), .Y(new_n4207));
  OAI21xp33_ASAP7_75t_L     g03951(.A1(new_n3987), .A2(new_n3997), .B(new_n4206), .Y(new_n4208));
  NOR2xp33_ASAP7_75t_L      g03952(.A(new_n4198), .B(new_n4208), .Y(new_n4209));
  OAI21xp33_ASAP7_75t_L     g03953(.A1(new_n4207), .A2(new_n4209), .B(new_n4021), .Y(new_n4210));
  A2O1A1Ixp33_ASAP7_75t_L   g03954(.A1(new_n3596), .A2(new_n3786), .B(new_n3818), .C(new_n4003), .Y(new_n4211));
  NAND4xp25_ASAP7_75t_L     g03955(.A(new_n4211), .B(new_n4205), .C(new_n3996), .D(new_n4210), .Y(new_n4212));
  AO22x1_ASAP7_75t_L        g03956(.A1(new_n4205), .A2(new_n4210), .B1(new_n3996), .B2(new_n4211), .Y(new_n4213));
  NAND2xp33_ASAP7_75t_L     g03957(.A(new_n4212), .B(new_n4213), .Y(new_n4214));
  NOR2xp33_ASAP7_75t_L      g03958(.A(\b[35] ), .B(\b[36] ), .Y(new_n4215));
  INVx1_ASAP7_75t_L         g03959(.A(\b[36] ), .Y(new_n4216));
  NOR2xp33_ASAP7_75t_L      g03960(.A(new_n3804), .B(new_n4216), .Y(new_n4217));
  NOR2xp33_ASAP7_75t_L      g03961(.A(new_n4215), .B(new_n4217), .Y(new_n4218));
  A2O1A1Ixp33_ASAP7_75t_L   g03962(.A1(\b[35] ), .A2(\b[34] ), .B(new_n3808), .C(new_n4218), .Y(new_n4219));
  O2A1O1Ixp33_ASAP7_75t_L   g03963(.A1(new_n3585), .A2(new_n3809), .B(new_n3806), .C(new_n3805), .Y(new_n4220));
  INVx1_ASAP7_75t_L         g03964(.A(new_n4218), .Y(new_n4221));
  NAND2xp33_ASAP7_75t_L     g03965(.A(new_n4221), .B(new_n4220), .Y(new_n4222));
  NAND2xp33_ASAP7_75t_L     g03966(.A(new_n4219), .B(new_n4222), .Y(new_n4223));
  AOI22xp33_ASAP7_75t_L     g03967(.A1(\b[34] ), .A2(new_n282), .B1(\b[36] ), .B2(new_n303), .Y(new_n4224));
  OAI221xp5_ASAP7_75t_L     g03968(.A1(new_n291), .A2(new_n3804), .B1(new_n268), .B2(new_n4223), .C(new_n4224), .Y(new_n4225));
  XNOR2x2_ASAP7_75t_L       g03969(.A(\a[2] ), .B(new_n4225), .Y(new_n4226));
  XOR2x2_ASAP7_75t_L        g03970(.A(new_n4226), .B(new_n4214), .Y(new_n4227));
  A2O1A1O1Ixp25_ASAP7_75t_L g03971(.A1(new_n3793), .A2(new_n3796), .B(new_n3791), .C(new_n4013), .D(new_n4011), .Y(new_n4228));
  XNOR2x2_ASAP7_75t_L       g03972(.A(new_n4228), .B(new_n4227), .Y(\f[36] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03973(.A1(new_n4016), .A2(new_n4013), .B(new_n4011), .C(new_n4227), .Y(new_n4230));
  AOI22xp33_ASAP7_75t_L     g03974(.A1(new_n444), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n471), .Y(new_n4231));
  OAI221xp5_ASAP7_75t_L     g03975(.A1(new_n468), .A2(new_n2982), .B1(new_n469), .B2(new_n3187), .C(new_n4231), .Y(new_n4232));
  XNOR2x2_ASAP7_75t_L       g03976(.A(new_n435), .B(new_n4232), .Y(new_n4233));
  NOR3xp33_ASAP7_75t_L      g03977(.A(new_n4186), .B(new_n4187), .C(new_n4184), .Y(new_n4234));
  INVx1_ASAP7_75t_L         g03978(.A(new_n4234), .Y(new_n4235));
  A2O1A1Ixp33_ASAP7_75t_L   g03979(.A1(new_n4185), .A2(new_n4189), .B(new_n4192), .C(new_n4235), .Y(new_n4236));
  INVx1_ASAP7_75t_L         g03980(.A(new_n2672), .Y(new_n4237));
  AOI22xp33_ASAP7_75t_L     g03981(.A1(\b[26] ), .A2(new_n651), .B1(\b[28] ), .B2(new_n581), .Y(new_n4238));
  INVx1_ASAP7_75t_L         g03982(.A(new_n4238), .Y(new_n4239));
  AOI221xp5_ASAP7_75t_L     g03983(.A1(\b[27] ), .A2(new_n584), .B1(new_n578), .B2(new_n4237), .C(new_n4239), .Y(new_n4240));
  XNOR2x2_ASAP7_75t_L       g03984(.A(new_n574), .B(new_n4240), .Y(new_n4241));
  OAI21xp33_ASAP7_75t_L     g03985(.A1(new_n4165), .A2(new_n4174), .B(new_n4176), .Y(new_n4242));
  AOI22xp33_ASAP7_75t_L     g03986(.A1(new_n2114), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n2259), .Y(new_n4243));
  OAI221xp5_ASAP7_75t_L     g03987(.A1(new_n2109), .A2(new_n760), .B1(new_n2257), .B2(new_n790), .C(new_n4243), .Y(new_n4244));
  XNOR2x2_ASAP7_75t_L       g03988(.A(\a[26] ), .B(new_n4244), .Y(new_n4245));
  INVx1_ASAP7_75t_L         g03989(.A(new_n4245), .Y(new_n4246));
  AOI22xp33_ASAP7_75t_L     g03990(.A1(new_n4099), .A2(new_n4100), .B1(new_n4094), .B2(new_n4098), .Y(new_n4247));
  A2O1A1O1Ixp25_ASAP7_75t_L g03991(.A1(new_n3882), .A2(new_n3880), .B(new_n3872), .C(new_n4101), .D(new_n4247), .Y(new_n4248));
  AOI22xp33_ASAP7_75t_L     g03992(.A1(new_n2552), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n2736), .Y(new_n4249));
  OAI221xp5_ASAP7_75t_L     g03993(.A1(new_n2547), .A2(new_n540), .B1(new_n2734), .B2(new_n624), .C(new_n4249), .Y(new_n4250));
  XNOR2x2_ASAP7_75t_L       g03994(.A(\a[29] ), .B(new_n4250), .Y(new_n4251));
  INVx1_ASAP7_75t_L         g03995(.A(new_n4251), .Y(new_n4252));
  NAND2xp33_ASAP7_75t_L     g03996(.A(new_n4077), .B(new_n4079), .Y(new_n4253));
  NAND3xp33_ASAP7_75t_L     g03997(.A(new_n4253), .B(new_n4073), .C(new_n4072), .Y(new_n4254));
  A2O1A1Ixp33_ASAP7_75t_L   g03998(.A1(new_n4081), .A2(new_n4080), .B(new_n4097), .C(new_n4254), .Y(new_n4255));
  AOI22xp33_ASAP7_75t_L     g03999(.A1(new_n3029), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n3258), .Y(new_n4256));
  OAI221xp5_ASAP7_75t_L     g04000(.A1(new_n3024), .A2(new_n418), .B1(new_n3256), .B2(new_n425), .C(new_n4256), .Y(new_n4257));
  OR2x4_ASAP7_75t_L         g04001(.A(new_n3015), .B(new_n4257), .Y(new_n4258));
  NAND2xp33_ASAP7_75t_L     g04002(.A(new_n3015), .B(new_n4257), .Y(new_n4259));
  NOR2xp33_ASAP7_75t_L      g04003(.A(new_n3862), .B(new_n3860), .Y(new_n4260));
  NAND2xp33_ASAP7_75t_L     g04004(.A(new_n4059), .B(new_n4260), .Y(new_n4261));
  NOR2xp33_ASAP7_75t_L      g04005(.A(new_n298), .B(new_n3853), .Y(new_n4262));
  NOR3xp33_ASAP7_75t_L      g04006(.A(new_n326), .B(new_n328), .C(new_n3856), .Y(new_n4263));
  OAI22xp33_ASAP7_75t_L     g04007(.A1(new_n4052), .A2(new_n276), .B1(new_n324), .B2(new_n4061), .Y(new_n4264));
  NOR4xp25_ASAP7_75t_L      g04008(.A(new_n4263), .B(new_n4264), .C(new_n3628), .D(new_n4262), .Y(new_n4265));
  OAI31xp33_ASAP7_75t_L     g04009(.A1(new_n4263), .A2(new_n4264), .A3(new_n4262), .B(new_n3628), .Y(new_n4266));
  INVx1_ASAP7_75t_L         g04010(.A(new_n4266), .Y(new_n4267));
  INVx1_ASAP7_75t_L         g04011(.A(\a[38] ), .Y(new_n4268));
  NOR2xp33_ASAP7_75t_L      g04012(.A(new_n4268), .B(new_n4058), .Y(new_n4269));
  AND2x2_ASAP7_75t_L        g04013(.A(new_n4055), .B(new_n4056), .Y(new_n4270));
  INVx1_ASAP7_75t_L         g04014(.A(\a[37] ), .Y(new_n4271));
  NAND2xp33_ASAP7_75t_L     g04015(.A(\a[38] ), .B(new_n4271), .Y(new_n4272));
  NAND2xp33_ASAP7_75t_L     g04016(.A(\a[37] ), .B(new_n4268), .Y(new_n4273));
  AOI21xp33_ASAP7_75t_L     g04017(.A1(new_n4273), .A2(new_n4272), .B(new_n4270), .Y(new_n4274));
  NAND3xp33_ASAP7_75t_L     g04018(.A(new_n4057), .B(new_n4272), .C(new_n4273), .Y(new_n4275));
  XNOR2x2_ASAP7_75t_L       g04019(.A(\a[37] ), .B(\a[36] ), .Y(new_n4276));
  OR2x4_ASAP7_75t_L         g04020(.A(new_n4276), .B(new_n4057), .Y(new_n4277));
  OAI22xp33_ASAP7_75t_L     g04021(.A1(new_n4277), .A2(new_n258), .B1(new_n261), .B2(new_n4275), .Y(new_n4278));
  A2O1A1Ixp33_ASAP7_75t_L   g04022(.A1(new_n269), .A2(new_n4274), .B(new_n4278), .C(new_n4269), .Y(new_n4279));
  INVx1_ASAP7_75t_L         g04023(.A(new_n4269), .Y(new_n4280));
  NAND2xp33_ASAP7_75t_L     g04024(.A(new_n269), .B(new_n4274), .Y(new_n4281));
  NAND2xp33_ASAP7_75t_L     g04025(.A(new_n4273), .B(new_n4272), .Y(new_n4282));
  NOR2xp33_ASAP7_75t_L      g04026(.A(new_n4282), .B(new_n4270), .Y(new_n4283));
  NAND2xp33_ASAP7_75t_L     g04027(.A(\b[1] ), .B(new_n4283), .Y(new_n4284));
  NOR2xp33_ASAP7_75t_L      g04028(.A(new_n4276), .B(new_n4057), .Y(new_n4285));
  NAND2xp33_ASAP7_75t_L     g04029(.A(\b[0] ), .B(new_n4285), .Y(new_n4286));
  NAND4xp25_ASAP7_75t_L     g04030(.A(new_n4280), .B(new_n4286), .C(new_n4284), .D(new_n4281), .Y(new_n4287));
  AND2x2_ASAP7_75t_L        g04031(.A(new_n4287), .B(new_n4279), .Y(new_n4288));
  NOR3xp33_ASAP7_75t_L      g04032(.A(new_n4288), .B(new_n4267), .C(new_n4265), .Y(new_n4289));
  INVx1_ASAP7_75t_L         g04033(.A(new_n4265), .Y(new_n4290));
  NAND2xp33_ASAP7_75t_L     g04034(.A(new_n4287), .B(new_n4279), .Y(new_n4291));
  AOI21xp33_ASAP7_75t_L     g04035(.A1(new_n4290), .A2(new_n4266), .B(new_n4291), .Y(new_n4292));
  AOI211xp5_ASAP7_75t_L     g04036(.A1(new_n4072), .A2(new_n4261), .B(new_n4289), .C(new_n4292), .Y(new_n4293));
  AOI22xp33_ASAP7_75t_L     g04037(.A1(new_n4060), .A2(new_n4065), .B1(new_n4069), .B2(new_n4071), .Y(new_n4294));
  NAND3xp33_ASAP7_75t_L     g04038(.A(new_n4291), .B(new_n4290), .C(new_n4266), .Y(new_n4295));
  OAI21xp33_ASAP7_75t_L     g04039(.A1(new_n4265), .A2(new_n4267), .B(new_n4288), .Y(new_n4296));
  AOI221xp5_ASAP7_75t_L     g04040(.A1(new_n4059), .A2(new_n4260), .B1(new_n4295), .B2(new_n4296), .C(new_n4294), .Y(new_n4297));
  OAI211xp5_ASAP7_75t_L     g04041(.A1(new_n4297), .A2(new_n4293), .B(new_n4259), .C(new_n4258), .Y(new_n4298));
  NAND2xp33_ASAP7_75t_L     g04042(.A(new_n4259), .B(new_n4258), .Y(new_n4299));
  NOR2xp33_ASAP7_75t_L      g04043(.A(new_n4292), .B(new_n4289), .Y(new_n4300));
  A2O1A1Ixp33_ASAP7_75t_L   g04044(.A1(new_n4260), .A2(new_n4059), .B(new_n4294), .C(new_n4300), .Y(new_n4301));
  INVx1_ASAP7_75t_L         g04045(.A(new_n4297), .Y(new_n4302));
  NAND3xp33_ASAP7_75t_L     g04046(.A(new_n4299), .B(new_n4301), .C(new_n4302), .Y(new_n4303));
  NAND3xp33_ASAP7_75t_L     g04047(.A(new_n4255), .B(new_n4298), .C(new_n4303), .Y(new_n4304));
  AND4x1_ASAP7_75t_L        g04048(.A(new_n4072), .B(new_n4079), .C(new_n4073), .D(new_n4077), .Y(new_n4305));
  AOI22xp33_ASAP7_75t_L     g04049(.A1(new_n4072), .A2(new_n4073), .B1(new_n4077), .B2(new_n4079), .Y(new_n4306));
  AND3x1_ASAP7_75t_L        g04050(.A(new_n4253), .B(new_n4073), .C(new_n4072), .Y(new_n4307));
  O2A1O1Ixp33_ASAP7_75t_L   g04051(.A1(new_n4305), .A2(new_n4306), .B(new_n4085), .C(new_n4307), .Y(new_n4308));
  AOI21xp33_ASAP7_75t_L     g04052(.A1(new_n4301), .A2(new_n4302), .B(new_n4299), .Y(new_n4309));
  AOI211xp5_ASAP7_75t_L     g04053(.A1(new_n4259), .A2(new_n4258), .B(new_n4297), .C(new_n4293), .Y(new_n4310));
  OAI21xp33_ASAP7_75t_L     g04054(.A1(new_n4309), .A2(new_n4310), .B(new_n4308), .Y(new_n4311));
  AOI21xp33_ASAP7_75t_L     g04055(.A1(new_n4304), .A2(new_n4311), .B(new_n4252), .Y(new_n4312));
  OAI221xp5_ASAP7_75t_L     g04056(.A1(new_n3845), .A2(new_n4096), .B1(new_n4305), .B2(new_n4306), .C(new_n3865), .Y(new_n4313));
  AOI211xp5_ASAP7_75t_L     g04057(.A1(new_n4313), .A2(new_n4254), .B(new_n4310), .C(new_n4309), .Y(new_n4314));
  AOI221xp5_ASAP7_75t_L     g04058(.A1(new_n4095), .A2(new_n4085), .B1(new_n4298), .B2(new_n4303), .C(new_n4307), .Y(new_n4315));
  NOR3xp33_ASAP7_75t_L      g04059(.A(new_n4315), .B(new_n4314), .C(new_n4251), .Y(new_n4316));
  OR3x1_ASAP7_75t_L         g04060(.A(new_n4248), .B(new_n4312), .C(new_n4316), .Y(new_n4317));
  OAI21xp33_ASAP7_75t_L     g04061(.A1(new_n4316), .A2(new_n4312), .B(new_n4248), .Y(new_n4318));
  AOI21xp33_ASAP7_75t_L     g04062(.A1(new_n4317), .A2(new_n4318), .B(new_n4246), .Y(new_n4319));
  NOR3xp33_ASAP7_75t_L      g04063(.A(new_n4248), .B(new_n4312), .C(new_n4316), .Y(new_n4320));
  OA21x2_ASAP7_75t_L        g04064(.A1(new_n4316), .A2(new_n4312), .B(new_n4248), .Y(new_n4321));
  NOR3xp33_ASAP7_75t_L      g04065(.A(new_n4321), .B(new_n4320), .C(new_n4245), .Y(new_n4322));
  NOR2xp33_ASAP7_75t_L      g04066(.A(new_n4322), .B(new_n4319), .Y(new_n4323));
  A2O1A1Ixp33_ASAP7_75t_L   g04067(.A1(new_n4131), .A2(new_n4112), .B(new_n4128), .C(new_n4323), .Y(new_n4324));
  A2O1A1O1Ixp25_ASAP7_75t_L g04068(.A1(new_n3891), .A2(new_n3892), .B(new_n4121), .C(new_n4112), .D(new_n4128), .Y(new_n4325));
  OAI21xp33_ASAP7_75t_L     g04069(.A1(new_n4320), .A2(new_n4321), .B(new_n4245), .Y(new_n4326));
  NAND3xp33_ASAP7_75t_L     g04070(.A(new_n4246), .B(new_n4317), .C(new_n4318), .Y(new_n4327));
  NAND2xp33_ASAP7_75t_L     g04071(.A(new_n4326), .B(new_n4327), .Y(new_n4328));
  NAND2xp33_ASAP7_75t_L     g04072(.A(new_n4325), .B(new_n4328), .Y(new_n4329));
  AOI22xp33_ASAP7_75t_L     g04073(.A1(new_n1704), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1837), .Y(new_n4330));
  OAI221xp5_ASAP7_75t_L     g04074(.A1(new_n1699), .A2(new_n942), .B1(new_n1827), .B2(new_n1035), .C(new_n4330), .Y(new_n4331));
  XNOR2x2_ASAP7_75t_L       g04075(.A(\a[23] ), .B(new_n4331), .Y(new_n4332));
  NAND3xp33_ASAP7_75t_L     g04076(.A(new_n4324), .B(new_n4329), .C(new_n4332), .Y(new_n4333));
  O2A1O1Ixp33_ASAP7_75t_L   g04077(.A1(new_n4127), .A2(new_n4119), .B(new_n4116), .C(new_n4328), .Y(new_n4334));
  OAI21xp33_ASAP7_75t_L     g04078(.A1(new_n4127), .A2(new_n4119), .B(new_n4116), .Y(new_n4335));
  NOR2xp33_ASAP7_75t_L      g04079(.A(new_n4335), .B(new_n4323), .Y(new_n4336));
  INVx1_ASAP7_75t_L         g04080(.A(new_n4332), .Y(new_n4337));
  OAI21xp33_ASAP7_75t_L     g04081(.A1(new_n4336), .A2(new_n4334), .B(new_n4337), .Y(new_n4338));
  NOR2xp33_ASAP7_75t_L      g04082(.A(new_n4122), .B(new_n4120), .Y(new_n4339));
  MAJIxp5_ASAP7_75t_L       g04083(.A(new_n4049), .B(new_n4125), .C(new_n4339), .Y(new_n4340));
  NAND3xp33_ASAP7_75t_L     g04084(.A(new_n4340), .B(new_n4338), .C(new_n4333), .Y(new_n4341));
  NOR3xp33_ASAP7_75t_L      g04085(.A(new_n4334), .B(new_n4336), .C(new_n4337), .Y(new_n4342));
  AOI21xp33_ASAP7_75t_L     g04086(.A1(new_n4324), .A2(new_n4329), .B(new_n4332), .Y(new_n4343));
  XNOR2x2_ASAP7_75t_L       g04087(.A(new_n4119), .B(new_n4117), .Y(new_n4344));
  MAJIxp5_ASAP7_75t_L       g04088(.A(new_n4137), .B(new_n4134), .C(new_n4344), .Y(new_n4345));
  OAI21xp33_ASAP7_75t_L     g04089(.A1(new_n4342), .A2(new_n4343), .B(new_n4345), .Y(new_n4346));
  AOI22xp33_ASAP7_75t_L     g04090(.A1(new_n1360), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1581), .Y(new_n4347));
  OAI221xp5_ASAP7_75t_L     g04091(.A1(new_n1373), .A2(new_n1313), .B1(new_n1359), .B2(new_n1438), .C(new_n4347), .Y(new_n4348));
  XNOR2x2_ASAP7_75t_L       g04092(.A(\a[20] ), .B(new_n4348), .Y(new_n4349));
  NAND3xp33_ASAP7_75t_L     g04093(.A(new_n4341), .B(new_n4346), .C(new_n4349), .Y(new_n4350));
  NOR3xp33_ASAP7_75t_L      g04094(.A(new_n4345), .B(new_n4343), .C(new_n4342), .Y(new_n4351));
  AOI21xp33_ASAP7_75t_L     g04095(.A1(new_n4338), .A2(new_n4333), .B(new_n4340), .Y(new_n4352));
  XNOR2x2_ASAP7_75t_L       g04096(.A(new_n1356), .B(new_n4348), .Y(new_n4353));
  OAI21xp33_ASAP7_75t_L     g04097(.A1(new_n4351), .A2(new_n4352), .B(new_n4353), .Y(new_n4354));
  NOR3xp33_ASAP7_75t_L      g04098(.A(new_n4144), .B(new_n4142), .C(new_n4143), .Y(new_n4355));
  A2O1A1O1Ixp25_ASAP7_75t_L g04099(.A1(new_n3925), .A2(new_n3934), .B(new_n4040), .C(new_n4145), .D(new_n4355), .Y(new_n4356));
  NAND3xp33_ASAP7_75t_L     g04100(.A(new_n4356), .B(new_n4354), .C(new_n4350), .Y(new_n4357));
  NAND2xp33_ASAP7_75t_L     g04101(.A(new_n4350), .B(new_n4354), .Y(new_n4358));
  A2O1A1Ixp33_ASAP7_75t_L   g04102(.A1(new_n4145), .A2(new_n4042), .B(new_n4355), .C(new_n4358), .Y(new_n4359));
  NAND2xp33_ASAP7_75t_L     g04103(.A(\b[21] ), .B(new_n1080), .Y(new_n4360));
  NAND2xp33_ASAP7_75t_L     g04104(.A(new_n1073), .B(new_n3728), .Y(new_n4361));
  AOI22xp33_ASAP7_75t_L     g04105(.A1(new_n1076), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1253), .Y(new_n4362));
  AND4x1_ASAP7_75t_L        g04106(.A(new_n4362), .B(new_n4361), .C(new_n4360), .D(\a[17] ), .Y(new_n4363));
  AOI31xp33_ASAP7_75t_L     g04107(.A1(new_n4361), .A2(new_n4360), .A3(new_n4362), .B(\a[17] ), .Y(new_n4364));
  NOR2xp33_ASAP7_75t_L      g04108(.A(new_n4364), .B(new_n4363), .Y(new_n4365));
  NAND3xp33_ASAP7_75t_L     g04109(.A(new_n4359), .B(new_n4357), .C(new_n4365), .Y(new_n4366));
  AND3x1_ASAP7_75t_L        g04110(.A(new_n4356), .B(new_n4354), .C(new_n4350), .Y(new_n4367));
  AOI21xp33_ASAP7_75t_L     g04111(.A1(new_n4354), .A2(new_n4350), .B(new_n4356), .Y(new_n4368));
  OR2x4_ASAP7_75t_L         g04112(.A(new_n4364), .B(new_n4363), .Y(new_n4369));
  OAI21xp33_ASAP7_75t_L     g04113(.A1(new_n4368), .A2(new_n4367), .B(new_n4369), .Y(new_n4370));
  NOR3xp33_ASAP7_75t_L      g04114(.A(new_n4148), .B(new_n4146), .C(new_n4158), .Y(new_n4371));
  INVx1_ASAP7_75t_L         g04115(.A(new_n4371), .Y(new_n4372));
  NAND4xp25_ASAP7_75t_L     g04116(.A(new_n4161), .B(new_n4372), .C(new_n4370), .D(new_n4366), .Y(new_n4373));
  NAND2xp33_ASAP7_75t_L     g04117(.A(new_n4370), .B(new_n4366), .Y(new_n4374));
  OAI21xp33_ASAP7_75t_L     g04118(.A1(new_n4371), .A2(new_n4169), .B(new_n4374), .Y(new_n4375));
  AOI22xp33_ASAP7_75t_L     g04119(.A1(new_n811), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n900), .Y(new_n4376));
  OAI31xp33_ASAP7_75t_L     g04120(.A1(new_n2074), .A2(new_n898), .A3(new_n2071), .B(new_n4376), .Y(new_n4377));
  AOI21xp33_ASAP7_75t_L     g04121(.A1(new_n815), .A2(\b[24] ), .B(new_n4377), .Y(new_n4378));
  NAND2xp33_ASAP7_75t_L     g04122(.A(\a[14] ), .B(new_n4378), .Y(new_n4379));
  A2O1A1Ixp33_ASAP7_75t_L   g04123(.A1(\b[24] ), .A2(new_n815), .B(new_n4377), .C(new_n806), .Y(new_n4380));
  NAND2xp33_ASAP7_75t_L     g04124(.A(new_n4380), .B(new_n4379), .Y(new_n4381));
  AO21x2_ASAP7_75t_L        g04125(.A1(new_n4373), .A2(new_n4375), .B(new_n4381), .Y(new_n4382));
  NAND3xp33_ASAP7_75t_L     g04126(.A(new_n4375), .B(new_n4373), .C(new_n4381), .Y(new_n4383));
  AOI21xp33_ASAP7_75t_L     g04127(.A1(new_n4383), .A2(new_n4382), .B(new_n4242), .Y(new_n4384));
  A2O1A1O1Ixp25_ASAP7_75t_L g04128(.A1(new_n3946), .A2(new_n3957), .B(new_n3959), .C(new_n4175), .D(new_n4171), .Y(new_n4385));
  NAND2xp33_ASAP7_75t_L     g04129(.A(new_n4383), .B(new_n4382), .Y(new_n4386));
  NOR2xp33_ASAP7_75t_L      g04130(.A(new_n4385), .B(new_n4386), .Y(new_n4387));
  OAI21xp33_ASAP7_75t_L     g04131(.A1(new_n4384), .A2(new_n4387), .B(new_n4241), .Y(new_n4388));
  AND2x2_ASAP7_75t_L        g04132(.A(\a[11] ), .B(new_n4240), .Y(new_n4389));
  NOR2xp33_ASAP7_75t_L      g04133(.A(\a[11] ), .B(new_n4240), .Y(new_n4390));
  NAND2xp33_ASAP7_75t_L     g04134(.A(new_n4385), .B(new_n4386), .Y(new_n4391));
  NAND3xp33_ASAP7_75t_L     g04135(.A(new_n4242), .B(new_n4382), .C(new_n4383), .Y(new_n4392));
  OAI211xp5_ASAP7_75t_L     g04136(.A1(new_n4390), .A2(new_n4389), .B(new_n4391), .C(new_n4392), .Y(new_n4393));
  NAND3xp33_ASAP7_75t_L     g04137(.A(new_n4236), .B(new_n4388), .C(new_n4393), .Y(new_n4394));
  AO221x2_ASAP7_75t_L       g04138(.A1(new_n4032), .A2(new_n4190), .B1(new_n4393), .B2(new_n4388), .C(new_n4234), .Y(new_n4395));
  AOI21xp33_ASAP7_75t_L     g04139(.A1(new_n4394), .A2(new_n4395), .B(new_n4233), .Y(new_n4396));
  AND3x1_ASAP7_75t_L        g04140(.A(new_n4394), .B(new_n4395), .C(new_n4233), .Y(new_n4397));
  NOR2xp33_ASAP7_75t_L      g04141(.A(new_n4396), .B(new_n4397), .Y(new_n4398));
  A2O1A1Ixp33_ASAP7_75t_L   g04142(.A1(new_n4201), .A2(new_n4208), .B(new_n4197), .C(new_n4398), .Y(new_n4399));
  A2O1A1O1Ixp25_ASAP7_75t_L g04143(.A1(new_n3980), .A2(new_n3983), .B(new_n4023), .C(new_n4201), .D(new_n4197), .Y(new_n4400));
  AO21x2_ASAP7_75t_L        g04144(.A1(new_n4395), .A2(new_n4394), .B(new_n4233), .Y(new_n4401));
  NAND3xp33_ASAP7_75t_L     g04145(.A(new_n4394), .B(new_n4395), .C(new_n4233), .Y(new_n4402));
  NAND2xp33_ASAP7_75t_L     g04146(.A(new_n4402), .B(new_n4401), .Y(new_n4403));
  NAND2xp33_ASAP7_75t_L     g04147(.A(new_n4400), .B(new_n4403), .Y(new_n4404));
  AOI22xp33_ASAP7_75t_L     g04148(.A1(new_n344), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n370), .Y(new_n4405));
  OAI221xp5_ASAP7_75t_L     g04149(.A1(new_n429), .A2(new_n3565), .B1(new_n366), .B2(new_n3591), .C(new_n4405), .Y(new_n4406));
  XNOR2x2_ASAP7_75t_L       g04150(.A(\a[5] ), .B(new_n4406), .Y(new_n4407));
  NAND3xp33_ASAP7_75t_L     g04151(.A(new_n4399), .B(new_n4404), .C(new_n4407), .Y(new_n4408));
  O2A1O1Ixp33_ASAP7_75t_L   g04152(.A1(new_n4200), .A2(new_n4194), .B(new_n4202), .C(new_n4403), .Y(new_n4409));
  NOR3xp33_ASAP7_75t_L      g04153(.A(new_n4398), .B(new_n4207), .C(new_n4197), .Y(new_n4410));
  INVx1_ASAP7_75t_L         g04154(.A(new_n4407), .Y(new_n4411));
  OAI21xp33_ASAP7_75t_L     g04155(.A1(new_n4409), .A2(new_n4410), .B(new_n4411), .Y(new_n4412));
  NAND2xp33_ASAP7_75t_L     g04156(.A(new_n4408), .B(new_n4412), .Y(new_n4413));
  NAND2xp33_ASAP7_75t_L     g04157(.A(new_n4210), .B(new_n4205), .Y(new_n4414));
  A2O1A1Ixp33_ASAP7_75t_L   g04158(.A1(new_n4009), .A2(new_n3780), .B(new_n4008), .C(new_n3996), .Y(new_n4415));
  OAI21xp33_ASAP7_75t_L     g04159(.A1(new_n4415), .A2(new_n4414), .B(new_n4205), .Y(new_n4416));
  NOR2xp33_ASAP7_75t_L      g04160(.A(new_n4416), .B(new_n4413), .Y(new_n4417));
  NOR3xp33_ASAP7_75t_L      g04161(.A(new_n4209), .B(new_n4207), .C(new_n4021), .Y(new_n4418));
  AOI31xp33_ASAP7_75t_L     g04162(.A1(new_n4211), .A2(new_n3996), .A3(new_n4210), .B(new_n4418), .Y(new_n4419));
  AOI21xp33_ASAP7_75t_L     g04163(.A1(new_n4412), .A2(new_n4408), .B(new_n4419), .Y(new_n4420));
  INVx1_ASAP7_75t_L         g04164(.A(new_n3805), .Y(new_n4421));
  A2O1A1Ixp33_ASAP7_75t_L   g04165(.A1(new_n3587), .A2(new_n3802), .B(new_n3807), .C(new_n4421), .Y(new_n4422));
  NOR2xp33_ASAP7_75t_L      g04166(.A(\b[36] ), .B(\b[37] ), .Y(new_n4423));
  INVx1_ASAP7_75t_L         g04167(.A(\b[37] ), .Y(new_n4424));
  NOR2xp33_ASAP7_75t_L      g04168(.A(new_n4216), .B(new_n4424), .Y(new_n4425));
  NOR2xp33_ASAP7_75t_L      g04169(.A(new_n4423), .B(new_n4425), .Y(new_n4426));
  A2O1A1Ixp33_ASAP7_75t_L   g04170(.A1(new_n4422), .A2(new_n4218), .B(new_n4217), .C(new_n4426), .Y(new_n4427));
  O2A1O1Ixp33_ASAP7_75t_L   g04171(.A1(new_n3805), .A2(new_n3808), .B(new_n4218), .C(new_n4217), .Y(new_n4428));
  INVx1_ASAP7_75t_L         g04172(.A(new_n4426), .Y(new_n4429));
  NAND2xp33_ASAP7_75t_L     g04173(.A(new_n4429), .B(new_n4428), .Y(new_n4430));
  NAND2xp33_ASAP7_75t_L     g04174(.A(new_n4430), .B(new_n4427), .Y(new_n4431));
  AOI22xp33_ASAP7_75t_L     g04175(.A1(\b[35] ), .A2(new_n282), .B1(\b[37] ), .B2(new_n303), .Y(new_n4432));
  OAI221xp5_ASAP7_75t_L     g04176(.A1(new_n291), .A2(new_n4216), .B1(new_n268), .B2(new_n4431), .C(new_n4432), .Y(new_n4433));
  XNOR2x2_ASAP7_75t_L       g04177(.A(\a[2] ), .B(new_n4433), .Y(new_n4434));
  OAI21xp33_ASAP7_75t_L     g04178(.A1(new_n4420), .A2(new_n4417), .B(new_n4434), .Y(new_n4435));
  NOR3xp33_ASAP7_75t_L      g04179(.A(new_n4417), .B(new_n4420), .C(new_n4434), .Y(new_n4436));
  INVx1_ASAP7_75t_L         g04180(.A(new_n4436), .Y(new_n4437));
  NAND2xp33_ASAP7_75t_L     g04181(.A(new_n4435), .B(new_n4437), .Y(new_n4438));
  O2A1O1Ixp33_ASAP7_75t_L   g04182(.A1(new_n4214), .A2(new_n4226), .B(new_n4230), .C(new_n4438), .Y(new_n4439));
  MAJIxp5_ASAP7_75t_L       g04183(.A(new_n4228), .B(new_n4226), .C(new_n4214), .Y(new_n4440));
  AOI21xp33_ASAP7_75t_L     g04184(.A1(new_n4437), .A2(new_n4435), .B(new_n4440), .Y(new_n4441));
  NOR2xp33_ASAP7_75t_L      g04185(.A(new_n4441), .B(new_n4439), .Y(\f[37] ));
  NAND2xp33_ASAP7_75t_L     g04186(.A(new_n4404), .B(new_n4399), .Y(new_n4443));
  MAJIxp5_ASAP7_75t_L       g04187(.A(new_n4419), .B(new_n4407), .C(new_n4443), .Y(new_n4444));
  NAND2xp33_ASAP7_75t_L     g04188(.A(\b[34] ), .B(new_n347), .Y(new_n4445));
  NAND2xp33_ASAP7_75t_L     g04189(.A(new_n341), .B(new_n3811), .Y(new_n4446));
  AOI22xp33_ASAP7_75t_L     g04190(.A1(new_n344), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n370), .Y(new_n4447));
  NAND3xp33_ASAP7_75t_L     g04191(.A(new_n4446), .B(new_n4445), .C(new_n4447), .Y(new_n4448));
  NOR2xp33_ASAP7_75t_L      g04192(.A(new_n338), .B(new_n4448), .Y(new_n4449));
  AOI31xp33_ASAP7_75t_L     g04193(.A1(new_n4446), .A2(new_n4445), .A3(new_n4447), .B(\a[5] ), .Y(new_n4450));
  NOR2xp33_ASAP7_75t_L      g04194(.A(new_n4450), .B(new_n4449), .Y(new_n4451));
  NOR2xp33_ASAP7_75t_L      g04195(.A(new_n3180), .B(new_n468), .Y(new_n4452));
  INVx1_ASAP7_75t_L         g04196(.A(new_n4452), .Y(new_n4453));
  NAND3xp33_ASAP7_75t_L     g04197(.A(new_n3210), .B(new_n441), .C(new_n3213), .Y(new_n4454));
  AOI22xp33_ASAP7_75t_L     g04198(.A1(new_n444), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n471), .Y(new_n4455));
  NAND4xp25_ASAP7_75t_L     g04199(.A(new_n4454), .B(\a[8] ), .C(new_n4453), .D(new_n4455), .Y(new_n4456));
  AOI31xp33_ASAP7_75t_L     g04200(.A1(new_n4454), .A2(new_n4453), .A3(new_n4455), .B(\a[8] ), .Y(new_n4457));
  INVx1_ASAP7_75t_L         g04201(.A(new_n4457), .Y(new_n4458));
  NAND2xp33_ASAP7_75t_L     g04202(.A(new_n4456), .B(new_n4458), .Y(new_n4459));
  INVx1_ASAP7_75t_L         g04203(.A(new_n4459), .Y(new_n4460));
  O2A1O1Ixp33_ASAP7_75t_L   g04204(.A1(new_n3968), .A2(new_n3976), .B(new_n4190), .C(new_n4234), .Y(new_n4461));
  INVx1_ASAP7_75t_L         g04205(.A(new_n4388), .Y(new_n4462));
  AOI22xp33_ASAP7_75t_L     g04206(.A1(\b[27] ), .A2(new_n651), .B1(\b[29] ), .B2(new_n581), .Y(new_n4463));
  OAI221xp5_ASAP7_75t_L     g04207(.A1(new_n821), .A2(new_n2666), .B1(new_n577), .B2(new_n2695), .C(new_n4463), .Y(new_n4464));
  XNOR2x2_ASAP7_75t_L       g04208(.A(new_n574), .B(new_n4464), .Y(new_n4465));
  AOI22xp33_ASAP7_75t_L     g04209(.A1(new_n811), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n900), .Y(new_n4466));
  OAI221xp5_ASAP7_75t_L     g04210(.A1(new_n904), .A2(new_n2067), .B1(new_n898), .B2(new_n2355), .C(new_n4466), .Y(new_n4467));
  NOR2xp33_ASAP7_75t_L      g04211(.A(new_n806), .B(new_n4467), .Y(new_n4468));
  AND2x2_ASAP7_75t_L        g04212(.A(new_n806), .B(new_n4467), .Y(new_n4469));
  NOR2xp33_ASAP7_75t_L      g04213(.A(new_n4468), .B(new_n4469), .Y(new_n4470));
  OAI31xp33_ASAP7_75t_L     g04214(.A1(new_n4162), .A2(new_n3933), .A3(new_n4163), .B(new_n4372), .Y(new_n4471));
  NOR3xp33_ASAP7_75t_L      g04215(.A(new_n4367), .B(new_n4368), .C(new_n4365), .Y(new_n4472));
  OAI21xp33_ASAP7_75t_L     g04216(.A1(new_n4319), .A2(new_n4325), .B(new_n4327), .Y(new_n4473));
  AOI22xp33_ASAP7_75t_L     g04217(.A1(new_n2114), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n2259), .Y(new_n4474));
  OAI221xp5_ASAP7_75t_L     g04218(.A1(new_n2109), .A2(new_n784), .B1(new_n2257), .B2(new_n875), .C(new_n4474), .Y(new_n4475));
  XNOR2x2_ASAP7_75t_L       g04219(.A(new_n2100), .B(new_n4475), .Y(new_n4476));
  NAND3xp33_ASAP7_75t_L     g04220(.A(new_n4252), .B(new_n4304), .C(new_n4311), .Y(new_n4477));
  OAI21xp33_ASAP7_75t_L     g04221(.A1(new_n4312), .A2(new_n4248), .B(new_n4477), .Y(new_n4478));
  NAND2xp33_ASAP7_75t_L     g04222(.A(\b[10] ), .B(new_n2553), .Y(new_n4479));
  NAND3xp33_ASAP7_75t_L     g04223(.A(new_n684), .B(new_n682), .C(new_n2544), .Y(new_n4480));
  AOI22xp33_ASAP7_75t_L     g04224(.A1(new_n2552), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n2736), .Y(new_n4481));
  NAND4xp25_ASAP7_75t_L     g04225(.A(new_n4480), .B(\a[29] ), .C(new_n4479), .D(new_n4481), .Y(new_n4482));
  NAND3xp33_ASAP7_75t_L     g04226(.A(new_n4480), .B(new_n4479), .C(new_n4481), .Y(new_n4483));
  NAND2xp33_ASAP7_75t_L     g04227(.A(new_n2538), .B(new_n4483), .Y(new_n4484));
  AND2x2_ASAP7_75t_L        g04228(.A(new_n4482), .B(new_n4484), .Y(new_n4485));
  A2O1A1Ixp33_ASAP7_75t_L   g04229(.A1(new_n4313), .A2(new_n4254), .B(new_n4309), .C(new_n4303), .Y(new_n4486));
  AOI22xp33_ASAP7_75t_L     g04230(.A1(new_n3029), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n3258), .Y(new_n4487));
  OAI221xp5_ASAP7_75t_L     g04231(.A1(new_n3024), .A2(new_n420), .B1(new_n3256), .B2(new_n494), .C(new_n4487), .Y(new_n4488));
  XNOR2x2_ASAP7_75t_L       g04232(.A(\a[32] ), .B(new_n4488), .Y(new_n4489));
  A2O1A1O1Ixp25_ASAP7_75t_L g04233(.A1(new_n4260), .A2(new_n4059), .B(new_n4294), .C(new_n4295), .D(new_n4292), .Y(new_n4490));
  NOR2xp33_ASAP7_75t_L      g04234(.A(new_n324), .B(new_n3853), .Y(new_n4491));
  NOR3xp33_ASAP7_75t_L      g04235(.A(new_n357), .B(new_n358), .C(new_n3856), .Y(new_n4492));
  OAI22xp33_ASAP7_75t_L     g04236(.A1(new_n4052), .A2(new_n298), .B1(new_n354), .B2(new_n4061), .Y(new_n4493));
  NOR3xp33_ASAP7_75t_L      g04237(.A(new_n4492), .B(new_n4493), .C(new_n4491), .Y(new_n4494));
  NAND2xp33_ASAP7_75t_L     g04238(.A(\a[35] ), .B(new_n4494), .Y(new_n4495));
  OAI31xp33_ASAP7_75t_L     g04239(.A1(new_n4492), .A2(new_n4491), .A3(new_n4493), .B(new_n3628), .Y(new_n4496));
  AOI21xp33_ASAP7_75t_L     g04240(.A1(new_n4274), .A2(new_n269), .B(new_n4278), .Y(new_n4497));
  NOR2xp33_ASAP7_75t_L      g04241(.A(new_n261), .B(new_n4277), .Y(new_n4498));
  NAND2xp33_ASAP7_75t_L     g04242(.A(new_n4282), .B(new_n4057), .Y(new_n4499));
  NAND2xp33_ASAP7_75t_L     g04243(.A(\b[2] ), .B(new_n4283), .Y(new_n4500));
  NAND3xp33_ASAP7_75t_L     g04244(.A(new_n4270), .B(new_n4282), .C(new_n4276), .Y(new_n4501));
  OAI221xp5_ASAP7_75t_L     g04245(.A1(new_n258), .A2(new_n4501), .B1(new_n280), .B2(new_n4499), .C(new_n4500), .Y(new_n4502));
  NOR2xp33_ASAP7_75t_L      g04246(.A(new_n4498), .B(new_n4502), .Y(new_n4503));
  A2O1A1Ixp33_ASAP7_75t_L   g04247(.A1(new_n4058), .A2(new_n4497), .B(new_n4268), .C(new_n4503), .Y(new_n4504));
  O2A1O1Ixp33_ASAP7_75t_L   g04248(.A1(new_n258), .A2(new_n4270), .B(new_n4497), .C(new_n4268), .Y(new_n4505));
  A2O1A1Ixp33_ASAP7_75t_L   g04249(.A1(\b[1] ), .A2(new_n4285), .B(new_n4502), .C(new_n4505), .Y(new_n4506));
  NAND4xp25_ASAP7_75t_L     g04250(.A(new_n4506), .B(new_n4495), .C(new_n4496), .D(new_n4504), .Y(new_n4507));
  NAND2xp33_ASAP7_75t_L     g04251(.A(new_n4496), .B(new_n4495), .Y(new_n4508));
  NAND3xp33_ASAP7_75t_L     g04252(.A(new_n4281), .B(new_n4284), .C(new_n4286), .Y(new_n4509));
  INVx1_ASAP7_75t_L         g04253(.A(new_n4498), .Y(new_n4510));
  NOR2xp33_ASAP7_75t_L      g04254(.A(new_n280), .B(new_n4499), .Y(new_n4511));
  AND3x1_ASAP7_75t_L        g04255(.A(new_n4270), .B(new_n4276), .C(new_n4282), .Y(new_n4512));
  AOI221xp5_ASAP7_75t_L     g04256(.A1(new_n4283), .A2(\b[2] ), .B1(new_n4512), .B2(\b[0] ), .C(new_n4511), .Y(new_n4513));
  NAND2xp33_ASAP7_75t_L     g04257(.A(new_n4510), .B(new_n4513), .Y(new_n4514));
  O2A1O1Ixp33_ASAP7_75t_L   g04258(.A1(new_n4059), .A2(new_n4509), .B(\a[38] ), .C(new_n4514), .Y(new_n4515));
  A2O1A1Ixp33_ASAP7_75t_L   g04259(.A1(\b[0] ), .A2(new_n4057), .B(new_n4509), .C(\a[38] ), .Y(new_n4516));
  O2A1O1Ixp33_ASAP7_75t_L   g04260(.A1(new_n4277), .A2(new_n261), .B(new_n4513), .C(new_n4516), .Y(new_n4517));
  OAI21xp33_ASAP7_75t_L     g04261(.A1(new_n4515), .A2(new_n4517), .B(new_n4508), .Y(new_n4518));
  AOI21xp33_ASAP7_75t_L     g04262(.A1(new_n4518), .A2(new_n4507), .B(new_n4490), .Y(new_n4519));
  AND3x1_ASAP7_75t_L        g04263(.A(new_n4490), .B(new_n4518), .C(new_n4507), .Y(new_n4520));
  OR3x1_ASAP7_75t_L         g04264(.A(new_n4520), .B(new_n4489), .C(new_n4519), .Y(new_n4521));
  OAI21xp33_ASAP7_75t_L     g04265(.A1(new_n4519), .A2(new_n4520), .B(new_n4489), .Y(new_n4522));
  NAND3xp33_ASAP7_75t_L     g04266(.A(new_n4486), .B(new_n4521), .C(new_n4522), .Y(new_n4523));
  A2O1A1O1Ixp25_ASAP7_75t_L g04267(.A1(new_n4085), .A2(new_n4095), .B(new_n4307), .C(new_n4298), .D(new_n4310), .Y(new_n4524));
  NOR3xp33_ASAP7_75t_L      g04268(.A(new_n4520), .B(new_n4489), .C(new_n4519), .Y(new_n4525));
  OA21x2_ASAP7_75t_L        g04269(.A1(new_n4519), .A2(new_n4520), .B(new_n4489), .Y(new_n4526));
  OAI21xp33_ASAP7_75t_L     g04270(.A1(new_n4525), .A2(new_n4526), .B(new_n4524), .Y(new_n4527));
  AOI21xp33_ASAP7_75t_L     g04271(.A1(new_n4523), .A2(new_n4527), .B(new_n4485), .Y(new_n4528));
  NAND2xp33_ASAP7_75t_L     g04272(.A(new_n4482), .B(new_n4484), .Y(new_n4529));
  NOR3xp33_ASAP7_75t_L      g04273(.A(new_n4524), .B(new_n4526), .C(new_n4525), .Y(new_n4530));
  AOI21xp33_ASAP7_75t_L     g04274(.A1(new_n4521), .A2(new_n4522), .B(new_n4486), .Y(new_n4531));
  NOR3xp33_ASAP7_75t_L      g04275(.A(new_n4530), .B(new_n4531), .C(new_n4529), .Y(new_n4532));
  OAI21xp33_ASAP7_75t_L     g04276(.A1(new_n4528), .A2(new_n4532), .B(new_n4478), .Y(new_n4533));
  OAI21xp33_ASAP7_75t_L     g04277(.A1(new_n4314), .A2(new_n4315), .B(new_n4251), .Y(new_n4534));
  A2O1A1O1Ixp25_ASAP7_75t_L g04278(.A1(new_n4101), .A2(new_n4050), .B(new_n4247), .C(new_n4534), .D(new_n4316), .Y(new_n4535));
  OAI21xp33_ASAP7_75t_L     g04279(.A1(new_n4531), .A2(new_n4530), .B(new_n4529), .Y(new_n4536));
  NAND3xp33_ASAP7_75t_L     g04280(.A(new_n4485), .B(new_n4523), .C(new_n4527), .Y(new_n4537));
  NAND3xp33_ASAP7_75t_L     g04281(.A(new_n4535), .B(new_n4536), .C(new_n4537), .Y(new_n4538));
  AO21x2_ASAP7_75t_L        g04282(.A1(new_n4538), .A2(new_n4533), .B(new_n4476), .Y(new_n4539));
  NAND3xp33_ASAP7_75t_L     g04283(.A(new_n4538), .B(new_n4533), .C(new_n4476), .Y(new_n4540));
  NAND3xp33_ASAP7_75t_L     g04284(.A(new_n4473), .B(new_n4539), .C(new_n4540), .Y(new_n4541));
  A2O1A1O1Ixp25_ASAP7_75t_L g04285(.A1(new_n4112), .A2(new_n4131), .B(new_n4128), .C(new_n4326), .D(new_n4322), .Y(new_n4542));
  NAND2xp33_ASAP7_75t_L     g04286(.A(new_n4540), .B(new_n4539), .Y(new_n4543));
  NAND2xp33_ASAP7_75t_L     g04287(.A(new_n4542), .B(new_n4543), .Y(new_n4544));
  NOR2xp33_ASAP7_75t_L      g04288(.A(new_n1030), .B(new_n1699), .Y(new_n4545));
  INVx1_ASAP7_75t_L         g04289(.A(new_n4545), .Y(new_n4546));
  NAND3xp33_ASAP7_75t_L     g04290(.A(new_n1206), .B(new_n1208), .C(new_n1695), .Y(new_n4547));
  AOI22xp33_ASAP7_75t_L     g04291(.A1(new_n1704), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1837), .Y(new_n4548));
  AND4x1_ASAP7_75t_L        g04292(.A(new_n4548), .B(new_n4547), .C(new_n4546), .D(\a[23] ), .Y(new_n4549));
  AOI31xp33_ASAP7_75t_L     g04293(.A1(new_n4547), .A2(new_n4546), .A3(new_n4548), .B(\a[23] ), .Y(new_n4550));
  NOR2xp33_ASAP7_75t_L      g04294(.A(new_n4550), .B(new_n4549), .Y(new_n4551));
  NAND3xp33_ASAP7_75t_L     g04295(.A(new_n4544), .B(new_n4541), .C(new_n4551), .Y(new_n4552));
  NOR2xp33_ASAP7_75t_L      g04296(.A(new_n4542), .B(new_n4543), .Y(new_n4553));
  AOI21xp33_ASAP7_75t_L     g04297(.A1(new_n4540), .A2(new_n4539), .B(new_n4473), .Y(new_n4554));
  INVx1_ASAP7_75t_L         g04298(.A(new_n4551), .Y(new_n4555));
  OAI21xp33_ASAP7_75t_L     g04299(.A1(new_n4554), .A2(new_n4553), .B(new_n4555), .Y(new_n4556));
  NAND2xp33_ASAP7_75t_L     g04300(.A(new_n4552), .B(new_n4556), .Y(new_n4557));
  XNOR2x2_ASAP7_75t_L       g04301(.A(new_n4325), .B(new_n4328), .Y(new_n4558));
  MAJIxp5_ASAP7_75t_L       g04302(.A(new_n4340), .B(new_n4558), .C(new_n4332), .Y(new_n4559));
  NOR2xp33_ASAP7_75t_L      g04303(.A(new_n4557), .B(new_n4559), .Y(new_n4560));
  NOR2xp33_ASAP7_75t_L      g04304(.A(new_n4336), .B(new_n4334), .Y(new_n4561));
  MAJIxp5_ASAP7_75t_L       g04305(.A(new_n4345), .B(new_n4337), .C(new_n4561), .Y(new_n4562));
  AOI21xp33_ASAP7_75t_L     g04306(.A1(new_n4556), .A2(new_n4552), .B(new_n4562), .Y(new_n4563));
  NAND2xp33_ASAP7_75t_L     g04307(.A(\b[19] ), .B(new_n1362), .Y(new_n4564));
  NAND2xp33_ASAP7_75t_L     g04308(.A(new_n1365), .B(new_n1886), .Y(new_n4565));
  AOI22xp33_ASAP7_75t_L     g04309(.A1(new_n1360), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1581), .Y(new_n4566));
  NAND4xp25_ASAP7_75t_L     g04310(.A(new_n4565), .B(\a[20] ), .C(new_n4564), .D(new_n4566), .Y(new_n4567));
  OAI21xp33_ASAP7_75t_L     g04311(.A1(new_n1359), .A2(new_n1547), .B(new_n4566), .Y(new_n4568));
  A2O1A1Ixp33_ASAP7_75t_L   g04312(.A1(\b[19] ), .A2(new_n1362), .B(new_n4568), .C(new_n1356), .Y(new_n4569));
  NAND2xp33_ASAP7_75t_L     g04313(.A(new_n4567), .B(new_n4569), .Y(new_n4570));
  NOR3xp33_ASAP7_75t_L      g04314(.A(new_n4560), .B(new_n4563), .C(new_n4570), .Y(new_n4571));
  NAND3xp33_ASAP7_75t_L     g04315(.A(new_n4562), .B(new_n4556), .C(new_n4552), .Y(new_n4572));
  NAND2xp33_ASAP7_75t_L     g04316(.A(new_n4557), .B(new_n4559), .Y(new_n4573));
  AND2x2_ASAP7_75t_L        g04317(.A(new_n4567), .B(new_n4569), .Y(new_n4574));
  AOI21xp33_ASAP7_75t_L     g04318(.A1(new_n4573), .A2(new_n4572), .B(new_n4574), .Y(new_n4575));
  NAND3xp33_ASAP7_75t_L     g04319(.A(new_n4341), .B(new_n4346), .C(new_n4353), .Y(new_n4576));
  A2O1A1Ixp33_ASAP7_75t_L   g04320(.A1(new_n4354), .A2(new_n4350), .B(new_n4356), .C(new_n4576), .Y(new_n4577));
  NOR3xp33_ASAP7_75t_L      g04321(.A(new_n4577), .B(new_n4575), .C(new_n4571), .Y(new_n4578));
  OA21x2_ASAP7_75t_L        g04322(.A1(new_n4571), .A2(new_n4575), .B(new_n4577), .Y(new_n4579));
  AOI22xp33_ASAP7_75t_L     g04323(.A1(new_n1076), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1253), .Y(new_n4580));
  OAI221xp5_ASAP7_75t_L     g04324(.A1(new_n1154), .A2(new_n1774), .B1(new_n1156), .B2(new_n1915), .C(new_n4580), .Y(new_n4581));
  XNOR2x2_ASAP7_75t_L       g04325(.A(\a[17] ), .B(new_n4581), .Y(new_n4582));
  OAI21xp33_ASAP7_75t_L     g04326(.A1(new_n4578), .A2(new_n4579), .B(new_n4582), .Y(new_n4583));
  NOR2xp33_ASAP7_75t_L      g04327(.A(new_n4575), .B(new_n4571), .Y(new_n4584));
  NAND2xp33_ASAP7_75t_L     g04328(.A(new_n4346), .B(new_n4341), .Y(new_n4585));
  MAJx2_ASAP7_75t_L         g04329(.A(new_n4356), .B(new_n4349), .C(new_n4585), .Y(new_n4586));
  NAND2xp33_ASAP7_75t_L     g04330(.A(new_n4584), .B(new_n4586), .Y(new_n4587));
  OAI21xp33_ASAP7_75t_L     g04331(.A1(new_n4571), .A2(new_n4575), .B(new_n4577), .Y(new_n4588));
  XNOR2x2_ASAP7_75t_L       g04332(.A(new_n1071), .B(new_n4581), .Y(new_n4589));
  NAND3xp33_ASAP7_75t_L     g04333(.A(new_n4587), .B(new_n4589), .C(new_n4588), .Y(new_n4590));
  AOI221xp5_ASAP7_75t_L     g04334(.A1(new_n4590), .A2(new_n4583), .B1(new_n4374), .B2(new_n4471), .C(new_n4472), .Y(new_n4591));
  INVx1_ASAP7_75t_L         g04335(.A(new_n4472), .Y(new_n4592));
  NAND2xp33_ASAP7_75t_L     g04336(.A(new_n4583), .B(new_n4590), .Y(new_n4593));
  AOI21xp33_ASAP7_75t_L     g04337(.A1(new_n4375), .A2(new_n4592), .B(new_n4593), .Y(new_n4594));
  OAI21xp33_ASAP7_75t_L     g04338(.A1(new_n4591), .A2(new_n4594), .B(new_n4470), .Y(new_n4595));
  O2A1O1Ixp33_ASAP7_75t_L   g04339(.A1(new_n4169), .A2(new_n4371), .B(new_n4374), .C(new_n4472), .Y(new_n4596));
  NAND2xp33_ASAP7_75t_L     g04340(.A(new_n4593), .B(new_n4596), .Y(new_n4597));
  AOI21xp33_ASAP7_75t_L     g04341(.A1(new_n4587), .A2(new_n4588), .B(new_n4589), .Y(new_n4598));
  NOR3xp33_ASAP7_75t_L      g04342(.A(new_n4579), .B(new_n4582), .C(new_n4578), .Y(new_n4599));
  NOR2xp33_ASAP7_75t_L      g04343(.A(new_n4599), .B(new_n4598), .Y(new_n4600));
  A2O1A1Ixp33_ASAP7_75t_L   g04344(.A1(new_n4471), .A2(new_n4374), .B(new_n4472), .C(new_n4600), .Y(new_n4601));
  OAI211xp5_ASAP7_75t_L     g04345(.A1(new_n4468), .A2(new_n4469), .B(new_n4601), .C(new_n4597), .Y(new_n4602));
  OAI211xp5_ASAP7_75t_L     g04346(.A1(new_n4177), .A2(new_n4174), .B(new_n4176), .C(new_n4383), .Y(new_n4603));
  NAND4xp25_ASAP7_75t_L     g04347(.A(new_n4602), .B(new_n4603), .C(new_n4382), .D(new_n4595), .Y(new_n4604));
  AO22x1_ASAP7_75t_L        g04348(.A1(new_n4382), .A2(new_n4603), .B1(new_n4595), .B2(new_n4602), .Y(new_n4605));
  AO21x2_ASAP7_75t_L        g04349(.A1(new_n4604), .A2(new_n4605), .B(new_n4465), .Y(new_n4606));
  NAND3xp33_ASAP7_75t_L     g04350(.A(new_n4605), .B(new_n4604), .C(new_n4465), .Y(new_n4607));
  NAND2xp33_ASAP7_75t_L     g04351(.A(new_n4607), .B(new_n4606), .Y(new_n4608));
  O2A1O1Ixp33_ASAP7_75t_L   g04352(.A1(new_n4461), .A2(new_n4462), .B(new_n4393), .C(new_n4608), .Y(new_n4609));
  NOR3xp33_ASAP7_75t_L      g04353(.A(new_n4387), .B(new_n4384), .C(new_n4241), .Y(new_n4610));
  A2O1A1O1Ixp25_ASAP7_75t_L g04354(.A1(new_n4032), .A2(new_n4190), .B(new_n4234), .C(new_n4388), .D(new_n4610), .Y(new_n4611));
  AND2x2_ASAP7_75t_L        g04355(.A(new_n4611), .B(new_n4608), .Y(new_n4612));
  OAI21xp33_ASAP7_75t_L     g04356(.A1(new_n4609), .A2(new_n4612), .B(new_n4460), .Y(new_n4613));
  AOI21xp33_ASAP7_75t_L     g04357(.A1(new_n4605), .A2(new_n4604), .B(new_n4465), .Y(new_n4614));
  AND3x1_ASAP7_75t_L        g04358(.A(new_n4605), .B(new_n4604), .C(new_n4465), .Y(new_n4615));
  NOR2xp33_ASAP7_75t_L      g04359(.A(new_n4614), .B(new_n4615), .Y(new_n4616));
  A2O1A1Ixp33_ASAP7_75t_L   g04360(.A1(new_n4388), .A2(new_n4236), .B(new_n4610), .C(new_n4616), .Y(new_n4617));
  NAND2xp33_ASAP7_75t_L     g04361(.A(new_n4611), .B(new_n4608), .Y(new_n4618));
  NAND3xp33_ASAP7_75t_L     g04362(.A(new_n4617), .B(new_n4459), .C(new_n4618), .Y(new_n4619));
  NAND2xp33_ASAP7_75t_L     g04363(.A(new_n4619), .B(new_n4613), .Y(new_n4620));
  O2A1O1Ixp33_ASAP7_75t_L   g04364(.A1(new_n4400), .A2(new_n4396), .B(new_n4402), .C(new_n4620), .Y(new_n4621));
  OAI21xp33_ASAP7_75t_L     g04365(.A1(new_n4396), .A2(new_n4400), .B(new_n4402), .Y(new_n4622));
  AOI21xp33_ASAP7_75t_L     g04366(.A1(new_n4619), .A2(new_n4613), .B(new_n4622), .Y(new_n4623));
  OAI21xp33_ASAP7_75t_L     g04367(.A1(new_n4623), .A2(new_n4621), .B(new_n4451), .Y(new_n4624));
  NAND3xp33_ASAP7_75t_L     g04368(.A(new_n4622), .B(new_n4613), .C(new_n4619), .Y(new_n4625));
  A2O1A1O1Ixp25_ASAP7_75t_L g04369(.A1(new_n4198), .A2(new_n4208), .B(new_n4197), .C(new_n4401), .D(new_n4397), .Y(new_n4626));
  NAND2xp33_ASAP7_75t_L     g04370(.A(new_n4626), .B(new_n4620), .Y(new_n4627));
  OAI211xp5_ASAP7_75t_L     g04371(.A1(new_n4449), .A2(new_n4450), .B(new_n4627), .C(new_n4625), .Y(new_n4628));
  NAND2xp33_ASAP7_75t_L     g04372(.A(new_n4628), .B(new_n4624), .Y(new_n4629));
  XNOR2x2_ASAP7_75t_L       g04373(.A(new_n4444), .B(new_n4629), .Y(new_n4630));
  NOR2xp33_ASAP7_75t_L      g04374(.A(\b[37] ), .B(\b[38] ), .Y(new_n4631));
  INVx1_ASAP7_75t_L         g04375(.A(\b[38] ), .Y(new_n4632));
  NOR2xp33_ASAP7_75t_L      g04376(.A(new_n4424), .B(new_n4632), .Y(new_n4633));
  NOR2xp33_ASAP7_75t_L      g04377(.A(new_n4631), .B(new_n4633), .Y(new_n4634));
  INVx1_ASAP7_75t_L         g04378(.A(new_n4634), .Y(new_n4635));
  O2A1O1Ixp33_ASAP7_75t_L   g04379(.A1(new_n4216), .A2(new_n4424), .B(new_n4427), .C(new_n4635), .Y(new_n4636));
  INVx1_ASAP7_75t_L         g04380(.A(new_n4217), .Y(new_n4637));
  O2A1O1Ixp33_ASAP7_75t_L   g04381(.A1(new_n4221), .A2(new_n4220), .B(new_n4637), .C(new_n4429), .Y(new_n4638));
  NOR3xp33_ASAP7_75t_L      g04382(.A(new_n4638), .B(new_n4634), .C(new_n4425), .Y(new_n4639));
  NOR2xp33_ASAP7_75t_L      g04383(.A(new_n4639), .B(new_n4636), .Y(new_n4640));
  INVx1_ASAP7_75t_L         g04384(.A(new_n4640), .Y(new_n4641));
  AOI22xp33_ASAP7_75t_L     g04385(.A1(\b[36] ), .A2(new_n282), .B1(\b[38] ), .B2(new_n303), .Y(new_n4642));
  OAI221xp5_ASAP7_75t_L     g04386(.A1(new_n291), .A2(new_n4424), .B1(new_n268), .B2(new_n4641), .C(new_n4642), .Y(new_n4643));
  XNOR2x2_ASAP7_75t_L       g04387(.A(\a[2] ), .B(new_n4643), .Y(new_n4644));
  INVx1_ASAP7_75t_L         g04388(.A(new_n4644), .Y(new_n4645));
  XNOR2x2_ASAP7_75t_L       g04389(.A(new_n4645), .B(new_n4630), .Y(new_n4646));
  AO21x2_ASAP7_75t_L        g04390(.A1(new_n4435), .A2(new_n4440), .B(new_n4436), .Y(new_n4647));
  XNOR2x2_ASAP7_75t_L       g04391(.A(new_n4647), .B(new_n4646), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g04392(.A(new_n4407), .B(new_n4443), .Y(new_n4649));
  NOR3xp33_ASAP7_75t_L      g04393(.A(new_n4621), .B(new_n4451), .C(new_n4623), .Y(new_n4650));
  A2O1A1O1Ixp25_ASAP7_75t_L g04394(.A1(new_n4416), .A2(new_n4413), .B(new_n4649), .C(new_n4624), .D(new_n4650), .Y(new_n4651));
  AOI22xp33_ASAP7_75t_L     g04395(.A1(new_n344), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n370), .Y(new_n4652));
  OAI221xp5_ASAP7_75t_L     g04396(.A1(new_n429), .A2(new_n3804), .B1(new_n366), .B2(new_n4223), .C(new_n4652), .Y(new_n4653));
  XNOR2x2_ASAP7_75t_L       g04397(.A(\a[5] ), .B(new_n4653), .Y(new_n4654));
  AOI21xp33_ASAP7_75t_L     g04398(.A1(new_n4617), .A2(new_n4618), .B(new_n4459), .Y(new_n4655));
  OAI21xp33_ASAP7_75t_L     g04399(.A1(new_n4614), .A2(new_n4611), .B(new_n4607), .Y(new_n4656));
  AOI22xp33_ASAP7_75t_L     g04400(.A1(\b[28] ), .A2(new_n651), .B1(\b[30] ), .B2(new_n581), .Y(new_n4657));
  OAI221xp5_ASAP7_75t_L     g04401(.A1(new_n821), .A2(new_n2688), .B1(new_n577), .B2(new_n2990), .C(new_n4657), .Y(new_n4658));
  XNOR2x2_ASAP7_75t_L       g04402(.A(\a[11] ), .B(new_n4658), .Y(new_n4659));
  INVx1_ASAP7_75t_L         g04403(.A(new_n4659), .Y(new_n4660));
  NOR3xp33_ASAP7_75t_L      g04404(.A(new_n4594), .B(new_n4591), .C(new_n4470), .Y(new_n4661));
  AOI31xp33_ASAP7_75t_L     g04405(.A1(new_n4603), .A2(new_n4595), .A3(new_n4382), .B(new_n4661), .Y(new_n4662));
  NOR3xp33_ASAP7_75t_L      g04406(.A(new_n4553), .B(new_n4554), .C(new_n4551), .Y(new_n4663));
  OAI22xp33_ASAP7_75t_L     g04407(.A1(new_n1829), .A2(new_n1030), .B1(new_n1313), .B2(new_n1696), .Y(new_n4664));
  AOI221xp5_ASAP7_75t_L     g04408(.A1(new_n1706), .A2(\b[17] ), .B1(new_n1695), .B2(new_n1319), .C(new_n4664), .Y(new_n4665));
  AND2x2_ASAP7_75t_L        g04409(.A(\a[23] ), .B(new_n4665), .Y(new_n4666));
  NOR2xp33_ASAP7_75t_L      g04410(.A(\a[23] ), .B(new_n4665), .Y(new_n4667));
  OAI21xp33_ASAP7_75t_L     g04411(.A1(new_n4542), .A2(new_n4543), .B(new_n4540), .Y(new_n4668));
  NAND5xp2_ASAP7_75t_L      g04412(.A(\a[38] ), .B(new_n4281), .C(new_n4284), .D(new_n4286), .E(new_n4058), .Y(new_n4669));
  INVx1_ASAP7_75t_L         g04413(.A(\a[39] ), .Y(new_n4670));
  NAND2xp33_ASAP7_75t_L     g04414(.A(\a[38] ), .B(new_n4670), .Y(new_n4671));
  NAND2xp33_ASAP7_75t_L     g04415(.A(\a[39] ), .B(new_n4268), .Y(new_n4672));
  AND2x2_ASAP7_75t_L        g04416(.A(new_n4671), .B(new_n4672), .Y(new_n4673));
  NOR2xp33_ASAP7_75t_L      g04417(.A(new_n258), .B(new_n4673), .Y(new_n4674));
  OAI31xp33_ASAP7_75t_L     g04418(.A1(new_n4669), .A2(new_n4502), .A3(new_n4498), .B(new_n4674), .Y(new_n4675));
  NOR2xp33_ASAP7_75t_L      g04419(.A(new_n4268), .B(new_n4059), .Y(new_n4676));
  INVx1_ASAP7_75t_L         g04420(.A(new_n4674), .Y(new_n4677));
  NAND5xp2_ASAP7_75t_L      g04421(.A(new_n4497), .B(new_n4677), .C(new_n4513), .D(new_n4676), .E(new_n4510), .Y(new_n4678));
  NOR2xp33_ASAP7_75t_L      g04422(.A(new_n276), .B(new_n4277), .Y(new_n4679));
  NAND2xp33_ASAP7_75t_L     g04423(.A(\b[3] ), .B(new_n4283), .Y(new_n4680));
  OAI221xp5_ASAP7_75t_L     g04424(.A1(new_n4501), .A2(new_n261), .B1(new_n4499), .B2(new_n302), .C(new_n4680), .Y(new_n4681));
  OR3x1_ASAP7_75t_L         g04425(.A(new_n4681), .B(new_n4268), .C(new_n4679), .Y(new_n4682));
  A2O1A1Ixp33_ASAP7_75t_L   g04426(.A1(\b[2] ), .A2(new_n4285), .B(new_n4681), .C(new_n4268), .Y(new_n4683));
  AO22x1_ASAP7_75t_L        g04427(.A1(new_n4675), .A2(new_n4678), .B1(new_n4683), .B2(new_n4682), .Y(new_n4684));
  NAND4xp25_ASAP7_75t_L     g04428(.A(new_n4682), .B(new_n4678), .C(new_n4675), .D(new_n4683), .Y(new_n4685));
  NAND2xp33_ASAP7_75t_L     g04429(.A(\b[5] ), .B(new_n3639), .Y(new_n4686));
  NAND2xp33_ASAP7_75t_L     g04430(.A(new_n3630), .B(new_n526), .Y(new_n4687));
  AOI22xp33_ASAP7_75t_L     g04431(.A1(new_n3633), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n3858), .Y(new_n4688));
  NAND4xp25_ASAP7_75t_L     g04432(.A(new_n4687), .B(\a[35] ), .C(new_n4686), .D(new_n4688), .Y(new_n4689));
  AOI31xp33_ASAP7_75t_L     g04433(.A1(new_n4687), .A2(new_n4686), .A3(new_n4688), .B(\a[35] ), .Y(new_n4690));
  INVx1_ASAP7_75t_L         g04434(.A(new_n4690), .Y(new_n4691));
  NAND4xp25_ASAP7_75t_L     g04435(.A(new_n4691), .B(new_n4684), .C(new_n4685), .D(new_n4689), .Y(new_n4692));
  AOI22xp33_ASAP7_75t_L     g04436(.A1(new_n4678), .A2(new_n4675), .B1(new_n4683), .B2(new_n4682), .Y(new_n4693));
  AND4x1_ASAP7_75t_L        g04437(.A(new_n4678), .B(new_n4682), .C(new_n4675), .D(new_n4683), .Y(new_n4694));
  INVx1_ASAP7_75t_L         g04438(.A(new_n4689), .Y(new_n4695));
  OAI22xp33_ASAP7_75t_L     g04439(.A1(new_n4695), .A2(new_n4690), .B1(new_n4693), .B2(new_n4694), .Y(new_n4696));
  NAND2xp33_ASAP7_75t_L     g04440(.A(new_n4696), .B(new_n4692), .Y(new_n4697));
  NOR2xp33_ASAP7_75t_L      g04441(.A(new_n4515), .B(new_n4517), .Y(new_n4698));
  NAND2xp33_ASAP7_75t_L     g04442(.A(new_n4508), .B(new_n4698), .Y(new_n4699));
  A2O1A1Ixp33_ASAP7_75t_L   g04443(.A1(new_n4507), .A2(new_n4518), .B(new_n4490), .C(new_n4699), .Y(new_n4700));
  NOR2xp33_ASAP7_75t_L      g04444(.A(new_n4697), .B(new_n4700), .Y(new_n4701));
  AND2x2_ASAP7_75t_L        g04445(.A(new_n4696), .B(new_n4692), .Y(new_n4702));
  A2O1A1Ixp33_ASAP7_75t_L   g04446(.A1(new_n4072), .A2(new_n4261), .B(new_n4289), .C(new_n4296), .Y(new_n4703));
  MAJIxp5_ASAP7_75t_L       g04447(.A(new_n4703), .B(new_n4508), .C(new_n4698), .Y(new_n4704));
  NOR2xp33_ASAP7_75t_L      g04448(.A(new_n4704), .B(new_n4702), .Y(new_n4705));
  NAND2xp33_ASAP7_75t_L     g04449(.A(\b[8] ), .B(new_n3030), .Y(new_n4706));
  NAND2xp33_ASAP7_75t_L     g04450(.A(new_n3021), .B(new_n731), .Y(new_n4707));
  AOI22xp33_ASAP7_75t_L     g04451(.A1(new_n3029), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n3258), .Y(new_n4708));
  NAND4xp25_ASAP7_75t_L     g04452(.A(new_n4707), .B(\a[32] ), .C(new_n4706), .D(new_n4708), .Y(new_n4709));
  OAI21xp33_ASAP7_75t_L     g04453(.A1(new_n3256), .A2(new_n548), .B(new_n4708), .Y(new_n4710));
  A2O1A1Ixp33_ASAP7_75t_L   g04454(.A1(\b[8] ), .A2(new_n3030), .B(new_n4710), .C(new_n3015), .Y(new_n4711));
  NAND2xp33_ASAP7_75t_L     g04455(.A(new_n4711), .B(new_n4709), .Y(new_n4712));
  NOR3xp33_ASAP7_75t_L      g04456(.A(new_n4712), .B(new_n4705), .C(new_n4701), .Y(new_n4713));
  NAND2xp33_ASAP7_75t_L     g04457(.A(new_n4704), .B(new_n4702), .Y(new_n4714));
  A2O1A1Ixp33_ASAP7_75t_L   g04458(.A1(new_n4698), .A2(new_n4508), .B(new_n4519), .C(new_n4697), .Y(new_n4715));
  AOI22xp33_ASAP7_75t_L     g04459(.A1(new_n4709), .A2(new_n4711), .B1(new_n4715), .B2(new_n4714), .Y(new_n4716));
  OAI21xp33_ASAP7_75t_L     g04460(.A1(new_n4526), .A2(new_n4524), .B(new_n4521), .Y(new_n4717));
  NOR3xp33_ASAP7_75t_L      g04461(.A(new_n4717), .B(new_n4716), .C(new_n4713), .Y(new_n4718));
  NAND4xp25_ASAP7_75t_L     g04462(.A(new_n4714), .B(new_n4715), .C(new_n4711), .D(new_n4709), .Y(new_n4719));
  OAI21xp33_ASAP7_75t_L     g04463(.A1(new_n4701), .A2(new_n4705), .B(new_n4712), .Y(new_n4720));
  A2O1A1O1Ixp25_ASAP7_75t_L g04464(.A1(new_n4298), .A2(new_n4255), .B(new_n4310), .C(new_n4522), .D(new_n4525), .Y(new_n4721));
  AOI21xp33_ASAP7_75t_L     g04465(.A1(new_n4720), .A2(new_n4719), .B(new_n4721), .Y(new_n4722));
  NOR2xp33_ASAP7_75t_L      g04466(.A(new_n679), .B(new_n2547), .Y(new_n4723));
  AOI22xp33_ASAP7_75t_L     g04467(.A1(new_n2552), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n2736), .Y(new_n4724));
  OAI31xp33_ASAP7_75t_L     g04468(.A1(new_n1231), .A2(new_n764), .A3(new_n2734), .B(new_n4724), .Y(new_n4725));
  OR3x1_ASAP7_75t_L         g04469(.A(new_n4725), .B(new_n2538), .C(new_n4723), .Y(new_n4726));
  A2O1A1Ixp33_ASAP7_75t_L   g04470(.A1(\b[11] ), .A2(new_n2553), .B(new_n4725), .C(new_n2538), .Y(new_n4727));
  AND2x2_ASAP7_75t_L        g04471(.A(new_n4727), .B(new_n4726), .Y(new_n4728));
  OAI21xp33_ASAP7_75t_L     g04472(.A1(new_n4722), .A2(new_n4718), .B(new_n4728), .Y(new_n4729));
  NAND3xp33_ASAP7_75t_L     g04473(.A(new_n4721), .B(new_n4720), .C(new_n4719), .Y(new_n4730));
  OAI21xp33_ASAP7_75t_L     g04474(.A1(new_n4713), .A2(new_n4716), .B(new_n4717), .Y(new_n4731));
  NAND2xp33_ASAP7_75t_L     g04475(.A(new_n4727), .B(new_n4726), .Y(new_n4732));
  NAND3xp33_ASAP7_75t_L     g04476(.A(new_n4730), .B(new_n4731), .C(new_n4732), .Y(new_n4733));
  NAND2xp33_ASAP7_75t_L     g04477(.A(new_n4527), .B(new_n4523), .Y(new_n4734));
  MAJIxp5_ASAP7_75t_L       g04478(.A(new_n4535), .B(new_n4485), .C(new_n4734), .Y(new_n4735));
  NAND3xp33_ASAP7_75t_L     g04479(.A(new_n4735), .B(new_n4733), .C(new_n4729), .Y(new_n4736));
  INVx1_ASAP7_75t_L         g04480(.A(new_n4729), .Y(new_n4737));
  NOR3xp33_ASAP7_75t_L      g04481(.A(new_n4718), .B(new_n4728), .C(new_n4722), .Y(new_n4738));
  NOR2xp33_ASAP7_75t_L      g04482(.A(new_n4485), .B(new_n4734), .Y(new_n4739));
  O2A1O1Ixp33_ASAP7_75t_L   g04483(.A1(new_n4528), .A2(new_n4532), .B(new_n4478), .C(new_n4739), .Y(new_n4740));
  OAI21xp33_ASAP7_75t_L     g04484(.A1(new_n4738), .A2(new_n4737), .B(new_n4740), .Y(new_n4741));
  AOI22xp33_ASAP7_75t_L     g04485(.A1(new_n2114), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n2259), .Y(new_n4742));
  OAI221xp5_ASAP7_75t_L     g04486(.A1(new_n2109), .A2(new_n869), .B1(new_n2257), .B2(new_n950), .C(new_n4742), .Y(new_n4743));
  XNOR2x2_ASAP7_75t_L       g04487(.A(\a[26] ), .B(new_n4743), .Y(new_n4744));
  NAND3xp33_ASAP7_75t_L     g04488(.A(new_n4741), .B(new_n4736), .C(new_n4744), .Y(new_n4745));
  NOR3xp33_ASAP7_75t_L      g04489(.A(new_n4740), .B(new_n4738), .C(new_n4737), .Y(new_n4746));
  AOI21xp33_ASAP7_75t_L     g04490(.A1(new_n4733), .A2(new_n4729), .B(new_n4735), .Y(new_n4747));
  XNOR2x2_ASAP7_75t_L       g04491(.A(new_n2100), .B(new_n4743), .Y(new_n4748));
  OAI21xp33_ASAP7_75t_L     g04492(.A1(new_n4747), .A2(new_n4746), .B(new_n4748), .Y(new_n4749));
  NAND2xp33_ASAP7_75t_L     g04493(.A(new_n4745), .B(new_n4749), .Y(new_n4750));
  NAND2xp33_ASAP7_75t_L     g04494(.A(new_n4668), .B(new_n4750), .Y(new_n4751));
  AND3x1_ASAP7_75t_L        g04495(.A(new_n4533), .B(new_n4538), .C(new_n4476), .Y(new_n4752));
  A2O1A1O1Ixp25_ASAP7_75t_L g04496(.A1(new_n4326), .A2(new_n4335), .B(new_n4322), .C(new_n4539), .D(new_n4752), .Y(new_n4753));
  NAND3xp33_ASAP7_75t_L     g04497(.A(new_n4753), .B(new_n4745), .C(new_n4749), .Y(new_n4754));
  OAI211xp5_ASAP7_75t_L     g04498(.A1(new_n4667), .A2(new_n4666), .B(new_n4751), .C(new_n4754), .Y(new_n4755));
  XNOR2x2_ASAP7_75t_L       g04499(.A(new_n1689), .B(new_n4665), .Y(new_n4756));
  AOI21xp33_ASAP7_75t_L     g04500(.A1(new_n4749), .A2(new_n4745), .B(new_n4753), .Y(new_n4757));
  NOR2xp33_ASAP7_75t_L      g04501(.A(new_n4668), .B(new_n4750), .Y(new_n4758));
  OAI21xp33_ASAP7_75t_L     g04502(.A1(new_n4757), .A2(new_n4758), .B(new_n4756), .Y(new_n4759));
  AO221x2_ASAP7_75t_L       g04503(.A1(new_n4559), .A2(new_n4557), .B1(new_n4755), .B2(new_n4759), .C(new_n4663), .Y(new_n4760));
  INVx1_ASAP7_75t_L         g04504(.A(new_n4663), .Y(new_n4761));
  A2O1A1Ixp33_ASAP7_75t_L   g04505(.A1(new_n4556), .A2(new_n4552), .B(new_n4562), .C(new_n4761), .Y(new_n4762));
  NAND3xp33_ASAP7_75t_L     g04506(.A(new_n4762), .B(new_n4755), .C(new_n4759), .Y(new_n4763));
  AOI22xp33_ASAP7_75t_L     g04507(.A1(new_n1360), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1581), .Y(new_n4764));
  OAI221xp5_ASAP7_75t_L     g04508(.A1(new_n1373), .A2(new_n1539), .B1(new_n1359), .B2(new_n1662), .C(new_n4764), .Y(new_n4765));
  XNOR2x2_ASAP7_75t_L       g04509(.A(\a[20] ), .B(new_n4765), .Y(new_n4766));
  NAND3xp33_ASAP7_75t_L     g04510(.A(new_n4763), .B(new_n4760), .C(new_n4766), .Y(new_n4767));
  AOI21xp33_ASAP7_75t_L     g04511(.A1(new_n4759), .A2(new_n4755), .B(new_n4762), .Y(new_n4768));
  NAND2xp33_ASAP7_75t_L     g04512(.A(new_n4759), .B(new_n4755), .Y(new_n4769));
  AOI21xp33_ASAP7_75t_L     g04513(.A1(new_n4573), .A2(new_n4761), .B(new_n4769), .Y(new_n4770));
  XNOR2x2_ASAP7_75t_L       g04514(.A(new_n1356), .B(new_n4765), .Y(new_n4771));
  OAI21xp33_ASAP7_75t_L     g04515(.A1(new_n4768), .A2(new_n4770), .B(new_n4771), .Y(new_n4772));
  NAND2xp33_ASAP7_75t_L     g04516(.A(new_n4767), .B(new_n4772), .Y(new_n4773));
  NOR3xp33_ASAP7_75t_L      g04517(.A(new_n4574), .B(new_n4560), .C(new_n4563), .Y(new_n4774));
  NOR3xp33_ASAP7_75t_L      g04518(.A(new_n4773), .B(new_n4579), .C(new_n4774), .Y(new_n4775));
  O2A1O1Ixp33_ASAP7_75t_L   g04519(.A1(new_n4571), .A2(new_n4575), .B(new_n4577), .C(new_n4774), .Y(new_n4776));
  AOI21xp33_ASAP7_75t_L     g04520(.A1(new_n4772), .A2(new_n4767), .B(new_n4776), .Y(new_n4777));
  OAI22xp33_ASAP7_75t_L     g04521(.A1(new_n1158), .A2(new_n1774), .B1(new_n1929), .B2(new_n1259), .Y(new_n4778));
  AOI221xp5_ASAP7_75t_L     g04522(.A1(\b[23] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n1935), .C(new_n4778), .Y(new_n4779));
  XNOR2x2_ASAP7_75t_L       g04523(.A(new_n1071), .B(new_n4779), .Y(new_n4780));
  OAI21xp33_ASAP7_75t_L     g04524(.A1(new_n4777), .A2(new_n4775), .B(new_n4780), .Y(new_n4781));
  NAND3xp33_ASAP7_75t_L     g04525(.A(new_n4776), .B(new_n4772), .C(new_n4767), .Y(new_n4782));
  OAI21xp33_ASAP7_75t_L     g04526(.A1(new_n4774), .A2(new_n4579), .B(new_n4773), .Y(new_n4783));
  XNOR2x2_ASAP7_75t_L       g04527(.A(\a[17] ), .B(new_n4779), .Y(new_n4784));
  NAND3xp33_ASAP7_75t_L     g04528(.A(new_n4783), .B(new_n4784), .C(new_n4782), .Y(new_n4785));
  NOR3xp33_ASAP7_75t_L      g04529(.A(new_n4369), .B(new_n4367), .C(new_n4368), .Y(new_n4786));
  AOI21xp33_ASAP7_75t_L     g04530(.A1(new_n4359), .A2(new_n4357), .B(new_n4365), .Y(new_n4787));
  NOR2xp33_ASAP7_75t_L      g04531(.A(new_n4786), .B(new_n4787), .Y(new_n4788));
  NAND2xp33_ASAP7_75t_L     g04532(.A(new_n4167), .B(new_n4168), .Y(new_n4789));
  AOI31xp33_ASAP7_75t_L     g04533(.A1(new_n4789), .A2(new_n3942), .A3(new_n4160), .B(new_n4371), .Y(new_n4790));
  OAI211xp5_ASAP7_75t_L     g04534(.A1(new_n4788), .A2(new_n4790), .B(new_n4592), .C(new_n4590), .Y(new_n4791));
  NAND4xp25_ASAP7_75t_L     g04535(.A(new_n4791), .B(new_n4781), .C(new_n4583), .D(new_n4785), .Y(new_n4792));
  AOI21xp33_ASAP7_75t_L     g04536(.A1(new_n4783), .A2(new_n4782), .B(new_n4784), .Y(new_n4793));
  NOR3xp33_ASAP7_75t_L      g04537(.A(new_n4775), .B(new_n4777), .C(new_n4780), .Y(new_n4794));
  AOI211xp5_ASAP7_75t_L     g04538(.A1(new_n4471), .A2(new_n4374), .B(new_n4472), .C(new_n4599), .Y(new_n4795));
  OAI22xp33_ASAP7_75t_L     g04539(.A1(new_n4795), .A2(new_n4598), .B1(new_n4793), .B2(new_n4794), .Y(new_n4796));
  NAND2xp33_ASAP7_75t_L     g04540(.A(\b[26] ), .B(new_n815), .Y(new_n4797));
  NAND2xp33_ASAP7_75t_L     g04541(.A(new_n808), .B(new_n2504), .Y(new_n4798));
  AOI22xp33_ASAP7_75t_L     g04542(.A1(new_n811), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n900), .Y(new_n4799));
  NAND4xp25_ASAP7_75t_L     g04543(.A(new_n4798), .B(\a[14] ), .C(new_n4797), .D(new_n4799), .Y(new_n4800));
  NAND2xp33_ASAP7_75t_L     g04544(.A(new_n4799), .B(new_n4798), .Y(new_n4801));
  A2O1A1Ixp33_ASAP7_75t_L   g04545(.A1(\b[26] ), .A2(new_n815), .B(new_n4801), .C(new_n806), .Y(new_n4802));
  AND2x2_ASAP7_75t_L        g04546(.A(new_n4800), .B(new_n4802), .Y(new_n4803));
  NAND3xp33_ASAP7_75t_L     g04547(.A(new_n4796), .B(new_n4792), .C(new_n4803), .Y(new_n4804));
  NOR4xp25_ASAP7_75t_L      g04548(.A(new_n4795), .B(new_n4598), .C(new_n4793), .D(new_n4794), .Y(new_n4805));
  AOI22xp33_ASAP7_75t_L     g04549(.A1(new_n4785), .A2(new_n4781), .B1(new_n4583), .B2(new_n4791), .Y(new_n4806));
  NAND2xp33_ASAP7_75t_L     g04550(.A(new_n4800), .B(new_n4802), .Y(new_n4807));
  OAI21xp33_ASAP7_75t_L     g04551(.A1(new_n4806), .A2(new_n4805), .B(new_n4807), .Y(new_n4808));
  AOI21xp33_ASAP7_75t_L     g04552(.A1(new_n4804), .A2(new_n4808), .B(new_n4662), .Y(new_n4809));
  INVx1_ASAP7_75t_L         g04553(.A(new_n4809), .Y(new_n4810));
  NAND3xp33_ASAP7_75t_L     g04554(.A(new_n4662), .B(new_n4804), .C(new_n4808), .Y(new_n4811));
  NAND3xp33_ASAP7_75t_L     g04555(.A(new_n4810), .B(new_n4660), .C(new_n4811), .Y(new_n4812));
  INVx1_ASAP7_75t_L         g04556(.A(new_n4811), .Y(new_n4813));
  OAI21xp33_ASAP7_75t_L     g04557(.A1(new_n4809), .A2(new_n4813), .B(new_n4659), .Y(new_n4814));
  NAND3xp33_ASAP7_75t_L     g04558(.A(new_n4656), .B(new_n4812), .C(new_n4814), .Y(new_n4815));
  A2O1A1O1Ixp25_ASAP7_75t_L g04559(.A1(new_n4388), .A2(new_n4236), .B(new_n4610), .C(new_n4606), .D(new_n4615), .Y(new_n4816));
  NOR3xp33_ASAP7_75t_L      g04560(.A(new_n4813), .B(new_n4809), .C(new_n4659), .Y(new_n4817));
  AOI21xp33_ASAP7_75t_L     g04561(.A1(new_n4810), .A2(new_n4811), .B(new_n4660), .Y(new_n4818));
  OAI21xp33_ASAP7_75t_L     g04562(.A1(new_n4818), .A2(new_n4817), .B(new_n4816), .Y(new_n4819));
  NAND2xp33_ASAP7_75t_L     g04563(.A(\b[32] ), .B(new_n447), .Y(new_n4820));
  NOR2xp33_ASAP7_75t_L      g04564(.A(new_n3570), .B(new_n3582), .Y(new_n4821));
  NAND2xp33_ASAP7_75t_L     g04565(.A(new_n441), .B(new_n4821), .Y(new_n4822));
  AOI22xp33_ASAP7_75t_L     g04566(.A1(new_n444), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n471), .Y(new_n4823));
  NAND4xp25_ASAP7_75t_L     g04567(.A(new_n4822), .B(\a[8] ), .C(new_n4820), .D(new_n4823), .Y(new_n4824));
  NAND2xp33_ASAP7_75t_L     g04568(.A(new_n4823), .B(new_n4822), .Y(new_n4825));
  A2O1A1Ixp33_ASAP7_75t_L   g04569(.A1(\b[32] ), .A2(new_n447), .B(new_n4825), .C(new_n435), .Y(new_n4826));
  AND2x2_ASAP7_75t_L        g04570(.A(new_n4824), .B(new_n4826), .Y(new_n4827));
  NAND3xp33_ASAP7_75t_L     g04571(.A(new_n4815), .B(new_n4827), .C(new_n4819), .Y(new_n4828));
  NOR3xp33_ASAP7_75t_L      g04572(.A(new_n4816), .B(new_n4817), .C(new_n4818), .Y(new_n4829));
  AOI21xp33_ASAP7_75t_L     g04573(.A1(new_n4814), .A2(new_n4812), .B(new_n4656), .Y(new_n4830));
  NAND2xp33_ASAP7_75t_L     g04574(.A(new_n4824), .B(new_n4826), .Y(new_n4831));
  OAI21xp33_ASAP7_75t_L     g04575(.A1(new_n4829), .A2(new_n4830), .B(new_n4831), .Y(new_n4832));
  AND2x2_ASAP7_75t_L        g04576(.A(new_n4828), .B(new_n4832), .Y(new_n4833));
  O2A1O1Ixp33_ASAP7_75t_L   g04577(.A1(new_n4626), .A2(new_n4655), .B(new_n4619), .C(new_n4833), .Y(new_n4834));
  OAI21xp33_ASAP7_75t_L     g04578(.A1(new_n4655), .A2(new_n4626), .B(new_n4619), .Y(new_n4835));
  NAND2xp33_ASAP7_75t_L     g04579(.A(new_n4828), .B(new_n4832), .Y(new_n4836));
  NOR2xp33_ASAP7_75t_L      g04580(.A(new_n4836), .B(new_n4835), .Y(new_n4837));
  OAI21xp33_ASAP7_75t_L     g04581(.A1(new_n4837), .A2(new_n4834), .B(new_n4654), .Y(new_n4838));
  INVx1_ASAP7_75t_L         g04582(.A(new_n4654), .Y(new_n4839));
  NAND2xp33_ASAP7_75t_L     g04583(.A(new_n4836), .B(new_n4835), .Y(new_n4840));
  INVx1_ASAP7_75t_L         g04584(.A(new_n4837), .Y(new_n4841));
  NAND3xp33_ASAP7_75t_L     g04585(.A(new_n4841), .B(new_n4839), .C(new_n4840), .Y(new_n4842));
  NAND2xp33_ASAP7_75t_L     g04586(.A(new_n4838), .B(new_n4842), .Y(new_n4843));
  XNOR2x2_ASAP7_75t_L       g04587(.A(new_n4651), .B(new_n4843), .Y(new_n4844));
  A2O1A1O1Ixp25_ASAP7_75t_L g04588(.A1(new_n4218), .A2(new_n4422), .B(new_n4217), .C(new_n4426), .D(new_n4425), .Y(new_n4845));
  INVx1_ASAP7_75t_L         g04589(.A(new_n4633), .Y(new_n4846));
  NOR2xp33_ASAP7_75t_L      g04590(.A(\b[38] ), .B(\b[39] ), .Y(new_n4847));
  INVx1_ASAP7_75t_L         g04591(.A(\b[39] ), .Y(new_n4848));
  NOR2xp33_ASAP7_75t_L      g04592(.A(new_n4632), .B(new_n4848), .Y(new_n4849));
  NOR2xp33_ASAP7_75t_L      g04593(.A(new_n4847), .B(new_n4849), .Y(new_n4850));
  INVx1_ASAP7_75t_L         g04594(.A(new_n4850), .Y(new_n4851));
  O2A1O1Ixp33_ASAP7_75t_L   g04595(.A1(new_n4635), .A2(new_n4845), .B(new_n4846), .C(new_n4851), .Y(new_n4852));
  INVx1_ASAP7_75t_L         g04596(.A(new_n4852), .Y(new_n4853));
  INVx1_ASAP7_75t_L         g04597(.A(new_n3808), .Y(new_n4854));
  A2O1A1Ixp33_ASAP7_75t_L   g04598(.A1(new_n4854), .A2(new_n4421), .B(new_n4215), .C(new_n4637), .Y(new_n4855));
  A2O1A1O1Ixp25_ASAP7_75t_L g04599(.A1(new_n4426), .A2(new_n4855), .B(new_n4425), .C(new_n4634), .D(new_n4633), .Y(new_n4856));
  NAND2xp33_ASAP7_75t_L     g04600(.A(new_n4851), .B(new_n4856), .Y(new_n4857));
  NAND2xp33_ASAP7_75t_L     g04601(.A(new_n4857), .B(new_n4853), .Y(new_n4858));
  AOI22xp33_ASAP7_75t_L     g04602(.A1(\b[37] ), .A2(new_n282), .B1(\b[39] ), .B2(new_n303), .Y(new_n4859));
  OAI221xp5_ASAP7_75t_L     g04603(.A1(new_n291), .A2(new_n4632), .B1(new_n268), .B2(new_n4858), .C(new_n4859), .Y(new_n4860));
  XNOR2x2_ASAP7_75t_L       g04604(.A(\a[2] ), .B(new_n4860), .Y(new_n4861));
  XOR2x2_ASAP7_75t_L        g04605(.A(new_n4861), .B(new_n4844), .Y(new_n4862));
  MAJIxp5_ASAP7_75t_L       g04606(.A(new_n4647), .B(new_n4645), .C(new_n4630), .Y(new_n4863));
  XNOR2x2_ASAP7_75t_L       g04607(.A(new_n4863), .B(new_n4862), .Y(\f[39] ));
  MAJIxp5_ASAP7_75t_L       g04608(.A(new_n4863), .B(new_n4844), .C(new_n4861), .Y(new_n4865));
  A2O1A1Ixp33_ASAP7_75t_L   g04609(.A1(new_n4855), .A2(new_n4426), .B(new_n4425), .C(new_n4634), .Y(new_n4866));
  INVx1_ASAP7_75t_L         g04610(.A(new_n4849), .Y(new_n4867));
  NOR2xp33_ASAP7_75t_L      g04611(.A(\b[39] ), .B(\b[40] ), .Y(new_n4868));
  INVx1_ASAP7_75t_L         g04612(.A(\b[40] ), .Y(new_n4869));
  NOR2xp33_ASAP7_75t_L      g04613(.A(new_n4848), .B(new_n4869), .Y(new_n4870));
  NOR2xp33_ASAP7_75t_L      g04614(.A(new_n4868), .B(new_n4870), .Y(new_n4871));
  INVx1_ASAP7_75t_L         g04615(.A(new_n4871), .Y(new_n4872));
  A2O1A1O1Ixp25_ASAP7_75t_L g04616(.A1(new_n4846), .A2(new_n4866), .B(new_n4847), .C(new_n4867), .D(new_n4872), .Y(new_n4873));
  A2O1A1Ixp33_ASAP7_75t_L   g04617(.A1(new_n4866), .A2(new_n4846), .B(new_n4847), .C(new_n4867), .Y(new_n4874));
  NOR2xp33_ASAP7_75t_L      g04618(.A(new_n4871), .B(new_n4874), .Y(new_n4875));
  NOR2xp33_ASAP7_75t_L      g04619(.A(new_n4873), .B(new_n4875), .Y(new_n4876));
  NAND2xp33_ASAP7_75t_L     g04620(.A(new_n267), .B(new_n4876), .Y(new_n4877));
  AOI22xp33_ASAP7_75t_L     g04621(.A1(\b[38] ), .A2(new_n282), .B1(\b[40] ), .B2(new_n303), .Y(new_n4878));
  NAND2xp33_ASAP7_75t_L     g04622(.A(new_n4878), .B(new_n4877), .Y(new_n4879));
  AOI211xp5_ASAP7_75t_L     g04623(.A1(\b[39] ), .A2(new_n272), .B(new_n262), .C(new_n4879), .Y(new_n4880));
  INVx1_ASAP7_75t_L         g04624(.A(new_n4879), .Y(new_n4881));
  O2A1O1Ixp33_ASAP7_75t_L   g04625(.A1(new_n4848), .A2(new_n291), .B(new_n4881), .C(\a[2] ), .Y(new_n4882));
  NOR2xp33_ASAP7_75t_L      g04626(.A(new_n4880), .B(new_n4882), .Y(new_n4883));
  INVx1_ASAP7_75t_L         g04627(.A(new_n4651), .Y(new_n4884));
  NOR3xp33_ASAP7_75t_L      g04628(.A(new_n4834), .B(new_n4837), .C(new_n4654), .Y(new_n4885));
  NOR3xp33_ASAP7_75t_L      g04629(.A(new_n4830), .B(new_n4829), .C(new_n4827), .Y(new_n4886));
  AOI22xp33_ASAP7_75t_L     g04630(.A1(new_n444), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n471), .Y(new_n4887));
  OAI221xp5_ASAP7_75t_L     g04631(.A1(new_n468), .A2(new_n3565), .B1(new_n469), .B2(new_n3591), .C(new_n4887), .Y(new_n4888));
  XNOR2x2_ASAP7_75t_L       g04632(.A(new_n435), .B(new_n4888), .Y(new_n4889));
  OAI21xp33_ASAP7_75t_L     g04633(.A1(new_n4818), .A2(new_n4816), .B(new_n4812), .Y(new_n4890));
  NAND2xp33_ASAP7_75t_L     g04634(.A(new_n4792), .B(new_n4796), .Y(new_n4891));
  MAJIxp5_ASAP7_75t_L       g04635(.A(new_n4662), .B(new_n4891), .C(new_n4803), .Y(new_n4892));
  AOI22xp33_ASAP7_75t_L     g04636(.A1(new_n811), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n900), .Y(new_n4893));
  INVx1_ASAP7_75t_L         g04637(.A(new_n4893), .Y(new_n4894));
  AOI221xp5_ASAP7_75t_L     g04638(.A1(\b[27] ), .A2(new_n815), .B1(new_n808), .B2(new_n4237), .C(new_n4894), .Y(new_n4895));
  XNOR2x2_ASAP7_75t_L       g04639(.A(\a[14] ), .B(new_n4895), .Y(new_n4896));
  NAND2xp33_ASAP7_75t_L     g04640(.A(new_n4536), .B(new_n4537), .Y(new_n4897));
  A2O1A1O1Ixp25_ASAP7_75t_L g04641(.A1(new_n4478), .A2(new_n4897), .B(new_n4739), .C(new_n4729), .D(new_n4738), .Y(new_n4898));
  AOI22xp33_ASAP7_75t_L     g04642(.A1(new_n2552), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n2736), .Y(new_n4899));
  OAI221xp5_ASAP7_75t_L     g04643(.A1(new_n2547), .A2(new_n760), .B1(new_n2734), .B2(new_n790), .C(new_n4899), .Y(new_n4900));
  XNOR2x2_ASAP7_75t_L       g04644(.A(\a[29] ), .B(new_n4900), .Y(new_n4901));
  INVx1_ASAP7_75t_L         g04645(.A(new_n4901), .Y(new_n4902));
  NOR2xp33_ASAP7_75t_L      g04646(.A(new_n4701), .B(new_n4705), .Y(new_n4903));
  MAJIxp5_ASAP7_75t_L       g04647(.A(new_n4717), .B(new_n4903), .C(new_n4712), .Y(new_n4904));
  NOR3xp33_ASAP7_75t_L      g04648(.A(new_n4514), .B(new_n4677), .C(new_n4669), .Y(new_n4905));
  NAND2xp33_ASAP7_75t_L     g04649(.A(\b[3] ), .B(new_n4285), .Y(new_n4906));
  NAND2xp33_ASAP7_75t_L     g04650(.A(new_n4274), .B(new_n329), .Y(new_n4907));
  AOI22xp33_ASAP7_75t_L     g04651(.A1(new_n4283), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n4512), .Y(new_n4908));
  NAND4xp25_ASAP7_75t_L     g04652(.A(new_n4907), .B(\a[38] ), .C(new_n4906), .D(new_n4908), .Y(new_n4909));
  AOI31xp33_ASAP7_75t_L     g04653(.A1(new_n4907), .A2(new_n4906), .A3(new_n4908), .B(\a[38] ), .Y(new_n4910));
  INVx1_ASAP7_75t_L         g04654(.A(new_n4910), .Y(new_n4911));
  NAND2xp33_ASAP7_75t_L     g04655(.A(\a[41] ), .B(new_n4674), .Y(new_n4912));
  INVx1_ASAP7_75t_L         g04656(.A(\a[40] ), .Y(new_n4913));
  NAND2xp33_ASAP7_75t_L     g04657(.A(\a[41] ), .B(new_n4913), .Y(new_n4914));
  INVx1_ASAP7_75t_L         g04658(.A(\a[41] ), .Y(new_n4915));
  NAND2xp33_ASAP7_75t_L     g04659(.A(\a[40] ), .B(new_n4915), .Y(new_n4916));
  AOI21xp33_ASAP7_75t_L     g04660(.A1(new_n4916), .A2(new_n4914), .B(new_n4673), .Y(new_n4917));
  NAND2xp33_ASAP7_75t_L     g04661(.A(new_n269), .B(new_n4917), .Y(new_n4918));
  NAND2xp33_ASAP7_75t_L     g04662(.A(new_n4916), .B(new_n4914), .Y(new_n4919));
  NOR2xp33_ASAP7_75t_L      g04663(.A(new_n4919), .B(new_n4673), .Y(new_n4920));
  NAND2xp33_ASAP7_75t_L     g04664(.A(\b[1] ), .B(new_n4920), .Y(new_n4921));
  NAND2xp33_ASAP7_75t_L     g04665(.A(new_n4672), .B(new_n4671), .Y(new_n4922));
  XNOR2x2_ASAP7_75t_L       g04666(.A(\a[40] ), .B(\a[39] ), .Y(new_n4923));
  NOR2xp33_ASAP7_75t_L      g04667(.A(new_n4923), .B(new_n4922), .Y(new_n4924));
  NAND2xp33_ASAP7_75t_L     g04668(.A(\b[0] ), .B(new_n4924), .Y(new_n4925));
  NAND3xp33_ASAP7_75t_L     g04669(.A(new_n4918), .B(new_n4921), .C(new_n4925), .Y(new_n4926));
  XOR2x2_ASAP7_75t_L        g04670(.A(new_n4912), .B(new_n4926), .Y(new_n4927));
  NAND3xp33_ASAP7_75t_L     g04671(.A(new_n4911), .B(new_n4927), .C(new_n4909), .Y(new_n4928));
  INVx1_ASAP7_75t_L         g04672(.A(new_n4909), .Y(new_n4929));
  XNOR2x2_ASAP7_75t_L       g04673(.A(new_n4912), .B(new_n4926), .Y(new_n4930));
  OAI21xp33_ASAP7_75t_L     g04674(.A1(new_n4910), .A2(new_n4929), .B(new_n4930), .Y(new_n4931));
  OAI211xp5_ASAP7_75t_L     g04675(.A1(new_n4905), .A2(new_n4693), .B(new_n4928), .C(new_n4931), .Y(new_n4932));
  INVx1_ASAP7_75t_L         g04676(.A(new_n4905), .Y(new_n4933));
  NOR3xp33_ASAP7_75t_L      g04677(.A(new_n4930), .B(new_n4929), .C(new_n4910), .Y(new_n4934));
  AOI21xp33_ASAP7_75t_L     g04678(.A1(new_n4911), .A2(new_n4909), .B(new_n4927), .Y(new_n4935));
  OAI211xp5_ASAP7_75t_L     g04679(.A1(new_n4934), .A2(new_n4935), .B(new_n4933), .C(new_n4684), .Y(new_n4936));
  NOR2xp33_ASAP7_75t_L      g04680(.A(new_n418), .B(new_n3853), .Y(new_n4937));
  AOI22xp33_ASAP7_75t_L     g04681(.A1(new_n3633), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n3858), .Y(new_n4938));
  OAI21xp33_ASAP7_75t_L     g04682(.A1(new_n3856), .A2(new_n425), .B(new_n4938), .Y(new_n4939));
  OR3x1_ASAP7_75t_L         g04683(.A(new_n4939), .B(new_n3628), .C(new_n4937), .Y(new_n4940));
  A2O1A1Ixp33_ASAP7_75t_L   g04684(.A1(\b[6] ), .A2(new_n3639), .B(new_n4939), .C(new_n3628), .Y(new_n4941));
  NAND4xp25_ASAP7_75t_L     g04685(.A(new_n4936), .B(new_n4940), .C(new_n4941), .D(new_n4932), .Y(new_n4942));
  AOI211xp5_ASAP7_75t_L     g04686(.A1(new_n4684), .A2(new_n4933), .B(new_n4934), .C(new_n4935), .Y(new_n4943));
  AOI211xp5_ASAP7_75t_L     g04687(.A1(new_n4928), .A2(new_n4931), .B(new_n4905), .C(new_n4693), .Y(new_n4944));
  NAND2xp33_ASAP7_75t_L     g04688(.A(new_n4941), .B(new_n4940), .Y(new_n4945));
  OAI21xp33_ASAP7_75t_L     g04689(.A1(new_n4943), .A2(new_n4944), .B(new_n4945), .Y(new_n4946));
  AOI211xp5_ASAP7_75t_L     g04690(.A1(new_n4691), .A2(new_n4689), .B(new_n4693), .C(new_n4694), .Y(new_n4947));
  AOI21xp33_ASAP7_75t_L     g04691(.A1(new_n4700), .A2(new_n4697), .B(new_n4947), .Y(new_n4948));
  NAND3xp33_ASAP7_75t_L     g04692(.A(new_n4948), .B(new_n4946), .C(new_n4942), .Y(new_n4949));
  NAND2xp33_ASAP7_75t_L     g04693(.A(new_n4942), .B(new_n4946), .Y(new_n4950));
  A2O1A1Ixp33_ASAP7_75t_L   g04694(.A1(new_n4697), .A2(new_n4700), .B(new_n4947), .C(new_n4950), .Y(new_n4951));
  NOR2xp33_ASAP7_75t_L      g04695(.A(new_n540), .B(new_n3024), .Y(new_n4952));
  INVx1_ASAP7_75t_L         g04696(.A(new_n4952), .Y(new_n4953));
  NAND2xp33_ASAP7_75t_L     g04697(.A(new_n3021), .B(new_n2143), .Y(new_n4954));
  AOI22xp33_ASAP7_75t_L     g04698(.A1(new_n3029), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n3258), .Y(new_n4955));
  AND4x1_ASAP7_75t_L        g04699(.A(new_n4955), .B(new_n4954), .C(new_n4953), .D(\a[32] ), .Y(new_n4956));
  AOI31xp33_ASAP7_75t_L     g04700(.A1(new_n4954), .A2(new_n4953), .A3(new_n4955), .B(\a[32] ), .Y(new_n4957));
  OR2x4_ASAP7_75t_L         g04701(.A(new_n4957), .B(new_n4956), .Y(new_n4958));
  AOI21xp33_ASAP7_75t_L     g04702(.A1(new_n4951), .A2(new_n4949), .B(new_n4958), .Y(new_n4959));
  INVx1_ASAP7_75t_L         g04703(.A(new_n4947), .Y(new_n4960));
  A2O1A1Ixp33_ASAP7_75t_L   g04704(.A1(new_n4696), .A2(new_n4692), .B(new_n4704), .C(new_n4960), .Y(new_n4961));
  NOR2xp33_ASAP7_75t_L      g04705(.A(new_n4950), .B(new_n4961), .Y(new_n4962));
  AOI21xp33_ASAP7_75t_L     g04706(.A1(new_n4946), .A2(new_n4942), .B(new_n4948), .Y(new_n4963));
  NOR2xp33_ASAP7_75t_L      g04707(.A(new_n4957), .B(new_n4956), .Y(new_n4964));
  NOR3xp33_ASAP7_75t_L      g04708(.A(new_n4962), .B(new_n4964), .C(new_n4963), .Y(new_n4965));
  OAI21xp33_ASAP7_75t_L     g04709(.A1(new_n4959), .A2(new_n4965), .B(new_n4904), .Y(new_n4966));
  AOI211xp5_ASAP7_75t_L     g04710(.A1(new_n4711), .A2(new_n4709), .B(new_n4701), .C(new_n4705), .Y(new_n4967));
  INVx1_ASAP7_75t_L         g04711(.A(new_n4967), .Y(new_n4968));
  A2O1A1Ixp33_ASAP7_75t_L   g04712(.A1(new_n4720), .A2(new_n4719), .B(new_n4721), .C(new_n4968), .Y(new_n4969));
  OAI21xp33_ASAP7_75t_L     g04713(.A1(new_n4963), .A2(new_n4962), .B(new_n4964), .Y(new_n4970));
  NAND3xp33_ASAP7_75t_L     g04714(.A(new_n4958), .B(new_n4951), .C(new_n4949), .Y(new_n4971));
  NAND3xp33_ASAP7_75t_L     g04715(.A(new_n4969), .B(new_n4970), .C(new_n4971), .Y(new_n4972));
  AOI21xp33_ASAP7_75t_L     g04716(.A1(new_n4972), .A2(new_n4966), .B(new_n4902), .Y(new_n4973));
  NAND2xp33_ASAP7_75t_L     g04717(.A(new_n4719), .B(new_n4720), .Y(new_n4974));
  AOI221xp5_ASAP7_75t_L     g04718(.A1(new_n4974), .A2(new_n4717), .B1(new_n4970), .B2(new_n4971), .C(new_n4967), .Y(new_n4975));
  NOR3xp33_ASAP7_75t_L      g04719(.A(new_n4904), .B(new_n4959), .C(new_n4965), .Y(new_n4976));
  NOR3xp33_ASAP7_75t_L      g04720(.A(new_n4976), .B(new_n4975), .C(new_n4901), .Y(new_n4977));
  NOR3xp33_ASAP7_75t_L      g04721(.A(new_n4898), .B(new_n4973), .C(new_n4977), .Y(new_n4978));
  OAI21xp33_ASAP7_75t_L     g04722(.A1(new_n4975), .A2(new_n4976), .B(new_n4901), .Y(new_n4979));
  NAND3xp33_ASAP7_75t_L     g04723(.A(new_n4972), .B(new_n4902), .C(new_n4966), .Y(new_n4980));
  AOI221xp5_ASAP7_75t_L     g04724(.A1(new_n4729), .A2(new_n4735), .B1(new_n4979), .B2(new_n4980), .C(new_n4738), .Y(new_n4981));
  AOI22xp33_ASAP7_75t_L     g04725(.A1(new_n2114), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n2259), .Y(new_n4982));
  OAI221xp5_ASAP7_75t_L     g04726(.A1(new_n2109), .A2(new_n942), .B1(new_n2257), .B2(new_n1035), .C(new_n4982), .Y(new_n4983));
  XNOR2x2_ASAP7_75t_L       g04727(.A(new_n2100), .B(new_n4983), .Y(new_n4984));
  NOR3xp33_ASAP7_75t_L      g04728(.A(new_n4981), .B(new_n4978), .C(new_n4984), .Y(new_n4985));
  INVx1_ASAP7_75t_L         g04729(.A(new_n4739), .Y(new_n4986));
  A2O1A1Ixp33_ASAP7_75t_L   g04730(.A1(new_n4533), .A2(new_n4986), .B(new_n4737), .C(new_n4733), .Y(new_n4987));
  NAND3xp33_ASAP7_75t_L     g04731(.A(new_n4987), .B(new_n4979), .C(new_n4980), .Y(new_n4988));
  OAI21xp33_ASAP7_75t_L     g04732(.A1(new_n4973), .A2(new_n4977), .B(new_n4898), .Y(new_n4989));
  XNOR2x2_ASAP7_75t_L       g04733(.A(\a[26] ), .B(new_n4983), .Y(new_n4990));
  AOI21xp33_ASAP7_75t_L     g04734(.A1(new_n4988), .A2(new_n4989), .B(new_n4990), .Y(new_n4991));
  NOR2xp33_ASAP7_75t_L      g04735(.A(new_n4985), .B(new_n4991), .Y(new_n4992));
  NOR3xp33_ASAP7_75t_L      g04736(.A(new_n4746), .B(new_n4747), .C(new_n4744), .Y(new_n4993));
  O2A1O1Ixp33_ASAP7_75t_L   g04737(.A1(new_n4752), .A2(new_n4553), .B(new_n4750), .C(new_n4993), .Y(new_n4994));
  NAND2xp33_ASAP7_75t_L     g04738(.A(new_n4992), .B(new_n4994), .Y(new_n4995));
  NAND3xp33_ASAP7_75t_L     g04739(.A(new_n4988), .B(new_n4989), .C(new_n4990), .Y(new_n4996));
  OAI21xp33_ASAP7_75t_L     g04740(.A1(new_n4978), .A2(new_n4981), .B(new_n4984), .Y(new_n4997));
  NAND2xp33_ASAP7_75t_L     g04741(.A(new_n4997), .B(new_n4996), .Y(new_n4998));
  A2O1A1Ixp33_ASAP7_75t_L   g04742(.A1(new_n4668), .A2(new_n4750), .B(new_n4993), .C(new_n4998), .Y(new_n4999));
  AOI22xp33_ASAP7_75t_L     g04743(.A1(new_n1704), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1837), .Y(new_n5000));
  OAI221xp5_ASAP7_75t_L     g04744(.A1(new_n1699), .A2(new_n1313), .B1(new_n1827), .B2(new_n1438), .C(new_n5000), .Y(new_n5001));
  XNOR2x2_ASAP7_75t_L       g04745(.A(\a[23] ), .B(new_n5001), .Y(new_n5002));
  NAND3xp33_ASAP7_75t_L     g04746(.A(new_n4995), .B(new_n4999), .C(new_n5002), .Y(new_n5003));
  NAND3xp33_ASAP7_75t_L     g04747(.A(new_n4741), .B(new_n4736), .C(new_n4748), .Y(new_n5004));
  A2O1A1Ixp33_ASAP7_75t_L   g04748(.A1(new_n4745), .A2(new_n4749), .B(new_n4753), .C(new_n5004), .Y(new_n5005));
  NOR2xp33_ASAP7_75t_L      g04749(.A(new_n5005), .B(new_n4998), .Y(new_n5006));
  A2O1A1O1Ixp25_ASAP7_75t_L g04750(.A1(new_n4745), .A2(new_n4749), .B(new_n4753), .C(new_n5004), .D(new_n4992), .Y(new_n5007));
  INVx1_ASAP7_75t_L         g04751(.A(new_n5002), .Y(new_n5008));
  OAI21xp33_ASAP7_75t_L     g04752(.A1(new_n5006), .A2(new_n5007), .B(new_n5008), .Y(new_n5009));
  NOR3xp33_ASAP7_75t_L      g04753(.A(new_n4758), .B(new_n4757), .C(new_n4756), .Y(new_n5010));
  A2O1A1O1Ixp25_ASAP7_75t_L g04754(.A1(new_n4557), .A2(new_n4559), .B(new_n4663), .C(new_n4759), .D(new_n5010), .Y(new_n5011));
  AND3x1_ASAP7_75t_L        g04755(.A(new_n5011), .B(new_n5009), .C(new_n5003), .Y(new_n5012));
  AOI21xp33_ASAP7_75t_L     g04756(.A1(new_n5003), .A2(new_n5009), .B(new_n5011), .Y(new_n5013));
  NOR2xp33_ASAP7_75t_L      g04757(.A(new_n1655), .B(new_n1373), .Y(new_n5014));
  AOI22xp33_ASAP7_75t_L     g04758(.A1(new_n1360), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1581), .Y(new_n5015));
  OAI21xp33_ASAP7_75t_L     g04759(.A1(new_n1359), .A2(new_n1780), .B(new_n5015), .Y(new_n5016));
  OR3x1_ASAP7_75t_L         g04760(.A(new_n5016), .B(new_n1356), .C(new_n5014), .Y(new_n5017));
  A2O1A1Ixp33_ASAP7_75t_L   g04761(.A1(\b[21] ), .A2(new_n1362), .B(new_n5016), .C(new_n1356), .Y(new_n5018));
  NAND2xp33_ASAP7_75t_L     g04762(.A(new_n5018), .B(new_n5017), .Y(new_n5019));
  NOR3xp33_ASAP7_75t_L      g04763(.A(new_n5012), .B(new_n5013), .C(new_n5019), .Y(new_n5020));
  NAND3xp33_ASAP7_75t_L     g04764(.A(new_n5011), .B(new_n5003), .C(new_n5009), .Y(new_n5021));
  AO21x2_ASAP7_75t_L        g04765(.A1(new_n5003), .A2(new_n5009), .B(new_n5011), .Y(new_n5022));
  AND2x2_ASAP7_75t_L        g04766(.A(new_n5018), .B(new_n5017), .Y(new_n5023));
  AOI21xp33_ASAP7_75t_L     g04767(.A1(new_n5022), .A2(new_n5021), .B(new_n5023), .Y(new_n5024));
  NOR2xp33_ASAP7_75t_L      g04768(.A(new_n5024), .B(new_n5020), .Y(new_n5025));
  NAND3xp33_ASAP7_75t_L     g04769(.A(new_n4763), .B(new_n4760), .C(new_n4771), .Y(new_n5026));
  NAND3xp33_ASAP7_75t_L     g04770(.A(new_n5025), .B(new_n4783), .C(new_n5026), .Y(new_n5027));
  NAND3xp33_ASAP7_75t_L     g04771(.A(new_n5022), .B(new_n5023), .C(new_n5021), .Y(new_n5028));
  OAI21xp33_ASAP7_75t_L     g04772(.A1(new_n5013), .A2(new_n5012), .B(new_n5019), .Y(new_n5029));
  NAND2xp33_ASAP7_75t_L     g04773(.A(new_n5028), .B(new_n5029), .Y(new_n5030));
  A2O1A1Ixp33_ASAP7_75t_L   g04774(.A1(new_n4772), .A2(new_n4767), .B(new_n4776), .C(new_n5026), .Y(new_n5031));
  NAND2xp33_ASAP7_75t_L     g04775(.A(new_n5030), .B(new_n5031), .Y(new_n5032));
  OAI22xp33_ASAP7_75t_L     g04776(.A1(new_n1158), .A2(new_n1909), .B1(new_n2067), .B2(new_n1259), .Y(new_n5033));
  AOI221xp5_ASAP7_75t_L     g04777(.A1(\b[24] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n2648), .C(new_n5033), .Y(new_n5034));
  XNOR2x2_ASAP7_75t_L       g04778(.A(new_n1071), .B(new_n5034), .Y(new_n5035));
  NAND3xp33_ASAP7_75t_L     g04779(.A(new_n5027), .B(new_n5035), .C(new_n5032), .Y(new_n5036));
  NOR2xp33_ASAP7_75t_L      g04780(.A(new_n5030), .B(new_n5031), .Y(new_n5037));
  AOI21xp33_ASAP7_75t_L     g04781(.A1(new_n4783), .A2(new_n5026), .B(new_n5025), .Y(new_n5038));
  XNOR2x2_ASAP7_75t_L       g04782(.A(\a[17] ), .B(new_n5034), .Y(new_n5039));
  OAI21xp33_ASAP7_75t_L     g04783(.A1(new_n5037), .A2(new_n5038), .B(new_n5039), .Y(new_n5040));
  AOI31xp33_ASAP7_75t_L     g04784(.A1(new_n4791), .A2(new_n4781), .A3(new_n4583), .B(new_n4794), .Y(new_n5041));
  AOI21xp33_ASAP7_75t_L     g04785(.A1(new_n5040), .A2(new_n5036), .B(new_n5041), .Y(new_n5042));
  AND3x1_ASAP7_75t_L        g04786(.A(new_n5041), .B(new_n5040), .C(new_n5036), .Y(new_n5043));
  OAI21xp33_ASAP7_75t_L     g04787(.A1(new_n5042), .A2(new_n5043), .B(new_n4896), .Y(new_n5044));
  XNOR2x2_ASAP7_75t_L       g04788(.A(new_n806), .B(new_n4895), .Y(new_n5045));
  AO21x2_ASAP7_75t_L        g04789(.A1(new_n5036), .A2(new_n5040), .B(new_n5041), .Y(new_n5046));
  NAND3xp33_ASAP7_75t_L     g04790(.A(new_n5041), .B(new_n5040), .C(new_n5036), .Y(new_n5047));
  NAND3xp33_ASAP7_75t_L     g04791(.A(new_n5046), .B(new_n5045), .C(new_n5047), .Y(new_n5048));
  NAND3xp33_ASAP7_75t_L     g04792(.A(new_n4892), .B(new_n5044), .C(new_n5048), .Y(new_n5049));
  AO31x2_ASAP7_75t_L        g04793(.A1(new_n4603), .A2(new_n4595), .A3(new_n4382), .B(new_n4661), .Y(new_n5050));
  NAND2xp33_ASAP7_75t_L     g04794(.A(new_n4804), .B(new_n4808), .Y(new_n5051));
  NOR2xp33_ASAP7_75t_L      g04795(.A(new_n4803), .B(new_n4891), .Y(new_n5052));
  AO221x2_ASAP7_75t_L       g04796(.A1(new_n5051), .A2(new_n5050), .B1(new_n5044), .B2(new_n5048), .C(new_n5052), .Y(new_n5053));
  AOI22xp33_ASAP7_75t_L     g04797(.A1(\b[29] ), .A2(new_n651), .B1(\b[31] ), .B2(new_n581), .Y(new_n5054));
  OAI221xp5_ASAP7_75t_L     g04798(.A1(new_n821), .A2(new_n2982), .B1(new_n577), .B2(new_n3187), .C(new_n5054), .Y(new_n5055));
  XNOR2x2_ASAP7_75t_L       g04799(.A(\a[11] ), .B(new_n5055), .Y(new_n5056));
  NAND3xp33_ASAP7_75t_L     g04800(.A(new_n5053), .B(new_n5049), .C(new_n5056), .Y(new_n5057));
  NOR2xp33_ASAP7_75t_L      g04801(.A(new_n4806), .B(new_n4805), .Y(new_n5058));
  MAJIxp5_ASAP7_75t_L       g04802(.A(new_n5050), .B(new_n5058), .C(new_n4807), .Y(new_n5059));
  NAND2xp33_ASAP7_75t_L     g04803(.A(new_n5048), .B(new_n5044), .Y(new_n5060));
  NOR2xp33_ASAP7_75t_L      g04804(.A(new_n5059), .B(new_n5060), .Y(new_n5061));
  AOI21xp33_ASAP7_75t_L     g04805(.A1(new_n5048), .A2(new_n5044), .B(new_n4892), .Y(new_n5062));
  INVx1_ASAP7_75t_L         g04806(.A(new_n5056), .Y(new_n5063));
  OAI21xp33_ASAP7_75t_L     g04807(.A1(new_n5062), .A2(new_n5061), .B(new_n5063), .Y(new_n5064));
  NAND3xp33_ASAP7_75t_L     g04808(.A(new_n4890), .B(new_n5057), .C(new_n5064), .Y(new_n5065));
  NOR3xp33_ASAP7_75t_L      g04809(.A(new_n5061), .B(new_n5063), .C(new_n5062), .Y(new_n5066));
  AOI21xp33_ASAP7_75t_L     g04810(.A1(new_n5053), .A2(new_n5049), .B(new_n5056), .Y(new_n5067));
  OAI221xp5_ASAP7_75t_L     g04811(.A1(new_n4818), .A2(new_n4816), .B1(new_n5067), .B2(new_n5066), .C(new_n4812), .Y(new_n5068));
  AOI21xp33_ASAP7_75t_L     g04812(.A1(new_n5065), .A2(new_n5068), .B(new_n4889), .Y(new_n5069));
  AND3x1_ASAP7_75t_L        g04813(.A(new_n5065), .B(new_n5068), .C(new_n4889), .Y(new_n5070));
  NOR2xp33_ASAP7_75t_L      g04814(.A(new_n5069), .B(new_n5070), .Y(new_n5071));
  A2O1A1Ixp33_ASAP7_75t_L   g04815(.A1(new_n4836), .A2(new_n4835), .B(new_n4886), .C(new_n5071), .Y(new_n5072));
  AOI21xp33_ASAP7_75t_L     g04816(.A1(new_n4835), .A2(new_n4836), .B(new_n4886), .Y(new_n5073));
  AO21x2_ASAP7_75t_L        g04817(.A1(new_n5068), .A2(new_n5065), .B(new_n4889), .Y(new_n5074));
  NAND3xp33_ASAP7_75t_L     g04818(.A(new_n5065), .B(new_n5068), .C(new_n4889), .Y(new_n5075));
  NAND2xp33_ASAP7_75t_L     g04819(.A(new_n5075), .B(new_n5074), .Y(new_n5076));
  NAND2xp33_ASAP7_75t_L     g04820(.A(new_n5076), .B(new_n5073), .Y(new_n5077));
  AOI22xp33_ASAP7_75t_L     g04821(.A1(new_n344), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n370), .Y(new_n5078));
  OAI221xp5_ASAP7_75t_L     g04822(.A1(new_n429), .A2(new_n4216), .B1(new_n366), .B2(new_n4431), .C(new_n5078), .Y(new_n5079));
  XNOR2x2_ASAP7_75t_L       g04823(.A(\a[5] ), .B(new_n5079), .Y(new_n5080));
  NAND3xp33_ASAP7_75t_L     g04824(.A(new_n5072), .B(new_n5077), .C(new_n5080), .Y(new_n5081));
  NOR2xp33_ASAP7_75t_L      g04825(.A(new_n5076), .B(new_n5073), .Y(new_n5082));
  AOI221xp5_ASAP7_75t_L     g04826(.A1(new_n4835), .A2(new_n4836), .B1(new_n5074), .B2(new_n5075), .C(new_n4886), .Y(new_n5083));
  INVx1_ASAP7_75t_L         g04827(.A(new_n5080), .Y(new_n5084));
  OAI21xp33_ASAP7_75t_L     g04828(.A1(new_n5083), .A2(new_n5082), .B(new_n5084), .Y(new_n5085));
  NAND2xp33_ASAP7_75t_L     g04829(.A(new_n5081), .B(new_n5085), .Y(new_n5086));
  A2O1A1Ixp33_ASAP7_75t_L   g04830(.A1(new_n4884), .A2(new_n4838), .B(new_n4885), .C(new_n5086), .Y(new_n5087));
  A2O1A1O1Ixp25_ASAP7_75t_L g04831(.A1(new_n4624), .A2(new_n4444), .B(new_n4650), .C(new_n4838), .D(new_n4885), .Y(new_n5088));
  NAND3xp33_ASAP7_75t_L     g04832(.A(new_n5088), .B(new_n5081), .C(new_n5085), .Y(new_n5089));
  NAND2xp33_ASAP7_75t_L     g04833(.A(new_n5089), .B(new_n5087), .Y(new_n5090));
  NOR2xp33_ASAP7_75t_L      g04834(.A(new_n4883), .B(new_n5090), .Y(new_n5091));
  INVx1_ASAP7_75t_L         g04835(.A(new_n5091), .Y(new_n5092));
  NAND2xp33_ASAP7_75t_L     g04836(.A(new_n4883), .B(new_n5090), .Y(new_n5093));
  NAND2xp33_ASAP7_75t_L     g04837(.A(new_n5093), .B(new_n5092), .Y(new_n5094));
  XNOR2x2_ASAP7_75t_L       g04838(.A(new_n4865), .B(new_n5094), .Y(\f[40] ));
  AOI21xp33_ASAP7_75t_L     g04839(.A1(new_n4865), .A2(new_n5093), .B(new_n5091), .Y(new_n5096));
  NAND3xp33_ASAP7_75t_L     g04840(.A(new_n5072), .B(new_n5077), .C(new_n5084), .Y(new_n5097));
  A2O1A1Ixp33_ASAP7_75t_L   g04841(.A1(new_n5081), .A2(new_n5085), .B(new_n5088), .C(new_n5097), .Y(new_n5098));
  OAI22xp33_ASAP7_75t_L     g04842(.A1(new_n407), .A2(new_n4216), .B1(new_n4632), .B2(new_n343), .Y(new_n5099));
  AOI221xp5_ASAP7_75t_L     g04843(.A1(\b[37] ), .A2(new_n347), .B1(new_n341), .B2(new_n4640), .C(new_n5099), .Y(new_n5100));
  XNOR2x2_ASAP7_75t_L       g04844(.A(new_n338), .B(new_n5100), .Y(new_n5101));
  INVx1_ASAP7_75t_L         g04845(.A(new_n5101), .Y(new_n5102));
  INVx1_ASAP7_75t_L         g04846(.A(new_n5073), .Y(new_n5103));
  A2O1A1O1Ixp25_ASAP7_75t_L g04847(.A1(new_n4814), .A2(new_n4656), .B(new_n4817), .C(new_n5057), .D(new_n5067), .Y(new_n5104));
  NOR2xp33_ASAP7_75t_L      g04848(.A(new_n3180), .B(new_n821), .Y(new_n5105));
  INVx1_ASAP7_75t_L         g04849(.A(new_n5105), .Y(new_n5106));
  NAND3xp33_ASAP7_75t_L     g04850(.A(new_n3210), .B(new_n578), .C(new_n3213), .Y(new_n5107));
  AOI22xp33_ASAP7_75t_L     g04851(.A1(\b[30] ), .A2(new_n651), .B1(\b[32] ), .B2(new_n581), .Y(new_n5108));
  AND4x1_ASAP7_75t_L        g04852(.A(new_n5108), .B(new_n5107), .C(new_n5106), .D(\a[11] ), .Y(new_n5109));
  AOI31xp33_ASAP7_75t_L     g04853(.A1(new_n5107), .A2(new_n5106), .A3(new_n5108), .B(\a[11] ), .Y(new_n5110));
  NOR2xp33_ASAP7_75t_L      g04854(.A(new_n5110), .B(new_n5109), .Y(new_n5111));
  INVx1_ASAP7_75t_L         g04855(.A(new_n5111), .Y(new_n5112));
  NOR3xp33_ASAP7_75t_L      g04856(.A(new_n5043), .B(new_n5042), .C(new_n5045), .Y(new_n5113));
  INVx1_ASAP7_75t_L         g04857(.A(new_n5113), .Y(new_n5114));
  A2O1A1Ixp33_ASAP7_75t_L   g04858(.A1(new_n5044), .A2(new_n5048), .B(new_n5059), .C(new_n5114), .Y(new_n5115));
  AOI22xp33_ASAP7_75t_L     g04859(.A1(new_n811), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n900), .Y(new_n5116));
  OAI221xp5_ASAP7_75t_L     g04860(.A1(new_n904), .A2(new_n2666), .B1(new_n898), .B2(new_n2695), .C(new_n5116), .Y(new_n5117));
  XNOR2x2_ASAP7_75t_L       g04861(.A(\a[14] ), .B(new_n5117), .Y(new_n5118));
  NOR2xp33_ASAP7_75t_L      g04862(.A(new_n5037), .B(new_n5038), .Y(new_n5119));
  OAI31xp33_ASAP7_75t_L     g04863(.A1(new_n4795), .A2(new_n4793), .A3(new_n4598), .B(new_n4785), .Y(new_n5120));
  MAJIxp5_ASAP7_75t_L       g04864(.A(new_n5120), .B(new_n5119), .C(new_n5039), .Y(new_n5121));
  AOI22xp33_ASAP7_75t_L     g04865(.A1(new_n1076), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1253), .Y(new_n5122));
  OAI221xp5_ASAP7_75t_L     g04866(.A1(new_n1154), .A2(new_n2067), .B1(new_n1156), .B2(new_n2355), .C(new_n5122), .Y(new_n5123));
  XNOR2x2_ASAP7_75t_L       g04867(.A(\a[17] ), .B(new_n5123), .Y(new_n5124));
  INVx1_ASAP7_75t_L         g04868(.A(new_n5124), .Y(new_n5125));
  NAND3xp33_ASAP7_75t_L     g04869(.A(new_n5022), .B(new_n5021), .C(new_n5019), .Y(new_n5126));
  INVx1_ASAP7_75t_L         g04870(.A(new_n5126), .Y(new_n5127));
  O2A1O1Ixp33_ASAP7_75t_L   g04871(.A1(new_n5020), .A2(new_n5024), .B(new_n5031), .C(new_n5127), .Y(new_n5128));
  NOR3xp33_ASAP7_75t_L      g04872(.A(new_n4981), .B(new_n4978), .C(new_n4990), .Y(new_n5129));
  NAND2xp33_ASAP7_75t_L     g04873(.A(\b[16] ), .B(new_n2115), .Y(new_n5130));
  NAND3xp33_ASAP7_75t_L     g04874(.A(new_n1206), .B(new_n1208), .C(new_n2106), .Y(new_n5131));
  AOI22xp33_ASAP7_75t_L     g04875(.A1(new_n2114), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n2259), .Y(new_n5132));
  NAND4xp25_ASAP7_75t_L     g04876(.A(new_n5131), .B(\a[26] ), .C(new_n5130), .D(new_n5132), .Y(new_n5133));
  OAI31xp33_ASAP7_75t_L     g04877(.A1(new_n1796), .A2(new_n1205), .A3(new_n2257), .B(new_n5132), .Y(new_n5134));
  A2O1A1Ixp33_ASAP7_75t_L   g04878(.A1(\b[16] ), .A2(new_n2115), .B(new_n5134), .C(new_n2100), .Y(new_n5135));
  NAND2xp33_ASAP7_75t_L     g04879(.A(new_n5133), .B(new_n5135), .Y(new_n5136));
  OAI21xp33_ASAP7_75t_L     g04880(.A1(new_n4973), .A2(new_n4898), .B(new_n4980), .Y(new_n5137));
  AOI22xp33_ASAP7_75t_L     g04881(.A1(new_n2552), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n2736), .Y(new_n5138));
  OAI221xp5_ASAP7_75t_L     g04882(.A1(new_n2547), .A2(new_n784), .B1(new_n2734), .B2(new_n875), .C(new_n5138), .Y(new_n5139));
  XNOR2x2_ASAP7_75t_L       g04883(.A(new_n2538), .B(new_n5139), .Y(new_n5140));
  NOR2xp33_ASAP7_75t_L      g04884(.A(new_n4944), .B(new_n4943), .Y(new_n5141));
  AOI22xp33_ASAP7_75t_L     g04885(.A1(new_n3633), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n3858), .Y(new_n5142));
  OAI221xp5_ASAP7_75t_L     g04886(.A1(new_n3853), .A2(new_n420), .B1(new_n3856), .B2(new_n494), .C(new_n5142), .Y(new_n5143));
  NOR2xp33_ASAP7_75t_L      g04887(.A(new_n3628), .B(new_n5143), .Y(new_n5144));
  AND2x2_ASAP7_75t_L        g04888(.A(new_n3628), .B(new_n5143), .Y(new_n5145));
  O2A1O1Ixp33_ASAP7_75t_L   g04889(.A1(new_n4905), .A2(new_n4693), .B(new_n4928), .C(new_n4935), .Y(new_n5146));
  NOR2xp33_ASAP7_75t_L      g04890(.A(new_n324), .B(new_n4277), .Y(new_n5147));
  NOR3xp33_ASAP7_75t_L      g04891(.A(new_n357), .B(new_n358), .C(new_n4499), .Y(new_n5148));
  OAI22xp33_ASAP7_75t_L     g04892(.A1(new_n4501), .A2(new_n298), .B1(new_n354), .B2(new_n4275), .Y(new_n5149));
  NOR4xp25_ASAP7_75t_L      g04893(.A(new_n5148), .B(new_n4268), .C(new_n5149), .D(new_n5147), .Y(new_n5150));
  INVx1_ASAP7_75t_L         g04894(.A(new_n5150), .Y(new_n5151));
  OAI31xp33_ASAP7_75t_L     g04895(.A1(new_n5148), .A2(new_n5147), .A3(new_n5149), .B(new_n4268), .Y(new_n5152));
  NAND3xp33_ASAP7_75t_L     g04896(.A(new_n4922), .B(new_n4914), .C(new_n4916), .Y(new_n5153));
  OR2x4_ASAP7_75t_L         g04897(.A(new_n4923), .B(new_n4922), .Y(new_n5154));
  OAI22xp33_ASAP7_75t_L     g04898(.A1(new_n5154), .A2(new_n258), .B1(new_n261), .B2(new_n5153), .Y(new_n5155));
  AOI21xp33_ASAP7_75t_L     g04899(.A1(new_n4917), .A2(new_n269), .B(new_n5155), .Y(new_n5156));
  NOR2xp33_ASAP7_75t_L      g04900(.A(new_n261), .B(new_n5154), .Y(new_n5157));
  NAND2xp33_ASAP7_75t_L     g04901(.A(new_n4919), .B(new_n4922), .Y(new_n5158));
  NAND2xp33_ASAP7_75t_L     g04902(.A(\b[2] ), .B(new_n4920), .Y(new_n5159));
  NAND3xp33_ASAP7_75t_L     g04903(.A(new_n4673), .B(new_n4919), .C(new_n4923), .Y(new_n5160));
  OAI221xp5_ASAP7_75t_L     g04904(.A1(new_n258), .A2(new_n5160), .B1(new_n280), .B2(new_n5158), .C(new_n5159), .Y(new_n5161));
  NOR2xp33_ASAP7_75t_L      g04905(.A(new_n5157), .B(new_n5161), .Y(new_n5162));
  A2O1A1Ixp33_ASAP7_75t_L   g04906(.A1(new_n4677), .A2(new_n5156), .B(new_n4915), .C(new_n5162), .Y(new_n5163));
  O2A1O1Ixp33_ASAP7_75t_L   g04907(.A1(new_n258), .A2(new_n4673), .B(new_n5156), .C(new_n4915), .Y(new_n5164));
  INVx1_ASAP7_75t_L         g04908(.A(new_n5157), .Y(new_n5165));
  NOR2xp33_ASAP7_75t_L      g04909(.A(new_n280), .B(new_n5158), .Y(new_n5166));
  AND3x1_ASAP7_75t_L        g04910(.A(new_n4673), .B(new_n4923), .C(new_n4919), .Y(new_n5167));
  AOI221xp5_ASAP7_75t_L     g04911(.A1(new_n4920), .A2(\b[2] ), .B1(new_n5167), .B2(\b[0] ), .C(new_n5166), .Y(new_n5168));
  NAND2xp33_ASAP7_75t_L     g04912(.A(new_n5165), .B(new_n5168), .Y(new_n5169));
  NAND2xp33_ASAP7_75t_L     g04913(.A(new_n5169), .B(new_n5164), .Y(new_n5170));
  NAND4xp25_ASAP7_75t_L     g04914(.A(new_n5170), .B(new_n5151), .C(new_n5152), .D(new_n5163), .Y(new_n5171));
  INVx1_ASAP7_75t_L         g04915(.A(new_n5152), .Y(new_n5172));
  O2A1O1Ixp33_ASAP7_75t_L   g04916(.A1(new_n4674), .A2(new_n4926), .B(\a[41] ), .C(new_n5169), .Y(new_n5173));
  A2O1A1Ixp33_ASAP7_75t_L   g04917(.A1(\b[0] ), .A2(new_n4922), .B(new_n4926), .C(\a[41] ), .Y(new_n5174));
  O2A1O1Ixp33_ASAP7_75t_L   g04918(.A1(new_n5154), .A2(new_n261), .B(new_n5168), .C(new_n5174), .Y(new_n5175));
  OAI22xp33_ASAP7_75t_L     g04919(.A1(new_n5175), .A2(new_n5173), .B1(new_n5172), .B2(new_n5150), .Y(new_n5176));
  AOI21xp33_ASAP7_75t_L     g04920(.A1(new_n5176), .A2(new_n5171), .B(new_n5146), .Y(new_n5177));
  A2O1A1Ixp33_ASAP7_75t_L   g04921(.A1(new_n4684), .A2(new_n4933), .B(new_n4934), .C(new_n4931), .Y(new_n5178));
  NAND2xp33_ASAP7_75t_L     g04922(.A(new_n5176), .B(new_n5171), .Y(new_n5179));
  NOR2xp33_ASAP7_75t_L      g04923(.A(new_n5178), .B(new_n5179), .Y(new_n5180));
  OAI22xp33_ASAP7_75t_L     g04924(.A1(new_n5180), .A2(new_n5177), .B1(new_n5145), .B2(new_n5144), .Y(new_n5181));
  XNOR2x2_ASAP7_75t_L       g04925(.A(\a[35] ), .B(new_n5143), .Y(new_n5182));
  NAND2xp33_ASAP7_75t_L     g04926(.A(new_n5178), .B(new_n5179), .Y(new_n5183));
  NAND3xp33_ASAP7_75t_L     g04927(.A(new_n5146), .B(new_n5171), .C(new_n5176), .Y(new_n5184));
  NAND3xp33_ASAP7_75t_L     g04928(.A(new_n5183), .B(new_n5182), .C(new_n5184), .Y(new_n5185));
  AND2x2_ASAP7_75t_L        g04929(.A(new_n5185), .B(new_n5181), .Y(new_n5186));
  A2O1A1Ixp33_ASAP7_75t_L   g04930(.A1(new_n4945), .A2(new_n5141), .B(new_n4963), .C(new_n5186), .Y(new_n5187));
  NAND2xp33_ASAP7_75t_L     g04931(.A(new_n4945), .B(new_n5141), .Y(new_n5188));
  NAND2xp33_ASAP7_75t_L     g04932(.A(new_n5185), .B(new_n5181), .Y(new_n5189));
  NAND3xp33_ASAP7_75t_L     g04933(.A(new_n4951), .B(new_n5188), .C(new_n5189), .Y(new_n5190));
  AOI22xp33_ASAP7_75t_L     g04934(.A1(new_n3029), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n3258), .Y(new_n5191));
  OAI221xp5_ASAP7_75t_L     g04935(.A1(new_n3024), .A2(new_n617), .B1(new_n3256), .B2(new_n685), .C(new_n5191), .Y(new_n5192));
  XNOR2x2_ASAP7_75t_L       g04936(.A(\a[32] ), .B(new_n5192), .Y(new_n5193));
  NAND3xp33_ASAP7_75t_L     g04937(.A(new_n5187), .B(new_n5190), .C(new_n5193), .Y(new_n5194));
  A2O1A1O1Ixp25_ASAP7_75t_L g04938(.A1(new_n4946), .A2(new_n4942), .B(new_n4948), .C(new_n5188), .D(new_n5189), .Y(new_n5195));
  A2O1A1Ixp33_ASAP7_75t_L   g04939(.A1(new_n4946), .A2(new_n4942), .B(new_n4948), .C(new_n5188), .Y(new_n5196));
  NOR2xp33_ASAP7_75t_L      g04940(.A(new_n5196), .B(new_n5186), .Y(new_n5197));
  XNOR2x2_ASAP7_75t_L       g04941(.A(new_n3015), .B(new_n5192), .Y(new_n5198));
  OAI21xp33_ASAP7_75t_L     g04942(.A1(new_n5195), .A2(new_n5197), .B(new_n5198), .Y(new_n5199));
  NAND3xp33_ASAP7_75t_L     g04943(.A(new_n4731), .B(new_n4968), .C(new_n4971), .Y(new_n5200));
  NAND4xp25_ASAP7_75t_L     g04944(.A(new_n5200), .B(new_n4970), .C(new_n5194), .D(new_n5199), .Y(new_n5201));
  NOR3xp33_ASAP7_75t_L      g04945(.A(new_n5197), .B(new_n5195), .C(new_n5198), .Y(new_n5202));
  AOI21xp33_ASAP7_75t_L     g04946(.A1(new_n5187), .A2(new_n5190), .B(new_n5193), .Y(new_n5203));
  AOI211xp5_ASAP7_75t_L     g04947(.A1(new_n4974), .A2(new_n4717), .B(new_n4967), .C(new_n4965), .Y(new_n5204));
  OAI22xp33_ASAP7_75t_L     g04948(.A1(new_n5203), .A2(new_n5202), .B1(new_n4959), .B2(new_n5204), .Y(new_n5205));
  AO21x2_ASAP7_75t_L        g04949(.A1(new_n5201), .A2(new_n5205), .B(new_n5140), .Y(new_n5206));
  NAND3xp33_ASAP7_75t_L     g04950(.A(new_n5205), .B(new_n5201), .C(new_n5140), .Y(new_n5207));
  NAND3xp33_ASAP7_75t_L     g04951(.A(new_n5137), .B(new_n5206), .C(new_n5207), .Y(new_n5208));
  A2O1A1O1Ixp25_ASAP7_75t_L g04952(.A1(new_n4729), .A2(new_n4735), .B(new_n4738), .C(new_n4979), .D(new_n4977), .Y(new_n5209));
  AOI21xp33_ASAP7_75t_L     g04953(.A1(new_n5205), .A2(new_n5201), .B(new_n5140), .Y(new_n5210));
  AND3x1_ASAP7_75t_L        g04954(.A(new_n5205), .B(new_n5201), .C(new_n5140), .Y(new_n5211));
  OAI21xp33_ASAP7_75t_L     g04955(.A1(new_n5210), .A2(new_n5211), .B(new_n5209), .Y(new_n5212));
  AOI21xp33_ASAP7_75t_L     g04956(.A1(new_n5208), .A2(new_n5212), .B(new_n5136), .Y(new_n5213));
  AND2x2_ASAP7_75t_L        g04957(.A(new_n5133), .B(new_n5135), .Y(new_n5214));
  NOR3xp33_ASAP7_75t_L      g04958(.A(new_n5209), .B(new_n5210), .C(new_n5211), .Y(new_n5215));
  AOI21xp33_ASAP7_75t_L     g04959(.A1(new_n5207), .A2(new_n5206), .B(new_n5137), .Y(new_n5216));
  NOR3xp33_ASAP7_75t_L      g04960(.A(new_n5216), .B(new_n5215), .C(new_n5214), .Y(new_n5217));
  NOR2xp33_ASAP7_75t_L      g04961(.A(new_n5213), .B(new_n5217), .Y(new_n5218));
  A2O1A1Ixp33_ASAP7_75t_L   g04962(.A1(new_n5005), .A2(new_n4998), .B(new_n5129), .C(new_n5218), .Y(new_n5219));
  O2A1O1Ixp33_ASAP7_75t_L   g04963(.A1(new_n4985), .A2(new_n4991), .B(new_n5005), .C(new_n5129), .Y(new_n5220));
  OAI21xp33_ASAP7_75t_L     g04964(.A1(new_n5215), .A2(new_n5216), .B(new_n5214), .Y(new_n5221));
  NAND3xp33_ASAP7_75t_L     g04965(.A(new_n5208), .B(new_n5136), .C(new_n5212), .Y(new_n5222));
  NAND2xp33_ASAP7_75t_L     g04966(.A(new_n5222), .B(new_n5221), .Y(new_n5223));
  NAND2xp33_ASAP7_75t_L     g04967(.A(new_n5223), .B(new_n5220), .Y(new_n5224));
  AOI22xp33_ASAP7_75t_L     g04968(.A1(new_n1704), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1837), .Y(new_n5225));
  OAI21xp33_ASAP7_75t_L     g04969(.A1(new_n1827), .A2(new_n1547), .B(new_n5225), .Y(new_n5226));
  AOI211xp5_ASAP7_75t_L     g04970(.A1(\b[19] ), .A2(new_n1706), .B(new_n1689), .C(new_n5226), .Y(new_n5227));
  NAND2xp33_ASAP7_75t_L     g04971(.A(\b[19] ), .B(new_n1706), .Y(new_n5228));
  NAND2xp33_ASAP7_75t_L     g04972(.A(new_n1695), .B(new_n1886), .Y(new_n5229));
  AOI31xp33_ASAP7_75t_L     g04973(.A1(new_n5229), .A2(new_n5228), .A3(new_n5225), .B(\a[23] ), .Y(new_n5230));
  NOR2xp33_ASAP7_75t_L      g04974(.A(new_n5230), .B(new_n5227), .Y(new_n5231));
  NAND3xp33_ASAP7_75t_L     g04975(.A(new_n5219), .B(new_n5224), .C(new_n5231), .Y(new_n5232));
  INVx1_ASAP7_75t_L         g04976(.A(new_n5129), .Y(new_n5233));
  O2A1O1Ixp33_ASAP7_75t_L   g04977(.A1(new_n4992), .A2(new_n4994), .B(new_n5233), .C(new_n5223), .Y(new_n5234));
  AOI221xp5_ASAP7_75t_L     g04978(.A1(new_n5222), .A2(new_n5221), .B1(new_n5005), .B2(new_n4998), .C(new_n5129), .Y(new_n5235));
  NAND4xp25_ASAP7_75t_L     g04979(.A(new_n5229), .B(\a[23] ), .C(new_n5228), .D(new_n5225), .Y(new_n5236));
  A2O1A1Ixp33_ASAP7_75t_L   g04980(.A1(\b[19] ), .A2(new_n1706), .B(new_n5226), .C(new_n1689), .Y(new_n5237));
  NAND2xp33_ASAP7_75t_L     g04981(.A(new_n5236), .B(new_n5237), .Y(new_n5238));
  OAI21xp33_ASAP7_75t_L     g04982(.A1(new_n5235), .A2(new_n5234), .B(new_n5238), .Y(new_n5239));
  NAND2xp33_ASAP7_75t_L     g04983(.A(new_n5239), .B(new_n5232), .Y(new_n5240));
  NAND3xp33_ASAP7_75t_L     g04984(.A(new_n5008), .B(new_n4995), .C(new_n4999), .Y(new_n5241));
  A2O1A1Ixp33_ASAP7_75t_L   g04985(.A1(new_n5009), .A2(new_n5003), .B(new_n5011), .C(new_n5241), .Y(new_n5242));
  NOR2xp33_ASAP7_75t_L      g04986(.A(new_n5242), .B(new_n5240), .Y(new_n5243));
  NOR3xp33_ASAP7_75t_L      g04987(.A(new_n5234), .B(new_n5235), .C(new_n5238), .Y(new_n5244));
  INVx1_ASAP7_75t_L         g04988(.A(new_n5239), .Y(new_n5245));
  OA21x2_ASAP7_75t_L        g04989(.A1(new_n5244), .A2(new_n5245), .B(new_n5242), .Y(new_n5246));
  NOR2xp33_ASAP7_75t_L      g04990(.A(new_n1774), .B(new_n1373), .Y(new_n5247));
  INVx1_ASAP7_75t_L         g04991(.A(new_n5247), .Y(new_n5248));
  NAND3xp33_ASAP7_75t_L     g04992(.A(new_n1912), .B(new_n1365), .C(new_n1914), .Y(new_n5249));
  AOI22xp33_ASAP7_75t_L     g04993(.A1(new_n1360), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1581), .Y(new_n5250));
  AND4x1_ASAP7_75t_L        g04994(.A(new_n5250), .B(new_n5249), .C(new_n5248), .D(\a[20] ), .Y(new_n5251));
  AOI31xp33_ASAP7_75t_L     g04995(.A1(new_n5249), .A2(new_n5248), .A3(new_n5250), .B(\a[20] ), .Y(new_n5252));
  NOR2xp33_ASAP7_75t_L      g04996(.A(new_n5252), .B(new_n5251), .Y(new_n5253));
  OAI21xp33_ASAP7_75t_L     g04997(.A1(new_n5243), .A2(new_n5246), .B(new_n5253), .Y(new_n5254));
  NAND4xp25_ASAP7_75t_L     g04998(.A(new_n5022), .B(new_n5241), .C(new_n5239), .D(new_n5232), .Y(new_n5255));
  NAND2xp33_ASAP7_75t_L     g04999(.A(new_n5242), .B(new_n5240), .Y(new_n5256));
  INVx1_ASAP7_75t_L         g05000(.A(new_n5253), .Y(new_n5257));
  NAND3xp33_ASAP7_75t_L     g05001(.A(new_n5255), .B(new_n5256), .C(new_n5257), .Y(new_n5258));
  NAND2xp33_ASAP7_75t_L     g05002(.A(new_n5258), .B(new_n5254), .Y(new_n5259));
  NAND2xp33_ASAP7_75t_L     g05003(.A(new_n5259), .B(new_n5128), .Y(new_n5260));
  AOI21xp33_ASAP7_75t_L     g05004(.A1(new_n5255), .A2(new_n5256), .B(new_n5257), .Y(new_n5261));
  NOR3xp33_ASAP7_75t_L      g05005(.A(new_n5246), .B(new_n5243), .C(new_n5253), .Y(new_n5262));
  NOR2xp33_ASAP7_75t_L      g05006(.A(new_n5261), .B(new_n5262), .Y(new_n5263));
  A2O1A1Ixp33_ASAP7_75t_L   g05007(.A1(new_n5031), .A2(new_n5030), .B(new_n5127), .C(new_n5263), .Y(new_n5264));
  AOI21xp33_ASAP7_75t_L     g05008(.A1(new_n5264), .A2(new_n5260), .B(new_n5125), .Y(new_n5265));
  AOI221xp5_ASAP7_75t_L     g05009(.A1(new_n5031), .A2(new_n5030), .B1(new_n5258), .B2(new_n5254), .C(new_n5127), .Y(new_n5266));
  INVx1_ASAP7_75t_L         g05010(.A(new_n5026), .Y(new_n5267));
  O2A1O1Ixp33_ASAP7_75t_L   g05011(.A1(new_n4774), .A2(new_n4579), .B(new_n4773), .C(new_n5267), .Y(new_n5268));
  O2A1O1Ixp33_ASAP7_75t_L   g05012(.A1(new_n5025), .A2(new_n5268), .B(new_n5126), .C(new_n5259), .Y(new_n5269));
  NOR3xp33_ASAP7_75t_L      g05013(.A(new_n5269), .B(new_n5266), .C(new_n5124), .Y(new_n5270));
  NOR3xp33_ASAP7_75t_L      g05014(.A(new_n5121), .B(new_n5265), .C(new_n5270), .Y(new_n5271));
  NAND2xp33_ASAP7_75t_L     g05015(.A(new_n5039), .B(new_n5119), .Y(new_n5272));
  A2O1A1Ixp33_ASAP7_75t_L   g05016(.A1(new_n5040), .A2(new_n5036), .B(new_n5041), .C(new_n5272), .Y(new_n5273));
  NOR2xp33_ASAP7_75t_L      g05017(.A(new_n5270), .B(new_n5265), .Y(new_n5274));
  NOR2xp33_ASAP7_75t_L      g05018(.A(new_n5273), .B(new_n5274), .Y(new_n5275));
  OAI21xp33_ASAP7_75t_L     g05019(.A1(new_n5271), .A2(new_n5275), .B(new_n5118), .Y(new_n5276));
  INVx1_ASAP7_75t_L         g05020(.A(new_n5118), .Y(new_n5277));
  A2O1A1Ixp33_ASAP7_75t_L   g05021(.A1(new_n5039), .A2(new_n5119), .B(new_n5042), .C(new_n5274), .Y(new_n5278));
  OAI21xp33_ASAP7_75t_L     g05022(.A1(new_n5265), .A2(new_n5270), .B(new_n5121), .Y(new_n5279));
  NAND3xp33_ASAP7_75t_L     g05023(.A(new_n5278), .B(new_n5277), .C(new_n5279), .Y(new_n5280));
  NAND3xp33_ASAP7_75t_L     g05024(.A(new_n5115), .B(new_n5276), .C(new_n5280), .Y(new_n5281));
  NOR2xp33_ASAP7_75t_L      g05025(.A(new_n5042), .B(new_n5043), .Y(new_n5282));
  MAJIxp5_ASAP7_75t_L       g05026(.A(new_n4892), .B(new_n4896), .C(new_n5282), .Y(new_n5283));
  AOI21xp33_ASAP7_75t_L     g05027(.A1(new_n5278), .A2(new_n5279), .B(new_n5277), .Y(new_n5284));
  NOR3xp33_ASAP7_75t_L      g05028(.A(new_n5275), .B(new_n5271), .C(new_n5118), .Y(new_n5285));
  OAI21xp33_ASAP7_75t_L     g05029(.A1(new_n5284), .A2(new_n5285), .B(new_n5283), .Y(new_n5286));
  AOI21xp33_ASAP7_75t_L     g05030(.A1(new_n5281), .A2(new_n5286), .B(new_n5112), .Y(new_n5287));
  NOR3xp33_ASAP7_75t_L      g05031(.A(new_n5283), .B(new_n5284), .C(new_n5285), .Y(new_n5288));
  AOI221xp5_ASAP7_75t_L     g05032(.A1(new_n4892), .A2(new_n5060), .B1(new_n5276), .B2(new_n5280), .C(new_n5113), .Y(new_n5289));
  NOR3xp33_ASAP7_75t_L      g05033(.A(new_n5288), .B(new_n5289), .C(new_n5111), .Y(new_n5290));
  OR3x1_ASAP7_75t_L         g05034(.A(new_n5104), .B(new_n5287), .C(new_n5290), .Y(new_n5291));
  OAI21xp33_ASAP7_75t_L     g05035(.A1(new_n5290), .A2(new_n5287), .B(new_n5104), .Y(new_n5292));
  NAND2xp33_ASAP7_75t_L     g05036(.A(\b[34] ), .B(new_n447), .Y(new_n5293));
  NAND2xp33_ASAP7_75t_L     g05037(.A(new_n441), .B(new_n3811), .Y(new_n5294));
  AOI22xp33_ASAP7_75t_L     g05038(.A1(new_n444), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n471), .Y(new_n5295));
  NAND4xp25_ASAP7_75t_L     g05039(.A(new_n5294), .B(\a[8] ), .C(new_n5293), .D(new_n5295), .Y(new_n5296));
  NAND2xp33_ASAP7_75t_L     g05040(.A(new_n5295), .B(new_n5294), .Y(new_n5297));
  A2O1A1Ixp33_ASAP7_75t_L   g05041(.A1(\b[34] ), .A2(new_n447), .B(new_n5297), .C(new_n435), .Y(new_n5298));
  NAND2xp33_ASAP7_75t_L     g05042(.A(new_n5296), .B(new_n5298), .Y(new_n5299));
  INVx1_ASAP7_75t_L         g05043(.A(new_n5299), .Y(new_n5300));
  NAND3xp33_ASAP7_75t_L     g05044(.A(new_n5291), .B(new_n5300), .C(new_n5292), .Y(new_n5301));
  NOR3xp33_ASAP7_75t_L      g05045(.A(new_n5104), .B(new_n5287), .C(new_n5290), .Y(new_n5302));
  INVx1_ASAP7_75t_L         g05046(.A(new_n5292), .Y(new_n5303));
  OAI21xp33_ASAP7_75t_L     g05047(.A1(new_n5302), .A2(new_n5303), .B(new_n5299), .Y(new_n5304));
  NAND2xp33_ASAP7_75t_L     g05048(.A(new_n5301), .B(new_n5304), .Y(new_n5305));
  A2O1A1Ixp33_ASAP7_75t_L   g05049(.A1(new_n5074), .A2(new_n5103), .B(new_n5070), .C(new_n5305), .Y(new_n5306));
  A2O1A1O1Ixp25_ASAP7_75t_L g05050(.A1(new_n4836), .A2(new_n4835), .B(new_n4886), .C(new_n5074), .D(new_n5070), .Y(new_n5307));
  NOR3xp33_ASAP7_75t_L      g05051(.A(new_n5303), .B(new_n5299), .C(new_n5302), .Y(new_n5308));
  AOI21xp33_ASAP7_75t_L     g05052(.A1(new_n5291), .A2(new_n5292), .B(new_n5300), .Y(new_n5309));
  NOR2xp33_ASAP7_75t_L      g05053(.A(new_n5309), .B(new_n5308), .Y(new_n5310));
  NAND2xp33_ASAP7_75t_L     g05054(.A(new_n5307), .B(new_n5310), .Y(new_n5311));
  NAND3xp33_ASAP7_75t_L     g05055(.A(new_n5306), .B(new_n5311), .C(new_n5102), .Y(new_n5312));
  O2A1O1Ixp33_ASAP7_75t_L   g05056(.A1(new_n5073), .A2(new_n5069), .B(new_n5075), .C(new_n5310), .Y(new_n5313));
  OAI21xp33_ASAP7_75t_L     g05057(.A1(new_n5076), .A2(new_n5073), .B(new_n5075), .Y(new_n5314));
  NOR2xp33_ASAP7_75t_L      g05058(.A(new_n5305), .B(new_n5314), .Y(new_n5315));
  OAI21xp33_ASAP7_75t_L     g05059(.A1(new_n5315), .A2(new_n5313), .B(new_n5101), .Y(new_n5316));
  AOI21xp33_ASAP7_75t_L     g05060(.A1(new_n5316), .A2(new_n5312), .B(new_n5098), .Y(new_n5317));
  NAND2xp33_ASAP7_75t_L     g05061(.A(new_n5312), .B(new_n5316), .Y(new_n5318));
  A2O1A1O1Ixp25_ASAP7_75t_L g05062(.A1(new_n5081), .A2(new_n5085), .B(new_n5088), .C(new_n5097), .D(new_n5318), .Y(new_n5319));
  NOR2xp33_ASAP7_75t_L      g05063(.A(\b[40] ), .B(\b[41] ), .Y(new_n5320));
  INVx1_ASAP7_75t_L         g05064(.A(\b[41] ), .Y(new_n5321));
  NOR2xp33_ASAP7_75t_L      g05065(.A(new_n4869), .B(new_n5321), .Y(new_n5322));
  NOR2xp33_ASAP7_75t_L      g05066(.A(new_n5320), .B(new_n5322), .Y(new_n5323));
  A2O1A1Ixp33_ASAP7_75t_L   g05067(.A1(new_n4874), .A2(new_n4871), .B(new_n4870), .C(new_n5323), .Y(new_n5324));
  O2A1O1Ixp33_ASAP7_75t_L   g05068(.A1(new_n4849), .A2(new_n4852), .B(new_n4871), .C(new_n4870), .Y(new_n5325));
  OAI21xp33_ASAP7_75t_L     g05069(.A1(new_n5320), .A2(new_n5322), .B(new_n5325), .Y(new_n5326));
  NAND2xp33_ASAP7_75t_L     g05070(.A(new_n5324), .B(new_n5326), .Y(new_n5327));
  AOI22xp33_ASAP7_75t_L     g05071(.A1(\b[39] ), .A2(new_n282), .B1(\b[41] ), .B2(new_n303), .Y(new_n5328));
  OAI221xp5_ASAP7_75t_L     g05072(.A1(new_n291), .A2(new_n4869), .B1(new_n268), .B2(new_n5327), .C(new_n5328), .Y(new_n5329));
  XNOR2x2_ASAP7_75t_L       g05073(.A(\a[2] ), .B(new_n5329), .Y(new_n5330));
  OAI21xp33_ASAP7_75t_L     g05074(.A1(new_n5317), .A2(new_n5319), .B(new_n5330), .Y(new_n5331));
  NOR3xp33_ASAP7_75t_L      g05075(.A(new_n5319), .B(new_n5330), .C(new_n5317), .Y(new_n5332));
  INVx1_ASAP7_75t_L         g05076(.A(new_n5332), .Y(new_n5333));
  NAND2xp33_ASAP7_75t_L     g05077(.A(new_n5331), .B(new_n5333), .Y(new_n5334));
  XOR2x2_ASAP7_75t_L        g05078(.A(new_n5096), .B(new_n5334), .Y(\f[41] ));
  INVx1_ASAP7_75t_L         g05079(.A(new_n5322), .Y(new_n5336));
  NOR2xp33_ASAP7_75t_L      g05080(.A(\b[41] ), .B(\b[42] ), .Y(new_n5337));
  INVx1_ASAP7_75t_L         g05081(.A(\b[42] ), .Y(new_n5338));
  NOR2xp33_ASAP7_75t_L      g05082(.A(new_n5321), .B(new_n5338), .Y(new_n5339));
  NOR2xp33_ASAP7_75t_L      g05083(.A(new_n5337), .B(new_n5339), .Y(new_n5340));
  INVx1_ASAP7_75t_L         g05084(.A(new_n5340), .Y(new_n5341));
  O2A1O1Ixp33_ASAP7_75t_L   g05085(.A1(new_n5320), .A2(new_n5325), .B(new_n5336), .C(new_n5341), .Y(new_n5342));
  INVx1_ASAP7_75t_L         g05086(.A(new_n5342), .Y(new_n5343));
  A2O1A1O1Ixp25_ASAP7_75t_L g05087(.A1(new_n4871), .A2(new_n4874), .B(new_n4870), .C(new_n5323), .D(new_n5322), .Y(new_n5344));
  NAND2xp33_ASAP7_75t_L     g05088(.A(new_n5341), .B(new_n5344), .Y(new_n5345));
  NAND2xp33_ASAP7_75t_L     g05089(.A(new_n5345), .B(new_n5343), .Y(new_n5346));
  AOI22xp33_ASAP7_75t_L     g05090(.A1(\b[40] ), .A2(new_n282), .B1(\b[42] ), .B2(new_n303), .Y(new_n5347));
  OAI221xp5_ASAP7_75t_L     g05091(.A1(new_n291), .A2(new_n5321), .B1(new_n268), .B2(new_n5346), .C(new_n5347), .Y(new_n5348));
  XNOR2x2_ASAP7_75t_L       g05092(.A(\a[2] ), .B(new_n5348), .Y(new_n5349));
  NOR3xp33_ASAP7_75t_L      g05093(.A(new_n5313), .B(new_n5315), .C(new_n5101), .Y(new_n5350));
  NAND2xp33_ASAP7_75t_L     g05094(.A(\b[38] ), .B(new_n347), .Y(new_n5351));
  INVx1_ASAP7_75t_L         g05095(.A(new_n4858), .Y(new_n5352));
  NAND2xp33_ASAP7_75t_L     g05096(.A(new_n341), .B(new_n5352), .Y(new_n5353));
  AOI22xp33_ASAP7_75t_L     g05097(.A1(new_n344), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n370), .Y(new_n5354));
  AND4x1_ASAP7_75t_L        g05098(.A(new_n5354), .B(new_n5353), .C(new_n5351), .D(\a[5] ), .Y(new_n5355));
  AOI31xp33_ASAP7_75t_L     g05099(.A1(new_n5353), .A2(new_n5351), .A3(new_n5354), .B(\a[5] ), .Y(new_n5356));
  NAND3xp33_ASAP7_75t_L     g05100(.A(new_n5291), .B(new_n5292), .C(new_n5299), .Y(new_n5357));
  AOI22xp33_ASAP7_75t_L     g05101(.A1(new_n444), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n471), .Y(new_n5358));
  OAI21xp33_ASAP7_75t_L     g05102(.A1(new_n469), .A2(new_n4223), .B(new_n5358), .Y(new_n5359));
  AOI21xp33_ASAP7_75t_L     g05103(.A1(new_n447), .A2(\b[35] ), .B(new_n5359), .Y(new_n5360));
  NAND2xp33_ASAP7_75t_L     g05104(.A(\a[8] ), .B(new_n5360), .Y(new_n5361));
  A2O1A1Ixp33_ASAP7_75t_L   g05105(.A1(\b[35] ), .A2(new_n447), .B(new_n5359), .C(new_n435), .Y(new_n5362));
  AND2x2_ASAP7_75t_L        g05106(.A(new_n5362), .B(new_n5361), .Y(new_n5363));
  OAI21xp33_ASAP7_75t_L     g05107(.A1(new_n5289), .A2(new_n5288), .B(new_n5111), .Y(new_n5364));
  A2O1A1O1Ixp25_ASAP7_75t_L g05108(.A1(new_n5057), .A2(new_n4890), .B(new_n5067), .C(new_n5364), .D(new_n5290), .Y(new_n5365));
  OAI21xp33_ASAP7_75t_L     g05109(.A1(new_n5284), .A2(new_n5283), .B(new_n5280), .Y(new_n5366));
  NOR2xp33_ASAP7_75t_L      g05110(.A(new_n2688), .B(new_n904), .Y(new_n5367));
  INVx1_ASAP7_75t_L         g05111(.A(new_n5367), .Y(new_n5368));
  NAND2xp33_ASAP7_75t_L     g05112(.A(new_n808), .B(new_n2989), .Y(new_n5369));
  AOI22xp33_ASAP7_75t_L     g05113(.A1(new_n811), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n900), .Y(new_n5370));
  AND4x1_ASAP7_75t_L        g05114(.A(new_n5370), .B(new_n5369), .C(new_n5368), .D(\a[14] ), .Y(new_n5371));
  AOI31xp33_ASAP7_75t_L     g05115(.A1(new_n5369), .A2(new_n5368), .A3(new_n5370), .B(\a[14] ), .Y(new_n5372));
  NOR2xp33_ASAP7_75t_L      g05116(.A(new_n5372), .B(new_n5371), .Y(new_n5373));
  INVx1_ASAP7_75t_L         g05117(.A(new_n5373), .Y(new_n5374));
  OAI21xp33_ASAP7_75t_L     g05118(.A1(new_n5266), .A2(new_n5269), .B(new_n5124), .Y(new_n5375));
  A2O1A1Ixp33_ASAP7_75t_L   g05119(.A1(new_n4751), .A2(new_n5004), .B(new_n4992), .C(new_n5233), .Y(new_n5376));
  OAI21xp33_ASAP7_75t_L     g05120(.A1(new_n5210), .A2(new_n5209), .B(new_n5207), .Y(new_n5377));
  AOI22xp33_ASAP7_75t_L     g05121(.A1(new_n2552), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n2736), .Y(new_n5378));
  OAI221xp5_ASAP7_75t_L     g05122(.A1(new_n2547), .A2(new_n869), .B1(new_n2734), .B2(new_n950), .C(new_n5378), .Y(new_n5379));
  XNOR2x2_ASAP7_75t_L       g05123(.A(new_n2538), .B(new_n5379), .Y(new_n5380));
  INVx1_ASAP7_75t_L         g05124(.A(new_n5380), .Y(new_n5381));
  OAI31xp33_ASAP7_75t_L     g05125(.A1(new_n5204), .A2(new_n5202), .A3(new_n4959), .B(new_n5199), .Y(new_n5382));
  AOI22xp33_ASAP7_75t_L     g05126(.A1(new_n3029), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n3258), .Y(new_n5383));
  INVx1_ASAP7_75t_L         g05127(.A(new_n5383), .Y(new_n5384));
  AOI221xp5_ASAP7_75t_L     g05128(.A1(new_n3030), .A2(\b[11] ), .B1(new_n3021), .B2(new_n1232), .C(new_n5384), .Y(new_n5385));
  XNOR2x2_ASAP7_75t_L       g05129(.A(new_n3015), .B(new_n5385), .Y(new_n5386));
  NOR3xp33_ASAP7_75t_L      g05130(.A(new_n5180), .B(new_n5182), .C(new_n5177), .Y(new_n5387));
  NAND5xp2_ASAP7_75t_L      g05131(.A(\a[41] ), .B(new_n4918), .C(new_n4921), .D(new_n4925), .E(new_n4677), .Y(new_n5388));
  INVx1_ASAP7_75t_L         g05132(.A(\a[42] ), .Y(new_n5389));
  NAND2xp33_ASAP7_75t_L     g05133(.A(\a[41] ), .B(new_n5389), .Y(new_n5390));
  NAND2xp33_ASAP7_75t_L     g05134(.A(\a[42] ), .B(new_n4915), .Y(new_n5391));
  AND2x2_ASAP7_75t_L        g05135(.A(new_n5390), .B(new_n5391), .Y(new_n5392));
  NOR2xp33_ASAP7_75t_L      g05136(.A(new_n258), .B(new_n5392), .Y(new_n5393));
  OAI31xp33_ASAP7_75t_L     g05137(.A1(new_n5388), .A2(new_n5161), .A3(new_n5157), .B(new_n5393), .Y(new_n5394));
  NOR2xp33_ASAP7_75t_L      g05138(.A(new_n4915), .B(new_n4674), .Y(new_n5395));
  INVx1_ASAP7_75t_L         g05139(.A(new_n5393), .Y(new_n5396));
  NAND5xp2_ASAP7_75t_L      g05140(.A(new_n5156), .B(new_n5396), .C(new_n5168), .D(new_n5395), .E(new_n5165), .Y(new_n5397));
  NOR2xp33_ASAP7_75t_L      g05141(.A(new_n276), .B(new_n5154), .Y(new_n5398));
  NAND2xp33_ASAP7_75t_L     g05142(.A(\b[3] ), .B(new_n4920), .Y(new_n5399));
  OAI221xp5_ASAP7_75t_L     g05143(.A1(new_n5160), .A2(new_n261), .B1(new_n5158), .B2(new_n302), .C(new_n5399), .Y(new_n5400));
  OR3x1_ASAP7_75t_L         g05144(.A(new_n5400), .B(new_n4915), .C(new_n5398), .Y(new_n5401));
  A2O1A1Ixp33_ASAP7_75t_L   g05145(.A1(\b[2] ), .A2(new_n4924), .B(new_n5400), .C(new_n4915), .Y(new_n5402));
  AO22x1_ASAP7_75t_L        g05146(.A1(new_n5394), .A2(new_n5397), .B1(new_n5402), .B2(new_n5401), .Y(new_n5403));
  NAND4xp25_ASAP7_75t_L     g05147(.A(new_n5401), .B(new_n5397), .C(new_n5394), .D(new_n5402), .Y(new_n5404));
  NAND2xp33_ASAP7_75t_L     g05148(.A(\b[5] ), .B(new_n4285), .Y(new_n5405));
  NAND2xp33_ASAP7_75t_L     g05149(.A(new_n4274), .B(new_n526), .Y(new_n5406));
  AOI22xp33_ASAP7_75t_L     g05150(.A1(new_n4283), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n4512), .Y(new_n5407));
  NAND4xp25_ASAP7_75t_L     g05151(.A(new_n5406), .B(\a[38] ), .C(new_n5405), .D(new_n5407), .Y(new_n5408));
  AOI31xp33_ASAP7_75t_L     g05152(.A1(new_n5406), .A2(new_n5405), .A3(new_n5407), .B(\a[38] ), .Y(new_n5409));
  INVx1_ASAP7_75t_L         g05153(.A(new_n5409), .Y(new_n5410));
  NAND4xp25_ASAP7_75t_L     g05154(.A(new_n5410), .B(new_n5403), .C(new_n5404), .D(new_n5408), .Y(new_n5411));
  AOI22xp33_ASAP7_75t_L     g05155(.A1(new_n5397), .A2(new_n5394), .B1(new_n5402), .B2(new_n5401), .Y(new_n5412));
  AND4x1_ASAP7_75t_L        g05156(.A(new_n5397), .B(new_n5401), .C(new_n5394), .D(new_n5402), .Y(new_n5413));
  INVx1_ASAP7_75t_L         g05157(.A(new_n5408), .Y(new_n5414));
  OAI22xp33_ASAP7_75t_L     g05158(.A1(new_n5414), .A2(new_n5409), .B1(new_n5412), .B2(new_n5413), .Y(new_n5415));
  AND2x2_ASAP7_75t_L        g05159(.A(new_n5415), .B(new_n5411), .Y(new_n5416));
  NAND2xp33_ASAP7_75t_L     g05160(.A(new_n5152), .B(new_n5151), .Y(new_n5417));
  NOR2xp33_ASAP7_75t_L      g05161(.A(new_n5173), .B(new_n5175), .Y(new_n5418));
  MAJIxp5_ASAP7_75t_L       g05162(.A(new_n5178), .B(new_n5417), .C(new_n5418), .Y(new_n5419));
  NAND2xp33_ASAP7_75t_L     g05163(.A(new_n5419), .B(new_n5416), .Y(new_n5420));
  NAND2xp33_ASAP7_75t_L     g05164(.A(new_n5415), .B(new_n5411), .Y(new_n5421));
  A2O1A1Ixp33_ASAP7_75t_L   g05165(.A1(new_n5418), .A2(new_n5417), .B(new_n5177), .C(new_n5421), .Y(new_n5422));
  NAND2xp33_ASAP7_75t_L     g05166(.A(\b[8] ), .B(new_n3639), .Y(new_n5423));
  NAND2xp33_ASAP7_75t_L     g05167(.A(new_n3630), .B(new_n731), .Y(new_n5424));
  AOI22xp33_ASAP7_75t_L     g05168(.A1(new_n3633), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n3858), .Y(new_n5425));
  NAND4xp25_ASAP7_75t_L     g05169(.A(new_n5424), .B(\a[35] ), .C(new_n5423), .D(new_n5425), .Y(new_n5426));
  OAI211xp5_ASAP7_75t_L     g05170(.A1(new_n3856), .A2(new_n548), .B(new_n5423), .C(new_n5425), .Y(new_n5427));
  NAND2xp33_ASAP7_75t_L     g05171(.A(new_n3628), .B(new_n5427), .Y(new_n5428));
  NAND2xp33_ASAP7_75t_L     g05172(.A(new_n5428), .B(new_n5426), .Y(new_n5429));
  AOI21xp33_ASAP7_75t_L     g05173(.A1(new_n5422), .A2(new_n5420), .B(new_n5429), .Y(new_n5430));
  NAND2xp33_ASAP7_75t_L     g05174(.A(new_n5417), .B(new_n5418), .Y(new_n5431));
  A2O1A1Ixp33_ASAP7_75t_L   g05175(.A1(new_n5171), .A2(new_n5176), .B(new_n5146), .C(new_n5431), .Y(new_n5432));
  NOR2xp33_ASAP7_75t_L      g05176(.A(new_n5421), .B(new_n5432), .Y(new_n5433));
  NOR2xp33_ASAP7_75t_L      g05177(.A(new_n5419), .B(new_n5416), .Y(new_n5434));
  AOI211xp5_ASAP7_75t_L     g05178(.A1(new_n5428), .A2(new_n5426), .B(new_n5433), .C(new_n5434), .Y(new_n5435));
  NOR2xp33_ASAP7_75t_L      g05179(.A(new_n5430), .B(new_n5435), .Y(new_n5436));
  A2O1A1Ixp33_ASAP7_75t_L   g05180(.A1(new_n5189), .A2(new_n5196), .B(new_n5387), .C(new_n5436), .Y(new_n5437));
  AOI21xp33_ASAP7_75t_L     g05181(.A1(new_n5196), .A2(new_n5189), .B(new_n5387), .Y(new_n5438));
  OAI211xp5_ASAP7_75t_L     g05182(.A1(new_n5433), .A2(new_n5434), .B(new_n5426), .C(new_n5428), .Y(new_n5439));
  NAND3xp33_ASAP7_75t_L     g05183(.A(new_n5429), .B(new_n5420), .C(new_n5422), .Y(new_n5440));
  NAND2xp33_ASAP7_75t_L     g05184(.A(new_n5440), .B(new_n5439), .Y(new_n5441));
  NAND2xp33_ASAP7_75t_L     g05185(.A(new_n5438), .B(new_n5441), .Y(new_n5442));
  AOI21xp33_ASAP7_75t_L     g05186(.A1(new_n5437), .A2(new_n5442), .B(new_n5386), .Y(new_n5443));
  XNOR2x2_ASAP7_75t_L       g05187(.A(\a[32] ), .B(new_n5385), .Y(new_n5444));
  NOR2xp33_ASAP7_75t_L      g05188(.A(new_n5438), .B(new_n5441), .Y(new_n5445));
  AOI221xp5_ASAP7_75t_L     g05189(.A1(new_n5196), .A2(new_n5189), .B1(new_n5440), .B2(new_n5439), .C(new_n5387), .Y(new_n5446));
  NOR3xp33_ASAP7_75t_L      g05190(.A(new_n5445), .B(new_n5446), .C(new_n5444), .Y(new_n5447));
  OAI21xp33_ASAP7_75t_L     g05191(.A1(new_n5443), .A2(new_n5447), .B(new_n5382), .Y(new_n5448));
  AOI31xp33_ASAP7_75t_L     g05192(.A1(new_n5200), .A2(new_n5194), .A3(new_n4970), .B(new_n5203), .Y(new_n5449));
  OAI21xp33_ASAP7_75t_L     g05193(.A1(new_n5446), .A2(new_n5445), .B(new_n5444), .Y(new_n5450));
  NAND3xp33_ASAP7_75t_L     g05194(.A(new_n5437), .B(new_n5442), .C(new_n5386), .Y(new_n5451));
  NAND3xp33_ASAP7_75t_L     g05195(.A(new_n5449), .B(new_n5450), .C(new_n5451), .Y(new_n5452));
  NAND3xp33_ASAP7_75t_L     g05196(.A(new_n5381), .B(new_n5448), .C(new_n5452), .Y(new_n5453));
  AOI21xp33_ASAP7_75t_L     g05197(.A1(new_n5451), .A2(new_n5450), .B(new_n5449), .Y(new_n5454));
  NOR3xp33_ASAP7_75t_L      g05198(.A(new_n5382), .B(new_n5443), .C(new_n5447), .Y(new_n5455));
  OAI21xp33_ASAP7_75t_L     g05199(.A1(new_n5454), .A2(new_n5455), .B(new_n5380), .Y(new_n5456));
  NAND3xp33_ASAP7_75t_L     g05200(.A(new_n5377), .B(new_n5453), .C(new_n5456), .Y(new_n5457));
  A2O1A1O1Ixp25_ASAP7_75t_L g05201(.A1(new_n4979), .A2(new_n4987), .B(new_n4977), .C(new_n5206), .D(new_n5211), .Y(new_n5458));
  NOR3xp33_ASAP7_75t_L      g05202(.A(new_n5455), .B(new_n5454), .C(new_n5380), .Y(new_n5459));
  AOI21xp33_ASAP7_75t_L     g05203(.A1(new_n5452), .A2(new_n5448), .B(new_n5381), .Y(new_n5460));
  OAI21xp33_ASAP7_75t_L     g05204(.A1(new_n5459), .A2(new_n5460), .B(new_n5458), .Y(new_n5461));
  AOI22xp33_ASAP7_75t_L     g05205(.A1(new_n2114), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n2259), .Y(new_n5462));
  OAI31xp33_ASAP7_75t_L     g05206(.A1(new_n1318), .A2(new_n1317), .A3(new_n2257), .B(new_n5462), .Y(new_n5463));
  AOI21xp33_ASAP7_75t_L     g05207(.A1(new_n2115), .A2(\b[17] ), .B(new_n5463), .Y(new_n5464));
  NAND2xp33_ASAP7_75t_L     g05208(.A(\a[26] ), .B(new_n5464), .Y(new_n5465));
  A2O1A1Ixp33_ASAP7_75t_L   g05209(.A1(\b[17] ), .A2(new_n2115), .B(new_n5463), .C(new_n2100), .Y(new_n5466));
  AND2x2_ASAP7_75t_L        g05210(.A(new_n5466), .B(new_n5465), .Y(new_n5467));
  AOI21xp33_ASAP7_75t_L     g05211(.A1(new_n5457), .A2(new_n5461), .B(new_n5467), .Y(new_n5468));
  NOR3xp33_ASAP7_75t_L      g05212(.A(new_n5458), .B(new_n5459), .C(new_n5460), .Y(new_n5469));
  AOI21xp33_ASAP7_75t_L     g05213(.A1(new_n5456), .A2(new_n5453), .B(new_n5377), .Y(new_n5470));
  NAND2xp33_ASAP7_75t_L     g05214(.A(new_n5466), .B(new_n5465), .Y(new_n5471));
  NOR3xp33_ASAP7_75t_L      g05215(.A(new_n5469), .B(new_n5470), .C(new_n5471), .Y(new_n5472));
  NOR2xp33_ASAP7_75t_L      g05216(.A(new_n5468), .B(new_n5472), .Y(new_n5473));
  A2O1A1Ixp33_ASAP7_75t_L   g05217(.A1(new_n5218), .A2(new_n5376), .B(new_n5217), .C(new_n5473), .Y(new_n5474));
  A2O1A1O1Ixp25_ASAP7_75t_L g05218(.A1(new_n5005), .A2(new_n4998), .B(new_n5129), .C(new_n5221), .D(new_n5217), .Y(new_n5475));
  OAI21xp33_ASAP7_75t_L     g05219(.A1(new_n5470), .A2(new_n5469), .B(new_n5471), .Y(new_n5476));
  NAND3xp33_ASAP7_75t_L     g05220(.A(new_n5467), .B(new_n5457), .C(new_n5461), .Y(new_n5477));
  NAND2xp33_ASAP7_75t_L     g05221(.A(new_n5476), .B(new_n5477), .Y(new_n5478));
  NAND2xp33_ASAP7_75t_L     g05222(.A(new_n5475), .B(new_n5478), .Y(new_n5479));
  AOI22xp33_ASAP7_75t_L     g05223(.A1(new_n1704), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1837), .Y(new_n5480));
  OAI31xp33_ASAP7_75t_L     g05224(.A1(new_n1660), .A2(new_n1659), .A3(new_n1827), .B(new_n5480), .Y(new_n5481));
  AOI211xp5_ASAP7_75t_L     g05225(.A1(\b[20] ), .A2(new_n1706), .B(new_n1689), .C(new_n5481), .Y(new_n5482));
  AOI21xp33_ASAP7_75t_L     g05226(.A1(new_n1706), .A2(\b[20] ), .B(new_n5481), .Y(new_n5483));
  NOR2xp33_ASAP7_75t_L      g05227(.A(\a[23] ), .B(new_n5483), .Y(new_n5484));
  NOR2xp33_ASAP7_75t_L      g05228(.A(new_n5482), .B(new_n5484), .Y(new_n5485));
  NAND3xp33_ASAP7_75t_L     g05229(.A(new_n5474), .B(new_n5479), .C(new_n5485), .Y(new_n5486));
  NOR2xp33_ASAP7_75t_L      g05230(.A(new_n5475), .B(new_n5478), .Y(new_n5487));
  AOI221xp5_ASAP7_75t_L     g05231(.A1(new_n5477), .A2(new_n5476), .B1(new_n5218), .B2(new_n5376), .C(new_n5217), .Y(new_n5488));
  OR2x4_ASAP7_75t_L         g05232(.A(new_n5482), .B(new_n5484), .Y(new_n5489));
  OAI21xp33_ASAP7_75t_L     g05233(.A1(new_n5487), .A2(new_n5488), .B(new_n5489), .Y(new_n5490));
  NAND2xp33_ASAP7_75t_L     g05234(.A(new_n5490), .B(new_n5486), .Y(new_n5491));
  NOR3xp33_ASAP7_75t_L      g05235(.A(new_n5234), .B(new_n5231), .C(new_n5235), .Y(new_n5492));
  NOR3xp33_ASAP7_75t_L      g05236(.A(new_n5246), .B(new_n5491), .C(new_n5492), .Y(new_n5493));
  NOR3xp33_ASAP7_75t_L      g05237(.A(new_n5488), .B(new_n5487), .C(new_n5489), .Y(new_n5494));
  AOI21xp33_ASAP7_75t_L     g05238(.A1(new_n5474), .A2(new_n5479), .B(new_n5485), .Y(new_n5495));
  NOR2xp33_ASAP7_75t_L      g05239(.A(new_n5494), .B(new_n5495), .Y(new_n5496));
  NOR2xp33_ASAP7_75t_L      g05240(.A(new_n5235), .B(new_n5234), .Y(new_n5497));
  MAJIxp5_ASAP7_75t_L       g05241(.A(new_n5242), .B(new_n5497), .C(new_n5238), .Y(new_n5498));
  NOR2xp33_ASAP7_75t_L      g05242(.A(new_n5498), .B(new_n5496), .Y(new_n5499));
  AOI22xp33_ASAP7_75t_L     g05243(.A1(new_n1360), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n1581), .Y(new_n5500));
  INVx1_ASAP7_75t_L         g05244(.A(new_n5500), .Y(new_n5501));
  AOI221xp5_ASAP7_75t_L     g05245(.A1(\b[23] ), .A2(new_n1362), .B1(new_n1365), .B2(new_n1935), .C(new_n5501), .Y(new_n5502));
  XNOR2x2_ASAP7_75t_L       g05246(.A(new_n1356), .B(new_n5502), .Y(new_n5503));
  OAI21xp33_ASAP7_75t_L     g05247(.A1(new_n5499), .A2(new_n5493), .B(new_n5503), .Y(new_n5504));
  NAND2xp33_ASAP7_75t_L     g05248(.A(new_n5498), .B(new_n5496), .Y(new_n5505));
  A2O1A1Ixp33_ASAP7_75t_L   g05249(.A1(new_n5240), .A2(new_n5242), .B(new_n5492), .C(new_n5491), .Y(new_n5506));
  XNOR2x2_ASAP7_75t_L       g05250(.A(\a[20] ), .B(new_n5502), .Y(new_n5507));
  NAND3xp33_ASAP7_75t_L     g05251(.A(new_n5506), .B(new_n5507), .C(new_n5505), .Y(new_n5508));
  OAI211xp5_ASAP7_75t_L     g05252(.A1(new_n5025), .A2(new_n5268), .B(new_n5126), .C(new_n5258), .Y(new_n5509));
  NAND4xp25_ASAP7_75t_L     g05253(.A(new_n5509), .B(new_n5254), .C(new_n5504), .D(new_n5508), .Y(new_n5510));
  AOI21xp33_ASAP7_75t_L     g05254(.A1(new_n5506), .A2(new_n5505), .B(new_n5507), .Y(new_n5511));
  NOR3xp33_ASAP7_75t_L      g05255(.A(new_n5493), .B(new_n5499), .C(new_n5503), .Y(new_n5512));
  AOI211xp5_ASAP7_75t_L     g05256(.A1(new_n5031), .A2(new_n5030), .B(new_n5127), .C(new_n5262), .Y(new_n5513));
  OAI22xp33_ASAP7_75t_L     g05257(.A1(new_n5513), .A2(new_n5261), .B1(new_n5511), .B2(new_n5512), .Y(new_n5514));
  NOR2xp33_ASAP7_75t_L      g05258(.A(new_n2348), .B(new_n1154), .Y(new_n5515));
  INVx1_ASAP7_75t_L         g05259(.A(new_n5515), .Y(new_n5516));
  NAND2xp33_ASAP7_75t_L     g05260(.A(new_n1073), .B(new_n2504), .Y(new_n5517));
  AOI22xp33_ASAP7_75t_L     g05261(.A1(new_n1076), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1253), .Y(new_n5518));
  AND4x1_ASAP7_75t_L        g05262(.A(new_n5518), .B(new_n5517), .C(new_n5516), .D(\a[17] ), .Y(new_n5519));
  AOI31xp33_ASAP7_75t_L     g05263(.A1(new_n5517), .A2(new_n5516), .A3(new_n5518), .B(\a[17] ), .Y(new_n5520));
  NOR2xp33_ASAP7_75t_L      g05264(.A(new_n5520), .B(new_n5519), .Y(new_n5521));
  NAND3xp33_ASAP7_75t_L     g05265(.A(new_n5510), .B(new_n5514), .C(new_n5521), .Y(new_n5522));
  NOR4xp25_ASAP7_75t_L      g05266(.A(new_n5513), .B(new_n5512), .C(new_n5261), .D(new_n5511), .Y(new_n5523));
  AOI22xp33_ASAP7_75t_L     g05267(.A1(new_n5508), .A2(new_n5504), .B1(new_n5254), .B2(new_n5509), .Y(new_n5524));
  INVx1_ASAP7_75t_L         g05268(.A(new_n5521), .Y(new_n5525));
  OAI21xp33_ASAP7_75t_L     g05269(.A1(new_n5523), .A2(new_n5524), .B(new_n5525), .Y(new_n5526));
  NAND2xp33_ASAP7_75t_L     g05270(.A(new_n5522), .B(new_n5526), .Y(new_n5527));
  A2O1A1Ixp33_ASAP7_75t_L   g05271(.A1(new_n5375), .A2(new_n5273), .B(new_n5270), .C(new_n5527), .Y(new_n5528));
  NAND2xp33_ASAP7_75t_L     g05272(.A(new_n5036), .B(new_n5040), .Y(new_n5529));
  NAND2xp33_ASAP7_75t_L     g05273(.A(new_n5032), .B(new_n5027), .Y(new_n5530));
  NOR2xp33_ASAP7_75t_L      g05274(.A(new_n5035), .B(new_n5530), .Y(new_n5531));
  A2O1A1O1Ixp25_ASAP7_75t_L g05275(.A1(new_n5120), .A2(new_n5529), .B(new_n5531), .C(new_n5375), .D(new_n5270), .Y(new_n5532));
  NAND3xp33_ASAP7_75t_L     g05276(.A(new_n5532), .B(new_n5522), .C(new_n5526), .Y(new_n5533));
  NAND3xp33_ASAP7_75t_L     g05277(.A(new_n5528), .B(new_n5533), .C(new_n5374), .Y(new_n5534));
  AOI21xp33_ASAP7_75t_L     g05278(.A1(new_n5526), .A2(new_n5522), .B(new_n5532), .Y(new_n5535));
  AOI211xp5_ASAP7_75t_L     g05279(.A1(new_n5273), .A2(new_n5375), .B(new_n5270), .C(new_n5527), .Y(new_n5536));
  OAI21xp33_ASAP7_75t_L     g05280(.A1(new_n5535), .A2(new_n5536), .B(new_n5373), .Y(new_n5537));
  NAND3xp33_ASAP7_75t_L     g05281(.A(new_n5366), .B(new_n5534), .C(new_n5537), .Y(new_n5538));
  A2O1A1O1Ixp25_ASAP7_75t_L g05282(.A1(new_n4892), .A2(new_n5060), .B(new_n5113), .C(new_n5276), .D(new_n5285), .Y(new_n5539));
  NOR3xp33_ASAP7_75t_L      g05283(.A(new_n5536), .B(new_n5373), .C(new_n5535), .Y(new_n5540));
  AOI21xp33_ASAP7_75t_L     g05284(.A1(new_n5528), .A2(new_n5533), .B(new_n5374), .Y(new_n5541));
  OAI21xp33_ASAP7_75t_L     g05285(.A1(new_n5540), .A2(new_n5541), .B(new_n5539), .Y(new_n5542));
  NAND2xp33_ASAP7_75t_L     g05286(.A(\b[31] ), .B(new_n651), .Y(new_n5543));
  OAI221xp5_ASAP7_75t_L     g05287(.A1(new_n580), .A2(new_n3565), .B1(new_n577), .B2(new_n3572), .C(new_n5543), .Y(new_n5544));
  AOI21xp33_ASAP7_75t_L     g05288(.A1(new_n584), .A2(\b[32] ), .B(new_n5544), .Y(new_n5545));
  NAND2xp33_ASAP7_75t_L     g05289(.A(\a[11] ), .B(new_n5545), .Y(new_n5546));
  A2O1A1Ixp33_ASAP7_75t_L   g05290(.A1(\b[32] ), .A2(new_n584), .B(new_n5544), .C(new_n574), .Y(new_n5547));
  AND2x2_ASAP7_75t_L        g05291(.A(new_n5547), .B(new_n5546), .Y(new_n5548));
  NAND3xp33_ASAP7_75t_L     g05292(.A(new_n5548), .B(new_n5542), .C(new_n5538), .Y(new_n5549));
  NOR3xp33_ASAP7_75t_L      g05293(.A(new_n5539), .B(new_n5540), .C(new_n5541), .Y(new_n5550));
  AOI21xp33_ASAP7_75t_L     g05294(.A1(new_n5537), .A2(new_n5534), .B(new_n5366), .Y(new_n5551));
  NAND2xp33_ASAP7_75t_L     g05295(.A(new_n5547), .B(new_n5546), .Y(new_n5552));
  OAI21xp33_ASAP7_75t_L     g05296(.A1(new_n5550), .A2(new_n5551), .B(new_n5552), .Y(new_n5553));
  AOI21xp33_ASAP7_75t_L     g05297(.A1(new_n5553), .A2(new_n5549), .B(new_n5365), .Y(new_n5554));
  NAND3xp33_ASAP7_75t_L     g05298(.A(new_n5281), .B(new_n5112), .C(new_n5286), .Y(new_n5555));
  OAI21xp33_ASAP7_75t_L     g05299(.A1(new_n5287), .A2(new_n5104), .B(new_n5555), .Y(new_n5556));
  NOR3xp33_ASAP7_75t_L      g05300(.A(new_n5551), .B(new_n5550), .C(new_n5552), .Y(new_n5557));
  AOI21xp33_ASAP7_75t_L     g05301(.A1(new_n5542), .A2(new_n5538), .B(new_n5548), .Y(new_n5558));
  NOR3xp33_ASAP7_75t_L      g05302(.A(new_n5556), .B(new_n5557), .C(new_n5558), .Y(new_n5559));
  OAI21xp33_ASAP7_75t_L     g05303(.A1(new_n5554), .A2(new_n5559), .B(new_n5363), .Y(new_n5560));
  NAND2xp33_ASAP7_75t_L     g05304(.A(new_n5362), .B(new_n5361), .Y(new_n5561));
  OAI21xp33_ASAP7_75t_L     g05305(.A1(new_n5557), .A2(new_n5558), .B(new_n5556), .Y(new_n5562));
  NAND3xp33_ASAP7_75t_L     g05306(.A(new_n5365), .B(new_n5549), .C(new_n5553), .Y(new_n5563));
  NAND3xp33_ASAP7_75t_L     g05307(.A(new_n5563), .B(new_n5562), .C(new_n5561), .Y(new_n5564));
  NAND2xp33_ASAP7_75t_L     g05308(.A(new_n5564), .B(new_n5560), .Y(new_n5565));
  O2A1O1Ixp33_ASAP7_75t_L   g05309(.A1(new_n5307), .A2(new_n5310), .B(new_n5357), .C(new_n5565), .Y(new_n5566));
  A2O1A1Ixp33_ASAP7_75t_L   g05310(.A1(new_n5301), .A2(new_n5304), .B(new_n5307), .C(new_n5357), .Y(new_n5567));
  AOI21xp33_ASAP7_75t_L     g05311(.A1(new_n5564), .A2(new_n5560), .B(new_n5567), .Y(new_n5568));
  OAI22xp33_ASAP7_75t_L     g05312(.A1(new_n5568), .A2(new_n5566), .B1(new_n5356), .B2(new_n5355), .Y(new_n5569));
  NOR2xp33_ASAP7_75t_L      g05313(.A(new_n5356), .B(new_n5355), .Y(new_n5570));
  NAND3xp33_ASAP7_75t_L     g05314(.A(new_n5567), .B(new_n5560), .C(new_n5564), .Y(new_n5571));
  OAI211xp5_ASAP7_75t_L     g05315(.A1(new_n5307), .A2(new_n5310), .B(new_n5565), .C(new_n5357), .Y(new_n5572));
  NAND3xp33_ASAP7_75t_L     g05316(.A(new_n5571), .B(new_n5572), .C(new_n5570), .Y(new_n5573));
  NAND2xp33_ASAP7_75t_L     g05317(.A(new_n5573), .B(new_n5569), .Y(new_n5574));
  A2O1A1Ixp33_ASAP7_75t_L   g05318(.A1(new_n5316), .A2(new_n5098), .B(new_n5350), .C(new_n5574), .Y(new_n5575));
  INVx1_ASAP7_75t_L         g05319(.A(new_n4838), .Y(new_n5576));
  OAI21xp33_ASAP7_75t_L     g05320(.A1(new_n5576), .A2(new_n4651), .B(new_n4842), .Y(new_n5577));
  INVx1_ASAP7_75t_L         g05321(.A(new_n5097), .Y(new_n5578));
  A2O1A1O1Ixp25_ASAP7_75t_L g05322(.A1(new_n5086), .A2(new_n5577), .B(new_n5578), .C(new_n5316), .D(new_n5350), .Y(new_n5579));
  NAND3xp33_ASAP7_75t_L     g05323(.A(new_n5579), .B(new_n5569), .C(new_n5573), .Y(new_n5580));
  NAND2xp33_ASAP7_75t_L     g05324(.A(new_n5580), .B(new_n5575), .Y(new_n5581));
  XOR2x2_ASAP7_75t_L        g05325(.A(new_n5349), .B(new_n5581), .Y(new_n5582));
  A2O1A1O1Ixp25_ASAP7_75t_L g05326(.A1(new_n5093), .A2(new_n4865), .B(new_n5091), .C(new_n5331), .D(new_n5332), .Y(new_n5583));
  XNOR2x2_ASAP7_75t_L       g05327(.A(new_n5583), .B(new_n5582), .Y(\f[42] ));
  OAI211xp5_ASAP7_75t_L     g05328(.A1(new_n5356), .A2(new_n5355), .B(new_n5571), .C(new_n5572), .Y(new_n5585));
  A2O1A1Ixp33_ASAP7_75t_L   g05329(.A1(new_n5569), .A2(new_n5573), .B(new_n5579), .C(new_n5585), .Y(new_n5586));
  NAND2xp33_ASAP7_75t_L     g05330(.A(\b[39] ), .B(new_n347), .Y(new_n5587));
  NAND2xp33_ASAP7_75t_L     g05331(.A(new_n341), .B(new_n4876), .Y(new_n5588));
  AOI22xp33_ASAP7_75t_L     g05332(.A1(new_n344), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n370), .Y(new_n5589));
  NAND4xp25_ASAP7_75t_L     g05333(.A(new_n5588), .B(\a[5] ), .C(new_n5587), .D(new_n5589), .Y(new_n5590));
  NAND2xp33_ASAP7_75t_L     g05334(.A(new_n5589), .B(new_n5588), .Y(new_n5591));
  A2O1A1Ixp33_ASAP7_75t_L   g05335(.A1(\b[39] ), .A2(new_n347), .B(new_n5591), .C(new_n338), .Y(new_n5592));
  NAND2xp33_ASAP7_75t_L     g05336(.A(new_n5590), .B(new_n5592), .Y(new_n5593));
  INVx1_ASAP7_75t_L         g05337(.A(new_n5593), .Y(new_n5594));
  INVx1_ASAP7_75t_L         g05338(.A(new_n5564), .Y(new_n5595));
  OAI21xp33_ASAP7_75t_L     g05339(.A1(new_n5541), .A2(new_n5539), .B(new_n5534), .Y(new_n5596));
  NAND3xp33_ASAP7_75t_L     g05340(.A(new_n5510), .B(new_n5514), .C(new_n5525), .Y(new_n5597));
  A2O1A1Ixp33_ASAP7_75t_L   g05341(.A1(new_n5522), .A2(new_n5526), .B(new_n5532), .C(new_n5597), .Y(new_n5598));
  AOI22xp33_ASAP7_75t_L     g05342(.A1(new_n1076), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n1253), .Y(new_n5599));
  INVx1_ASAP7_75t_L         g05343(.A(new_n5599), .Y(new_n5600));
  AOI221xp5_ASAP7_75t_L     g05344(.A1(\b[27] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n4237), .C(new_n5600), .Y(new_n5601));
  XNOR2x2_ASAP7_75t_L       g05345(.A(new_n1071), .B(new_n5601), .Y(new_n5602));
  NAND2xp33_ASAP7_75t_L     g05346(.A(new_n5442), .B(new_n5437), .Y(new_n5603));
  MAJIxp5_ASAP7_75t_L       g05347(.A(new_n5449), .B(new_n5386), .C(new_n5603), .Y(new_n5604));
  AOI22xp33_ASAP7_75t_L     g05348(.A1(new_n3029), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n3258), .Y(new_n5605));
  OAI221xp5_ASAP7_75t_L     g05349(.A1(new_n3024), .A2(new_n760), .B1(new_n3256), .B2(new_n790), .C(new_n5605), .Y(new_n5606));
  XNOR2x2_ASAP7_75t_L       g05350(.A(\a[32] ), .B(new_n5606), .Y(new_n5607));
  A2O1A1O1Ixp25_ASAP7_75t_L g05351(.A1(new_n5189), .A2(new_n5196), .B(new_n5387), .C(new_n5439), .D(new_n5435), .Y(new_n5608));
  NOR3xp33_ASAP7_75t_L      g05352(.A(new_n5169), .B(new_n5396), .C(new_n5388), .Y(new_n5609));
  NAND2xp33_ASAP7_75t_L     g05353(.A(\b[3] ), .B(new_n4924), .Y(new_n5610));
  NAND2xp33_ASAP7_75t_L     g05354(.A(new_n4917), .B(new_n329), .Y(new_n5611));
  AOI22xp33_ASAP7_75t_L     g05355(.A1(new_n4920), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n5167), .Y(new_n5612));
  NAND4xp25_ASAP7_75t_L     g05356(.A(new_n5611), .B(\a[41] ), .C(new_n5610), .D(new_n5612), .Y(new_n5613));
  AOI31xp33_ASAP7_75t_L     g05357(.A1(new_n5611), .A2(new_n5610), .A3(new_n5612), .B(\a[41] ), .Y(new_n5614));
  INVx1_ASAP7_75t_L         g05358(.A(new_n5614), .Y(new_n5615));
  NAND2xp33_ASAP7_75t_L     g05359(.A(\a[44] ), .B(new_n5393), .Y(new_n5616));
  INVx1_ASAP7_75t_L         g05360(.A(\a[43] ), .Y(new_n5617));
  NAND2xp33_ASAP7_75t_L     g05361(.A(\a[44] ), .B(new_n5617), .Y(new_n5618));
  INVx1_ASAP7_75t_L         g05362(.A(\a[44] ), .Y(new_n5619));
  NAND2xp33_ASAP7_75t_L     g05363(.A(\a[43] ), .B(new_n5619), .Y(new_n5620));
  AOI21xp33_ASAP7_75t_L     g05364(.A1(new_n5620), .A2(new_n5618), .B(new_n5392), .Y(new_n5621));
  NAND2xp33_ASAP7_75t_L     g05365(.A(new_n269), .B(new_n5621), .Y(new_n5622));
  NAND2xp33_ASAP7_75t_L     g05366(.A(new_n5620), .B(new_n5618), .Y(new_n5623));
  NOR2xp33_ASAP7_75t_L      g05367(.A(new_n5623), .B(new_n5392), .Y(new_n5624));
  NAND2xp33_ASAP7_75t_L     g05368(.A(\b[1] ), .B(new_n5624), .Y(new_n5625));
  NAND2xp33_ASAP7_75t_L     g05369(.A(new_n5391), .B(new_n5390), .Y(new_n5626));
  XNOR2x2_ASAP7_75t_L       g05370(.A(\a[43] ), .B(\a[42] ), .Y(new_n5627));
  NOR2xp33_ASAP7_75t_L      g05371(.A(new_n5627), .B(new_n5626), .Y(new_n5628));
  NAND2xp33_ASAP7_75t_L     g05372(.A(\b[0] ), .B(new_n5628), .Y(new_n5629));
  NAND3xp33_ASAP7_75t_L     g05373(.A(new_n5622), .B(new_n5625), .C(new_n5629), .Y(new_n5630));
  XOR2x2_ASAP7_75t_L        g05374(.A(new_n5616), .B(new_n5630), .Y(new_n5631));
  NAND3xp33_ASAP7_75t_L     g05375(.A(new_n5615), .B(new_n5631), .C(new_n5613), .Y(new_n5632));
  INVx1_ASAP7_75t_L         g05376(.A(new_n5613), .Y(new_n5633));
  XNOR2x2_ASAP7_75t_L       g05377(.A(new_n5616), .B(new_n5630), .Y(new_n5634));
  OAI21xp33_ASAP7_75t_L     g05378(.A1(new_n5614), .A2(new_n5633), .B(new_n5634), .Y(new_n5635));
  OAI211xp5_ASAP7_75t_L     g05379(.A1(new_n5609), .A2(new_n5412), .B(new_n5632), .C(new_n5635), .Y(new_n5636));
  INVx1_ASAP7_75t_L         g05380(.A(new_n5609), .Y(new_n5637));
  NOR3xp33_ASAP7_75t_L      g05381(.A(new_n5634), .B(new_n5633), .C(new_n5614), .Y(new_n5638));
  AOI21xp33_ASAP7_75t_L     g05382(.A1(new_n5615), .A2(new_n5613), .B(new_n5631), .Y(new_n5639));
  OAI211xp5_ASAP7_75t_L     g05383(.A1(new_n5638), .A2(new_n5639), .B(new_n5637), .C(new_n5403), .Y(new_n5640));
  NAND2xp33_ASAP7_75t_L     g05384(.A(\b[6] ), .B(new_n4285), .Y(new_n5641));
  NAND2xp33_ASAP7_75t_L     g05385(.A(new_n4274), .B(new_n2084), .Y(new_n5642));
  AOI22xp33_ASAP7_75t_L     g05386(.A1(new_n4283), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n4512), .Y(new_n5643));
  NAND4xp25_ASAP7_75t_L     g05387(.A(new_n5642), .B(\a[38] ), .C(new_n5641), .D(new_n5643), .Y(new_n5644));
  OAI211xp5_ASAP7_75t_L     g05388(.A1(new_n4499), .A2(new_n425), .B(new_n5641), .C(new_n5643), .Y(new_n5645));
  NAND2xp33_ASAP7_75t_L     g05389(.A(new_n4268), .B(new_n5645), .Y(new_n5646));
  NAND4xp25_ASAP7_75t_L     g05390(.A(new_n5640), .B(new_n5644), .C(new_n5646), .D(new_n5636), .Y(new_n5647));
  AO22x1_ASAP7_75t_L        g05391(.A1(new_n5646), .A2(new_n5644), .B1(new_n5636), .B2(new_n5640), .Y(new_n5648));
  AND2x2_ASAP7_75t_L        g05392(.A(new_n5647), .B(new_n5648), .Y(new_n5649));
  AOI211xp5_ASAP7_75t_L     g05393(.A1(new_n5410), .A2(new_n5408), .B(new_n5412), .C(new_n5413), .Y(new_n5650));
  AOI21xp33_ASAP7_75t_L     g05394(.A1(new_n5432), .A2(new_n5421), .B(new_n5650), .Y(new_n5651));
  NAND2xp33_ASAP7_75t_L     g05395(.A(new_n5651), .B(new_n5649), .Y(new_n5652));
  NAND2xp33_ASAP7_75t_L     g05396(.A(new_n5647), .B(new_n5648), .Y(new_n5653));
  A2O1A1Ixp33_ASAP7_75t_L   g05397(.A1(new_n5421), .A2(new_n5432), .B(new_n5650), .C(new_n5653), .Y(new_n5654));
  AOI22xp33_ASAP7_75t_L     g05398(.A1(new_n3633), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n3858), .Y(new_n5655));
  OAI221xp5_ASAP7_75t_L     g05399(.A1(new_n3853), .A2(new_n540), .B1(new_n3856), .B2(new_n624), .C(new_n5655), .Y(new_n5656));
  XNOR2x2_ASAP7_75t_L       g05400(.A(\a[35] ), .B(new_n5656), .Y(new_n5657));
  INVx1_ASAP7_75t_L         g05401(.A(new_n5657), .Y(new_n5658));
  AOI21xp33_ASAP7_75t_L     g05402(.A1(new_n5652), .A2(new_n5654), .B(new_n5658), .Y(new_n5659));
  AND3x1_ASAP7_75t_L        g05403(.A(new_n5652), .B(new_n5658), .C(new_n5654), .Y(new_n5660));
  OA21x2_ASAP7_75t_L        g05404(.A1(new_n5659), .A2(new_n5660), .B(new_n5608), .Y(new_n5661));
  NOR3xp33_ASAP7_75t_L      g05405(.A(new_n5660), .B(new_n5608), .C(new_n5659), .Y(new_n5662));
  OAI21xp33_ASAP7_75t_L     g05406(.A1(new_n5662), .A2(new_n5661), .B(new_n5607), .Y(new_n5663));
  OR3x1_ASAP7_75t_L         g05407(.A(new_n5661), .B(new_n5607), .C(new_n5662), .Y(new_n5664));
  NAND3xp33_ASAP7_75t_L     g05408(.A(new_n5604), .B(new_n5663), .C(new_n5664), .Y(new_n5665));
  NOR2xp33_ASAP7_75t_L      g05409(.A(new_n5446), .B(new_n5445), .Y(new_n5666));
  MAJIxp5_ASAP7_75t_L       g05410(.A(new_n5382), .B(new_n5444), .C(new_n5666), .Y(new_n5667));
  OA21x2_ASAP7_75t_L        g05411(.A1(new_n5662), .A2(new_n5661), .B(new_n5607), .Y(new_n5668));
  NOR3xp33_ASAP7_75t_L      g05412(.A(new_n5661), .B(new_n5662), .C(new_n5607), .Y(new_n5669));
  OAI21xp33_ASAP7_75t_L     g05413(.A1(new_n5668), .A2(new_n5669), .B(new_n5667), .Y(new_n5670));
  AOI22xp33_ASAP7_75t_L     g05414(.A1(new_n2552), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n2736), .Y(new_n5671));
  OAI221xp5_ASAP7_75t_L     g05415(.A1(new_n2547), .A2(new_n942), .B1(new_n2734), .B2(new_n1035), .C(new_n5671), .Y(new_n5672));
  XNOR2x2_ASAP7_75t_L       g05416(.A(\a[29] ), .B(new_n5672), .Y(new_n5673));
  NAND3xp33_ASAP7_75t_L     g05417(.A(new_n5665), .B(new_n5670), .C(new_n5673), .Y(new_n5674));
  NOR3xp33_ASAP7_75t_L      g05418(.A(new_n5667), .B(new_n5668), .C(new_n5669), .Y(new_n5675));
  AOI21xp33_ASAP7_75t_L     g05419(.A1(new_n5664), .A2(new_n5663), .B(new_n5604), .Y(new_n5676));
  INVx1_ASAP7_75t_L         g05420(.A(new_n5673), .Y(new_n5677));
  OAI21xp33_ASAP7_75t_L     g05421(.A1(new_n5676), .A2(new_n5675), .B(new_n5677), .Y(new_n5678));
  NOR2xp33_ASAP7_75t_L      g05422(.A(new_n5454), .B(new_n5455), .Y(new_n5679));
  MAJIxp5_ASAP7_75t_L       g05423(.A(new_n5377), .B(new_n5380), .C(new_n5679), .Y(new_n5680));
  NAND3xp33_ASAP7_75t_L     g05424(.A(new_n5680), .B(new_n5678), .C(new_n5674), .Y(new_n5681));
  NOR3xp33_ASAP7_75t_L      g05425(.A(new_n5675), .B(new_n5676), .C(new_n5677), .Y(new_n5682));
  AOI21xp33_ASAP7_75t_L     g05426(.A1(new_n5665), .A2(new_n5670), .B(new_n5673), .Y(new_n5683));
  NAND2xp33_ASAP7_75t_L     g05427(.A(new_n5448), .B(new_n5452), .Y(new_n5684));
  MAJIxp5_ASAP7_75t_L       g05428(.A(new_n5458), .B(new_n5381), .C(new_n5684), .Y(new_n5685));
  OAI21xp33_ASAP7_75t_L     g05429(.A1(new_n5682), .A2(new_n5683), .B(new_n5685), .Y(new_n5686));
  AOI22xp33_ASAP7_75t_L     g05430(.A1(new_n2114), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n2259), .Y(new_n5687));
  OAI221xp5_ASAP7_75t_L     g05431(.A1(new_n2109), .A2(new_n1313), .B1(new_n2257), .B2(new_n1438), .C(new_n5687), .Y(new_n5688));
  XNOR2x2_ASAP7_75t_L       g05432(.A(\a[26] ), .B(new_n5688), .Y(new_n5689));
  NAND3xp33_ASAP7_75t_L     g05433(.A(new_n5681), .B(new_n5689), .C(new_n5686), .Y(new_n5690));
  AOI21xp33_ASAP7_75t_L     g05434(.A1(new_n5681), .A2(new_n5686), .B(new_n5689), .Y(new_n5691));
  INVx1_ASAP7_75t_L         g05435(.A(new_n5691), .Y(new_n5692));
  A2O1A1O1Ixp25_ASAP7_75t_L g05436(.A1(new_n5218), .A2(new_n5376), .B(new_n5217), .C(new_n5477), .D(new_n5468), .Y(new_n5693));
  NAND3xp33_ASAP7_75t_L     g05437(.A(new_n5693), .B(new_n5692), .C(new_n5690), .Y(new_n5694));
  AND3x1_ASAP7_75t_L        g05438(.A(new_n5681), .B(new_n5689), .C(new_n5686), .Y(new_n5695));
  OAI21xp33_ASAP7_75t_L     g05439(.A1(new_n5472), .A2(new_n5475), .B(new_n5476), .Y(new_n5696));
  OAI21xp33_ASAP7_75t_L     g05440(.A1(new_n5695), .A2(new_n5691), .B(new_n5696), .Y(new_n5697));
  NAND2xp33_ASAP7_75t_L     g05441(.A(\b[21] ), .B(new_n1706), .Y(new_n5698));
  NAND2xp33_ASAP7_75t_L     g05442(.A(new_n1695), .B(new_n3728), .Y(new_n5699));
  AOI22xp33_ASAP7_75t_L     g05443(.A1(new_n1704), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1837), .Y(new_n5700));
  NAND4xp25_ASAP7_75t_L     g05444(.A(new_n5699), .B(\a[23] ), .C(new_n5698), .D(new_n5700), .Y(new_n5701));
  OAI21xp33_ASAP7_75t_L     g05445(.A1(new_n1827), .A2(new_n1780), .B(new_n5700), .Y(new_n5702));
  A2O1A1Ixp33_ASAP7_75t_L   g05446(.A1(\b[21] ), .A2(new_n1706), .B(new_n5702), .C(new_n1689), .Y(new_n5703));
  NAND2xp33_ASAP7_75t_L     g05447(.A(new_n5701), .B(new_n5703), .Y(new_n5704));
  INVx1_ASAP7_75t_L         g05448(.A(new_n5704), .Y(new_n5705));
  NAND3xp33_ASAP7_75t_L     g05449(.A(new_n5694), .B(new_n5705), .C(new_n5697), .Y(new_n5706));
  NOR3xp33_ASAP7_75t_L      g05450(.A(new_n5696), .B(new_n5691), .C(new_n5695), .Y(new_n5707));
  AOI21xp33_ASAP7_75t_L     g05451(.A1(new_n5692), .A2(new_n5690), .B(new_n5693), .Y(new_n5708));
  OAI21xp33_ASAP7_75t_L     g05452(.A1(new_n5707), .A2(new_n5708), .B(new_n5704), .Y(new_n5709));
  NAND2xp33_ASAP7_75t_L     g05453(.A(new_n5706), .B(new_n5709), .Y(new_n5710));
  NOR3xp33_ASAP7_75t_L      g05454(.A(new_n5488), .B(new_n5487), .C(new_n5485), .Y(new_n5711));
  INVx1_ASAP7_75t_L         g05455(.A(new_n5711), .Y(new_n5712));
  OAI21xp33_ASAP7_75t_L     g05456(.A1(new_n5498), .A2(new_n5496), .B(new_n5712), .Y(new_n5713));
  NOR2xp33_ASAP7_75t_L      g05457(.A(new_n5710), .B(new_n5713), .Y(new_n5714));
  NOR3xp33_ASAP7_75t_L      g05458(.A(new_n5708), .B(new_n5707), .C(new_n5704), .Y(new_n5715));
  AOI21xp33_ASAP7_75t_L     g05459(.A1(new_n5694), .A2(new_n5697), .B(new_n5705), .Y(new_n5716));
  NOR2xp33_ASAP7_75t_L      g05460(.A(new_n5715), .B(new_n5716), .Y(new_n5717));
  AOI21xp33_ASAP7_75t_L     g05461(.A1(new_n5506), .A2(new_n5712), .B(new_n5717), .Y(new_n5718));
  AOI22xp33_ASAP7_75t_L     g05462(.A1(new_n1360), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n1581), .Y(new_n5719));
  INVx1_ASAP7_75t_L         g05463(.A(new_n5719), .Y(new_n5720));
  AOI221xp5_ASAP7_75t_L     g05464(.A1(\b[24] ), .A2(new_n1362), .B1(new_n1365), .B2(new_n2648), .C(new_n5720), .Y(new_n5721));
  XNOR2x2_ASAP7_75t_L       g05465(.A(\a[20] ), .B(new_n5721), .Y(new_n5722));
  NOR3xp33_ASAP7_75t_L      g05466(.A(new_n5718), .B(new_n5714), .C(new_n5722), .Y(new_n5723));
  A2O1A1O1Ixp25_ASAP7_75t_L g05467(.A1(new_n5242), .A2(new_n5240), .B(new_n5492), .C(new_n5491), .D(new_n5711), .Y(new_n5724));
  NAND2xp33_ASAP7_75t_L     g05468(.A(new_n5717), .B(new_n5724), .Y(new_n5725));
  NAND2xp33_ASAP7_75t_L     g05469(.A(new_n5710), .B(new_n5713), .Y(new_n5726));
  XNOR2x2_ASAP7_75t_L       g05470(.A(new_n1356), .B(new_n5721), .Y(new_n5727));
  AOI21xp33_ASAP7_75t_L     g05471(.A1(new_n5725), .A2(new_n5726), .B(new_n5727), .Y(new_n5728));
  OAI31xp33_ASAP7_75t_L     g05472(.A1(new_n5513), .A2(new_n5511), .A3(new_n5261), .B(new_n5508), .Y(new_n5729));
  OAI21xp33_ASAP7_75t_L     g05473(.A1(new_n5723), .A2(new_n5728), .B(new_n5729), .Y(new_n5730));
  NAND3xp33_ASAP7_75t_L     g05474(.A(new_n5725), .B(new_n5726), .C(new_n5727), .Y(new_n5731));
  OAI21xp33_ASAP7_75t_L     g05475(.A1(new_n5714), .A2(new_n5718), .B(new_n5722), .Y(new_n5732));
  NAND4xp25_ASAP7_75t_L     g05476(.A(new_n5510), .B(new_n5731), .C(new_n5732), .D(new_n5508), .Y(new_n5733));
  AOI21xp33_ASAP7_75t_L     g05477(.A1(new_n5733), .A2(new_n5730), .B(new_n5602), .Y(new_n5734));
  XNOR2x2_ASAP7_75t_L       g05478(.A(\a[17] ), .B(new_n5601), .Y(new_n5735));
  AOI31xp33_ASAP7_75t_L     g05479(.A1(new_n5509), .A2(new_n5504), .A3(new_n5254), .B(new_n5512), .Y(new_n5736));
  AOI21xp33_ASAP7_75t_L     g05480(.A1(new_n5732), .A2(new_n5731), .B(new_n5736), .Y(new_n5737));
  NOR3xp33_ASAP7_75t_L      g05481(.A(new_n5729), .B(new_n5728), .C(new_n5723), .Y(new_n5738));
  NOR3xp33_ASAP7_75t_L      g05482(.A(new_n5737), .B(new_n5738), .C(new_n5735), .Y(new_n5739));
  NOR2xp33_ASAP7_75t_L      g05483(.A(new_n5734), .B(new_n5739), .Y(new_n5740));
  NAND2xp33_ASAP7_75t_L     g05484(.A(new_n5598), .B(new_n5740), .Y(new_n5741));
  INVx1_ASAP7_75t_L         g05485(.A(new_n5597), .Y(new_n5742));
  A2O1A1O1Ixp25_ASAP7_75t_L g05486(.A1(new_n5273), .A2(new_n5274), .B(new_n5270), .C(new_n5527), .D(new_n5742), .Y(new_n5743));
  OAI21xp33_ASAP7_75t_L     g05487(.A1(new_n5738), .A2(new_n5737), .B(new_n5735), .Y(new_n5744));
  NAND3xp33_ASAP7_75t_L     g05488(.A(new_n5733), .B(new_n5602), .C(new_n5730), .Y(new_n5745));
  NAND2xp33_ASAP7_75t_L     g05489(.A(new_n5745), .B(new_n5744), .Y(new_n5746));
  NAND2xp33_ASAP7_75t_L     g05490(.A(new_n5746), .B(new_n5743), .Y(new_n5747));
  AOI22xp33_ASAP7_75t_L     g05491(.A1(new_n811), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n900), .Y(new_n5748));
  OAI221xp5_ASAP7_75t_L     g05492(.A1(new_n904), .A2(new_n2982), .B1(new_n898), .B2(new_n3187), .C(new_n5748), .Y(new_n5749));
  XNOR2x2_ASAP7_75t_L       g05493(.A(\a[14] ), .B(new_n5749), .Y(new_n5750));
  NAND3xp33_ASAP7_75t_L     g05494(.A(new_n5747), .B(new_n5741), .C(new_n5750), .Y(new_n5751));
  NOR2xp33_ASAP7_75t_L      g05495(.A(new_n5746), .B(new_n5743), .Y(new_n5752));
  NOR2xp33_ASAP7_75t_L      g05496(.A(new_n5598), .B(new_n5740), .Y(new_n5753));
  INVx1_ASAP7_75t_L         g05497(.A(new_n5750), .Y(new_n5754));
  OAI21xp33_ASAP7_75t_L     g05498(.A1(new_n5753), .A2(new_n5752), .B(new_n5754), .Y(new_n5755));
  NAND3xp33_ASAP7_75t_L     g05499(.A(new_n5596), .B(new_n5751), .C(new_n5755), .Y(new_n5756));
  A2O1A1O1Ixp25_ASAP7_75t_L g05500(.A1(new_n5276), .A2(new_n5115), .B(new_n5285), .C(new_n5537), .D(new_n5540), .Y(new_n5757));
  NAND2xp33_ASAP7_75t_L     g05501(.A(new_n5751), .B(new_n5755), .Y(new_n5758));
  NAND2xp33_ASAP7_75t_L     g05502(.A(new_n5757), .B(new_n5758), .Y(new_n5759));
  AOI22xp33_ASAP7_75t_L     g05503(.A1(\b[32] ), .A2(new_n651), .B1(\b[34] ), .B2(new_n581), .Y(new_n5760));
  OAI221xp5_ASAP7_75t_L     g05504(.A1(new_n821), .A2(new_n3565), .B1(new_n577), .B2(new_n3591), .C(new_n5760), .Y(new_n5761));
  XNOR2x2_ASAP7_75t_L       g05505(.A(\a[11] ), .B(new_n5761), .Y(new_n5762));
  NAND3xp33_ASAP7_75t_L     g05506(.A(new_n5759), .B(new_n5756), .C(new_n5762), .Y(new_n5763));
  O2A1O1Ixp33_ASAP7_75t_L   g05507(.A1(new_n5539), .A2(new_n5541), .B(new_n5534), .C(new_n5758), .Y(new_n5764));
  AOI21xp33_ASAP7_75t_L     g05508(.A1(new_n5755), .A2(new_n5751), .B(new_n5596), .Y(new_n5765));
  INVx1_ASAP7_75t_L         g05509(.A(new_n5762), .Y(new_n5766));
  OAI21xp33_ASAP7_75t_L     g05510(.A1(new_n5765), .A2(new_n5764), .B(new_n5766), .Y(new_n5767));
  NOR2xp33_ASAP7_75t_L      g05511(.A(new_n5550), .B(new_n5551), .Y(new_n5768));
  MAJIxp5_ASAP7_75t_L       g05512(.A(new_n5556), .B(new_n5552), .C(new_n5768), .Y(new_n5769));
  NAND3xp33_ASAP7_75t_L     g05513(.A(new_n5769), .B(new_n5767), .C(new_n5763), .Y(new_n5770));
  NOR3xp33_ASAP7_75t_L      g05514(.A(new_n5764), .B(new_n5766), .C(new_n5765), .Y(new_n5771));
  AOI21xp33_ASAP7_75t_L     g05515(.A1(new_n5759), .A2(new_n5756), .B(new_n5762), .Y(new_n5772));
  NAND2xp33_ASAP7_75t_L     g05516(.A(new_n5542), .B(new_n5538), .Y(new_n5773));
  MAJIxp5_ASAP7_75t_L       g05517(.A(new_n5365), .B(new_n5548), .C(new_n5773), .Y(new_n5774));
  OAI21xp33_ASAP7_75t_L     g05518(.A1(new_n5772), .A2(new_n5771), .B(new_n5774), .Y(new_n5775));
  AOI22xp33_ASAP7_75t_L     g05519(.A1(new_n444), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n471), .Y(new_n5776));
  OAI221xp5_ASAP7_75t_L     g05520(.A1(new_n468), .A2(new_n4216), .B1(new_n469), .B2(new_n4431), .C(new_n5776), .Y(new_n5777));
  XNOR2x2_ASAP7_75t_L       g05521(.A(\a[8] ), .B(new_n5777), .Y(new_n5778));
  INVx1_ASAP7_75t_L         g05522(.A(new_n5778), .Y(new_n5779));
  AOI21xp33_ASAP7_75t_L     g05523(.A1(new_n5770), .A2(new_n5775), .B(new_n5779), .Y(new_n5780));
  NOR3xp33_ASAP7_75t_L      g05524(.A(new_n5774), .B(new_n5772), .C(new_n5771), .Y(new_n5781));
  AOI21xp33_ASAP7_75t_L     g05525(.A1(new_n5767), .A2(new_n5763), .B(new_n5769), .Y(new_n5782));
  NOR3xp33_ASAP7_75t_L      g05526(.A(new_n5781), .B(new_n5778), .C(new_n5782), .Y(new_n5783));
  NOR2xp33_ASAP7_75t_L      g05527(.A(new_n5780), .B(new_n5783), .Y(new_n5784));
  NOR3xp33_ASAP7_75t_L      g05528(.A(new_n5784), .B(new_n5566), .C(new_n5595), .Y(new_n5785));
  INVx1_ASAP7_75t_L         g05529(.A(new_n5567), .Y(new_n5786));
  OAI21xp33_ASAP7_75t_L     g05530(.A1(new_n5782), .A2(new_n5781), .B(new_n5778), .Y(new_n5787));
  NAND3xp33_ASAP7_75t_L     g05531(.A(new_n5770), .B(new_n5775), .C(new_n5779), .Y(new_n5788));
  NAND2xp33_ASAP7_75t_L     g05532(.A(new_n5788), .B(new_n5787), .Y(new_n5789));
  O2A1O1Ixp33_ASAP7_75t_L   g05533(.A1(new_n5565), .A2(new_n5786), .B(new_n5564), .C(new_n5789), .Y(new_n5790));
  OAI21xp33_ASAP7_75t_L     g05534(.A1(new_n5790), .A2(new_n5785), .B(new_n5594), .Y(new_n5791));
  INVx1_ASAP7_75t_L         g05535(.A(new_n5357), .Y(new_n5792));
  A2O1A1O1Ixp25_ASAP7_75t_L g05536(.A1(new_n5305), .A2(new_n5314), .B(new_n5792), .C(new_n5560), .D(new_n5595), .Y(new_n5793));
  NAND2xp33_ASAP7_75t_L     g05537(.A(new_n5793), .B(new_n5789), .Y(new_n5794));
  A2O1A1Ixp33_ASAP7_75t_L   g05538(.A1(new_n5560), .A2(new_n5567), .B(new_n5595), .C(new_n5784), .Y(new_n5795));
  NAND3xp33_ASAP7_75t_L     g05539(.A(new_n5795), .B(new_n5794), .C(new_n5593), .Y(new_n5796));
  NAND3xp33_ASAP7_75t_L     g05540(.A(new_n5586), .B(new_n5791), .C(new_n5796), .Y(new_n5797));
  INVx1_ASAP7_75t_L         g05541(.A(new_n5585), .Y(new_n5798));
  A2O1A1O1Ixp25_ASAP7_75t_L g05542(.A1(new_n5098), .A2(new_n5316), .B(new_n5350), .C(new_n5574), .D(new_n5798), .Y(new_n5799));
  NAND2xp33_ASAP7_75t_L     g05543(.A(new_n5796), .B(new_n5791), .Y(new_n5800));
  NAND2xp33_ASAP7_75t_L     g05544(.A(new_n5800), .B(new_n5799), .Y(new_n5801));
  NAND2xp33_ASAP7_75t_L     g05545(.A(\b[42] ), .B(new_n272), .Y(new_n5802));
  INVx1_ASAP7_75t_L         g05546(.A(new_n5339), .Y(new_n5803));
  NOR2xp33_ASAP7_75t_L      g05547(.A(\b[42] ), .B(\b[43] ), .Y(new_n5804));
  INVx1_ASAP7_75t_L         g05548(.A(\b[43] ), .Y(new_n5805));
  NOR2xp33_ASAP7_75t_L      g05549(.A(new_n5338), .B(new_n5805), .Y(new_n5806));
  NOR2xp33_ASAP7_75t_L      g05550(.A(new_n5804), .B(new_n5806), .Y(new_n5807));
  INVx1_ASAP7_75t_L         g05551(.A(new_n5807), .Y(new_n5808));
  A2O1A1O1Ixp25_ASAP7_75t_L g05552(.A1(new_n5336), .A2(new_n5324), .B(new_n5337), .C(new_n5803), .D(new_n5808), .Y(new_n5809));
  A2O1A1Ixp33_ASAP7_75t_L   g05553(.A1(new_n5324), .A2(new_n5336), .B(new_n5337), .C(new_n5803), .Y(new_n5810));
  NOR2xp33_ASAP7_75t_L      g05554(.A(new_n5807), .B(new_n5810), .Y(new_n5811));
  NOR2xp33_ASAP7_75t_L      g05555(.A(new_n5809), .B(new_n5811), .Y(new_n5812));
  NAND2xp33_ASAP7_75t_L     g05556(.A(new_n267), .B(new_n5812), .Y(new_n5813));
  AOI22xp33_ASAP7_75t_L     g05557(.A1(\b[41] ), .A2(new_n282), .B1(\b[43] ), .B2(new_n303), .Y(new_n5814));
  AND4x1_ASAP7_75t_L        g05558(.A(new_n5814), .B(new_n5813), .C(new_n5802), .D(\a[2] ), .Y(new_n5815));
  AOI31xp33_ASAP7_75t_L     g05559(.A1(new_n5813), .A2(new_n5802), .A3(new_n5814), .B(\a[2] ), .Y(new_n5816));
  NOR2xp33_ASAP7_75t_L      g05560(.A(new_n5816), .B(new_n5815), .Y(new_n5817));
  NAND3xp33_ASAP7_75t_L     g05561(.A(new_n5801), .B(new_n5797), .C(new_n5817), .Y(new_n5818));
  NOR2xp33_ASAP7_75t_L      g05562(.A(new_n5800), .B(new_n5799), .Y(new_n5819));
  AOI21xp33_ASAP7_75t_L     g05563(.A1(new_n5796), .A2(new_n5791), .B(new_n5586), .Y(new_n5820));
  INVx1_ASAP7_75t_L         g05564(.A(new_n5817), .Y(new_n5821));
  OAI21xp33_ASAP7_75t_L     g05565(.A1(new_n5820), .A2(new_n5819), .B(new_n5821), .Y(new_n5822));
  NAND2xp33_ASAP7_75t_L     g05566(.A(new_n5818), .B(new_n5822), .Y(new_n5823));
  MAJIxp5_ASAP7_75t_L       g05567(.A(new_n5583), .B(new_n5349), .C(new_n5581), .Y(new_n5824));
  XOR2x2_ASAP7_75t_L        g05568(.A(new_n5824), .B(new_n5823), .Y(\f[43] ));
  NOR3xp33_ASAP7_75t_L      g05569(.A(new_n5819), .B(new_n5820), .C(new_n5817), .Y(new_n5826));
  AOI21xp33_ASAP7_75t_L     g05570(.A1(new_n5823), .A2(new_n5824), .B(new_n5826), .Y(new_n5827));
  NOR2xp33_ASAP7_75t_L      g05571(.A(\b[43] ), .B(\b[44] ), .Y(new_n5828));
  INVx1_ASAP7_75t_L         g05572(.A(\b[44] ), .Y(new_n5829));
  NOR2xp33_ASAP7_75t_L      g05573(.A(new_n5805), .B(new_n5829), .Y(new_n5830));
  NOR2xp33_ASAP7_75t_L      g05574(.A(new_n5828), .B(new_n5830), .Y(new_n5831));
  A2O1A1Ixp33_ASAP7_75t_L   g05575(.A1(new_n5810), .A2(new_n5807), .B(new_n5806), .C(new_n5831), .Y(new_n5832));
  O2A1O1Ixp33_ASAP7_75t_L   g05576(.A1(new_n5339), .A2(new_n5342), .B(new_n5807), .C(new_n5806), .Y(new_n5833));
  OAI21xp33_ASAP7_75t_L     g05577(.A1(new_n5828), .A2(new_n5830), .B(new_n5833), .Y(new_n5834));
  NAND2xp33_ASAP7_75t_L     g05578(.A(new_n5832), .B(new_n5834), .Y(new_n5835));
  AOI22xp33_ASAP7_75t_L     g05579(.A1(\b[42] ), .A2(new_n282), .B1(\b[44] ), .B2(new_n303), .Y(new_n5836));
  OAI221xp5_ASAP7_75t_L     g05580(.A1(new_n291), .A2(new_n5805), .B1(new_n268), .B2(new_n5835), .C(new_n5836), .Y(new_n5837));
  XNOR2x2_ASAP7_75t_L       g05581(.A(\a[2] ), .B(new_n5837), .Y(new_n5838));
  AO21x2_ASAP7_75t_L        g05582(.A1(new_n5316), .A2(new_n5098), .B(new_n5350), .Y(new_n5839));
  NOR3xp33_ASAP7_75t_L      g05583(.A(new_n5785), .B(new_n5790), .C(new_n5594), .Y(new_n5840));
  A2O1A1O1Ixp25_ASAP7_75t_L g05584(.A1(new_n5574), .A2(new_n5839), .B(new_n5798), .C(new_n5791), .D(new_n5840), .Y(new_n5841));
  NAND2xp33_ASAP7_75t_L     g05585(.A(\b[40] ), .B(new_n347), .Y(new_n5842));
  NAND3xp33_ASAP7_75t_L     g05586(.A(new_n5326), .B(new_n5324), .C(new_n341), .Y(new_n5843));
  AOI22xp33_ASAP7_75t_L     g05587(.A1(new_n344), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n370), .Y(new_n5844));
  AND4x1_ASAP7_75t_L        g05588(.A(new_n5844), .B(new_n5843), .C(new_n5842), .D(\a[5] ), .Y(new_n5845));
  AOI31xp33_ASAP7_75t_L     g05589(.A1(new_n5843), .A2(new_n5842), .A3(new_n5844), .B(\a[5] ), .Y(new_n5846));
  NOR3xp33_ASAP7_75t_L      g05590(.A(new_n5752), .B(new_n5753), .C(new_n5754), .Y(new_n5847));
  OAI21xp33_ASAP7_75t_L     g05591(.A1(new_n5847), .A2(new_n5757), .B(new_n5755), .Y(new_n5848));
  NAND2xp33_ASAP7_75t_L     g05592(.A(\b[31] ), .B(new_n815), .Y(new_n5849));
  NAND3xp33_ASAP7_75t_L     g05593(.A(new_n3210), .B(new_n808), .C(new_n3213), .Y(new_n5850));
  AOI22xp33_ASAP7_75t_L     g05594(.A1(new_n811), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n900), .Y(new_n5851));
  AND4x1_ASAP7_75t_L        g05595(.A(new_n5851), .B(new_n5850), .C(new_n5849), .D(\a[14] ), .Y(new_n5852));
  AOI31xp33_ASAP7_75t_L     g05596(.A1(new_n5850), .A2(new_n5849), .A3(new_n5851), .B(\a[14] ), .Y(new_n5853));
  NOR2xp33_ASAP7_75t_L      g05597(.A(new_n5853), .B(new_n5852), .Y(new_n5854));
  NOR3xp33_ASAP7_75t_L      g05598(.A(new_n5737), .B(new_n5738), .C(new_n5602), .Y(new_n5855));
  AOI21xp33_ASAP7_75t_L     g05599(.A1(new_n5598), .A2(new_n5746), .B(new_n5855), .Y(new_n5856));
  AOI22xp33_ASAP7_75t_L     g05600(.A1(new_n1076), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1253), .Y(new_n5857));
  OAI221xp5_ASAP7_75t_L     g05601(.A1(new_n1154), .A2(new_n2666), .B1(new_n1156), .B2(new_n2695), .C(new_n5857), .Y(new_n5858));
  XNOR2x2_ASAP7_75t_L       g05602(.A(\a[17] ), .B(new_n5858), .Y(new_n5859));
  NOR2xp33_ASAP7_75t_L      g05603(.A(new_n5714), .B(new_n5718), .Y(new_n5860));
  MAJIxp5_ASAP7_75t_L       g05604(.A(new_n5729), .B(new_n5860), .C(new_n5722), .Y(new_n5861));
  AOI22xp33_ASAP7_75t_L     g05605(.A1(new_n1360), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1581), .Y(new_n5862));
  OAI221xp5_ASAP7_75t_L     g05606(.A1(new_n1373), .A2(new_n2067), .B1(new_n1359), .B2(new_n2355), .C(new_n5862), .Y(new_n5863));
  XNOR2x2_ASAP7_75t_L       g05607(.A(\a[20] ), .B(new_n5863), .Y(new_n5864));
  INVx1_ASAP7_75t_L         g05608(.A(new_n5864), .Y(new_n5865));
  NOR3xp33_ASAP7_75t_L      g05609(.A(new_n5708), .B(new_n5707), .C(new_n5705), .Y(new_n5866));
  NAND2xp33_ASAP7_75t_L     g05610(.A(new_n5670), .B(new_n5665), .Y(new_n5867));
  MAJIxp5_ASAP7_75t_L       g05611(.A(new_n5680), .B(new_n5673), .C(new_n5867), .Y(new_n5868));
  AOI22xp33_ASAP7_75t_L     g05612(.A1(new_n2552), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n2736), .Y(new_n5869));
  OAI221xp5_ASAP7_75t_L     g05613(.A1(new_n2547), .A2(new_n1030), .B1(new_n2734), .B2(new_n1209), .C(new_n5869), .Y(new_n5870));
  XNOR2x2_ASAP7_75t_L       g05614(.A(\a[29] ), .B(new_n5870), .Y(new_n5871));
  AOI22xp33_ASAP7_75t_L     g05615(.A1(new_n3029), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n3258), .Y(new_n5872));
  OAI221xp5_ASAP7_75t_L     g05616(.A1(new_n3024), .A2(new_n784), .B1(new_n3256), .B2(new_n875), .C(new_n5872), .Y(new_n5873));
  XNOR2x2_ASAP7_75t_L       g05617(.A(\a[32] ), .B(new_n5873), .Y(new_n5874));
  INVx1_ASAP7_75t_L         g05618(.A(new_n5659), .Y(new_n5875));
  INVx1_ASAP7_75t_L         g05619(.A(new_n5650), .Y(new_n5876));
  A2O1A1Ixp33_ASAP7_75t_L   g05620(.A1(new_n5415), .A2(new_n5411), .B(new_n5419), .C(new_n5876), .Y(new_n5877));
  NAND2xp33_ASAP7_75t_L     g05621(.A(new_n5644), .B(new_n5646), .Y(new_n5878));
  NAND3xp33_ASAP7_75t_L     g05622(.A(new_n5878), .B(new_n5640), .C(new_n5636), .Y(new_n5879));
  INVx1_ASAP7_75t_L         g05623(.A(new_n5879), .Y(new_n5880));
  AOI22xp33_ASAP7_75t_L     g05624(.A1(new_n4283), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n4512), .Y(new_n5881));
  OAI221xp5_ASAP7_75t_L     g05625(.A1(new_n4277), .A2(new_n420), .B1(new_n4499), .B2(new_n494), .C(new_n5881), .Y(new_n5882));
  XNOR2x2_ASAP7_75t_L       g05626(.A(\a[38] ), .B(new_n5882), .Y(new_n5883));
  A2O1A1Ixp33_ASAP7_75t_L   g05627(.A1(new_n5403), .A2(new_n5637), .B(new_n5638), .C(new_n5635), .Y(new_n5884));
  NOR2xp33_ASAP7_75t_L      g05628(.A(new_n324), .B(new_n5154), .Y(new_n5885));
  NOR3xp33_ASAP7_75t_L      g05629(.A(new_n357), .B(new_n358), .C(new_n5158), .Y(new_n5886));
  OAI22xp33_ASAP7_75t_L     g05630(.A1(new_n5160), .A2(new_n298), .B1(new_n354), .B2(new_n5153), .Y(new_n5887));
  NOR3xp33_ASAP7_75t_L      g05631(.A(new_n5886), .B(new_n5887), .C(new_n5885), .Y(new_n5888));
  NAND2xp33_ASAP7_75t_L     g05632(.A(\a[41] ), .B(new_n5888), .Y(new_n5889));
  OAI31xp33_ASAP7_75t_L     g05633(.A1(new_n5886), .A2(new_n5885), .A3(new_n5887), .B(new_n4915), .Y(new_n5890));
  AND3x1_ASAP7_75t_L        g05634(.A(new_n5622), .B(new_n5625), .C(new_n5629), .Y(new_n5891));
  NAND2xp33_ASAP7_75t_L     g05635(.A(new_n5623), .B(new_n5626), .Y(new_n5892));
  NOR2xp33_ASAP7_75t_L      g05636(.A(new_n280), .B(new_n5892), .Y(new_n5893));
  NAND3xp33_ASAP7_75t_L     g05637(.A(new_n5626), .B(new_n5618), .C(new_n5620), .Y(new_n5894));
  NAND3xp33_ASAP7_75t_L     g05638(.A(new_n5392), .B(new_n5623), .C(new_n5627), .Y(new_n5895));
  OAI22xp33_ASAP7_75t_L     g05639(.A1(new_n5895), .A2(new_n258), .B1(new_n276), .B2(new_n5894), .Y(new_n5896));
  AOI211xp5_ASAP7_75t_L     g05640(.A1(\b[1] ), .A2(new_n5628), .B(new_n5893), .C(new_n5896), .Y(new_n5897));
  A2O1A1Ixp33_ASAP7_75t_L   g05641(.A1(new_n5891), .A2(new_n5396), .B(new_n5619), .C(new_n5897), .Y(new_n5898));
  O2A1O1Ixp33_ASAP7_75t_L   g05642(.A1(new_n258), .A2(new_n5392), .B(new_n5891), .C(new_n5619), .Y(new_n5899));
  INVx1_ASAP7_75t_L         g05643(.A(new_n5628), .Y(new_n5900));
  AND3x1_ASAP7_75t_L        g05644(.A(new_n5392), .B(new_n5627), .C(new_n5623), .Y(new_n5901));
  AOI221xp5_ASAP7_75t_L     g05645(.A1(new_n5624), .A2(\b[2] ), .B1(new_n5901), .B2(\b[0] ), .C(new_n5893), .Y(new_n5902));
  OAI21xp33_ASAP7_75t_L     g05646(.A1(new_n261), .A2(new_n5900), .B(new_n5902), .Y(new_n5903));
  NAND2xp33_ASAP7_75t_L     g05647(.A(new_n5903), .B(new_n5899), .Y(new_n5904));
  NAND4xp25_ASAP7_75t_L     g05648(.A(new_n5904), .B(new_n5889), .C(new_n5890), .D(new_n5898), .Y(new_n5905));
  NAND2xp33_ASAP7_75t_L     g05649(.A(new_n5890), .B(new_n5889), .Y(new_n5906));
  INVx1_ASAP7_75t_L         g05650(.A(new_n5898), .Y(new_n5907));
  A2O1A1Ixp33_ASAP7_75t_L   g05651(.A1(\b[0] ), .A2(new_n5626), .B(new_n5630), .C(\a[44] ), .Y(new_n5908));
  O2A1O1Ixp33_ASAP7_75t_L   g05652(.A1(new_n5900), .A2(new_n261), .B(new_n5902), .C(new_n5908), .Y(new_n5909));
  OAI21xp33_ASAP7_75t_L     g05653(.A1(new_n5907), .A2(new_n5909), .B(new_n5906), .Y(new_n5910));
  NAND2xp33_ASAP7_75t_L     g05654(.A(new_n5905), .B(new_n5910), .Y(new_n5911));
  NAND2xp33_ASAP7_75t_L     g05655(.A(new_n5884), .B(new_n5911), .Y(new_n5912));
  O2A1O1Ixp33_ASAP7_75t_L   g05656(.A1(new_n5609), .A2(new_n5412), .B(new_n5632), .C(new_n5639), .Y(new_n5913));
  NAND3xp33_ASAP7_75t_L     g05657(.A(new_n5913), .B(new_n5905), .C(new_n5910), .Y(new_n5914));
  AOI21xp33_ASAP7_75t_L     g05658(.A1(new_n5912), .A2(new_n5914), .B(new_n5883), .Y(new_n5915));
  XNOR2x2_ASAP7_75t_L       g05659(.A(new_n4268), .B(new_n5882), .Y(new_n5916));
  AOI21xp33_ASAP7_75t_L     g05660(.A1(new_n5910), .A2(new_n5905), .B(new_n5913), .Y(new_n5917));
  NOR2xp33_ASAP7_75t_L      g05661(.A(new_n5884), .B(new_n5911), .Y(new_n5918));
  NOR3xp33_ASAP7_75t_L      g05662(.A(new_n5918), .B(new_n5917), .C(new_n5916), .Y(new_n5919));
  NOR2xp33_ASAP7_75t_L      g05663(.A(new_n5915), .B(new_n5919), .Y(new_n5920));
  A2O1A1Ixp33_ASAP7_75t_L   g05664(.A1(new_n5877), .A2(new_n5653), .B(new_n5880), .C(new_n5920), .Y(new_n5921));
  AOI21xp33_ASAP7_75t_L     g05665(.A1(new_n5653), .A2(new_n5877), .B(new_n5880), .Y(new_n5922));
  OAI21xp33_ASAP7_75t_L     g05666(.A1(new_n5917), .A2(new_n5918), .B(new_n5916), .Y(new_n5923));
  NAND3xp33_ASAP7_75t_L     g05667(.A(new_n5912), .B(new_n5883), .C(new_n5914), .Y(new_n5924));
  NAND2xp33_ASAP7_75t_L     g05668(.A(new_n5924), .B(new_n5923), .Y(new_n5925));
  NAND2xp33_ASAP7_75t_L     g05669(.A(new_n5925), .B(new_n5922), .Y(new_n5926));
  AOI22xp33_ASAP7_75t_L     g05670(.A1(new_n3633), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n3858), .Y(new_n5927));
  OAI221xp5_ASAP7_75t_L     g05671(.A1(new_n3853), .A2(new_n617), .B1(new_n3856), .B2(new_n685), .C(new_n5927), .Y(new_n5928));
  XNOR2x2_ASAP7_75t_L       g05672(.A(\a[35] ), .B(new_n5928), .Y(new_n5929));
  NAND3xp33_ASAP7_75t_L     g05673(.A(new_n5921), .B(new_n5926), .C(new_n5929), .Y(new_n5930));
  AO21x2_ASAP7_75t_L        g05674(.A1(new_n5926), .A2(new_n5921), .B(new_n5929), .Y(new_n5931));
  NAND3xp33_ASAP7_75t_L     g05675(.A(new_n5652), .B(new_n5658), .C(new_n5654), .Y(new_n5932));
  NAND2xp33_ASAP7_75t_L     g05676(.A(new_n5932), .B(new_n5608), .Y(new_n5933));
  AND4x1_ASAP7_75t_L        g05677(.A(new_n5933), .B(new_n5931), .C(new_n5930), .D(new_n5875), .Y(new_n5934));
  AOI22xp33_ASAP7_75t_L     g05678(.A1(new_n5931), .A2(new_n5930), .B1(new_n5875), .B2(new_n5933), .Y(new_n5935));
  OAI21xp33_ASAP7_75t_L     g05679(.A1(new_n5935), .A2(new_n5934), .B(new_n5874), .Y(new_n5936));
  INVx1_ASAP7_75t_L         g05680(.A(new_n5874), .Y(new_n5937));
  NAND4xp25_ASAP7_75t_L     g05681(.A(new_n5933), .B(new_n5931), .C(new_n5875), .D(new_n5930), .Y(new_n5938));
  AO22x1_ASAP7_75t_L        g05682(.A1(new_n5930), .A2(new_n5931), .B1(new_n5875), .B2(new_n5933), .Y(new_n5939));
  NAND3xp33_ASAP7_75t_L     g05683(.A(new_n5939), .B(new_n5937), .C(new_n5938), .Y(new_n5940));
  NAND2xp33_ASAP7_75t_L     g05684(.A(new_n5936), .B(new_n5940), .Y(new_n5941));
  O2A1O1Ixp33_ASAP7_75t_L   g05685(.A1(new_n5667), .A2(new_n5668), .B(new_n5664), .C(new_n5941), .Y(new_n5942));
  NAND2xp33_ASAP7_75t_L     g05686(.A(new_n5444), .B(new_n5666), .Y(new_n5943));
  A2O1A1Ixp33_ASAP7_75t_L   g05687(.A1(new_n5448), .A2(new_n5943), .B(new_n5668), .C(new_n5664), .Y(new_n5944));
  AOI21xp33_ASAP7_75t_L     g05688(.A1(new_n5939), .A2(new_n5938), .B(new_n5937), .Y(new_n5945));
  NOR3xp33_ASAP7_75t_L      g05689(.A(new_n5934), .B(new_n5935), .C(new_n5874), .Y(new_n5946));
  NOR2xp33_ASAP7_75t_L      g05690(.A(new_n5946), .B(new_n5945), .Y(new_n5947));
  NOR2xp33_ASAP7_75t_L      g05691(.A(new_n5944), .B(new_n5947), .Y(new_n5948));
  OAI21xp33_ASAP7_75t_L     g05692(.A1(new_n5948), .A2(new_n5942), .B(new_n5871), .Y(new_n5949));
  INVx1_ASAP7_75t_L         g05693(.A(new_n5871), .Y(new_n5950));
  A2O1A1Ixp33_ASAP7_75t_L   g05694(.A1(new_n5663), .A2(new_n5604), .B(new_n5669), .C(new_n5947), .Y(new_n5951));
  NAND2xp33_ASAP7_75t_L     g05695(.A(new_n5450), .B(new_n5451), .Y(new_n5952));
  NOR2xp33_ASAP7_75t_L      g05696(.A(new_n5386), .B(new_n5603), .Y(new_n5953));
  A2O1A1O1Ixp25_ASAP7_75t_L g05697(.A1(new_n5382), .A2(new_n5952), .B(new_n5953), .C(new_n5663), .D(new_n5669), .Y(new_n5954));
  NAND2xp33_ASAP7_75t_L     g05698(.A(new_n5954), .B(new_n5941), .Y(new_n5955));
  NAND3xp33_ASAP7_75t_L     g05699(.A(new_n5950), .B(new_n5951), .C(new_n5955), .Y(new_n5956));
  NAND3xp33_ASAP7_75t_L     g05700(.A(new_n5868), .B(new_n5949), .C(new_n5956), .Y(new_n5957));
  NOR2xp33_ASAP7_75t_L      g05701(.A(new_n5676), .B(new_n5675), .Y(new_n5958));
  NAND2xp33_ASAP7_75t_L     g05702(.A(new_n5677), .B(new_n5958), .Y(new_n5959));
  AOI21xp33_ASAP7_75t_L     g05703(.A1(new_n5951), .A2(new_n5955), .B(new_n5950), .Y(new_n5960));
  NOR3xp33_ASAP7_75t_L      g05704(.A(new_n5942), .B(new_n5948), .C(new_n5871), .Y(new_n5961));
  OAI211xp5_ASAP7_75t_L     g05705(.A1(new_n5961), .A2(new_n5960), .B(new_n5959), .C(new_n5686), .Y(new_n5962));
  AOI22xp33_ASAP7_75t_L     g05706(.A1(new_n2114), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n2259), .Y(new_n5963));
  OAI221xp5_ASAP7_75t_L     g05707(.A1(new_n2109), .A2(new_n1432), .B1(new_n2257), .B2(new_n1547), .C(new_n5963), .Y(new_n5964));
  XNOR2x2_ASAP7_75t_L       g05708(.A(\a[26] ), .B(new_n5964), .Y(new_n5965));
  NAND3xp33_ASAP7_75t_L     g05709(.A(new_n5962), .B(new_n5957), .C(new_n5965), .Y(new_n5966));
  AO21x2_ASAP7_75t_L        g05710(.A1(new_n5957), .A2(new_n5962), .B(new_n5965), .Y(new_n5967));
  NAND2xp33_ASAP7_75t_L     g05711(.A(new_n5686), .B(new_n5681), .Y(new_n5968));
  NOR2xp33_ASAP7_75t_L      g05712(.A(new_n5689), .B(new_n5968), .Y(new_n5969));
  INVx1_ASAP7_75t_L         g05713(.A(new_n5969), .Y(new_n5970));
  AND4x1_ASAP7_75t_L        g05714(.A(new_n5697), .B(new_n5970), .C(new_n5966), .D(new_n5967), .Y(new_n5971));
  O2A1O1Ixp33_ASAP7_75t_L   g05715(.A1(new_n5695), .A2(new_n5691), .B(new_n5696), .C(new_n5969), .Y(new_n5972));
  AOI21xp33_ASAP7_75t_L     g05716(.A1(new_n5967), .A2(new_n5966), .B(new_n5972), .Y(new_n5973));
  NOR2xp33_ASAP7_75t_L      g05717(.A(new_n1774), .B(new_n1699), .Y(new_n5974));
  INVx1_ASAP7_75t_L         g05718(.A(new_n5974), .Y(new_n5975));
  NAND3xp33_ASAP7_75t_L     g05719(.A(new_n1912), .B(new_n1695), .C(new_n1914), .Y(new_n5976));
  AOI22xp33_ASAP7_75t_L     g05720(.A1(new_n1704), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1837), .Y(new_n5977));
  AND4x1_ASAP7_75t_L        g05721(.A(new_n5977), .B(new_n5976), .C(new_n5975), .D(\a[23] ), .Y(new_n5978));
  AOI31xp33_ASAP7_75t_L     g05722(.A1(new_n5976), .A2(new_n5975), .A3(new_n5977), .B(\a[23] ), .Y(new_n5979));
  NOR2xp33_ASAP7_75t_L      g05723(.A(new_n5979), .B(new_n5978), .Y(new_n5980));
  OAI21xp33_ASAP7_75t_L     g05724(.A1(new_n5973), .A2(new_n5971), .B(new_n5980), .Y(new_n5981));
  NAND3xp33_ASAP7_75t_L     g05725(.A(new_n5972), .B(new_n5967), .C(new_n5966), .Y(new_n5982));
  INVx1_ASAP7_75t_L         g05726(.A(new_n5966), .Y(new_n5983));
  AOI21xp33_ASAP7_75t_L     g05727(.A1(new_n5962), .A2(new_n5957), .B(new_n5965), .Y(new_n5984));
  MAJIxp5_ASAP7_75t_L       g05728(.A(new_n5693), .B(new_n5689), .C(new_n5968), .Y(new_n5985));
  OAI21xp33_ASAP7_75t_L     g05729(.A1(new_n5984), .A2(new_n5983), .B(new_n5985), .Y(new_n5986));
  INVx1_ASAP7_75t_L         g05730(.A(new_n5980), .Y(new_n5987));
  NAND3xp33_ASAP7_75t_L     g05731(.A(new_n5986), .B(new_n5982), .C(new_n5987), .Y(new_n5988));
  AOI221xp5_ASAP7_75t_L     g05732(.A1(new_n5981), .A2(new_n5988), .B1(new_n5710), .B2(new_n5713), .C(new_n5866), .Y(new_n5989));
  INVx1_ASAP7_75t_L         g05733(.A(new_n5989), .Y(new_n5990));
  AOI21xp33_ASAP7_75t_L     g05734(.A1(new_n5986), .A2(new_n5982), .B(new_n5987), .Y(new_n5991));
  NOR3xp33_ASAP7_75t_L      g05735(.A(new_n5971), .B(new_n5973), .C(new_n5980), .Y(new_n5992));
  NOR2xp33_ASAP7_75t_L      g05736(.A(new_n5992), .B(new_n5991), .Y(new_n5993));
  A2O1A1Ixp33_ASAP7_75t_L   g05737(.A1(new_n5713), .A2(new_n5710), .B(new_n5866), .C(new_n5993), .Y(new_n5994));
  AOI21xp33_ASAP7_75t_L     g05738(.A1(new_n5990), .A2(new_n5994), .B(new_n5865), .Y(new_n5995));
  INVx1_ASAP7_75t_L         g05739(.A(new_n5866), .Y(new_n5996));
  NAND2xp33_ASAP7_75t_L     g05740(.A(new_n5988), .B(new_n5981), .Y(new_n5997));
  O2A1O1Ixp33_ASAP7_75t_L   g05741(.A1(new_n5717), .A2(new_n5724), .B(new_n5996), .C(new_n5997), .Y(new_n5998));
  NOR3xp33_ASAP7_75t_L      g05742(.A(new_n5998), .B(new_n5989), .C(new_n5864), .Y(new_n5999));
  NOR3xp33_ASAP7_75t_L      g05743(.A(new_n5861), .B(new_n5995), .C(new_n5999), .Y(new_n6000));
  NAND2xp33_ASAP7_75t_L     g05744(.A(new_n5731), .B(new_n5732), .Y(new_n6001));
  NAND2xp33_ASAP7_75t_L     g05745(.A(new_n5726), .B(new_n5725), .Y(new_n6002));
  NOR2xp33_ASAP7_75t_L      g05746(.A(new_n5727), .B(new_n6002), .Y(new_n6003));
  OAI21xp33_ASAP7_75t_L     g05747(.A1(new_n5989), .A2(new_n5998), .B(new_n5864), .Y(new_n6004));
  NAND3xp33_ASAP7_75t_L     g05748(.A(new_n5990), .B(new_n5994), .C(new_n5865), .Y(new_n6005));
  AOI221xp5_ASAP7_75t_L     g05749(.A1(new_n6001), .A2(new_n5729), .B1(new_n6004), .B2(new_n6005), .C(new_n6003), .Y(new_n6006));
  OAI21xp33_ASAP7_75t_L     g05750(.A1(new_n6006), .A2(new_n6000), .B(new_n5859), .Y(new_n6007));
  INVx1_ASAP7_75t_L         g05751(.A(new_n5859), .Y(new_n6008));
  MAJIxp5_ASAP7_75t_L       g05752(.A(new_n5736), .B(new_n6002), .C(new_n5727), .Y(new_n6009));
  NAND3xp33_ASAP7_75t_L     g05753(.A(new_n6009), .B(new_n6004), .C(new_n6005), .Y(new_n6010));
  OAI21xp33_ASAP7_75t_L     g05754(.A1(new_n5995), .A2(new_n5999), .B(new_n5861), .Y(new_n6011));
  NAND3xp33_ASAP7_75t_L     g05755(.A(new_n6010), .B(new_n6008), .C(new_n6011), .Y(new_n6012));
  NAND2xp33_ASAP7_75t_L     g05756(.A(new_n6007), .B(new_n6012), .Y(new_n6013));
  NOR2xp33_ASAP7_75t_L      g05757(.A(new_n5856), .B(new_n6013), .Y(new_n6014));
  AOI221xp5_ASAP7_75t_L     g05758(.A1(new_n5598), .A2(new_n5746), .B1(new_n6007), .B2(new_n6012), .C(new_n5855), .Y(new_n6015));
  OAI21xp33_ASAP7_75t_L     g05759(.A1(new_n6015), .A2(new_n6014), .B(new_n5854), .Y(new_n6016));
  INVx1_ASAP7_75t_L         g05760(.A(new_n5854), .Y(new_n6017));
  INVx1_ASAP7_75t_L         g05761(.A(new_n5855), .Y(new_n6018));
  A2O1A1Ixp33_ASAP7_75t_L   g05762(.A1(new_n5528), .A2(new_n5597), .B(new_n5740), .C(new_n6018), .Y(new_n6019));
  AOI21xp33_ASAP7_75t_L     g05763(.A1(new_n6010), .A2(new_n6011), .B(new_n6008), .Y(new_n6020));
  NOR3xp33_ASAP7_75t_L      g05764(.A(new_n6000), .B(new_n6006), .C(new_n5859), .Y(new_n6021));
  NOR2xp33_ASAP7_75t_L      g05765(.A(new_n6021), .B(new_n6020), .Y(new_n6022));
  NAND2xp33_ASAP7_75t_L     g05766(.A(new_n6022), .B(new_n6019), .Y(new_n6023));
  NAND2xp33_ASAP7_75t_L     g05767(.A(new_n5856), .B(new_n6013), .Y(new_n6024));
  NAND3xp33_ASAP7_75t_L     g05768(.A(new_n6023), .B(new_n6017), .C(new_n6024), .Y(new_n6025));
  NAND3xp33_ASAP7_75t_L     g05769(.A(new_n5848), .B(new_n6016), .C(new_n6025), .Y(new_n6026));
  AOI21xp33_ASAP7_75t_L     g05770(.A1(new_n5747), .A2(new_n5741), .B(new_n5750), .Y(new_n6027));
  A2O1A1O1Ixp25_ASAP7_75t_L g05771(.A1(new_n5537), .A2(new_n5366), .B(new_n5540), .C(new_n5751), .D(new_n6027), .Y(new_n6028));
  AOI21xp33_ASAP7_75t_L     g05772(.A1(new_n6023), .A2(new_n6024), .B(new_n6017), .Y(new_n6029));
  NOR3xp33_ASAP7_75t_L      g05773(.A(new_n6014), .B(new_n6015), .C(new_n5854), .Y(new_n6030));
  OAI21xp33_ASAP7_75t_L     g05774(.A1(new_n6030), .A2(new_n6029), .B(new_n6028), .Y(new_n6031));
  NOR2xp33_ASAP7_75t_L      g05775(.A(new_n3584), .B(new_n821), .Y(new_n6032));
  INVx1_ASAP7_75t_L         g05776(.A(new_n6032), .Y(new_n6033));
  NAND2xp33_ASAP7_75t_L     g05777(.A(new_n578), .B(new_n3811), .Y(new_n6034));
  AOI22xp33_ASAP7_75t_L     g05778(.A1(\b[33] ), .A2(new_n651), .B1(\b[35] ), .B2(new_n581), .Y(new_n6035));
  AND4x1_ASAP7_75t_L        g05779(.A(new_n6035), .B(new_n6034), .C(new_n6033), .D(\a[11] ), .Y(new_n6036));
  AOI31xp33_ASAP7_75t_L     g05780(.A1(new_n6034), .A2(new_n6033), .A3(new_n6035), .B(\a[11] ), .Y(new_n6037));
  NOR2xp33_ASAP7_75t_L      g05781(.A(new_n6037), .B(new_n6036), .Y(new_n6038));
  NAND3xp33_ASAP7_75t_L     g05782(.A(new_n6026), .B(new_n6031), .C(new_n6038), .Y(new_n6039));
  NOR3xp33_ASAP7_75t_L      g05783(.A(new_n6028), .B(new_n6029), .C(new_n6030), .Y(new_n6040));
  AOI21xp33_ASAP7_75t_L     g05784(.A1(new_n6025), .A2(new_n6016), .B(new_n5848), .Y(new_n6041));
  INVx1_ASAP7_75t_L         g05785(.A(new_n6038), .Y(new_n6042));
  OAI21xp33_ASAP7_75t_L     g05786(.A1(new_n6040), .A2(new_n6041), .B(new_n6042), .Y(new_n6043));
  NAND3xp33_ASAP7_75t_L     g05787(.A(new_n5759), .B(new_n5756), .C(new_n5766), .Y(new_n6044));
  NAND4xp25_ASAP7_75t_L     g05788(.A(new_n5775), .B(new_n6044), .C(new_n6043), .D(new_n6039), .Y(new_n6045));
  NAND2xp33_ASAP7_75t_L     g05789(.A(new_n6039), .B(new_n6043), .Y(new_n6046));
  A2O1A1Ixp33_ASAP7_75t_L   g05790(.A1(new_n5767), .A2(new_n5763), .B(new_n5769), .C(new_n6044), .Y(new_n6047));
  NAND2xp33_ASAP7_75t_L     g05791(.A(new_n6047), .B(new_n6046), .Y(new_n6048));
  NAND2xp33_ASAP7_75t_L     g05792(.A(\b[37] ), .B(new_n447), .Y(new_n6049));
  NAND2xp33_ASAP7_75t_L     g05793(.A(new_n441), .B(new_n4640), .Y(new_n6050));
  AOI22xp33_ASAP7_75t_L     g05794(.A1(new_n444), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n471), .Y(new_n6051));
  NAND4xp25_ASAP7_75t_L     g05795(.A(new_n6050), .B(\a[8] ), .C(new_n6049), .D(new_n6051), .Y(new_n6052));
  NAND2xp33_ASAP7_75t_L     g05796(.A(new_n6051), .B(new_n6050), .Y(new_n6053));
  A2O1A1Ixp33_ASAP7_75t_L   g05797(.A1(\b[37] ), .A2(new_n447), .B(new_n6053), .C(new_n435), .Y(new_n6054));
  AND2x2_ASAP7_75t_L        g05798(.A(new_n6052), .B(new_n6054), .Y(new_n6055));
  NAND3xp33_ASAP7_75t_L     g05799(.A(new_n6048), .B(new_n6045), .C(new_n6055), .Y(new_n6056));
  NOR2xp33_ASAP7_75t_L      g05800(.A(new_n6047), .B(new_n6046), .Y(new_n6057));
  AOI22xp33_ASAP7_75t_L     g05801(.A1(new_n6039), .A2(new_n6043), .B1(new_n6044), .B2(new_n5775), .Y(new_n6058));
  NAND2xp33_ASAP7_75t_L     g05802(.A(new_n6052), .B(new_n6054), .Y(new_n6059));
  OAI21xp33_ASAP7_75t_L     g05803(.A1(new_n6058), .A2(new_n6057), .B(new_n6059), .Y(new_n6060));
  AOI221xp5_ASAP7_75t_L     g05804(.A1(new_n5793), .A2(new_n5788), .B1(new_n6056), .B2(new_n6060), .C(new_n5780), .Y(new_n6061));
  INVx1_ASAP7_75t_L         g05805(.A(new_n5793), .Y(new_n6062));
  NAND2xp33_ASAP7_75t_L     g05806(.A(new_n6056), .B(new_n6060), .Y(new_n6063));
  O2A1O1Ixp33_ASAP7_75t_L   g05807(.A1(new_n5783), .A2(new_n6062), .B(new_n5787), .C(new_n6063), .Y(new_n6064));
  OAI22xp33_ASAP7_75t_L     g05808(.A1(new_n6064), .A2(new_n6061), .B1(new_n5846), .B2(new_n5845), .Y(new_n6065));
  NOR2xp33_ASAP7_75t_L      g05809(.A(new_n5846), .B(new_n5845), .Y(new_n6066));
  INVx1_ASAP7_75t_L         g05810(.A(new_n6061), .Y(new_n6067));
  NOR3xp33_ASAP7_75t_L      g05811(.A(new_n6057), .B(new_n6058), .C(new_n6059), .Y(new_n6068));
  AOI21xp33_ASAP7_75t_L     g05812(.A1(new_n6048), .A2(new_n6045), .B(new_n6055), .Y(new_n6069));
  NOR2xp33_ASAP7_75t_L      g05813(.A(new_n6069), .B(new_n6068), .Y(new_n6070));
  A2O1A1Ixp33_ASAP7_75t_L   g05814(.A1(new_n5788), .A2(new_n5793), .B(new_n5780), .C(new_n6070), .Y(new_n6071));
  NAND3xp33_ASAP7_75t_L     g05815(.A(new_n6067), .B(new_n6071), .C(new_n6066), .Y(new_n6072));
  AOI21xp33_ASAP7_75t_L     g05816(.A1(new_n6072), .A2(new_n6065), .B(new_n5841), .Y(new_n6073));
  A2O1A1Ixp33_ASAP7_75t_L   g05817(.A1(new_n5575), .A2(new_n5585), .B(new_n5800), .C(new_n5796), .Y(new_n6074));
  NAND2xp33_ASAP7_75t_L     g05818(.A(new_n6065), .B(new_n6072), .Y(new_n6075));
  NOR2xp33_ASAP7_75t_L      g05819(.A(new_n6075), .B(new_n6074), .Y(new_n6076));
  NOR3xp33_ASAP7_75t_L      g05820(.A(new_n6076), .B(new_n6073), .C(new_n5838), .Y(new_n6077));
  INVx1_ASAP7_75t_L         g05821(.A(new_n6077), .Y(new_n6078));
  OAI21xp33_ASAP7_75t_L     g05822(.A1(new_n6073), .A2(new_n6076), .B(new_n5838), .Y(new_n6079));
  NAND2xp33_ASAP7_75t_L     g05823(.A(new_n6079), .B(new_n6078), .Y(new_n6080));
  XOR2x2_ASAP7_75t_L        g05824(.A(new_n5827), .B(new_n6080), .Y(\f[44] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g05825(.A1(new_n5824), .A2(new_n5823), .B(new_n5826), .C(new_n6079), .D(new_n6077), .Y(new_n6082));
  A2O1A1Ixp33_ASAP7_75t_L   g05826(.A1(new_n5791), .A2(new_n5586), .B(new_n5840), .C(new_n6075), .Y(new_n6083));
  NOR3xp33_ASAP7_75t_L      g05827(.A(new_n6041), .B(new_n6040), .C(new_n6038), .Y(new_n6084));
  NAND2xp33_ASAP7_75t_L     g05828(.A(\b[34] ), .B(new_n651), .Y(new_n6085));
  OAI221xp5_ASAP7_75t_L     g05829(.A1(new_n580), .A2(new_n4216), .B1(new_n577), .B2(new_n4223), .C(new_n6085), .Y(new_n6086));
  AOI21xp33_ASAP7_75t_L     g05830(.A1(new_n584), .A2(\b[35] ), .B(new_n6086), .Y(new_n6087));
  NAND2xp33_ASAP7_75t_L     g05831(.A(\a[11] ), .B(new_n6087), .Y(new_n6088));
  A2O1A1Ixp33_ASAP7_75t_L   g05832(.A1(\b[35] ), .A2(new_n584), .B(new_n6086), .C(new_n574), .Y(new_n6089));
  NAND2xp33_ASAP7_75t_L     g05833(.A(new_n6089), .B(new_n6088), .Y(new_n6090));
  OAI21xp33_ASAP7_75t_L     g05834(.A1(new_n6029), .A2(new_n6028), .B(new_n6025), .Y(new_n6091));
  NOR2xp33_ASAP7_75t_L      g05835(.A(new_n2688), .B(new_n1154), .Y(new_n6092));
  INVx1_ASAP7_75t_L         g05836(.A(new_n6092), .Y(new_n6093));
  NAND2xp33_ASAP7_75t_L     g05837(.A(new_n1073), .B(new_n2989), .Y(new_n6094));
  AOI22xp33_ASAP7_75t_L     g05838(.A1(new_n1076), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1253), .Y(new_n6095));
  AND4x1_ASAP7_75t_L        g05839(.A(new_n6095), .B(new_n6094), .C(new_n6093), .D(\a[17] ), .Y(new_n6096));
  AOI31xp33_ASAP7_75t_L     g05840(.A1(new_n6094), .A2(new_n6093), .A3(new_n6095), .B(\a[17] ), .Y(new_n6097));
  NOR2xp33_ASAP7_75t_L      g05841(.A(new_n6097), .B(new_n6096), .Y(new_n6098));
  INVx1_ASAP7_75t_L         g05842(.A(new_n6098), .Y(new_n6099));
  INVx1_ASAP7_75t_L         g05843(.A(new_n6003), .Y(new_n6100));
  A2O1A1Ixp33_ASAP7_75t_L   g05844(.A1(new_n6100), .A2(new_n5730), .B(new_n5995), .C(new_n6005), .Y(new_n6101));
  A2O1A1Ixp33_ASAP7_75t_L   g05845(.A1(new_n5686), .A2(new_n5959), .B(new_n5960), .C(new_n5956), .Y(new_n6102));
  A2O1A1O1Ixp25_ASAP7_75t_L g05846(.A1(new_n5663), .A2(new_n5604), .B(new_n5669), .C(new_n5936), .D(new_n5946), .Y(new_n6103));
  AOI22xp33_ASAP7_75t_L     g05847(.A1(new_n3029), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n3258), .Y(new_n6104));
  OAI221xp5_ASAP7_75t_L     g05848(.A1(new_n3024), .A2(new_n869), .B1(new_n3256), .B2(new_n950), .C(new_n6104), .Y(new_n6105));
  XNOR2x2_ASAP7_75t_L       g05849(.A(\a[32] ), .B(new_n6105), .Y(new_n6106));
  AOI21xp33_ASAP7_75t_L     g05850(.A1(new_n5921), .A2(new_n5926), .B(new_n5929), .Y(new_n6107));
  AO31x2_ASAP7_75t_L        g05851(.A1(new_n5933), .A2(new_n5930), .A3(new_n5875), .B(new_n6107), .Y(new_n6108));
  OAI22xp33_ASAP7_75t_L     g05852(.A1(new_n4052), .A2(new_n617), .B1(new_n760), .B2(new_n4061), .Y(new_n6109));
  AOI221xp5_ASAP7_75t_L     g05853(.A1(new_n3639), .A2(\b[11] ), .B1(new_n3630), .B2(new_n1232), .C(new_n6109), .Y(new_n6110));
  XNOR2x2_ASAP7_75t_L       g05854(.A(new_n3628), .B(new_n6110), .Y(new_n6111));
  A2O1A1Ixp33_ASAP7_75t_L   g05855(.A1(new_n5648), .A2(new_n5647), .B(new_n5651), .C(new_n5879), .Y(new_n6112));
  NOR3xp33_ASAP7_75t_L      g05856(.A(new_n5918), .B(new_n5917), .C(new_n5883), .Y(new_n6113));
  NAND5xp2_ASAP7_75t_L      g05857(.A(\a[44] ), .B(new_n5622), .C(new_n5625), .D(new_n5629), .E(new_n5396), .Y(new_n6114));
  INVx1_ASAP7_75t_L         g05858(.A(new_n6114), .Y(new_n6115));
  INVx1_ASAP7_75t_L         g05859(.A(\a[45] ), .Y(new_n6116));
  NAND2xp33_ASAP7_75t_L     g05860(.A(\a[44] ), .B(new_n6116), .Y(new_n6117));
  NAND2xp33_ASAP7_75t_L     g05861(.A(\a[45] ), .B(new_n5619), .Y(new_n6118));
  AND2x2_ASAP7_75t_L        g05862(.A(new_n6117), .B(new_n6118), .Y(new_n6119));
  NOR2xp33_ASAP7_75t_L      g05863(.A(new_n258), .B(new_n6119), .Y(new_n6120));
  INVx1_ASAP7_75t_L         g05864(.A(new_n6120), .Y(new_n6121));
  AOI21xp33_ASAP7_75t_L     g05865(.A1(new_n6115), .A2(new_n5897), .B(new_n6121), .Y(new_n6122));
  NOR3xp33_ASAP7_75t_L      g05866(.A(new_n5903), .B(new_n6120), .C(new_n6114), .Y(new_n6123));
  OAI22xp33_ASAP7_75t_L     g05867(.A1(new_n5895), .A2(new_n261), .B1(new_n298), .B2(new_n5894), .Y(new_n6124));
  AOI221xp5_ASAP7_75t_L     g05868(.A1(\b[2] ), .A2(new_n5628), .B1(new_n406), .B2(new_n5621), .C(new_n6124), .Y(new_n6125));
  NAND2xp33_ASAP7_75t_L     g05869(.A(\a[44] ), .B(new_n6125), .Y(new_n6126));
  NAND2xp33_ASAP7_75t_L     g05870(.A(\b[3] ), .B(new_n5624), .Y(new_n6127));
  OAI221xp5_ASAP7_75t_L     g05871(.A1(new_n5895), .A2(new_n261), .B1(new_n5892), .B2(new_n302), .C(new_n6127), .Y(new_n6128));
  A2O1A1Ixp33_ASAP7_75t_L   g05872(.A1(\b[2] ), .A2(new_n5628), .B(new_n6128), .C(new_n5619), .Y(new_n6129));
  NAND2xp33_ASAP7_75t_L     g05873(.A(new_n6129), .B(new_n6126), .Y(new_n6130));
  OAI21xp33_ASAP7_75t_L     g05874(.A1(new_n6122), .A2(new_n6123), .B(new_n6130), .Y(new_n6131));
  OAI21xp33_ASAP7_75t_L     g05875(.A1(new_n6114), .A2(new_n5903), .B(new_n6120), .Y(new_n6132));
  NAND3xp33_ASAP7_75t_L     g05876(.A(new_n6115), .B(new_n5897), .C(new_n6121), .Y(new_n6133));
  XNOR2x2_ASAP7_75t_L       g05877(.A(new_n5619), .B(new_n6125), .Y(new_n6134));
  NAND3xp33_ASAP7_75t_L     g05878(.A(new_n6134), .B(new_n6133), .C(new_n6132), .Y(new_n6135));
  NOR2xp33_ASAP7_75t_L      g05879(.A(new_n354), .B(new_n5154), .Y(new_n6136));
  INVx1_ASAP7_75t_L         g05880(.A(new_n6136), .Y(new_n6137));
  NAND2xp33_ASAP7_75t_L     g05881(.A(new_n4917), .B(new_n526), .Y(new_n6138));
  AOI22xp33_ASAP7_75t_L     g05882(.A1(new_n4920), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n5167), .Y(new_n6139));
  NAND4xp25_ASAP7_75t_L     g05883(.A(new_n6138), .B(\a[41] ), .C(new_n6137), .D(new_n6139), .Y(new_n6140));
  AOI31xp33_ASAP7_75t_L     g05884(.A1(new_n6138), .A2(new_n6137), .A3(new_n6139), .B(\a[41] ), .Y(new_n6141));
  INVx1_ASAP7_75t_L         g05885(.A(new_n6141), .Y(new_n6142));
  NAND4xp25_ASAP7_75t_L     g05886(.A(new_n6135), .B(new_n6140), .C(new_n6142), .D(new_n6131), .Y(new_n6143));
  AOI21xp33_ASAP7_75t_L     g05887(.A1(new_n6133), .A2(new_n6132), .B(new_n6134), .Y(new_n6144));
  AND4x1_ASAP7_75t_L        g05888(.A(new_n6133), .B(new_n6132), .C(new_n6129), .D(new_n6126), .Y(new_n6145));
  INVx1_ASAP7_75t_L         g05889(.A(new_n6140), .Y(new_n6146));
  OAI22xp33_ASAP7_75t_L     g05890(.A1(new_n6144), .A2(new_n6145), .B1(new_n6141), .B2(new_n6146), .Y(new_n6147));
  NOR2xp33_ASAP7_75t_L      g05891(.A(new_n5909), .B(new_n5907), .Y(new_n6148));
  MAJIxp5_ASAP7_75t_L       g05892(.A(new_n5884), .B(new_n5906), .C(new_n6148), .Y(new_n6149));
  NAND3xp33_ASAP7_75t_L     g05893(.A(new_n6149), .B(new_n6147), .C(new_n6143), .Y(new_n6150));
  NAND2xp33_ASAP7_75t_L     g05894(.A(new_n6143), .B(new_n6147), .Y(new_n6151));
  A2O1A1Ixp33_ASAP7_75t_L   g05895(.A1(new_n6148), .A2(new_n5906), .B(new_n5917), .C(new_n6151), .Y(new_n6152));
  NAND2xp33_ASAP7_75t_L     g05896(.A(\b[8] ), .B(new_n4285), .Y(new_n6153));
  NAND2xp33_ASAP7_75t_L     g05897(.A(new_n4274), .B(new_n731), .Y(new_n6154));
  AOI22xp33_ASAP7_75t_L     g05898(.A1(new_n4283), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n4512), .Y(new_n6155));
  NAND4xp25_ASAP7_75t_L     g05899(.A(new_n6154), .B(\a[38] ), .C(new_n6153), .D(new_n6155), .Y(new_n6156));
  OAI211xp5_ASAP7_75t_L     g05900(.A1(new_n4499), .A2(new_n548), .B(new_n6153), .C(new_n6155), .Y(new_n6157));
  NAND2xp33_ASAP7_75t_L     g05901(.A(new_n4268), .B(new_n6157), .Y(new_n6158));
  NAND2xp33_ASAP7_75t_L     g05902(.A(new_n6158), .B(new_n6156), .Y(new_n6159));
  AOI21xp33_ASAP7_75t_L     g05903(.A1(new_n6152), .A2(new_n6150), .B(new_n6159), .Y(new_n6160));
  NAND2xp33_ASAP7_75t_L     g05904(.A(new_n5906), .B(new_n6148), .Y(new_n6161));
  A2O1A1Ixp33_ASAP7_75t_L   g05905(.A1(new_n5905), .A2(new_n5910), .B(new_n5913), .C(new_n6161), .Y(new_n6162));
  NOR2xp33_ASAP7_75t_L      g05906(.A(new_n6162), .B(new_n6151), .Y(new_n6163));
  AOI21xp33_ASAP7_75t_L     g05907(.A1(new_n6147), .A2(new_n6143), .B(new_n6149), .Y(new_n6164));
  AOI211xp5_ASAP7_75t_L     g05908(.A1(new_n6158), .A2(new_n6156), .B(new_n6163), .C(new_n6164), .Y(new_n6165));
  NOR2xp33_ASAP7_75t_L      g05909(.A(new_n6160), .B(new_n6165), .Y(new_n6166));
  A2O1A1Ixp33_ASAP7_75t_L   g05910(.A1(new_n5925), .A2(new_n6112), .B(new_n6113), .C(new_n6166), .Y(new_n6167));
  O2A1O1Ixp33_ASAP7_75t_L   g05911(.A1(new_n5915), .A2(new_n5919), .B(new_n6112), .C(new_n6113), .Y(new_n6168));
  OAI211xp5_ASAP7_75t_L     g05912(.A1(new_n6163), .A2(new_n6164), .B(new_n6156), .C(new_n6158), .Y(new_n6169));
  NAND3xp33_ASAP7_75t_L     g05913(.A(new_n6159), .B(new_n6152), .C(new_n6150), .Y(new_n6170));
  NAND2xp33_ASAP7_75t_L     g05914(.A(new_n6170), .B(new_n6169), .Y(new_n6171));
  NAND2xp33_ASAP7_75t_L     g05915(.A(new_n6171), .B(new_n6168), .Y(new_n6172));
  AOI21xp33_ASAP7_75t_L     g05916(.A1(new_n6167), .A2(new_n6172), .B(new_n6111), .Y(new_n6173));
  XNOR2x2_ASAP7_75t_L       g05917(.A(\a[35] ), .B(new_n6110), .Y(new_n6174));
  INVx1_ASAP7_75t_L         g05918(.A(new_n6113), .Y(new_n6175));
  O2A1O1Ixp33_ASAP7_75t_L   g05919(.A1(new_n5922), .A2(new_n5920), .B(new_n6175), .C(new_n6171), .Y(new_n6176));
  AOI221xp5_ASAP7_75t_L     g05920(.A1(new_n6112), .A2(new_n5925), .B1(new_n6170), .B2(new_n6169), .C(new_n6113), .Y(new_n6177));
  NOR3xp33_ASAP7_75t_L      g05921(.A(new_n6176), .B(new_n6177), .C(new_n6174), .Y(new_n6178));
  OAI21xp33_ASAP7_75t_L     g05922(.A1(new_n6173), .A2(new_n6178), .B(new_n6108), .Y(new_n6179));
  AOI31xp33_ASAP7_75t_L     g05923(.A1(new_n5933), .A2(new_n5930), .A3(new_n5875), .B(new_n6107), .Y(new_n6180));
  OAI21xp33_ASAP7_75t_L     g05924(.A1(new_n6177), .A2(new_n6176), .B(new_n6174), .Y(new_n6181));
  NAND3xp33_ASAP7_75t_L     g05925(.A(new_n6167), .B(new_n6172), .C(new_n6111), .Y(new_n6182));
  NAND3xp33_ASAP7_75t_L     g05926(.A(new_n6180), .B(new_n6181), .C(new_n6182), .Y(new_n6183));
  AND3x1_ASAP7_75t_L        g05927(.A(new_n6179), .B(new_n6183), .C(new_n6106), .Y(new_n6184));
  AOI21xp33_ASAP7_75t_L     g05928(.A1(new_n6179), .A2(new_n6183), .B(new_n6106), .Y(new_n6185));
  NOR3xp33_ASAP7_75t_L      g05929(.A(new_n6103), .B(new_n6184), .C(new_n6185), .Y(new_n6186));
  NAND3xp33_ASAP7_75t_L     g05930(.A(new_n6179), .B(new_n6183), .C(new_n6106), .Y(new_n6187));
  AO21x2_ASAP7_75t_L        g05931(.A1(new_n6183), .A2(new_n6179), .B(new_n6106), .Y(new_n6188));
  AOI221xp5_ASAP7_75t_L     g05932(.A1(new_n5944), .A2(new_n5936), .B1(new_n6187), .B2(new_n6188), .C(new_n5946), .Y(new_n6189));
  OAI22xp33_ASAP7_75t_L     g05933(.A1(new_n2747), .A2(new_n1030), .B1(new_n1313), .B2(new_n2545), .Y(new_n6190));
  AOI221xp5_ASAP7_75t_L     g05934(.A1(new_n2553), .A2(\b[17] ), .B1(new_n2544), .B2(new_n1319), .C(new_n6190), .Y(new_n6191));
  XNOR2x2_ASAP7_75t_L       g05935(.A(\a[29] ), .B(new_n6191), .Y(new_n6192));
  OAI21xp33_ASAP7_75t_L     g05936(.A1(new_n6189), .A2(new_n6186), .B(new_n6192), .Y(new_n6193));
  OAI21xp33_ASAP7_75t_L     g05937(.A1(new_n5945), .A2(new_n5954), .B(new_n5940), .Y(new_n6194));
  NAND3xp33_ASAP7_75t_L     g05938(.A(new_n6194), .B(new_n6187), .C(new_n6188), .Y(new_n6195));
  OAI21xp33_ASAP7_75t_L     g05939(.A1(new_n6184), .A2(new_n6185), .B(new_n6103), .Y(new_n6196));
  XNOR2x2_ASAP7_75t_L       g05940(.A(new_n2538), .B(new_n6191), .Y(new_n6197));
  NAND3xp33_ASAP7_75t_L     g05941(.A(new_n6195), .B(new_n6196), .C(new_n6197), .Y(new_n6198));
  NAND3xp33_ASAP7_75t_L     g05942(.A(new_n6102), .B(new_n6193), .C(new_n6198), .Y(new_n6199));
  NAND2xp33_ASAP7_75t_L     g05943(.A(new_n5674), .B(new_n5678), .Y(new_n6200));
  NOR2xp33_ASAP7_75t_L      g05944(.A(new_n5673), .B(new_n5867), .Y(new_n6201));
  A2O1A1O1Ixp25_ASAP7_75t_L g05945(.A1(new_n5685), .A2(new_n6200), .B(new_n6201), .C(new_n5949), .D(new_n5961), .Y(new_n6202));
  AOI21xp33_ASAP7_75t_L     g05946(.A1(new_n6195), .A2(new_n6196), .B(new_n6197), .Y(new_n6203));
  NOR3xp33_ASAP7_75t_L      g05947(.A(new_n6186), .B(new_n6189), .C(new_n6192), .Y(new_n6204));
  OAI21xp33_ASAP7_75t_L     g05948(.A1(new_n6203), .A2(new_n6204), .B(new_n6202), .Y(new_n6205));
  AOI22xp33_ASAP7_75t_L     g05949(.A1(new_n2114), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n2259), .Y(new_n6206));
  OAI221xp5_ASAP7_75t_L     g05950(.A1(new_n2109), .A2(new_n1539), .B1(new_n2257), .B2(new_n1662), .C(new_n6206), .Y(new_n6207));
  XNOR2x2_ASAP7_75t_L       g05951(.A(\a[26] ), .B(new_n6207), .Y(new_n6208));
  NAND3xp33_ASAP7_75t_L     g05952(.A(new_n6199), .B(new_n6208), .C(new_n6205), .Y(new_n6209));
  NOR3xp33_ASAP7_75t_L      g05953(.A(new_n6202), .B(new_n6203), .C(new_n6204), .Y(new_n6210));
  AOI21xp33_ASAP7_75t_L     g05954(.A1(new_n6198), .A2(new_n6193), .B(new_n6102), .Y(new_n6211));
  XNOR2x2_ASAP7_75t_L       g05955(.A(new_n2100), .B(new_n6207), .Y(new_n6212));
  OAI21xp33_ASAP7_75t_L     g05956(.A1(new_n6211), .A2(new_n6210), .B(new_n6212), .Y(new_n6213));
  NAND2xp33_ASAP7_75t_L     g05957(.A(new_n6209), .B(new_n6213), .Y(new_n6214));
  NAND2xp33_ASAP7_75t_L     g05958(.A(new_n5957), .B(new_n5962), .Y(new_n6215));
  MAJIxp5_ASAP7_75t_L       g05959(.A(new_n5972), .B(new_n6215), .C(new_n5965), .Y(new_n6216));
  NOR2xp33_ASAP7_75t_L      g05960(.A(new_n6216), .B(new_n6214), .Y(new_n6217));
  NOR3xp33_ASAP7_75t_L      g05961(.A(new_n6210), .B(new_n6211), .C(new_n6212), .Y(new_n6218));
  AOI21xp33_ASAP7_75t_L     g05962(.A1(new_n6199), .A2(new_n6205), .B(new_n6208), .Y(new_n6219));
  NOR2xp33_ASAP7_75t_L      g05963(.A(new_n6219), .B(new_n6218), .Y(new_n6220));
  O2A1O1Ixp33_ASAP7_75t_L   g05964(.A1(new_n6215), .A2(new_n5965), .B(new_n5986), .C(new_n6220), .Y(new_n6221));
  OAI22xp33_ASAP7_75t_L     g05965(.A1(new_n1829), .A2(new_n1774), .B1(new_n1929), .B2(new_n1696), .Y(new_n6222));
  AOI221xp5_ASAP7_75t_L     g05966(.A1(\b[23] ), .A2(new_n1706), .B1(new_n1695), .B2(new_n1935), .C(new_n6222), .Y(new_n6223));
  XNOR2x2_ASAP7_75t_L       g05967(.A(new_n1689), .B(new_n6223), .Y(new_n6224));
  OAI21xp33_ASAP7_75t_L     g05968(.A1(new_n6217), .A2(new_n6221), .B(new_n6224), .Y(new_n6225));
  OAI211xp5_ASAP7_75t_L     g05969(.A1(new_n6215), .A2(new_n5965), .B(new_n6220), .C(new_n5986), .Y(new_n6226));
  NAND2xp33_ASAP7_75t_L     g05970(.A(new_n6216), .B(new_n6214), .Y(new_n6227));
  XNOR2x2_ASAP7_75t_L       g05971(.A(\a[23] ), .B(new_n6223), .Y(new_n6228));
  NAND3xp33_ASAP7_75t_L     g05972(.A(new_n6226), .B(new_n6228), .C(new_n6227), .Y(new_n6229));
  OAI211xp5_ASAP7_75t_L     g05973(.A1(new_n5717), .A2(new_n5724), .B(new_n5996), .C(new_n5988), .Y(new_n6230));
  NAND4xp25_ASAP7_75t_L     g05974(.A(new_n6230), .B(new_n6225), .C(new_n6229), .D(new_n5981), .Y(new_n6231));
  AOI21xp33_ASAP7_75t_L     g05975(.A1(new_n6226), .A2(new_n6227), .B(new_n6228), .Y(new_n6232));
  NOR3xp33_ASAP7_75t_L      g05976(.A(new_n6221), .B(new_n6224), .C(new_n6217), .Y(new_n6233));
  AOI211xp5_ASAP7_75t_L     g05977(.A1(new_n5713), .A2(new_n5710), .B(new_n5866), .C(new_n5992), .Y(new_n6234));
  OAI22xp33_ASAP7_75t_L     g05978(.A1(new_n6234), .A2(new_n5991), .B1(new_n6233), .B2(new_n6232), .Y(new_n6235));
  NOR2xp33_ASAP7_75t_L      g05979(.A(new_n2348), .B(new_n1373), .Y(new_n6236));
  INVx1_ASAP7_75t_L         g05980(.A(new_n6236), .Y(new_n6237));
  NAND2xp33_ASAP7_75t_L     g05981(.A(new_n1365), .B(new_n2504), .Y(new_n6238));
  AOI22xp33_ASAP7_75t_L     g05982(.A1(new_n1360), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1581), .Y(new_n6239));
  AND4x1_ASAP7_75t_L        g05983(.A(new_n6239), .B(new_n6238), .C(new_n6237), .D(\a[20] ), .Y(new_n6240));
  AOI31xp33_ASAP7_75t_L     g05984(.A1(new_n6238), .A2(new_n6237), .A3(new_n6239), .B(\a[20] ), .Y(new_n6241));
  NOR2xp33_ASAP7_75t_L      g05985(.A(new_n6241), .B(new_n6240), .Y(new_n6242));
  NAND3xp33_ASAP7_75t_L     g05986(.A(new_n6235), .B(new_n6231), .C(new_n6242), .Y(new_n6243));
  AO21x2_ASAP7_75t_L        g05987(.A1(new_n6231), .A2(new_n6235), .B(new_n6242), .Y(new_n6244));
  NAND2xp33_ASAP7_75t_L     g05988(.A(new_n6243), .B(new_n6244), .Y(new_n6245));
  NAND2xp33_ASAP7_75t_L     g05989(.A(new_n6245), .B(new_n6101), .Y(new_n6246));
  A2O1A1O1Ixp25_ASAP7_75t_L g05990(.A1(new_n5729), .A2(new_n6001), .B(new_n6003), .C(new_n6004), .D(new_n5999), .Y(new_n6247));
  NAND3xp33_ASAP7_75t_L     g05991(.A(new_n6247), .B(new_n6243), .C(new_n6244), .Y(new_n6248));
  NAND3xp33_ASAP7_75t_L     g05992(.A(new_n6246), .B(new_n6099), .C(new_n6248), .Y(new_n6249));
  AOI21xp33_ASAP7_75t_L     g05993(.A1(new_n6244), .A2(new_n6243), .B(new_n6247), .Y(new_n6250));
  NOR2xp33_ASAP7_75t_L      g05994(.A(new_n6245), .B(new_n6101), .Y(new_n6251));
  OAI21xp33_ASAP7_75t_L     g05995(.A1(new_n6250), .A2(new_n6251), .B(new_n6098), .Y(new_n6252));
  NAND2xp33_ASAP7_75t_L     g05996(.A(new_n6249), .B(new_n6252), .Y(new_n6253));
  O2A1O1Ixp33_ASAP7_75t_L   g05997(.A1(new_n5856), .A2(new_n6020), .B(new_n6012), .C(new_n6253), .Y(new_n6254));
  OAI21xp33_ASAP7_75t_L     g05998(.A1(new_n6020), .A2(new_n5856), .B(new_n6012), .Y(new_n6255));
  NOR3xp33_ASAP7_75t_L      g05999(.A(new_n6251), .B(new_n6250), .C(new_n6098), .Y(new_n6256));
  AOI21xp33_ASAP7_75t_L     g06000(.A1(new_n6246), .A2(new_n6248), .B(new_n6099), .Y(new_n6257));
  NOR2xp33_ASAP7_75t_L      g06001(.A(new_n6257), .B(new_n6256), .Y(new_n6258));
  NOR2xp33_ASAP7_75t_L      g06002(.A(new_n6258), .B(new_n6255), .Y(new_n6259));
  AOI22xp33_ASAP7_75t_L     g06003(.A1(new_n811), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n900), .Y(new_n6260));
  OAI221xp5_ASAP7_75t_L     g06004(.A1(new_n904), .A2(new_n3207), .B1(new_n898), .B2(new_n3572), .C(new_n6260), .Y(new_n6261));
  XNOR2x2_ASAP7_75t_L       g06005(.A(\a[14] ), .B(new_n6261), .Y(new_n6262));
  INVx1_ASAP7_75t_L         g06006(.A(new_n6262), .Y(new_n6263));
  NOR3xp33_ASAP7_75t_L      g06007(.A(new_n6259), .B(new_n6254), .C(new_n6263), .Y(new_n6264));
  A2O1A1Ixp33_ASAP7_75t_L   g06008(.A1(new_n6007), .A2(new_n6019), .B(new_n6021), .C(new_n6258), .Y(new_n6265));
  A2O1A1O1Ixp25_ASAP7_75t_L g06009(.A1(new_n5746), .A2(new_n5598), .B(new_n5855), .C(new_n6007), .D(new_n6021), .Y(new_n6266));
  NAND2xp33_ASAP7_75t_L     g06010(.A(new_n6266), .B(new_n6253), .Y(new_n6267));
  AOI21xp33_ASAP7_75t_L     g06011(.A1(new_n6265), .A2(new_n6267), .B(new_n6262), .Y(new_n6268));
  OAI21xp33_ASAP7_75t_L     g06012(.A1(new_n6264), .A2(new_n6268), .B(new_n6091), .Y(new_n6269));
  A2O1A1O1Ixp25_ASAP7_75t_L g06013(.A1(new_n5751), .A2(new_n5596), .B(new_n6027), .C(new_n6016), .D(new_n6030), .Y(new_n6270));
  NAND3xp33_ASAP7_75t_L     g06014(.A(new_n6265), .B(new_n6267), .C(new_n6262), .Y(new_n6271));
  OAI21xp33_ASAP7_75t_L     g06015(.A1(new_n6254), .A2(new_n6259), .B(new_n6263), .Y(new_n6272));
  NAND3xp33_ASAP7_75t_L     g06016(.A(new_n6270), .B(new_n6271), .C(new_n6272), .Y(new_n6273));
  NAND3xp33_ASAP7_75t_L     g06017(.A(new_n6090), .B(new_n6273), .C(new_n6269), .Y(new_n6274));
  AO21x2_ASAP7_75t_L        g06018(.A1(new_n6269), .A2(new_n6273), .B(new_n6090), .Y(new_n6275));
  AOI221xp5_ASAP7_75t_L     g06019(.A1(new_n6046), .A2(new_n6047), .B1(new_n6274), .B2(new_n6275), .C(new_n6084), .Y(new_n6276));
  AOI21xp33_ASAP7_75t_L     g06020(.A1(new_n6046), .A2(new_n6047), .B(new_n6084), .Y(new_n6277));
  NAND2xp33_ASAP7_75t_L     g06021(.A(new_n6274), .B(new_n6275), .Y(new_n6278));
  NOR2xp33_ASAP7_75t_L      g06022(.A(new_n6278), .B(new_n6277), .Y(new_n6279));
  AOI22xp33_ASAP7_75t_L     g06023(.A1(new_n444), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n471), .Y(new_n6280));
  OAI21xp33_ASAP7_75t_L     g06024(.A1(new_n469), .A2(new_n4858), .B(new_n6280), .Y(new_n6281));
  AOI21xp33_ASAP7_75t_L     g06025(.A1(new_n447), .A2(\b[38] ), .B(new_n6281), .Y(new_n6282));
  NAND2xp33_ASAP7_75t_L     g06026(.A(\a[8] ), .B(new_n6282), .Y(new_n6283));
  A2O1A1Ixp33_ASAP7_75t_L   g06027(.A1(\b[38] ), .A2(new_n447), .B(new_n6281), .C(new_n435), .Y(new_n6284));
  NAND2xp33_ASAP7_75t_L     g06028(.A(new_n6284), .B(new_n6283), .Y(new_n6285));
  NOR3xp33_ASAP7_75t_L      g06029(.A(new_n6279), .B(new_n6285), .C(new_n6276), .Y(new_n6286));
  NAND2xp33_ASAP7_75t_L     g06030(.A(new_n6278), .B(new_n6277), .Y(new_n6287));
  AND3x1_ASAP7_75t_L        g06031(.A(new_n6273), .B(new_n6090), .C(new_n6269), .Y(new_n6288));
  AOI21xp33_ASAP7_75t_L     g06032(.A1(new_n6273), .A2(new_n6269), .B(new_n6090), .Y(new_n6289));
  NOR2xp33_ASAP7_75t_L      g06033(.A(new_n6289), .B(new_n6288), .Y(new_n6290));
  OAI21xp33_ASAP7_75t_L     g06034(.A1(new_n6084), .A2(new_n6058), .B(new_n6290), .Y(new_n6291));
  AND2x2_ASAP7_75t_L        g06035(.A(new_n6284), .B(new_n6283), .Y(new_n6292));
  AOI21xp33_ASAP7_75t_L     g06036(.A1(new_n6291), .A2(new_n6287), .B(new_n6292), .Y(new_n6293));
  NOR2xp33_ASAP7_75t_L      g06037(.A(new_n6293), .B(new_n6286), .Y(new_n6294));
  AOI21xp33_ASAP7_75t_L     g06038(.A1(new_n5793), .A2(new_n5788), .B(new_n5780), .Y(new_n6295));
  NOR3xp33_ASAP7_75t_L      g06039(.A(new_n6057), .B(new_n6058), .C(new_n6055), .Y(new_n6296));
  AOI21xp33_ASAP7_75t_L     g06040(.A1(new_n6295), .A2(new_n6063), .B(new_n6296), .Y(new_n6297));
  NAND2xp33_ASAP7_75t_L     g06041(.A(new_n6297), .B(new_n6294), .Y(new_n6298));
  NAND3xp33_ASAP7_75t_L     g06042(.A(new_n6291), .B(new_n6287), .C(new_n6292), .Y(new_n6299));
  OAI21xp33_ASAP7_75t_L     g06043(.A1(new_n6276), .A2(new_n6279), .B(new_n6285), .Y(new_n6300));
  NAND2xp33_ASAP7_75t_L     g06044(.A(new_n6299), .B(new_n6300), .Y(new_n6301));
  OAI21xp33_ASAP7_75t_L     g06045(.A1(new_n6296), .A2(new_n6061), .B(new_n6301), .Y(new_n6302));
  NOR2xp33_ASAP7_75t_L      g06046(.A(new_n5321), .B(new_n429), .Y(new_n6303));
  INVx1_ASAP7_75t_L         g06047(.A(new_n6303), .Y(new_n6304));
  NAND3xp33_ASAP7_75t_L     g06048(.A(new_n5343), .B(new_n341), .C(new_n5345), .Y(new_n6305));
  AOI22xp33_ASAP7_75t_L     g06049(.A1(new_n344), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n370), .Y(new_n6306));
  AND4x1_ASAP7_75t_L        g06050(.A(new_n6306), .B(new_n6305), .C(new_n6304), .D(\a[5] ), .Y(new_n6307));
  AOI31xp33_ASAP7_75t_L     g06051(.A1(new_n6305), .A2(new_n6304), .A3(new_n6306), .B(\a[5] ), .Y(new_n6308));
  NOR2xp33_ASAP7_75t_L      g06052(.A(new_n6308), .B(new_n6307), .Y(new_n6309));
  NAND3xp33_ASAP7_75t_L     g06053(.A(new_n6298), .B(new_n6302), .C(new_n6309), .Y(new_n6310));
  NOR4xp25_ASAP7_75t_L      g06054(.A(new_n6061), .B(new_n6296), .C(new_n6293), .D(new_n6286), .Y(new_n6311));
  NOR2xp33_ASAP7_75t_L      g06055(.A(new_n6297), .B(new_n6294), .Y(new_n6312));
  INVx1_ASAP7_75t_L         g06056(.A(new_n6309), .Y(new_n6313));
  OAI21xp33_ASAP7_75t_L     g06057(.A1(new_n6311), .A2(new_n6312), .B(new_n6313), .Y(new_n6314));
  OAI211xp5_ASAP7_75t_L     g06058(.A1(new_n5845), .A2(new_n5846), .B(new_n6071), .C(new_n6067), .Y(new_n6315));
  NAND4xp25_ASAP7_75t_L     g06059(.A(new_n6083), .B(new_n6315), .C(new_n6314), .D(new_n6310), .Y(new_n6316));
  NAND2xp33_ASAP7_75t_L     g06060(.A(new_n6310), .B(new_n6314), .Y(new_n6317));
  A2O1A1Ixp33_ASAP7_75t_L   g06061(.A1(new_n6065), .A2(new_n6072), .B(new_n5841), .C(new_n6315), .Y(new_n6318));
  NAND2xp33_ASAP7_75t_L     g06062(.A(new_n6318), .B(new_n6317), .Y(new_n6319));
  NOR2xp33_ASAP7_75t_L      g06063(.A(\b[44] ), .B(\b[45] ), .Y(new_n6320));
  INVx1_ASAP7_75t_L         g06064(.A(\b[45] ), .Y(new_n6321));
  NOR2xp33_ASAP7_75t_L      g06065(.A(new_n5829), .B(new_n6321), .Y(new_n6322));
  NOR2xp33_ASAP7_75t_L      g06066(.A(new_n6320), .B(new_n6322), .Y(new_n6323));
  INVx1_ASAP7_75t_L         g06067(.A(new_n6323), .Y(new_n6324));
  O2A1O1Ixp33_ASAP7_75t_L   g06068(.A1(new_n5805), .A2(new_n5829), .B(new_n5832), .C(new_n6324), .Y(new_n6325));
  INVx1_ASAP7_75t_L         g06069(.A(new_n6325), .Y(new_n6326));
  A2O1A1O1Ixp25_ASAP7_75t_L g06070(.A1(new_n5807), .A2(new_n5810), .B(new_n5806), .C(new_n5831), .D(new_n5830), .Y(new_n6327));
  NAND2xp33_ASAP7_75t_L     g06071(.A(new_n6324), .B(new_n6327), .Y(new_n6328));
  NAND2xp33_ASAP7_75t_L     g06072(.A(new_n6328), .B(new_n6326), .Y(new_n6329));
  AOI22xp33_ASAP7_75t_L     g06073(.A1(\b[43] ), .A2(new_n282), .B1(\b[45] ), .B2(new_n303), .Y(new_n6330));
  OAI221xp5_ASAP7_75t_L     g06074(.A1(new_n291), .A2(new_n5829), .B1(new_n268), .B2(new_n6329), .C(new_n6330), .Y(new_n6331));
  XNOR2x2_ASAP7_75t_L       g06075(.A(new_n262), .B(new_n6331), .Y(new_n6332));
  AOI21xp33_ASAP7_75t_L     g06076(.A1(new_n6316), .A2(new_n6319), .B(new_n6332), .Y(new_n6333));
  NAND3xp33_ASAP7_75t_L     g06077(.A(new_n6316), .B(new_n6319), .C(new_n6332), .Y(new_n6334));
  INVx1_ASAP7_75t_L         g06078(.A(new_n6334), .Y(new_n6335));
  NOR2xp33_ASAP7_75t_L      g06079(.A(new_n6333), .B(new_n6335), .Y(new_n6336));
  XNOR2x2_ASAP7_75t_L       g06080(.A(new_n6082), .B(new_n6336), .Y(\f[45] ));
  INVx1_ASAP7_75t_L         g06081(.A(new_n5812), .Y(new_n6338));
  AOI22xp33_ASAP7_75t_L     g06082(.A1(new_n344), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n370), .Y(new_n6339));
  OAI21xp33_ASAP7_75t_L     g06083(.A1(new_n366), .A2(new_n6338), .B(new_n6339), .Y(new_n6340));
  AOI21xp33_ASAP7_75t_L     g06084(.A1(new_n347), .A2(\b[42] ), .B(new_n6340), .Y(new_n6341));
  NAND2xp33_ASAP7_75t_L     g06085(.A(\a[5] ), .B(new_n6341), .Y(new_n6342));
  A2O1A1Ixp33_ASAP7_75t_L   g06086(.A1(\b[42] ), .A2(new_n347), .B(new_n6340), .C(new_n338), .Y(new_n6343));
  AND2x2_ASAP7_75t_L        g06087(.A(new_n6343), .B(new_n6342), .Y(new_n6344));
  NOR3xp33_ASAP7_75t_L      g06088(.A(new_n6279), .B(new_n6292), .C(new_n6276), .Y(new_n6345));
  O2A1O1Ixp33_ASAP7_75t_L   g06089(.A1(new_n6061), .A2(new_n6296), .B(new_n6301), .C(new_n6345), .Y(new_n6346));
  OAI21xp33_ASAP7_75t_L     g06090(.A1(new_n6257), .A2(new_n6266), .B(new_n6249), .Y(new_n6347));
  OAI211xp5_ASAP7_75t_L     g06091(.A1(new_n6240), .A2(new_n6241), .B(new_n6235), .C(new_n6231), .Y(new_n6348));
  INVx1_ASAP7_75t_L         g06092(.A(new_n6348), .Y(new_n6349));
  AOI22xp33_ASAP7_75t_L     g06093(.A1(new_n1360), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n1581), .Y(new_n6350));
  INVx1_ASAP7_75t_L         g06094(.A(new_n6350), .Y(new_n6351));
  AOI221xp5_ASAP7_75t_L     g06095(.A1(\b[27] ), .A2(new_n1362), .B1(new_n1365), .B2(new_n4237), .C(new_n6351), .Y(new_n6352));
  XNOR2x2_ASAP7_75t_L       g06096(.A(new_n1356), .B(new_n6352), .Y(new_n6353));
  NAND2xp33_ASAP7_75t_L     g06097(.A(new_n6182), .B(new_n6181), .Y(new_n6354));
  NAND2xp33_ASAP7_75t_L     g06098(.A(new_n6172), .B(new_n6167), .Y(new_n6355));
  NOR2xp33_ASAP7_75t_L      g06099(.A(new_n6111), .B(new_n6355), .Y(new_n6356));
  AOI22xp33_ASAP7_75t_L     g06100(.A1(new_n3633), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n3858), .Y(new_n6357));
  OAI221xp5_ASAP7_75t_L     g06101(.A1(new_n3853), .A2(new_n760), .B1(new_n3856), .B2(new_n790), .C(new_n6357), .Y(new_n6358));
  XNOR2x2_ASAP7_75t_L       g06102(.A(\a[35] ), .B(new_n6358), .Y(new_n6359));
  A2O1A1Ixp33_ASAP7_75t_L   g06103(.A1(new_n5923), .A2(new_n5924), .B(new_n5922), .C(new_n6175), .Y(new_n6360));
  NOR3xp33_ASAP7_75t_L      g06104(.A(new_n5903), .B(new_n6121), .C(new_n6114), .Y(new_n6361));
  NAND2xp33_ASAP7_75t_L     g06105(.A(\b[3] ), .B(new_n5628), .Y(new_n6362));
  NAND2xp33_ASAP7_75t_L     g06106(.A(new_n5621), .B(new_n329), .Y(new_n6363));
  AOI22xp33_ASAP7_75t_L     g06107(.A1(new_n5624), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n5901), .Y(new_n6364));
  NAND4xp25_ASAP7_75t_L     g06108(.A(new_n6363), .B(\a[44] ), .C(new_n6362), .D(new_n6364), .Y(new_n6365));
  AOI31xp33_ASAP7_75t_L     g06109(.A1(new_n6363), .A2(new_n6362), .A3(new_n6364), .B(\a[44] ), .Y(new_n6366));
  INVx1_ASAP7_75t_L         g06110(.A(new_n6366), .Y(new_n6367));
  NAND2xp33_ASAP7_75t_L     g06111(.A(\a[47] ), .B(new_n6120), .Y(new_n6368));
  INVx1_ASAP7_75t_L         g06112(.A(\a[46] ), .Y(new_n6369));
  NAND2xp33_ASAP7_75t_L     g06113(.A(\a[47] ), .B(new_n6369), .Y(new_n6370));
  INVx1_ASAP7_75t_L         g06114(.A(\a[47] ), .Y(new_n6371));
  NAND2xp33_ASAP7_75t_L     g06115(.A(\a[46] ), .B(new_n6371), .Y(new_n6372));
  AOI21xp33_ASAP7_75t_L     g06116(.A1(new_n6372), .A2(new_n6370), .B(new_n6119), .Y(new_n6373));
  NAND2xp33_ASAP7_75t_L     g06117(.A(new_n269), .B(new_n6373), .Y(new_n6374));
  NAND2xp33_ASAP7_75t_L     g06118(.A(new_n6372), .B(new_n6370), .Y(new_n6375));
  NOR2xp33_ASAP7_75t_L      g06119(.A(new_n6375), .B(new_n6119), .Y(new_n6376));
  NAND2xp33_ASAP7_75t_L     g06120(.A(\b[1] ), .B(new_n6376), .Y(new_n6377));
  NAND2xp33_ASAP7_75t_L     g06121(.A(new_n6118), .B(new_n6117), .Y(new_n6378));
  XNOR2x2_ASAP7_75t_L       g06122(.A(\a[46] ), .B(\a[45] ), .Y(new_n6379));
  NOR2xp33_ASAP7_75t_L      g06123(.A(new_n6379), .B(new_n6378), .Y(new_n6380));
  NAND2xp33_ASAP7_75t_L     g06124(.A(\b[0] ), .B(new_n6380), .Y(new_n6381));
  NAND3xp33_ASAP7_75t_L     g06125(.A(new_n6374), .B(new_n6377), .C(new_n6381), .Y(new_n6382));
  XOR2x2_ASAP7_75t_L        g06126(.A(new_n6368), .B(new_n6382), .Y(new_n6383));
  NAND3xp33_ASAP7_75t_L     g06127(.A(new_n6367), .B(new_n6383), .C(new_n6365), .Y(new_n6384));
  INVx1_ASAP7_75t_L         g06128(.A(new_n6365), .Y(new_n6385));
  XNOR2x2_ASAP7_75t_L       g06129(.A(new_n6368), .B(new_n6382), .Y(new_n6386));
  OAI21xp33_ASAP7_75t_L     g06130(.A1(new_n6366), .A2(new_n6385), .B(new_n6386), .Y(new_n6387));
  OAI211xp5_ASAP7_75t_L     g06131(.A1(new_n6361), .A2(new_n6144), .B(new_n6384), .C(new_n6387), .Y(new_n6388));
  O2A1O1Ixp33_ASAP7_75t_L   g06132(.A1(new_n6122), .A2(new_n6123), .B(new_n6130), .C(new_n6361), .Y(new_n6389));
  NOR3xp33_ASAP7_75t_L      g06133(.A(new_n6386), .B(new_n6385), .C(new_n6366), .Y(new_n6390));
  AOI21xp33_ASAP7_75t_L     g06134(.A1(new_n6367), .A2(new_n6365), .B(new_n6383), .Y(new_n6391));
  OAI21xp33_ASAP7_75t_L     g06135(.A1(new_n6390), .A2(new_n6391), .B(new_n6389), .Y(new_n6392));
  AOI22xp33_ASAP7_75t_L     g06136(.A1(new_n4920), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n5167), .Y(new_n6393));
  OAI221xp5_ASAP7_75t_L     g06137(.A1(new_n5154), .A2(new_n418), .B1(new_n5158), .B2(new_n425), .C(new_n6393), .Y(new_n6394));
  XNOR2x2_ASAP7_75t_L       g06138(.A(\a[41] ), .B(new_n6394), .Y(new_n6395));
  NAND3xp33_ASAP7_75t_L     g06139(.A(new_n6388), .B(new_n6392), .C(new_n6395), .Y(new_n6396));
  NOR3xp33_ASAP7_75t_L      g06140(.A(new_n6389), .B(new_n6390), .C(new_n6391), .Y(new_n6397));
  AOI211xp5_ASAP7_75t_L     g06141(.A1(new_n6384), .A2(new_n6387), .B(new_n6361), .C(new_n6144), .Y(new_n6398));
  XNOR2x2_ASAP7_75t_L       g06142(.A(new_n4915), .B(new_n6394), .Y(new_n6399));
  OAI21xp33_ASAP7_75t_L     g06143(.A1(new_n6397), .A2(new_n6398), .B(new_n6399), .Y(new_n6400));
  NAND2xp33_ASAP7_75t_L     g06144(.A(new_n6400), .B(new_n6396), .Y(new_n6401));
  AOI211xp5_ASAP7_75t_L     g06145(.A1(new_n6140), .A2(new_n6142), .B(new_n6145), .C(new_n6144), .Y(new_n6402));
  INVx1_ASAP7_75t_L         g06146(.A(new_n6402), .Y(new_n6403));
  A2O1A1Ixp33_ASAP7_75t_L   g06147(.A1(new_n6147), .A2(new_n6143), .B(new_n6149), .C(new_n6403), .Y(new_n6404));
  NOR2xp33_ASAP7_75t_L      g06148(.A(new_n6404), .B(new_n6401), .Y(new_n6405));
  AOI21xp33_ASAP7_75t_L     g06149(.A1(new_n6151), .A2(new_n6162), .B(new_n6402), .Y(new_n6406));
  AOI21xp33_ASAP7_75t_L     g06150(.A1(new_n6400), .A2(new_n6396), .B(new_n6406), .Y(new_n6407));
  AOI22xp33_ASAP7_75t_L     g06151(.A1(new_n4283), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n4512), .Y(new_n6408));
  OAI221xp5_ASAP7_75t_L     g06152(.A1(new_n4277), .A2(new_n540), .B1(new_n4499), .B2(new_n624), .C(new_n6408), .Y(new_n6409));
  XNOR2x2_ASAP7_75t_L       g06153(.A(\a[38] ), .B(new_n6409), .Y(new_n6410));
  OAI21xp33_ASAP7_75t_L     g06154(.A1(new_n6407), .A2(new_n6405), .B(new_n6410), .Y(new_n6411));
  NAND3xp33_ASAP7_75t_L     g06155(.A(new_n6406), .B(new_n6400), .C(new_n6396), .Y(new_n6412));
  A2O1A1Ixp33_ASAP7_75t_L   g06156(.A1(new_n6151), .A2(new_n6162), .B(new_n6402), .C(new_n6401), .Y(new_n6413));
  INVx1_ASAP7_75t_L         g06157(.A(new_n6410), .Y(new_n6414));
  NAND3xp33_ASAP7_75t_L     g06158(.A(new_n6414), .B(new_n6413), .C(new_n6412), .Y(new_n6415));
  AOI221xp5_ASAP7_75t_L     g06159(.A1(new_n6415), .A2(new_n6411), .B1(new_n6166), .B2(new_n6360), .C(new_n6165), .Y(new_n6416));
  A2O1A1O1Ixp25_ASAP7_75t_L g06160(.A1(new_n5925), .A2(new_n6112), .B(new_n6113), .C(new_n6169), .D(new_n6165), .Y(new_n6417));
  AOI21xp33_ASAP7_75t_L     g06161(.A1(new_n6413), .A2(new_n6412), .B(new_n6414), .Y(new_n6418));
  NOR3xp33_ASAP7_75t_L      g06162(.A(new_n6405), .B(new_n6407), .C(new_n6410), .Y(new_n6419));
  NOR3xp33_ASAP7_75t_L      g06163(.A(new_n6417), .B(new_n6418), .C(new_n6419), .Y(new_n6420));
  OA21x2_ASAP7_75t_L        g06164(.A1(new_n6420), .A2(new_n6416), .B(new_n6359), .Y(new_n6421));
  NOR3xp33_ASAP7_75t_L      g06165(.A(new_n6416), .B(new_n6420), .C(new_n6359), .Y(new_n6422));
  NOR2xp33_ASAP7_75t_L      g06166(.A(new_n6422), .B(new_n6421), .Y(new_n6423));
  A2O1A1Ixp33_ASAP7_75t_L   g06167(.A1(new_n6354), .A2(new_n6108), .B(new_n6356), .C(new_n6423), .Y(new_n6424));
  OAI21xp33_ASAP7_75t_L     g06168(.A1(new_n6420), .A2(new_n6416), .B(new_n6359), .Y(new_n6425));
  OR3x1_ASAP7_75t_L         g06169(.A(new_n6416), .B(new_n6359), .C(new_n6420), .Y(new_n6426));
  NAND2xp33_ASAP7_75t_L     g06170(.A(new_n6425), .B(new_n6426), .Y(new_n6427));
  OAI211xp5_ASAP7_75t_L     g06171(.A1(new_n6111), .A2(new_n6355), .B(new_n6427), .C(new_n6179), .Y(new_n6428));
  AOI22xp33_ASAP7_75t_L     g06172(.A1(new_n3029), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n3258), .Y(new_n6429));
  OAI221xp5_ASAP7_75t_L     g06173(.A1(new_n3024), .A2(new_n942), .B1(new_n3256), .B2(new_n1035), .C(new_n6429), .Y(new_n6430));
  XNOR2x2_ASAP7_75t_L       g06174(.A(\a[32] ), .B(new_n6430), .Y(new_n6431));
  NAND3xp33_ASAP7_75t_L     g06175(.A(new_n6428), .B(new_n6424), .C(new_n6431), .Y(new_n6432));
  O2A1O1Ixp33_ASAP7_75t_L   g06176(.A1(new_n6111), .A2(new_n6355), .B(new_n6179), .C(new_n6427), .Y(new_n6433));
  MAJIxp5_ASAP7_75t_L       g06177(.A(new_n6180), .B(new_n6111), .C(new_n6355), .Y(new_n6434));
  NOR2xp33_ASAP7_75t_L      g06178(.A(new_n6434), .B(new_n6423), .Y(new_n6435));
  INVx1_ASAP7_75t_L         g06179(.A(new_n6431), .Y(new_n6436));
  OAI21xp33_ASAP7_75t_L     g06180(.A1(new_n6435), .A2(new_n6433), .B(new_n6436), .Y(new_n6437));
  NAND2xp33_ASAP7_75t_L     g06181(.A(new_n6183), .B(new_n6179), .Y(new_n6438));
  NOR2xp33_ASAP7_75t_L      g06182(.A(new_n6106), .B(new_n6438), .Y(new_n6439));
  INVx1_ASAP7_75t_L         g06183(.A(new_n6439), .Y(new_n6440));
  OAI21xp33_ASAP7_75t_L     g06184(.A1(new_n6184), .A2(new_n6185), .B(new_n6194), .Y(new_n6441));
  NAND4xp25_ASAP7_75t_L     g06185(.A(new_n6441), .B(new_n6432), .C(new_n6437), .D(new_n6440), .Y(new_n6442));
  NOR3xp33_ASAP7_75t_L      g06186(.A(new_n6433), .B(new_n6435), .C(new_n6436), .Y(new_n6443));
  AOI21xp33_ASAP7_75t_L     g06187(.A1(new_n6428), .A2(new_n6424), .B(new_n6431), .Y(new_n6444));
  MAJIxp5_ASAP7_75t_L       g06188(.A(new_n6103), .B(new_n6106), .C(new_n6438), .Y(new_n6445));
  OAI21xp33_ASAP7_75t_L     g06189(.A1(new_n6443), .A2(new_n6444), .B(new_n6445), .Y(new_n6446));
  AOI22xp33_ASAP7_75t_L     g06190(.A1(new_n2552), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n2736), .Y(new_n6447));
  OAI221xp5_ASAP7_75t_L     g06191(.A1(new_n2547), .A2(new_n1313), .B1(new_n2734), .B2(new_n1438), .C(new_n6447), .Y(new_n6448));
  XNOR2x2_ASAP7_75t_L       g06192(.A(\a[29] ), .B(new_n6448), .Y(new_n6449));
  NAND3xp33_ASAP7_75t_L     g06193(.A(new_n6442), .B(new_n6446), .C(new_n6449), .Y(new_n6450));
  AO21x2_ASAP7_75t_L        g06194(.A1(new_n6446), .A2(new_n6442), .B(new_n6449), .Y(new_n6451));
  A2O1A1O1Ixp25_ASAP7_75t_L g06195(.A1(new_n5949), .A2(new_n5868), .B(new_n5961), .C(new_n6198), .D(new_n6203), .Y(new_n6452));
  NAND3xp33_ASAP7_75t_L     g06196(.A(new_n6452), .B(new_n6451), .C(new_n6450), .Y(new_n6453));
  AO21x2_ASAP7_75t_L        g06197(.A1(new_n6450), .A2(new_n6451), .B(new_n6452), .Y(new_n6454));
  NAND2xp33_ASAP7_75t_L     g06198(.A(\b[21] ), .B(new_n2115), .Y(new_n6455));
  NAND2xp33_ASAP7_75t_L     g06199(.A(new_n2106), .B(new_n3728), .Y(new_n6456));
  AOI22xp33_ASAP7_75t_L     g06200(.A1(new_n2114), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n2259), .Y(new_n6457));
  AND4x1_ASAP7_75t_L        g06201(.A(new_n6457), .B(new_n6456), .C(new_n6455), .D(\a[26] ), .Y(new_n6458));
  AOI31xp33_ASAP7_75t_L     g06202(.A1(new_n6456), .A2(new_n6455), .A3(new_n6457), .B(\a[26] ), .Y(new_n6459));
  NOR2xp33_ASAP7_75t_L      g06203(.A(new_n6459), .B(new_n6458), .Y(new_n6460));
  NAND3xp33_ASAP7_75t_L     g06204(.A(new_n6454), .B(new_n6453), .C(new_n6460), .Y(new_n6461));
  AND3x1_ASAP7_75t_L        g06205(.A(new_n6452), .B(new_n6451), .C(new_n6450), .Y(new_n6462));
  AOI21xp33_ASAP7_75t_L     g06206(.A1(new_n6451), .A2(new_n6450), .B(new_n6452), .Y(new_n6463));
  OR2x4_ASAP7_75t_L         g06207(.A(new_n6459), .B(new_n6458), .Y(new_n6464));
  OAI21xp33_ASAP7_75t_L     g06208(.A1(new_n6463), .A2(new_n6462), .B(new_n6464), .Y(new_n6465));
  NAND2xp33_ASAP7_75t_L     g06209(.A(new_n6461), .B(new_n6465), .Y(new_n6466));
  NOR3xp33_ASAP7_75t_L      g06210(.A(new_n6210), .B(new_n6211), .C(new_n6208), .Y(new_n6467));
  AOI211xp5_ASAP7_75t_L     g06211(.A1(new_n6216), .A2(new_n6214), .B(new_n6467), .C(new_n6466), .Y(new_n6468));
  NOR3xp33_ASAP7_75t_L      g06212(.A(new_n6462), .B(new_n6464), .C(new_n6463), .Y(new_n6469));
  AOI21xp33_ASAP7_75t_L     g06213(.A1(new_n6454), .A2(new_n6453), .B(new_n6460), .Y(new_n6470));
  NOR2xp33_ASAP7_75t_L      g06214(.A(new_n6470), .B(new_n6469), .Y(new_n6471));
  O2A1O1Ixp33_ASAP7_75t_L   g06215(.A1(new_n6218), .A2(new_n6219), .B(new_n6216), .C(new_n6467), .Y(new_n6472));
  NOR2xp33_ASAP7_75t_L      g06216(.A(new_n6471), .B(new_n6472), .Y(new_n6473));
  OAI22xp33_ASAP7_75t_L     g06217(.A1(new_n1829), .A2(new_n1909), .B1(new_n2067), .B2(new_n1696), .Y(new_n6474));
  AOI221xp5_ASAP7_75t_L     g06218(.A1(\b[24] ), .A2(new_n1706), .B1(new_n1695), .B2(new_n2648), .C(new_n6474), .Y(new_n6475));
  XNOR2x2_ASAP7_75t_L       g06219(.A(\a[23] ), .B(new_n6475), .Y(new_n6476));
  NOR3xp33_ASAP7_75t_L      g06220(.A(new_n6468), .B(new_n6473), .C(new_n6476), .Y(new_n6477));
  NAND2xp33_ASAP7_75t_L     g06221(.A(new_n6471), .B(new_n6472), .Y(new_n6478));
  A2O1A1Ixp33_ASAP7_75t_L   g06222(.A1(new_n6214), .A2(new_n6216), .B(new_n6467), .C(new_n6466), .Y(new_n6479));
  XNOR2x2_ASAP7_75t_L       g06223(.A(new_n1689), .B(new_n6475), .Y(new_n6480));
  AOI21xp33_ASAP7_75t_L     g06224(.A1(new_n6478), .A2(new_n6479), .B(new_n6480), .Y(new_n6481));
  OAI31xp33_ASAP7_75t_L     g06225(.A1(new_n6234), .A2(new_n6232), .A3(new_n5991), .B(new_n6229), .Y(new_n6482));
  OAI21xp33_ASAP7_75t_L     g06226(.A1(new_n6477), .A2(new_n6481), .B(new_n6482), .Y(new_n6483));
  NAND3xp33_ASAP7_75t_L     g06227(.A(new_n6478), .B(new_n6479), .C(new_n6480), .Y(new_n6484));
  OAI21xp33_ASAP7_75t_L     g06228(.A1(new_n6473), .A2(new_n6468), .B(new_n6476), .Y(new_n6485));
  AOI31xp33_ASAP7_75t_L     g06229(.A1(new_n6230), .A2(new_n6225), .A3(new_n5981), .B(new_n6233), .Y(new_n6486));
  NAND3xp33_ASAP7_75t_L     g06230(.A(new_n6486), .B(new_n6485), .C(new_n6484), .Y(new_n6487));
  AOI21xp33_ASAP7_75t_L     g06231(.A1(new_n6487), .A2(new_n6483), .B(new_n6353), .Y(new_n6488));
  XNOR2x2_ASAP7_75t_L       g06232(.A(\a[20] ), .B(new_n6352), .Y(new_n6489));
  AOI21xp33_ASAP7_75t_L     g06233(.A1(new_n6485), .A2(new_n6484), .B(new_n6486), .Y(new_n6490));
  NOR3xp33_ASAP7_75t_L      g06234(.A(new_n6482), .B(new_n6481), .C(new_n6477), .Y(new_n6491));
  NOR3xp33_ASAP7_75t_L      g06235(.A(new_n6491), .B(new_n6489), .C(new_n6490), .Y(new_n6492));
  NOR2xp33_ASAP7_75t_L      g06236(.A(new_n6488), .B(new_n6492), .Y(new_n6493));
  A2O1A1Ixp33_ASAP7_75t_L   g06237(.A1(new_n6245), .A2(new_n6101), .B(new_n6349), .C(new_n6493), .Y(new_n6494));
  A2O1A1O1Ixp25_ASAP7_75t_L g06238(.A1(new_n6004), .A2(new_n6009), .B(new_n5999), .C(new_n6245), .D(new_n6349), .Y(new_n6495));
  OAI21xp33_ASAP7_75t_L     g06239(.A1(new_n6490), .A2(new_n6491), .B(new_n6489), .Y(new_n6496));
  NAND3xp33_ASAP7_75t_L     g06240(.A(new_n6487), .B(new_n6483), .C(new_n6353), .Y(new_n6497));
  NAND2xp33_ASAP7_75t_L     g06241(.A(new_n6497), .B(new_n6496), .Y(new_n6498));
  NAND2xp33_ASAP7_75t_L     g06242(.A(new_n6498), .B(new_n6495), .Y(new_n6499));
  AOI22xp33_ASAP7_75t_L     g06243(.A1(new_n1076), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1253), .Y(new_n6500));
  OAI221xp5_ASAP7_75t_L     g06244(.A1(new_n1154), .A2(new_n2982), .B1(new_n1156), .B2(new_n3187), .C(new_n6500), .Y(new_n6501));
  XNOR2x2_ASAP7_75t_L       g06245(.A(\a[17] ), .B(new_n6501), .Y(new_n6502));
  NAND3xp33_ASAP7_75t_L     g06246(.A(new_n6499), .B(new_n6494), .C(new_n6502), .Y(new_n6503));
  NAND2xp33_ASAP7_75t_L     g06247(.A(new_n6231), .B(new_n6235), .Y(new_n6504));
  O2A1O1Ixp33_ASAP7_75t_L   g06248(.A1(new_n6504), .A2(new_n6242), .B(new_n6246), .C(new_n6498), .Y(new_n6505));
  A2O1A1Ixp33_ASAP7_75t_L   g06249(.A1(new_n6243), .A2(new_n6244), .B(new_n6247), .C(new_n6348), .Y(new_n6506));
  NOR2xp33_ASAP7_75t_L      g06250(.A(new_n6506), .B(new_n6493), .Y(new_n6507));
  INVx1_ASAP7_75t_L         g06251(.A(new_n6502), .Y(new_n6508));
  OAI21xp33_ASAP7_75t_L     g06252(.A1(new_n6507), .A2(new_n6505), .B(new_n6508), .Y(new_n6509));
  NAND3xp33_ASAP7_75t_L     g06253(.A(new_n6347), .B(new_n6503), .C(new_n6509), .Y(new_n6510));
  A2O1A1O1Ixp25_ASAP7_75t_L g06254(.A1(new_n6022), .A2(new_n6019), .B(new_n6021), .C(new_n6252), .D(new_n6256), .Y(new_n6511));
  NAND2xp33_ASAP7_75t_L     g06255(.A(new_n6509), .B(new_n6503), .Y(new_n6512));
  NAND2xp33_ASAP7_75t_L     g06256(.A(new_n6511), .B(new_n6512), .Y(new_n6513));
  AOI22xp33_ASAP7_75t_L     g06257(.A1(new_n811), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n900), .Y(new_n6514));
  OAI221xp5_ASAP7_75t_L     g06258(.A1(new_n904), .A2(new_n3565), .B1(new_n898), .B2(new_n3591), .C(new_n6514), .Y(new_n6515));
  XNOR2x2_ASAP7_75t_L       g06259(.A(\a[14] ), .B(new_n6515), .Y(new_n6516));
  NAND3xp33_ASAP7_75t_L     g06260(.A(new_n6513), .B(new_n6510), .C(new_n6516), .Y(new_n6517));
  O2A1O1Ixp33_ASAP7_75t_L   g06261(.A1(new_n6266), .A2(new_n6257), .B(new_n6249), .C(new_n6512), .Y(new_n6518));
  AOI21xp33_ASAP7_75t_L     g06262(.A1(new_n6509), .A2(new_n6503), .B(new_n6347), .Y(new_n6519));
  INVx1_ASAP7_75t_L         g06263(.A(new_n6516), .Y(new_n6520));
  OAI21xp33_ASAP7_75t_L     g06264(.A1(new_n6519), .A2(new_n6518), .B(new_n6520), .Y(new_n6521));
  NOR2xp33_ASAP7_75t_L      g06265(.A(new_n6254), .B(new_n6259), .Y(new_n6522));
  NAND2xp33_ASAP7_75t_L     g06266(.A(new_n6263), .B(new_n6522), .Y(new_n6523));
  NAND4xp25_ASAP7_75t_L     g06267(.A(new_n6269), .B(new_n6521), .C(new_n6523), .D(new_n6517), .Y(new_n6524));
  NOR3xp33_ASAP7_75t_L      g06268(.A(new_n6518), .B(new_n6519), .C(new_n6520), .Y(new_n6525));
  AOI21xp33_ASAP7_75t_L     g06269(.A1(new_n6513), .A2(new_n6510), .B(new_n6516), .Y(new_n6526));
  NAND2xp33_ASAP7_75t_L     g06270(.A(new_n6267), .B(new_n6265), .Y(new_n6527));
  MAJIxp5_ASAP7_75t_L       g06271(.A(new_n6270), .B(new_n6262), .C(new_n6527), .Y(new_n6528));
  OAI21xp33_ASAP7_75t_L     g06272(.A1(new_n6525), .A2(new_n6526), .B(new_n6528), .Y(new_n6529));
  AOI22xp33_ASAP7_75t_L     g06273(.A1(\b[35] ), .A2(new_n651), .B1(\b[37] ), .B2(new_n581), .Y(new_n6530));
  OAI221xp5_ASAP7_75t_L     g06274(.A1(new_n821), .A2(new_n4216), .B1(new_n577), .B2(new_n4431), .C(new_n6530), .Y(new_n6531));
  XNOR2x2_ASAP7_75t_L       g06275(.A(\a[11] ), .B(new_n6531), .Y(new_n6532));
  NAND3xp33_ASAP7_75t_L     g06276(.A(new_n6529), .B(new_n6524), .C(new_n6532), .Y(new_n6533));
  AO21x2_ASAP7_75t_L        g06277(.A1(new_n6524), .A2(new_n6529), .B(new_n6532), .Y(new_n6534));
  A2O1A1O1Ixp25_ASAP7_75t_L g06278(.A1(new_n6047), .A2(new_n6046), .B(new_n6084), .C(new_n6275), .D(new_n6288), .Y(new_n6535));
  NAND3xp33_ASAP7_75t_L     g06279(.A(new_n6535), .B(new_n6534), .C(new_n6533), .Y(new_n6536));
  AO21x2_ASAP7_75t_L        g06280(.A1(new_n6533), .A2(new_n6534), .B(new_n6535), .Y(new_n6537));
  NAND2xp33_ASAP7_75t_L     g06281(.A(\b[39] ), .B(new_n447), .Y(new_n6538));
  NAND2xp33_ASAP7_75t_L     g06282(.A(new_n441), .B(new_n4876), .Y(new_n6539));
  AOI22xp33_ASAP7_75t_L     g06283(.A1(new_n444), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n471), .Y(new_n6540));
  NAND4xp25_ASAP7_75t_L     g06284(.A(new_n6539), .B(\a[8] ), .C(new_n6538), .D(new_n6540), .Y(new_n6541));
  NAND2xp33_ASAP7_75t_L     g06285(.A(new_n6540), .B(new_n6539), .Y(new_n6542));
  A2O1A1Ixp33_ASAP7_75t_L   g06286(.A1(\b[39] ), .A2(new_n447), .B(new_n6542), .C(new_n435), .Y(new_n6543));
  NAND2xp33_ASAP7_75t_L     g06287(.A(new_n6541), .B(new_n6543), .Y(new_n6544));
  NAND3xp33_ASAP7_75t_L     g06288(.A(new_n6537), .B(new_n6536), .C(new_n6544), .Y(new_n6545));
  AO21x2_ASAP7_75t_L        g06289(.A1(new_n6536), .A2(new_n6537), .B(new_n6544), .Y(new_n6546));
  NAND2xp33_ASAP7_75t_L     g06290(.A(new_n6545), .B(new_n6546), .Y(new_n6547));
  NAND2xp33_ASAP7_75t_L     g06291(.A(new_n6547), .B(new_n6346), .Y(new_n6548));
  OAI31xp33_ASAP7_75t_L     g06292(.A1(new_n5566), .A2(new_n5595), .A3(new_n5783), .B(new_n5787), .Y(new_n6549));
  INVx1_ASAP7_75t_L         g06293(.A(new_n6296), .Y(new_n6550));
  OAI21xp33_ASAP7_75t_L     g06294(.A1(new_n6070), .A2(new_n6549), .B(new_n6550), .Y(new_n6551));
  AND3x1_ASAP7_75t_L        g06295(.A(new_n6537), .B(new_n6544), .C(new_n6536), .Y(new_n6552));
  AOI21xp33_ASAP7_75t_L     g06296(.A1(new_n6537), .A2(new_n6536), .B(new_n6544), .Y(new_n6553));
  NOR2xp33_ASAP7_75t_L      g06297(.A(new_n6553), .B(new_n6552), .Y(new_n6554));
  A2O1A1Ixp33_ASAP7_75t_L   g06298(.A1(new_n6551), .A2(new_n6301), .B(new_n6345), .C(new_n6554), .Y(new_n6555));
  NAND3xp33_ASAP7_75t_L     g06299(.A(new_n6555), .B(new_n6548), .C(new_n6344), .Y(new_n6556));
  NAND2xp33_ASAP7_75t_L     g06300(.A(new_n6343), .B(new_n6342), .Y(new_n6557));
  INVx1_ASAP7_75t_L         g06301(.A(new_n6345), .Y(new_n6558));
  OAI21xp33_ASAP7_75t_L     g06302(.A1(new_n6297), .A2(new_n6294), .B(new_n6558), .Y(new_n6559));
  NOR2xp33_ASAP7_75t_L      g06303(.A(new_n6554), .B(new_n6559), .Y(new_n6560));
  O2A1O1Ixp33_ASAP7_75t_L   g06304(.A1(new_n6294), .A2(new_n6297), .B(new_n6558), .C(new_n6547), .Y(new_n6561));
  OAI21xp33_ASAP7_75t_L     g06305(.A1(new_n6560), .A2(new_n6561), .B(new_n6557), .Y(new_n6562));
  NAND2xp33_ASAP7_75t_L     g06306(.A(new_n6556), .B(new_n6562), .Y(new_n6563));
  NOR3xp33_ASAP7_75t_L      g06307(.A(new_n6312), .B(new_n6309), .C(new_n6311), .Y(new_n6564));
  AOI21xp33_ASAP7_75t_L     g06308(.A1(new_n6317), .A2(new_n6318), .B(new_n6564), .Y(new_n6565));
  XNOR2x2_ASAP7_75t_L       g06309(.A(new_n6565), .B(new_n6563), .Y(new_n6566));
  NOR2xp33_ASAP7_75t_L      g06310(.A(\b[45] ), .B(\b[46] ), .Y(new_n6567));
  INVx1_ASAP7_75t_L         g06311(.A(\b[46] ), .Y(new_n6568));
  NOR2xp33_ASAP7_75t_L      g06312(.A(new_n6321), .B(new_n6568), .Y(new_n6569));
  NOR2xp33_ASAP7_75t_L      g06313(.A(new_n6567), .B(new_n6569), .Y(new_n6570));
  A2O1A1Ixp33_ASAP7_75t_L   g06314(.A1(\b[45] ), .A2(\b[44] ), .B(new_n6325), .C(new_n6570), .Y(new_n6571));
  OR3x1_ASAP7_75t_L         g06315(.A(new_n6325), .B(new_n6322), .C(new_n6570), .Y(new_n6572));
  NAND2xp33_ASAP7_75t_L     g06316(.A(new_n6571), .B(new_n6572), .Y(new_n6573));
  AOI22xp33_ASAP7_75t_L     g06317(.A1(\b[44] ), .A2(new_n282), .B1(\b[46] ), .B2(new_n303), .Y(new_n6574));
  OAI221xp5_ASAP7_75t_L     g06318(.A1(new_n291), .A2(new_n6321), .B1(new_n268), .B2(new_n6573), .C(new_n6574), .Y(new_n6575));
  XNOR2x2_ASAP7_75t_L       g06319(.A(new_n262), .B(new_n6575), .Y(new_n6576));
  XNOR2x2_ASAP7_75t_L       g06320(.A(new_n6576), .B(new_n6566), .Y(new_n6577));
  O2A1O1Ixp33_ASAP7_75t_L   g06321(.A1(new_n6082), .A2(new_n6333), .B(new_n6334), .C(new_n6577), .Y(new_n6578));
  INVx1_ASAP7_75t_L         g06322(.A(new_n6577), .Y(new_n6579));
  OAI21xp33_ASAP7_75t_L     g06323(.A1(new_n6333), .A2(new_n6082), .B(new_n6334), .Y(new_n6580));
  NOR2xp33_ASAP7_75t_L      g06324(.A(new_n6580), .B(new_n6579), .Y(new_n6581));
  NOR2xp33_ASAP7_75t_L      g06325(.A(new_n6578), .B(new_n6581), .Y(\f[46] ));
  NAND3xp33_ASAP7_75t_L     g06326(.A(new_n6555), .B(new_n6548), .C(new_n6557), .Y(new_n6583));
  A2O1A1Ixp33_ASAP7_75t_L   g06327(.A1(new_n6562), .A2(new_n6556), .B(new_n6565), .C(new_n6583), .Y(new_n6584));
  AOI22xp33_ASAP7_75t_L     g06328(.A1(new_n344), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n370), .Y(new_n6585));
  OAI221xp5_ASAP7_75t_L     g06329(.A1(new_n429), .A2(new_n5805), .B1(new_n366), .B2(new_n5835), .C(new_n6585), .Y(new_n6586));
  XNOR2x2_ASAP7_75t_L       g06330(.A(\a[5] ), .B(new_n6586), .Y(new_n6587));
  INVx1_ASAP7_75t_L         g06331(.A(new_n6587), .Y(new_n6588));
  NOR3xp33_ASAP7_75t_L      g06332(.A(new_n6505), .B(new_n6507), .C(new_n6508), .Y(new_n6589));
  OAI21xp33_ASAP7_75t_L     g06333(.A1(new_n6589), .A2(new_n6511), .B(new_n6509), .Y(new_n6590));
  NAND2xp33_ASAP7_75t_L     g06334(.A(\b[31] ), .B(new_n1080), .Y(new_n6591));
  NAND3xp33_ASAP7_75t_L     g06335(.A(new_n3210), .B(new_n1073), .C(new_n3213), .Y(new_n6592));
  AOI22xp33_ASAP7_75t_L     g06336(.A1(new_n1076), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1253), .Y(new_n6593));
  AND4x1_ASAP7_75t_L        g06337(.A(new_n6593), .B(new_n6592), .C(new_n6591), .D(\a[17] ), .Y(new_n6594));
  AOI31xp33_ASAP7_75t_L     g06338(.A1(new_n6592), .A2(new_n6591), .A3(new_n6593), .B(\a[17] ), .Y(new_n6595));
  NOR2xp33_ASAP7_75t_L      g06339(.A(new_n6595), .B(new_n6594), .Y(new_n6596));
  NOR2xp33_ASAP7_75t_L      g06340(.A(new_n6490), .B(new_n6491), .Y(new_n6597));
  MAJIxp5_ASAP7_75t_L       g06341(.A(new_n6506), .B(new_n6489), .C(new_n6597), .Y(new_n6598));
  AOI22xp33_ASAP7_75t_L     g06342(.A1(new_n1360), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1581), .Y(new_n6599));
  OAI221xp5_ASAP7_75t_L     g06343(.A1(new_n1373), .A2(new_n2666), .B1(new_n1359), .B2(new_n2695), .C(new_n6599), .Y(new_n6600));
  XNOR2x2_ASAP7_75t_L       g06344(.A(\a[20] ), .B(new_n6600), .Y(new_n6601));
  NOR2xp33_ASAP7_75t_L      g06345(.A(new_n6473), .B(new_n6468), .Y(new_n6602));
  MAJIxp5_ASAP7_75t_L       g06346(.A(new_n6482), .B(new_n6476), .C(new_n6602), .Y(new_n6603));
  AOI22xp33_ASAP7_75t_L     g06347(.A1(new_n1704), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1837), .Y(new_n6604));
  OAI221xp5_ASAP7_75t_L     g06348(.A1(new_n1699), .A2(new_n2067), .B1(new_n1827), .B2(new_n2355), .C(new_n6604), .Y(new_n6605));
  XNOR2x2_ASAP7_75t_L       g06349(.A(\a[23] ), .B(new_n6605), .Y(new_n6606));
  INVx1_ASAP7_75t_L         g06350(.A(new_n6606), .Y(new_n6607));
  NOR3xp33_ASAP7_75t_L      g06351(.A(new_n6462), .B(new_n6463), .C(new_n6460), .Y(new_n6608));
  A2O1A1O1Ixp25_ASAP7_75t_L g06352(.A1(new_n6216), .A2(new_n6214), .B(new_n6467), .C(new_n6466), .D(new_n6608), .Y(new_n6609));
  NAND2xp33_ASAP7_75t_L     g06353(.A(new_n6446), .B(new_n6442), .Y(new_n6610));
  MAJIxp5_ASAP7_75t_L       g06354(.A(new_n6452), .B(new_n6449), .C(new_n6610), .Y(new_n6611));
  O2A1O1Ixp33_ASAP7_75t_L   g06355(.A1(new_n6184), .A2(new_n6185), .B(new_n6194), .C(new_n6439), .Y(new_n6612));
  XOR2x2_ASAP7_75t_L        g06356(.A(new_n6434), .B(new_n6423), .Y(new_n6613));
  NAND2xp33_ASAP7_75t_L     g06357(.A(new_n6436), .B(new_n6613), .Y(new_n6614));
  A2O1A1Ixp33_ASAP7_75t_L   g06358(.A1(new_n6437), .A2(new_n6432), .B(new_n6612), .C(new_n6614), .Y(new_n6615));
  AOI22xp33_ASAP7_75t_L     g06359(.A1(new_n3029), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n3258), .Y(new_n6616));
  OAI221xp5_ASAP7_75t_L     g06360(.A1(new_n3024), .A2(new_n1030), .B1(new_n3256), .B2(new_n1209), .C(new_n6616), .Y(new_n6617));
  XNOR2x2_ASAP7_75t_L       g06361(.A(\a[32] ), .B(new_n6617), .Y(new_n6618));
  NOR3xp33_ASAP7_75t_L      g06362(.A(new_n6398), .B(new_n6397), .C(new_n6395), .Y(new_n6619));
  INVx1_ASAP7_75t_L         g06363(.A(new_n6619), .Y(new_n6620));
  A2O1A1Ixp33_ASAP7_75t_L   g06364(.A1(new_n6400), .A2(new_n6396), .B(new_n6406), .C(new_n6620), .Y(new_n6621));
  AOI22xp33_ASAP7_75t_L     g06365(.A1(new_n4920), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n5167), .Y(new_n6622));
  OAI221xp5_ASAP7_75t_L     g06366(.A1(new_n5154), .A2(new_n420), .B1(new_n5158), .B2(new_n494), .C(new_n6622), .Y(new_n6623));
  NOR2xp33_ASAP7_75t_L      g06367(.A(new_n4915), .B(new_n6623), .Y(new_n6624));
  AND2x2_ASAP7_75t_L        g06368(.A(new_n4915), .B(new_n6623), .Y(new_n6625));
  NAND2xp33_ASAP7_75t_L     g06369(.A(new_n6132), .B(new_n6133), .Y(new_n6626));
  A2O1A1O1Ixp25_ASAP7_75t_L g06370(.A1(new_n6130), .A2(new_n6626), .B(new_n6361), .C(new_n6384), .D(new_n6391), .Y(new_n6627));
  NAND2xp33_ASAP7_75t_L     g06371(.A(\b[4] ), .B(new_n5628), .Y(new_n6628));
  NOR3xp33_ASAP7_75t_L      g06372(.A(new_n357), .B(new_n358), .C(new_n5892), .Y(new_n6629));
  OAI22xp33_ASAP7_75t_L     g06373(.A1(new_n5895), .A2(new_n298), .B1(new_n354), .B2(new_n5894), .Y(new_n6630));
  NOR2xp33_ASAP7_75t_L      g06374(.A(new_n6630), .B(new_n6629), .Y(new_n6631));
  NAND3xp33_ASAP7_75t_L     g06375(.A(new_n6631), .B(new_n6628), .C(\a[44] ), .Y(new_n6632));
  INVx1_ASAP7_75t_L         g06376(.A(new_n6628), .Y(new_n6633));
  OAI31xp33_ASAP7_75t_L     g06377(.A1(new_n6629), .A2(new_n6633), .A3(new_n6630), .B(new_n5619), .Y(new_n6634));
  AND3x1_ASAP7_75t_L        g06378(.A(new_n6374), .B(new_n6377), .C(new_n6381), .Y(new_n6635));
  NAND2xp33_ASAP7_75t_L     g06379(.A(new_n6375), .B(new_n6378), .Y(new_n6636));
  NAND2xp33_ASAP7_75t_L     g06380(.A(\b[2] ), .B(new_n6376), .Y(new_n6637));
  NAND3xp33_ASAP7_75t_L     g06381(.A(new_n6119), .B(new_n6375), .C(new_n6379), .Y(new_n6638));
  OAI221xp5_ASAP7_75t_L     g06382(.A1(new_n258), .A2(new_n6638), .B1(new_n280), .B2(new_n6636), .C(new_n6637), .Y(new_n6639));
  AOI21xp33_ASAP7_75t_L     g06383(.A1(new_n6380), .A2(\b[1] ), .B(new_n6639), .Y(new_n6640));
  A2O1A1Ixp33_ASAP7_75t_L   g06384(.A1(new_n6121), .A2(new_n6635), .B(new_n6371), .C(new_n6640), .Y(new_n6641));
  O2A1O1Ixp33_ASAP7_75t_L   g06385(.A1(new_n258), .A2(new_n6119), .B(new_n6635), .C(new_n6371), .Y(new_n6642));
  A2O1A1Ixp33_ASAP7_75t_L   g06386(.A1(\b[1] ), .A2(new_n6380), .B(new_n6639), .C(new_n6642), .Y(new_n6643));
  NAND4xp25_ASAP7_75t_L     g06387(.A(new_n6643), .B(new_n6632), .C(new_n6634), .D(new_n6641), .Y(new_n6644));
  NAND2xp33_ASAP7_75t_L     g06388(.A(new_n6634), .B(new_n6632), .Y(new_n6645));
  INVx1_ASAP7_75t_L         g06389(.A(new_n6380), .Y(new_n6646));
  NOR2xp33_ASAP7_75t_L      g06390(.A(new_n280), .B(new_n6636), .Y(new_n6647));
  AND3x1_ASAP7_75t_L        g06391(.A(new_n6119), .B(new_n6379), .C(new_n6375), .Y(new_n6648));
  AOI221xp5_ASAP7_75t_L     g06392(.A1(new_n6376), .A2(\b[2] ), .B1(new_n6648), .B2(\b[0] ), .C(new_n6647), .Y(new_n6649));
  OAI21xp33_ASAP7_75t_L     g06393(.A1(new_n261), .A2(new_n6646), .B(new_n6649), .Y(new_n6650));
  O2A1O1Ixp33_ASAP7_75t_L   g06394(.A1(new_n6120), .A2(new_n6382), .B(\a[47] ), .C(new_n6650), .Y(new_n6651));
  A2O1A1Ixp33_ASAP7_75t_L   g06395(.A1(\b[0] ), .A2(new_n6378), .B(new_n6382), .C(\a[47] ), .Y(new_n6652));
  O2A1O1Ixp33_ASAP7_75t_L   g06396(.A1(new_n6646), .A2(new_n261), .B(new_n6649), .C(new_n6652), .Y(new_n6653));
  OAI21xp33_ASAP7_75t_L     g06397(.A1(new_n6651), .A2(new_n6653), .B(new_n6645), .Y(new_n6654));
  AOI21xp33_ASAP7_75t_L     g06398(.A1(new_n6654), .A2(new_n6644), .B(new_n6627), .Y(new_n6655));
  NAND3xp33_ASAP7_75t_L     g06399(.A(new_n6115), .B(new_n5897), .C(new_n6120), .Y(new_n6656));
  A2O1A1Ixp33_ASAP7_75t_L   g06400(.A1(new_n6131), .A2(new_n6656), .B(new_n6390), .C(new_n6387), .Y(new_n6657));
  NAND2xp33_ASAP7_75t_L     g06401(.A(new_n6644), .B(new_n6654), .Y(new_n6658));
  NOR2xp33_ASAP7_75t_L      g06402(.A(new_n6657), .B(new_n6658), .Y(new_n6659));
  OAI22xp33_ASAP7_75t_L     g06403(.A1(new_n6659), .A2(new_n6655), .B1(new_n6625), .B2(new_n6624), .Y(new_n6660));
  XNOR2x2_ASAP7_75t_L       g06404(.A(\a[41] ), .B(new_n6623), .Y(new_n6661));
  A2O1A1Ixp33_ASAP7_75t_L   g06405(.A1(new_n6133), .A2(new_n6132), .B(new_n6134), .C(new_n6656), .Y(new_n6662));
  A2O1A1Ixp33_ASAP7_75t_L   g06406(.A1(new_n6384), .A2(new_n6662), .B(new_n6391), .C(new_n6658), .Y(new_n6663));
  NAND3xp33_ASAP7_75t_L     g06407(.A(new_n6627), .B(new_n6644), .C(new_n6654), .Y(new_n6664));
  NAND3xp33_ASAP7_75t_L     g06408(.A(new_n6663), .B(new_n6664), .C(new_n6661), .Y(new_n6665));
  AND2x2_ASAP7_75t_L        g06409(.A(new_n6665), .B(new_n6660), .Y(new_n6666));
  NAND2xp33_ASAP7_75t_L     g06410(.A(new_n6621), .B(new_n6666), .Y(new_n6667));
  O2A1O1Ixp33_ASAP7_75t_L   g06411(.A1(new_n6402), .A2(new_n6164), .B(new_n6401), .C(new_n6619), .Y(new_n6668));
  NAND2xp33_ASAP7_75t_L     g06412(.A(new_n6665), .B(new_n6660), .Y(new_n6669));
  NAND2xp33_ASAP7_75t_L     g06413(.A(new_n6669), .B(new_n6668), .Y(new_n6670));
  AOI22xp33_ASAP7_75t_L     g06414(.A1(new_n4283), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n4512), .Y(new_n6671));
  OAI221xp5_ASAP7_75t_L     g06415(.A1(new_n4277), .A2(new_n617), .B1(new_n4499), .B2(new_n685), .C(new_n6671), .Y(new_n6672));
  XNOR2x2_ASAP7_75t_L       g06416(.A(\a[38] ), .B(new_n6672), .Y(new_n6673));
  NAND3xp33_ASAP7_75t_L     g06417(.A(new_n6667), .B(new_n6670), .C(new_n6673), .Y(new_n6674));
  A2O1A1O1Ixp25_ASAP7_75t_L g06418(.A1(new_n6400), .A2(new_n6396), .B(new_n6406), .C(new_n6620), .D(new_n6669), .Y(new_n6675));
  NOR2xp33_ASAP7_75t_L      g06419(.A(new_n6621), .B(new_n6666), .Y(new_n6676));
  INVx1_ASAP7_75t_L         g06420(.A(new_n6673), .Y(new_n6677));
  OAI21xp33_ASAP7_75t_L     g06421(.A1(new_n6675), .A2(new_n6676), .B(new_n6677), .Y(new_n6678));
  NAND2xp33_ASAP7_75t_L     g06422(.A(new_n6415), .B(new_n6417), .Y(new_n6679));
  NAND4xp25_ASAP7_75t_L     g06423(.A(new_n6679), .B(new_n6678), .C(new_n6674), .D(new_n6411), .Y(new_n6680));
  NOR3xp33_ASAP7_75t_L      g06424(.A(new_n6677), .B(new_n6676), .C(new_n6675), .Y(new_n6681));
  AOI21xp33_ASAP7_75t_L     g06425(.A1(new_n6667), .A2(new_n6670), .B(new_n6673), .Y(new_n6682));
  AOI211xp5_ASAP7_75t_L     g06426(.A1(new_n6360), .A2(new_n6166), .B(new_n6419), .C(new_n6165), .Y(new_n6683));
  OAI22xp33_ASAP7_75t_L     g06427(.A1(new_n6683), .A2(new_n6418), .B1(new_n6681), .B2(new_n6682), .Y(new_n6684));
  AOI22xp33_ASAP7_75t_L     g06428(.A1(new_n3633), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n3858), .Y(new_n6685));
  OAI221xp5_ASAP7_75t_L     g06429(.A1(new_n3853), .A2(new_n784), .B1(new_n3856), .B2(new_n875), .C(new_n6685), .Y(new_n6686));
  XNOR2x2_ASAP7_75t_L       g06430(.A(\a[35] ), .B(new_n6686), .Y(new_n6687));
  NAND3xp33_ASAP7_75t_L     g06431(.A(new_n6684), .B(new_n6680), .C(new_n6687), .Y(new_n6688));
  AND4x1_ASAP7_75t_L        g06432(.A(new_n6679), .B(new_n6678), .C(new_n6674), .D(new_n6411), .Y(new_n6689));
  AOI22xp33_ASAP7_75t_L     g06433(.A1(new_n6678), .A2(new_n6674), .B1(new_n6411), .B2(new_n6679), .Y(new_n6690));
  INVx1_ASAP7_75t_L         g06434(.A(new_n6687), .Y(new_n6691));
  OAI21xp33_ASAP7_75t_L     g06435(.A1(new_n6690), .A2(new_n6689), .B(new_n6691), .Y(new_n6692));
  NAND2xp33_ASAP7_75t_L     g06436(.A(new_n6692), .B(new_n6688), .Y(new_n6693));
  A2O1A1Ixp33_ASAP7_75t_L   g06437(.A1(new_n6423), .A2(new_n6434), .B(new_n6422), .C(new_n6693), .Y(new_n6694));
  A2O1A1O1Ixp25_ASAP7_75t_L g06438(.A1(new_n6108), .A2(new_n6354), .B(new_n6356), .C(new_n6425), .D(new_n6422), .Y(new_n6695));
  NAND3xp33_ASAP7_75t_L     g06439(.A(new_n6695), .B(new_n6688), .C(new_n6692), .Y(new_n6696));
  AOI21xp33_ASAP7_75t_L     g06440(.A1(new_n6694), .A2(new_n6696), .B(new_n6618), .Y(new_n6697));
  AND3x1_ASAP7_75t_L        g06441(.A(new_n6694), .B(new_n6696), .C(new_n6618), .Y(new_n6698));
  NOR2xp33_ASAP7_75t_L      g06442(.A(new_n6697), .B(new_n6698), .Y(new_n6699));
  NAND2xp33_ASAP7_75t_L     g06443(.A(new_n6615), .B(new_n6699), .Y(new_n6700));
  MAJIxp5_ASAP7_75t_L       g06444(.A(new_n6445), .B(new_n6436), .C(new_n6613), .Y(new_n6701));
  OAI21xp33_ASAP7_75t_L     g06445(.A1(new_n6697), .A2(new_n6698), .B(new_n6701), .Y(new_n6702));
  AOI22xp33_ASAP7_75t_L     g06446(.A1(new_n2552), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n2736), .Y(new_n6703));
  OAI221xp5_ASAP7_75t_L     g06447(.A1(new_n2547), .A2(new_n1432), .B1(new_n2734), .B2(new_n1547), .C(new_n6703), .Y(new_n6704));
  NOR2xp33_ASAP7_75t_L      g06448(.A(new_n2538), .B(new_n6704), .Y(new_n6705));
  AND2x2_ASAP7_75t_L        g06449(.A(new_n2538), .B(new_n6704), .Y(new_n6706));
  NOR2xp33_ASAP7_75t_L      g06450(.A(new_n6705), .B(new_n6706), .Y(new_n6707));
  AO21x2_ASAP7_75t_L        g06451(.A1(new_n6702), .A2(new_n6700), .B(new_n6707), .Y(new_n6708));
  NAND3xp33_ASAP7_75t_L     g06452(.A(new_n6700), .B(new_n6702), .C(new_n6707), .Y(new_n6709));
  AO21x2_ASAP7_75t_L        g06453(.A1(new_n6709), .A2(new_n6708), .B(new_n6611), .Y(new_n6710));
  NAND3xp33_ASAP7_75t_L     g06454(.A(new_n6708), .B(new_n6611), .C(new_n6709), .Y(new_n6711));
  AOI22xp33_ASAP7_75t_L     g06455(.A1(new_n2114), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n2259), .Y(new_n6712));
  OAI221xp5_ASAP7_75t_L     g06456(.A1(new_n2109), .A2(new_n1774), .B1(new_n2257), .B2(new_n1915), .C(new_n6712), .Y(new_n6713));
  XNOR2x2_ASAP7_75t_L       g06457(.A(new_n2100), .B(new_n6713), .Y(new_n6714));
  AO21x2_ASAP7_75t_L        g06458(.A1(new_n6711), .A2(new_n6710), .B(new_n6714), .Y(new_n6715));
  NAND3xp33_ASAP7_75t_L     g06459(.A(new_n6710), .B(new_n6714), .C(new_n6711), .Y(new_n6716));
  NAND2xp33_ASAP7_75t_L     g06460(.A(new_n6716), .B(new_n6715), .Y(new_n6717));
  NAND2xp33_ASAP7_75t_L     g06461(.A(new_n6609), .B(new_n6717), .Y(new_n6718));
  INVx1_ASAP7_75t_L         g06462(.A(new_n6467), .Y(new_n6719));
  INVx1_ASAP7_75t_L         g06463(.A(new_n6608), .Y(new_n6720));
  A2O1A1Ixp33_ASAP7_75t_L   g06464(.A1(new_n6227), .A2(new_n6719), .B(new_n6471), .C(new_n6720), .Y(new_n6721));
  NAND3xp33_ASAP7_75t_L     g06465(.A(new_n6721), .B(new_n6715), .C(new_n6716), .Y(new_n6722));
  AOI21xp33_ASAP7_75t_L     g06466(.A1(new_n6718), .A2(new_n6722), .B(new_n6607), .Y(new_n6723));
  AOI21xp33_ASAP7_75t_L     g06467(.A1(new_n6716), .A2(new_n6715), .B(new_n6721), .Y(new_n6724));
  NOR2xp33_ASAP7_75t_L      g06468(.A(new_n6609), .B(new_n6717), .Y(new_n6725));
  NOR3xp33_ASAP7_75t_L      g06469(.A(new_n6725), .B(new_n6724), .C(new_n6606), .Y(new_n6726));
  NOR3xp33_ASAP7_75t_L      g06470(.A(new_n6603), .B(new_n6723), .C(new_n6726), .Y(new_n6727));
  NAND2xp33_ASAP7_75t_L     g06471(.A(new_n6479), .B(new_n6478), .Y(new_n6728));
  MAJIxp5_ASAP7_75t_L       g06472(.A(new_n6486), .B(new_n6480), .C(new_n6728), .Y(new_n6729));
  OAI21xp33_ASAP7_75t_L     g06473(.A1(new_n6724), .A2(new_n6725), .B(new_n6606), .Y(new_n6730));
  NAND3xp33_ASAP7_75t_L     g06474(.A(new_n6718), .B(new_n6722), .C(new_n6607), .Y(new_n6731));
  AOI21xp33_ASAP7_75t_L     g06475(.A1(new_n6731), .A2(new_n6730), .B(new_n6729), .Y(new_n6732));
  OAI21xp33_ASAP7_75t_L     g06476(.A1(new_n6732), .A2(new_n6727), .B(new_n6601), .Y(new_n6733));
  INVx1_ASAP7_75t_L         g06477(.A(new_n6601), .Y(new_n6734));
  NAND3xp33_ASAP7_75t_L     g06478(.A(new_n6729), .B(new_n6730), .C(new_n6731), .Y(new_n6735));
  OAI21xp33_ASAP7_75t_L     g06479(.A1(new_n6723), .A2(new_n6726), .B(new_n6603), .Y(new_n6736));
  NAND3xp33_ASAP7_75t_L     g06480(.A(new_n6735), .B(new_n6736), .C(new_n6734), .Y(new_n6737));
  NAND2xp33_ASAP7_75t_L     g06481(.A(new_n6737), .B(new_n6733), .Y(new_n6738));
  NOR2xp33_ASAP7_75t_L      g06482(.A(new_n6598), .B(new_n6738), .Y(new_n6739));
  NOR3xp33_ASAP7_75t_L      g06483(.A(new_n6491), .B(new_n6490), .C(new_n6353), .Y(new_n6740));
  AOI221xp5_ASAP7_75t_L     g06484(.A1(new_n6506), .A2(new_n6498), .B1(new_n6737), .B2(new_n6733), .C(new_n6740), .Y(new_n6741));
  OAI21xp33_ASAP7_75t_L     g06485(.A1(new_n6741), .A2(new_n6739), .B(new_n6596), .Y(new_n6742));
  INVx1_ASAP7_75t_L         g06486(.A(new_n6596), .Y(new_n6743));
  AOI21xp33_ASAP7_75t_L     g06487(.A1(new_n6735), .A2(new_n6736), .B(new_n6734), .Y(new_n6744));
  NOR3xp33_ASAP7_75t_L      g06488(.A(new_n6727), .B(new_n6732), .C(new_n6601), .Y(new_n6745));
  NOR2xp33_ASAP7_75t_L      g06489(.A(new_n6744), .B(new_n6745), .Y(new_n6746));
  A2O1A1Ixp33_ASAP7_75t_L   g06490(.A1(new_n6498), .A2(new_n6506), .B(new_n6740), .C(new_n6746), .Y(new_n6747));
  NAND2xp33_ASAP7_75t_L     g06491(.A(new_n6598), .B(new_n6738), .Y(new_n6748));
  NAND3xp33_ASAP7_75t_L     g06492(.A(new_n6747), .B(new_n6743), .C(new_n6748), .Y(new_n6749));
  NAND3xp33_ASAP7_75t_L     g06493(.A(new_n6590), .B(new_n6742), .C(new_n6749), .Y(new_n6750));
  AOI21xp33_ASAP7_75t_L     g06494(.A1(new_n6499), .A2(new_n6494), .B(new_n6502), .Y(new_n6751));
  A2O1A1O1Ixp25_ASAP7_75t_L g06495(.A1(new_n6258), .A2(new_n6255), .B(new_n6256), .C(new_n6503), .D(new_n6751), .Y(new_n6752));
  AOI21xp33_ASAP7_75t_L     g06496(.A1(new_n6747), .A2(new_n6748), .B(new_n6743), .Y(new_n6753));
  NOR3xp33_ASAP7_75t_L      g06497(.A(new_n6739), .B(new_n6596), .C(new_n6741), .Y(new_n6754));
  OAI21xp33_ASAP7_75t_L     g06498(.A1(new_n6753), .A2(new_n6754), .B(new_n6752), .Y(new_n6755));
  NAND2xp33_ASAP7_75t_L     g06499(.A(\b[34] ), .B(new_n815), .Y(new_n6756));
  NAND2xp33_ASAP7_75t_L     g06500(.A(new_n808), .B(new_n3811), .Y(new_n6757));
  AOI22xp33_ASAP7_75t_L     g06501(.A1(new_n811), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n900), .Y(new_n6758));
  AND4x1_ASAP7_75t_L        g06502(.A(new_n6758), .B(new_n6757), .C(new_n6756), .D(\a[14] ), .Y(new_n6759));
  AOI31xp33_ASAP7_75t_L     g06503(.A1(new_n6757), .A2(new_n6756), .A3(new_n6758), .B(\a[14] ), .Y(new_n6760));
  NOR2xp33_ASAP7_75t_L      g06504(.A(new_n6760), .B(new_n6759), .Y(new_n6761));
  NAND3xp33_ASAP7_75t_L     g06505(.A(new_n6750), .B(new_n6755), .C(new_n6761), .Y(new_n6762));
  NOR3xp33_ASAP7_75t_L      g06506(.A(new_n6752), .B(new_n6753), .C(new_n6754), .Y(new_n6763));
  AOI221xp5_ASAP7_75t_L     g06507(.A1(new_n6347), .A2(new_n6503), .B1(new_n6742), .B2(new_n6749), .C(new_n6751), .Y(new_n6764));
  INVx1_ASAP7_75t_L         g06508(.A(new_n6761), .Y(new_n6765));
  OAI21xp33_ASAP7_75t_L     g06509(.A1(new_n6764), .A2(new_n6763), .B(new_n6765), .Y(new_n6766));
  NAND2xp33_ASAP7_75t_L     g06510(.A(new_n6766), .B(new_n6762), .Y(new_n6767));
  NAND2xp33_ASAP7_75t_L     g06511(.A(new_n6510), .B(new_n6513), .Y(new_n6768));
  MAJIxp5_ASAP7_75t_L       g06512(.A(new_n6091), .B(new_n6263), .C(new_n6522), .Y(new_n6769));
  MAJIxp5_ASAP7_75t_L       g06513(.A(new_n6769), .B(new_n6768), .C(new_n6516), .Y(new_n6770));
  NOR2xp33_ASAP7_75t_L      g06514(.A(new_n6770), .B(new_n6767), .Y(new_n6771));
  NOR2xp33_ASAP7_75t_L      g06515(.A(new_n6519), .B(new_n6518), .Y(new_n6772));
  MAJIxp5_ASAP7_75t_L       g06516(.A(new_n6528), .B(new_n6520), .C(new_n6772), .Y(new_n6773));
  AOI21xp33_ASAP7_75t_L     g06517(.A1(new_n6766), .A2(new_n6762), .B(new_n6773), .Y(new_n6774));
  AOI22xp33_ASAP7_75t_L     g06518(.A1(\b[36] ), .A2(new_n651), .B1(\b[38] ), .B2(new_n581), .Y(new_n6775));
  OAI221xp5_ASAP7_75t_L     g06519(.A1(new_n821), .A2(new_n4424), .B1(new_n577), .B2(new_n4641), .C(new_n6775), .Y(new_n6776));
  XNOR2x2_ASAP7_75t_L       g06520(.A(new_n574), .B(new_n6776), .Y(new_n6777));
  NOR3xp33_ASAP7_75t_L      g06521(.A(new_n6771), .B(new_n6774), .C(new_n6777), .Y(new_n6778));
  OA21x2_ASAP7_75t_L        g06522(.A1(new_n6774), .A2(new_n6771), .B(new_n6777), .Y(new_n6779));
  INVx1_ASAP7_75t_L         g06523(.A(new_n6532), .Y(new_n6780));
  NAND3xp33_ASAP7_75t_L     g06524(.A(new_n6524), .B(new_n6529), .C(new_n6780), .Y(new_n6781));
  A2O1A1Ixp33_ASAP7_75t_L   g06525(.A1(new_n6534), .A2(new_n6533), .B(new_n6535), .C(new_n6781), .Y(new_n6782));
  NOR3xp33_ASAP7_75t_L      g06526(.A(new_n6782), .B(new_n6779), .C(new_n6778), .Y(new_n6783));
  OA21x2_ASAP7_75t_L        g06527(.A1(new_n6778), .A2(new_n6779), .B(new_n6782), .Y(new_n6784));
  NOR2xp33_ASAP7_75t_L      g06528(.A(new_n4869), .B(new_n468), .Y(new_n6785));
  INVx1_ASAP7_75t_L         g06529(.A(new_n6785), .Y(new_n6786));
  NAND3xp33_ASAP7_75t_L     g06530(.A(new_n5326), .B(new_n5324), .C(new_n441), .Y(new_n6787));
  AOI22xp33_ASAP7_75t_L     g06531(.A1(new_n444), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n471), .Y(new_n6788));
  AND4x1_ASAP7_75t_L        g06532(.A(new_n6788), .B(new_n6787), .C(new_n6786), .D(\a[8] ), .Y(new_n6789));
  AOI31xp33_ASAP7_75t_L     g06533(.A1(new_n6787), .A2(new_n6786), .A3(new_n6788), .B(\a[8] ), .Y(new_n6790));
  NOR2xp33_ASAP7_75t_L      g06534(.A(new_n6790), .B(new_n6789), .Y(new_n6791));
  NOR3xp33_ASAP7_75t_L      g06535(.A(new_n6784), .B(new_n6791), .C(new_n6783), .Y(new_n6792));
  OR3x1_ASAP7_75t_L         g06536(.A(new_n6782), .B(new_n6778), .C(new_n6779), .Y(new_n6793));
  OAI21xp33_ASAP7_75t_L     g06537(.A1(new_n6778), .A2(new_n6779), .B(new_n6782), .Y(new_n6794));
  INVx1_ASAP7_75t_L         g06538(.A(new_n6791), .Y(new_n6795));
  AOI21xp33_ASAP7_75t_L     g06539(.A1(new_n6793), .A2(new_n6794), .B(new_n6795), .Y(new_n6796));
  NOR2xp33_ASAP7_75t_L      g06540(.A(new_n6792), .B(new_n6796), .Y(new_n6797));
  A2O1A1Ixp33_ASAP7_75t_L   g06541(.A1(new_n6546), .A2(new_n6559), .B(new_n6552), .C(new_n6797), .Y(new_n6798));
  NAND3xp33_ASAP7_75t_L     g06542(.A(new_n6793), .B(new_n6794), .C(new_n6795), .Y(new_n6799));
  OAI21xp33_ASAP7_75t_L     g06543(.A1(new_n6783), .A2(new_n6784), .B(new_n6791), .Y(new_n6800));
  NAND2xp33_ASAP7_75t_L     g06544(.A(new_n6800), .B(new_n6799), .Y(new_n6801));
  A2O1A1O1Ixp25_ASAP7_75t_L g06545(.A1(new_n6301), .A2(new_n6551), .B(new_n6345), .C(new_n6546), .D(new_n6552), .Y(new_n6802));
  NAND2xp33_ASAP7_75t_L     g06546(.A(new_n6802), .B(new_n6801), .Y(new_n6803));
  AOI21xp33_ASAP7_75t_L     g06547(.A1(new_n6798), .A2(new_n6803), .B(new_n6588), .Y(new_n6804));
  O2A1O1Ixp33_ASAP7_75t_L   g06548(.A1(new_n6346), .A2(new_n6553), .B(new_n6545), .C(new_n6801), .Y(new_n6805));
  A2O1A1Ixp33_ASAP7_75t_L   g06549(.A1(new_n6302), .A2(new_n6558), .B(new_n6547), .C(new_n6545), .Y(new_n6806));
  NOR2xp33_ASAP7_75t_L      g06550(.A(new_n6806), .B(new_n6797), .Y(new_n6807));
  NOR3xp33_ASAP7_75t_L      g06551(.A(new_n6805), .B(new_n6807), .C(new_n6587), .Y(new_n6808));
  NOR2xp33_ASAP7_75t_L      g06552(.A(new_n6804), .B(new_n6808), .Y(new_n6809));
  XNOR2x2_ASAP7_75t_L       g06553(.A(new_n6584), .B(new_n6809), .Y(new_n6810));
  NOR2xp33_ASAP7_75t_L      g06554(.A(\b[46] ), .B(\b[47] ), .Y(new_n6811));
  INVx1_ASAP7_75t_L         g06555(.A(\b[47] ), .Y(new_n6812));
  NOR2xp33_ASAP7_75t_L      g06556(.A(new_n6568), .B(new_n6812), .Y(new_n6813));
  NOR2xp33_ASAP7_75t_L      g06557(.A(new_n6811), .B(new_n6813), .Y(new_n6814));
  INVx1_ASAP7_75t_L         g06558(.A(new_n6814), .Y(new_n6815));
  O2A1O1Ixp33_ASAP7_75t_L   g06559(.A1(new_n6321), .A2(new_n6568), .B(new_n6571), .C(new_n6815), .Y(new_n6816));
  INVx1_ASAP7_75t_L         g06560(.A(new_n6816), .Y(new_n6817));
  O2A1O1Ixp33_ASAP7_75t_L   g06561(.A1(new_n6322), .A2(new_n6325), .B(new_n6570), .C(new_n6569), .Y(new_n6818));
  NAND2xp33_ASAP7_75t_L     g06562(.A(new_n6815), .B(new_n6818), .Y(new_n6819));
  NAND2xp33_ASAP7_75t_L     g06563(.A(new_n6819), .B(new_n6817), .Y(new_n6820));
  AOI22xp33_ASAP7_75t_L     g06564(.A1(\b[45] ), .A2(new_n282), .B1(\b[47] ), .B2(new_n303), .Y(new_n6821));
  OAI221xp5_ASAP7_75t_L     g06565(.A1(new_n291), .A2(new_n6568), .B1(new_n268), .B2(new_n6820), .C(new_n6821), .Y(new_n6822));
  XNOR2x2_ASAP7_75t_L       g06566(.A(\a[2] ), .B(new_n6822), .Y(new_n6823));
  XOR2x2_ASAP7_75t_L        g06567(.A(new_n6823), .B(new_n6810), .Y(new_n6824));
  MAJIxp5_ASAP7_75t_L       g06568(.A(new_n6580), .B(new_n6566), .C(new_n6576), .Y(new_n6825));
  XNOR2x2_ASAP7_75t_L       g06569(.A(new_n6825), .B(new_n6824), .Y(\f[47] ));
  A2O1A1Ixp33_ASAP7_75t_L   g06570(.A1(new_n6576), .A2(new_n6566), .B(new_n6578), .C(new_n6824), .Y(new_n6827));
  INVx1_ASAP7_75t_L         g06571(.A(new_n6813), .Y(new_n6828));
  NOR2xp33_ASAP7_75t_L      g06572(.A(\b[47] ), .B(\b[48] ), .Y(new_n6829));
  INVx1_ASAP7_75t_L         g06573(.A(\b[48] ), .Y(new_n6830));
  NOR2xp33_ASAP7_75t_L      g06574(.A(new_n6812), .B(new_n6830), .Y(new_n6831));
  NOR2xp33_ASAP7_75t_L      g06575(.A(new_n6829), .B(new_n6831), .Y(new_n6832));
  INVx1_ASAP7_75t_L         g06576(.A(new_n6832), .Y(new_n6833));
  O2A1O1Ixp33_ASAP7_75t_L   g06577(.A1(new_n6815), .A2(new_n6818), .B(new_n6828), .C(new_n6833), .Y(new_n6834));
  INVx1_ASAP7_75t_L         g06578(.A(new_n6834), .Y(new_n6835));
  NAND3xp33_ASAP7_75t_L     g06579(.A(new_n6817), .B(new_n6828), .C(new_n6833), .Y(new_n6836));
  NAND2xp33_ASAP7_75t_L     g06580(.A(new_n6835), .B(new_n6836), .Y(new_n6837));
  AOI22xp33_ASAP7_75t_L     g06581(.A1(\b[46] ), .A2(new_n282), .B1(\b[48] ), .B2(new_n303), .Y(new_n6838));
  OAI221xp5_ASAP7_75t_L     g06582(.A1(new_n291), .A2(new_n6812), .B1(new_n268), .B2(new_n6837), .C(new_n6838), .Y(new_n6839));
  XNOR2x2_ASAP7_75t_L       g06583(.A(\a[2] ), .B(new_n6839), .Y(new_n6840));
  AO21x2_ASAP7_75t_L        g06584(.A1(new_n6318), .A2(new_n6317), .B(new_n6564), .Y(new_n6841));
  NAND2xp33_ASAP7_75t_L     g06585(.A(new_n6548), .B(new_n6555), .Y(new_n6842));
  NOR2xp33_ASAP7_75t_L      g06586(.A(new_n6344), .B(new_n6842), .Y(new_n6843));
  OAI21xp33_ASAP7_75t_L     g06587(.A1(new_n6807), .A2(new_n6805), .B(new_n6587), .Y(new_n6844));
  A2O1A1O1Ixp25_ASAP7_75t_L g06588(.A1(new_n6563), .A2(new_n6841), .B(new_n6843), .C(new_n6844), .D(new_n6808), .Y(new_n6845));
  NAND2xp33_ASAP7_75t_L     g06589(.A(new_n6770), .B(new_n6767), .Y(new_n6846));
  NAND3xp33_ASAP7_75t_L     g06590(.A(new_n6750), .B(new_n6755), .C(new_n6765), .Y(new_n6847));
  INVx1_ASAP7_75t_L         g06591(.A(new_n4223), .Y(new_n6848));
  OAI22xp33_ASAP7_75t_L     g06592(.A1(new_n978), .A2(new_n3584), .B1(new_n4216), .B2(new_n977), .Y(new_n6849));
  AOI221xp5_ASAP7_75t_L     g06593(.A1(\b[35] ), .A2(new_n815), .B1(new_n808), .B2(new_n6848), .C(new_n6849), .Y(new_n6850));
  XNOR2x2_ASAP7_75t_L       g06594(.A(\a[14] ), .B(new_n6850), .Y(new_n6851));
  A2O1A1O1Ixp25_ASAP7_75t_L g06595(.A1(new_n6503), .A2(new_n6347), .B(new_n6751), .C(new_n6742), .D(new_n6754), .Y(new_n6852));
  OAI21xp33_ASAP7_75t_L     g06596(.A1(new_n6744), .A2(new_n6598), .B(new_n6737), .Y(new_n6853));
  AOI22xp33_ASAP7_75t_L     g06597(.A1(new_n1360), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1581), .Y(new_n6854));
  OAI221xp5_ASAP7_75t_L     g06598(.A1(new_n1373), .A2(new_n2688), .B1(new_n1359), .B2(new_n2990), .C(new_n6854), .Y(new_n6855));
  XNOR2x2_ASAP7_75t_L       g06599(.A(\a[20] ), .B(new_n6855), .Y(new_n6856));
  INVx1_ASAP7_75t_L         g06600(.A(new_n6856), .Y(new_n6857));
  NOR3xp33_ASAP7_75t_L      g06601(.A(new_n6689), .B(new_n6690), .C(new_n6687), .Y(new_n6858));
  INVx1_ASAP7_75t_L         g06602(.A(new_n6858), .Y(new_n6859));
  A2O1A1Ixp33_ASAP7_75t_L   g06603(.A1(new_n6688), .A2(new_n6692), .B(new_n6695), .C(new_n6859), .Y(new_n6860));
  AOI22xp33_ASAP7_75t_L     g06604(.A1(new_n3633), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n3858), .Y(new_n6861));
  OAI221xp5_ASAP7_75t_L     g06605(.A1(new_n3853), .A2(new_n869), .B1(new_n3856), .B2(new_n950), .C(new_n6861), .Y(new_n6862));
  XNOR2x2_ASAP7_75t_L       g06606(.A(\a[35] ), .B(new_n6862), .Y(new_n6863));
  INVx1_ASAP7_75t_L         g06607(.A(new_n6863), .Y(new_n6864));
  OAI31xp33_ASAP7_75t_L     g06608(.A1(new_n6683), .A2(new_n6681), .A3(new_n6418), .B(new_n6678), .Y(new_n6865));
  AOI22xp33_ASAP7_75t_L     g06609(.A1(new_n4283), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n4512), .Y(new_n6866));
  OAI221xp5_ASAP7_75t_L     g06610(.A1(new_n4277), .A2(new_n679), .B1(new_n4499), .B2(new_n768), .C(new_n6866), .Y(new_n6867));
  XNOR2x2_ASAP7_75t_L       g06611(.A(\a[38] ), .B(new_n6867), .Y(new_n6868));
  NOR3xp33_ASAP7_75t_L      g06612(.A(new_n6659), .B(new_n6655), .C(new_n6661), .Y(new_n6869));
  NAND5xp2_ASAP7_75t_L      g06613(.A(\a[47] ), .B(new_n6374), .C(new_n6377), .D(new_n6381), .E(new_n6121), .Y(new_n6870));
  INVx1_ASAP7_75t_L         g06614(.A(\a[48] ), .Y(new_n6871));
  NAND2xp33_ASAP7_75t_L     g06615(.A(\a[47] ), .B(new_n6871), .Y(new_n6872));
  NAND2xp33_ASAP7_75t_L     g06616(.A(\a[48] ), .B(new_n6371), .Y(new_n6873));
  AND2x2_ASAP7_75t_L        g06617(.A(new_n6872), .B(new_n6873), .Y(new_n6874));
  NOR2xp33_ASAP7_75t_L      g06618(.A(new_n258), .B(new_n6874), .Y(new_n6875));
  OAI21xp33_ASAP7_75t_L     g06619(.A1(new_n6870), .A2(new_n6650), .B(new_n6875), .Y(new_n6876));
  INVx1_ASAP7_75t_L         g06620(.A(new_n6870), .Y(new_n6877));
  INVx1_ASAP7_75t_L         g06621(.A(new_n6875), .Y(new_n6878));
  NAND3xp33_ASAP7_75t_L     g06622(.A(new_n6640), .B(new_n6877), .C(new_n6878), .Y(new_n6879));
  NAND3xp33_ASAP7_75t_L     g06623(.A(new_n6378), .B(new_n6370), .C(new_n6372), .Y(new_n6880));
  OAI22xp33_ASAP7_75t_L     g06624(.A1(new_n6638), .A2(new_n261), .B1(new_n298), .B2(new_n6880), .Y(new_n6881));
  AOI221xp5_ASAP7_75t_L     g06625(.A1(\b[2] ), .A2(new_n6380), .B1(new_n406), .B2(new_n6373), .C(new_n6881), .Y(new_n6882));
  NAND2xp33_ASAP7_75t_L     g06626(.A(\a[47] ), .B(new_n6882), .Y(new_n6883));
  NAND2xp33_ASAP7_75t_L     g06627(.A(\b[3] ), .B(new_n6376), .Y(new_n6884));
  OAI221xp5_ASAP7_75t_L     g06628(.A1(new_n6638), .A2(new_n261), .B1(new_n6636), .B2(new_n302), .C(new_n6884), .Y(new_n6885));
  A2O1A1Ixp33_ASAP7_75t_L   g06629(.A1(\b[2] ), .A2(new_n6380), .B(new_n6885), .C(new_n6371), .Y(new_n6886));
  AO22x1_ASAP7_75t_L        g06630(.A1(new_n6886), .A2(new_n6883), .B1(new_n6876), .B2(new_n6879), .Y(new_n6887));
  XNOR2x2_ASAP7_75t_L       g06631(.A(new_n6371), .B(new_n6882), .Y(new_n6888));
  NAND3xp33_ASAP7_75t_L     g06632(.A(new_n6888), .B(new_n6879), .C(new_n6876), .Y(new_n6889));
  NAND2xp33_ASAP7_75t_L     g06633(.A(\b[5] ), .B(new_n5628), .Y(new_n6890));
  NAND2xp33_ASAP7_75t_L     g06634(.A(new_n5621), .B(new_n526), .Y(new_n6891));
  AOI22xp33_ASAP7_75t_L     g06635(.A1(new_n5624), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n5901), .Y(new_n6892));
  NAND4xp25_ASAP7_75t_L     g06636(.A(new_n6891), .B(\a[44] ), .C(new_n6890), .D(new_n6892), .Y(new_n6893));
  AOI31xp33_ASAP7_75t_L     g06637(.A1(new_n6891), .A2(new_n6890), .A3(new_n6892), .B(\a[44] ), .Y(new_n6894));
  INVx1_ASAP7_75t_L         g06638(.A(new_n6894), .Y(new_n6895));
  NAND4xp25_ASAP7_75t_L     g06639(.A(new_n6887), .B(new_n6889), .C(new_n6895), .D(new_n6893), .Y(new_n6896));
  AOI21xp33_ASAP7_75t_L     g06640(.A1(new_n6879), .A2(new_n6876), .B(new_n6888), .Y(new_n6897));
  AND4x1_ASAP7_75t_L        g06641(.A(new_n6879), .B(new_n6876), .C(new_n6886), .D(new_n6883), .Y(new_n6898));
  INVx1_ASAP7_75t_L         g06642(.A(new_n6893), .Y(new_n6899));
  OAI22xp33_ASAP7_75t_L     g06643(.A1(new_n6898), .A2(new_n6897), .B1(new_n6894), .B2(new_n6899), .Y(new_n6900));
  AND2x2_ASAP7_75t_L        g06644(.A(new_n6896), .B(new_n6900), .Y(new_n6901));
  AOI211xp5_ASAP7_75t_L     g06645(.A1(new_n6632), .A2(new_n6634), .B(new_n6651), .C(new_n6653), .Y(new_n6902));
  A2O1A1O1Ixp25_ASAP7_75t_L g06646(.A1(new_n6384), .A2(new_n6662), .B(new_n6391), .C(new_n6658), .D(new_n6902), .Y(new_n6903));
  NAND2xp33_ASAP7_75t_L     g06647(.A(new_n6903), .B(new_n6901), .Y(new_n6904));
  NAND2xp33_ASAP7_75t_L     g06648(.A(new_n6896), .B(new_n6900), .Y(new_n6905));
  A2O1A1Ixp33_ASAP7_75t_L   g06649(.A1(new_n6657), .A2(new_n6658), .B(new_n6902), .C(new_n6905), .Y(new_n6906));
  AOI22xp33_ASAP7_75t_L     g06650(.A1(new_n4920), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n5167), .Y(new_n6907));
  OAI221xp5_ASAP7_75t_L     g06651(.A1(new_n5154), .A2(new_n488), .B1(new_n5158), .B2(new_n548), .C(new_n6907), .Y(new_n6908));
  XNOR2x2_ASAP7_75t_L       g06652(.A(new_n4915), .B(new_n6908), .Y(new_n6909));
  AOI21xp33_ASAP7_75t_L     g06653(.A1(new_n6904), .A2(new_n6906), .B(new_n6909), .Y(new_n6910));
  NOR2xp33_ASAP7_75t_L      g06654(.A(new_n6651), .B(new_n6653), .Y(new_n6911));
  NAND2xp33_ASAP7_75t_L     g06655(.A(new_n6645), .B(new_n6911), .Y(new_n6912));
  A2O1A1Ixp33_ASAP7_75t_L   g06656(.A1(new_n6644), .A2(new_n6654), .B(new_n6627), .C(new_n6912), .Y(new_n6913));
  NOR2xp33_ASAP7_75t_L      g06657(.A(new_n6905), .B(new_n6913), .Y(new_n6914));
  NOR2xp33_ASAP7_75t_L      g06658(.A(new_n6903), .B(new_n6901), .Y(new_n6915));
  XNOR2x2_ASAP7_75t_L       g06659(.A(\a[41] ), .B(new_n6908), .Y(new_n6916));
  NOR3xp33_ASAP7_75t_L      g06660(.A(new_n6915), .B(new_n6916), .C(new_n6914), .Y(new_n6917));
  NOR2xp33_ASAP7_75t_L      g06661(.A(new_n6910), .B(new_n6917), .Y(new_n6918));
  A2O1A1Ixp33_ASAP7_75t_L   g06662(.A1(new_n6669), .A2(new_n6621), .B(new_n6869), .C(new_n6918), .Y(new_n6919));
  A2O1A1O1Ixp25_ASAP7_75t_L g06663(.A1(new_n6404), .A2(new_n6401), .B(new_n6619), .C(new_n6669), .D(new_n6869), .Y(new_n6920));
  OAI21xp33_ASAP7_75t_L     g06664(.A1(new_n6914), .A2(new_n6915), .B(new_n6916), .Y(new_n6921));
  NAND3xp33_ASAP7_75t_L     g06665(.A(new_n6904), .B(new_n6906), .C(new_n6909), .Y(new_n6922));
  NAND2xp33_ASAP7_75t_L     g06666(.A(new_n6922), .B(new_n6921), .Y(new_n6923));
  NAND2xp33_ASAP7_75t_L     g06667(.A(new_n6923), .B(new_n6920), .Y(new_n6924));
  AOI21xp33_ASAP7_75t_L     g06668(.A1(new_n6919), .A2(new_n6924), .B(new_n6868), .Y(new_n6925));
  INVx1_ASAP7_75t_L         g06669(.A(new_n6868), .Y(new_n6926));
  OAI211xp5_ASAP7_75t_L     g06670(.A1(new_n6625), .A2(new_n6624), .B(new_n6663), .C(new_n6664), .Y(new_n6927));
  O2A1O1Ixp33_ASAP7_75t_L   g06671(.A1(new_n6668), .A2(new_n6666), .B(new_n6927), .C(new_n6923), .Y(new_n6928));
  A2O1A1Ixp33_ASAP7_75t_L   g06672(.A1(new_n6660), .A2(new_n6665), .B(new_n6668), .C(new_n6927), .Y(new_n6929));
  NOR2xp33_ASAP7_75t_L      g06673(.A(new_n6918), .B(new_n6929), .Y(new_n6930));
  NOR3xp33_ASAP7_75t_L      g06674(.A(new_n6930), .B(new_n6926), .C(new_n6928), .Y(new_n6931));
  OAI21xp33_ASAP7_75t_L     g06675(.A1(new_n6925), .A2(new_n6931), .B(new_n6865), .Y(new_n6932));
  AOI31xp33_ASAP7_75t_L     g06676(.A1(new_n6679), .A2(new_n6674), .A3(new_n6411), .B(new_n6682), .Y(new_n6933));
  OAI21xp33_ASAP7_75t_L     g06677(.A1(new_n6928), .A2(new_n6930), .B(new_n6926), .Y(new_n6934));
  NAND3xp33_ASAP7_75t_L     g06678(.A(new_n6919), .B(new_n6868), .C(new_n6924), .Y(new_n6935));
  NAND3xp33_ASAP7_75t_L     g06679(.A(new_n6933), .B(new_n6934), .C(new_n6935), .Y(new_n6936));
  NAND3xp33_ASAP7_75t_L     g06680(.A(new_n6864), .B(new_n6932), .C(new_n6936), .Y(new_n6937));
  AOI21xp33_ASAP7_75t_L     g06681(.A1(new_n6935), .A2(new_n6934), .B(new_n6933), .Y(new_n6938));
  NOR3xp33_ASAP7_75t_L      g06682(.A(new_n6865), .B(new_n6925), .C(new_n6931), .Y(new_n6939));
  OAI21xp33_ASAP7_75t_L     g06683(.A1(new_n6938), .A2(new_n6939), .B(new_n6863), .Y(new_n6940));
  NAND3xp33_ASAP7_75t_L     g06684(.A(new_n6860), .B(new_n6937), .C(new_n6940), .Y(new_n6941));
  A2O1A1O1Ixp25_ASAP7_75t_L g06685(.A1(new_n6434), .A2(new_n6423), .B(new_n6422), .C(new_n6693), .D(new_n6858), .Y(new_n6942));
  NAND2xp33_ASAP7_75t_L     g06686(.A(new_n6937), .B(new_n6940), .Y(new_n6943));
  NAND2xp33_ASAP7_75t_L     g06687(.A(new_n6943), .B(new_n6942), .Y(new_n6944));
  OAI22xp33_ASAP7_75t_L     g06688(.A1(new_n3402), .A2(new_n1030), .B1(new_n1313), .B2(new_n3022), .Y(new_n6945));
  AOI221xp5_ASAP7_75t_L     g06689(.A1(new_n3030), .A2(\b[17] ), .B1(new_n3021), .B2(new_n1319), .C(new_n6945), .Y(new_n6946));
  XNOR2x2_ASAP7_75t_L       g06690(.A(new_n3015), .B(new_n6946), .Y(new_n6947));
  NAND3xp33_ASAP7_75t_L     g06691(.A(new_n6944), .B(new_n6941), .C(new_n6947), .Y(new_n6948));
  NOR2xp33_ASAP7_75t_L      g06692(.A(new_n6943), .B(new_n6942), .Y(new_n6949));
  AOI21xp33_ASAP7_75t_L     g06693(.A1(new_n6940), .A2(new_n6937), .B(new_n6860), .Y(new_n6950));
  INVx1_ASAP7_75t_L         g06694(.A(new_n6947), .Y(new_n6951));
  OAI21xp33_ASAP7_75t_L     g06695(.A1(new_n6950), .A2(new_n6949), .B(new_n6951), .Y(new_n6952));
  NAND2xp33_ASAP7_75t_L     g06696(.A(new_n6948), .B(new_n6952), .Y(new_n6953));
  NAND2xp33_ASAP7_75t_L     g06697(.A(new_n6696), .B(new_n6694), .Y(new_n6954));
  MAJIxp5_ASAP7_75t_L       g06698(.A(new_n6701), .B(new_n6618), .C(new_n6954), .Y(new_n6955));
  NOR2xp33_ASAP7_75t_L      g06699(.A(new_n6955), .B(new_n6953), .Y(new_n6956));
  NOR3xp33_ASAP7_75t_L      g06700(.A(new_n6949), .B(new_n6950), .C(new_n6951), .Y(new_n6957));
  AOI21xp33_ASAP7_75t_L     g06701(.A1(new_n6944), .A2(new_n6941), .B(new_n6947), .Y(new_n6958));
  NOR2xp33_ASAP7_75t_L      g06702(.A(new_n6958), .B(new_n6957), .Y(new_n6959));
  NOR2xp33_ASAP7_75t_L      g06703(.A(new_n6618), .B(new_n6954), .Y(new_n6960));
  O2A1O1Ixp33_ASAP7_75t_L   g06704(.A1(new_n6697), .A2(new_n6698), .B(new_n6615), .C(new_n6960), .Y(new_n6961));
  NOR2xp33_ASAP7_75t_L      g06705(.A(new_n6959), .B(new_n6961), .Y(new_n6962));
  AOI22xp33_ASAP7_75t_L     g06706(.A1(new_n2552), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n2736), .Y(new_n6963));
  OAI221xp5_ASAP7_75t_L     g06707(.A1(new_n2547), .A2(new_n1539), .B1(new_n2734), .B2(new_n1662), .C(new_n6963), .Y(new_n6964));
  XNOR2x2_ASAP7_75t_L       g06708(.A(\a[29] ), .B(new_n6964), .Y(new_n6965));
  INVx1_ASAP7_75t_L         g06709(.A(new_n6965), .Y(new_n6966));
  NOR3xp33_ASAP7_75t_L      g06710(.A(new_n6962), .B(new_n6966), .C(new_n6956), .Y(new_n6967));
  NAND2xp33_ASAP7_75t_L     g06711(.A(new_n6959), .B(new_n6961), .Y(new_n6968));
  OAI21xp33_ASAP7_75t_L     g06712(.A1(new_n6957), .A2(new_n6958), .B(new_n6955), .Y(new_n6969));
  AOI21xp33_ASAP7_75t_L     g06713(.A1(new_n6968), .A2(new_n6969), .B(new_n6965), .Y(new_n6970));
  AOI21xp33_ASAP7_75t_L     g06714(.A1(new_n6700), .A2(new_n6702), .B(new_n6707), .Y(new_n6971));
  AO21x2_ASAP7_75t_L        g06715(.A1(new_n6709), .A2(new_n6611), .B(new_n6971), .Y(new_n6972));
  NOR3xp33_ASAP7_75t_L      g06716(.A(new_n6972), .B(new_n6970), .C(new_n6967), .Y(new_n6973));
  NAND3xp33_ASAP7_75t_L     g06717(.A(new_n6968), .B(new_n6969), .C(new_n6965), .Y(new_n6974));
  OAI21xp33_ASAP7_75t_L     g06718(.A1(new_n6956), .A2(new_n6962), .B(new_n6966), .Y(new_n6975));
  AOI21xp33_ASAP7_75t_L     g06719(.A1(new_n6611), .A2(new_n6709), .B(new_n6971), .Y(new_n6976));
  AOI21xp33_ASAP7_75t_L     g06720(.A1(new_n6975), .A2(new_n6974), .B(new_n6976), .Y(new_n6977));
  OAI22xp33_ASAP7_75t_L     g06721(.A1(new_n2269), .A2(new_n1774), .B1(new_n1929), .B2(new_n2107), .Y(new_n6978));
  AOI221xp5_ASAP7_75t_L     g06722(.A1(new_n2115), .A2(\b[23] ), .B1(new_n2106), .B2(new_n1935), .C(new_n6978), .Y(new_n6979));
  AND2x2_ASAP7_75t_L        g06723(.A(\a[26] ), .B(new_n6979), .Y(new_n6980));
  NOR2xp33_ASAP7_75t_L      g06724(.A(\a[26] ), .B(new_n6979), .Y(new_n6981));
  NOR2xp33_ASAP7_75t_L      g06725(.A(new_n6981), .B(new_n6980), .Y(new_n6982));
  OAI21xp33_ASAP7_75t_L     g06726(.A1(new_n6977), .A2(new_n6973), .B(new_n6982), .Y(new_n6983));
  NAND3xp33_ASAP7_75t_L     g06727(.A(new_n6976), .B(new_n6975), .C(new_n6974), .Y(new_n6984));
  OAI21xp33_ASAP7_75t_L     g06728(.A1(new_n6967), .A2(new_n6970), .B(new_n6972), .Y(new_n6985));
  OAI211xp5_ASAP7_75t_L     g06729(.A1(new_n6980), .A2(new_n6981), .B(new_n6985), .C(new_n6984), .Y(new_n6986));
  OAI211xp5_ASAP7_75t_L     g06730(.A1(new_n6471), .A2(new_n6472), .B(new_n6720), .C(new_n6716), .Y(new_n6987));
  NAND4xp25_ASAP7_75t_L     g06731(.A(new_n6987), .B(new_n6715), .C(new_n6983), .D(new_n6986), .Y(new_n6988));
  AO22x1_ASAP7_75t_L        g06732(.A1(new_n6983), .A2(new_n6986), .B1(new_n6715), .B2(new_n6987), .Y(new_n6989));
  NAND2xp33_ASAP7_75t_L     g06733(.A(\b[26] ), .B(new_n1706), .Y(new_n6990));
  NAND2xp33_ASAP7_75t_L     g06734(.A(new_n1695), .B(new_n2504), .Y(new_n6991));
  AOI22xp33_ASAP7_75t_L     g06735(.A1(new_n1704), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1837), .Y(new_n6992));
  AND4x1_ASAP7_75t_L        g06736(.A(new_n6992), .B(new_n6991), .C(new_n6990), .D(\a[23] ), .Y(new_n6993));
  AOI31xp33_ASAP7_75t_L     g06737(.A1(new_n6991), .A2(new_n6990), .A3(new_n6992), .B(\a[23] ), .Y(new_n6994));
  NOR2xp33_ASAP7_75t_L      g06738(.A(new_n6994), .B(new_n6993), .Y(new_n6995));
  NAND3xp33_ASAP7_75t_L     g06739(.A(new_n6989), .B(new_n6988), .C(new_n6995), .Y(new_n6996));
  AND4x1_ASAP7_75t_L        g06740(.A(new_n6987), .B(new_n6986), .C(new_n6983), .D(new_n6715), .Y(new_n6997));
  AOI22xp33_ASAP7_75t_L     g06741(.A1(new_n6986), .A2(new_n6983), .B1(new_n6715), .B2(new_n6987), .Y(new_n6998));
  OAI22xp33_ASAP7_75t_L     g06742(.A1(new_n6997), .A2(new_n6998), .B1(new_n6994), .B2(new_n6993), .Y(new_n6999));
  NAND2xp33_ASAP7_75t_L     g06743(.A(new_n6996), .B(new_n6999), .Y(new_n7000));
  A2O1A1Ixp33_ASAP7_75t_L   g06744(.A1(new_n6730), .A2(new_n6729), .B(new_n6726), .C(new_n7000), .Y(new_n7001));
  NAND2xp33_ASAP7_75t_L     g06745(.A(new_n6484), .B(new_n6485), .Y(new_n7002));
  NOR2xp33_ASAP7_75t_L      g06746(.A(new_n6480), .B(new_n6728), .Y(new_n7003));
  A2O1A1O1Ixp25_ASAP7_75t_L g06747(.A1(new_n6482), .A2(new_n7002), .B(new_n7003), .C(new_n6730), .D(new_n6726), .Y(new_n7004));
  NAND3xp33_ASAP7_75t_L     g06748(.A(new_n7004), .B(new_n6996), .C(new_n6999), .Y(new_n7005));
  NAND3xp33_ASAP7_75t_L     g06749(.A(new_n7001), .B(new_n7005), .C(new_n6857), .Y(new_n7006));
  AOI21xp33_ASAP7_75t_L     g06750(.A1(new_n6999), .A2(new_n6996), .B(new_n7004), .Y(new_n7007));
  NAND2xp33_ASAP7_75t_L     g06751(.A(new_n6476), .B(new_n6602), .Y(new_n7008));
  A2O1A1Ixp33_ASAP7_75t_L   g06752(.A1(new_n6483), .A2(new_n7008), .B(new_n6723), .C(new_n6731), .Y(new_n7009));
  NOR2xp33_ASAP7_75t_L      g06753(.A(new_n7000), .B(new_n7009), .Y(new_n7010));
  OAI21xp33_ASAP7_75t_L     g06754(.A1(new_n7007), .A2(new_n7010), .B(new_n6856), .Y(new_n7011));
  NAND3xp33_ASAP7_75t_L     g06755(.A(new_n6853), .B(new_n7006), .C(new_n7011), .Y(new_n7012));
  A2O1A1O1Ixp25_ASAP7_75t_L g06756(.A1(new_n6506), .A2(new_n6498), .B(new_n6740), .C(new_n6733), .D(new_n6745), .Y(new_n7013));
  NAND2xp33_ASAP7_75t_L     g06757(.A(new_n7011), .B(new_n7006), .Y(new_n7014));
  NAND2xp33_ASAP7_75t_L     g06758(.A(new_n7013), .B(new_n7014), .Y(new_n7015));
  AOI22xp33_ASAP7_75t_L     g06759(.A1(new_n1076), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1253), .Y(new_n7016));
  OAI221xp5_ASAP7_75t_L     g06760(.A1(new_n1154), .A2(new_n3207), .B1(new_n1156), .B2(new_n3572), .C(new_n7016), .Y(new_n7017));
  XNOR2x2_ASAP7_75t_L       g06761(.A(\a[17] ), .B(new_n7017), .Y(new_n7018));
  NAND3xp33_ASAP7_75t_L     g06762(.A(new_n7012), .B(new_n7015), .C(new_n7018), .Y(new_n7019));
  O2A1O1Ixp33_ASAP7_75t_L   g06763(.A1(new_n6598), .A2(new_n6744), .B(new_n6737), .C(new_n7014), .Y(new_n7020));
  AOI21xp33_ASAP7_75t_L     g06764(.A1(new_n7011), .A2(new_n7006), .B(new_n6853), .Y(new_n7021));
  INVx1_ASAP7_75t_L         g06765(.A(new_n7018), .Y(new_n7022));
  OAI21xp33_ASAP7_75t_L     g06766(.A1(new_n7021), .A2(new_n7020), .B(new_n7022), .Y(new_n7023));
  AO21x2_ASAP7_75t_L        g06767(.A1(new_n7023), .A2(new_n7019), .B(new_n6852), .Y(new_n7024));
  NAND3xp33_ASAP7_75t_L     g06768(.A(new_n6852), .B(new_n7019), .C(new_n7023), .Y(new_n7025));
  NAND3xp33_ASAP7_75t_L     g06769(.A(new_n7024), .B(new_n6851), .C(new_n7025), .Y(new_n7026));
  XNOR2x2_ASAP7_75t_L       g06770(.A(new_n806), .B(new_n6850), .Y(new_n7027));
  AOI21xp33_ASAP7_75t_L     g06771(.A1(new_n7019), .A2(new_n7023), .B(new_n6852), .Y(new_n7028));
  AND3x1_ASAP7_75t_L        g06772(.A(new_n6852), .B(new_n7023), .C(new_n7019), .Y(new_n7029));
  OAI21xp33_ASAP7_75t_L     g06773(.A1(new_n7028), .A2(new_n7029), .B(new_n7027), .Y(new_n7030));
  NAND2xp33_ASAP7_75t_L     g06774(.A(new_n7026), .B(new_n7030), .Y(new_n7031));
  NAND3xp33_ASAP7_75t_L     g06775(.A(new_n6846), .B(new_n7031), .C(new_n6847), .Y(new_n7032));
  INVx1_ASAP7_75t_L         g06776(.A(new_n6847), .Y(new_n7033));
  NOR3xp33_ASAP7_75t_L      g06777(.A(new_n7029), .B(new_n7028), .C(new_n7027), .Y(new_n7034));
  AOI21xp33_ASAP7_75t_L     g06778(.A1(new_n7024), .A2(new_n7025), .B(new_n6851), .Y(new_n7035));
  NOR2xp33_ASAP7_75t_L      g06779(.A(new_n7035), .B(new_n7034), .Y(new_n7036));
  A2O1A1Ixp33_ASAP7_75t_L   g06780(.A1(new_n6770), .A2(new_n6767), .B(new_n7033), .C(new_n7036), .Y(new_n7037));
  AOI22xp33_ASAP7_75t_L     g06781(.A1(\b[37] ), .A2(new_n651), .B1(\b[39] ), .B2(new_n581), .Y(new_n7038));
  OAI221xp5_ASAP7_75t_L     g06782(.A1(new_n821), .A2(new_n4632), .B1(new_n577), .B2(new_n4858), .C(new_n7038), .Y(new_n7039));
  XNOR2x2_ASAP7_75t_L       g06783(.A(\a[11] ), .B(new_n7039), .Y(new_n7040));
  NAND3xp33_ASAP7_75t_L     g06784(.A(new_n7037), .B(new_n7032), .C(new_n7040), .Y(new_n7041));
  A2O1A1Ixp33_ASAP7_75t_L   g06785(.A1(new_n6766), .A2(new_n6762), .B(new_n6773), .C(new_n6847), .Y(new_n7042));
  NOR2xp33_ASAP7_75t_L      g06786(.A(new_n7036), .B(new_n7042), .Y(new_n7043));
  A2O1A1O1Ixp25_ASAP7_75t_L g06787(.A1(new_n6766), .A2(new_n6762), .B(new_n6773), .C(new_n6847), .D(new_n7031), .Y(new_n7044));
  INVx1_ASAP7_75t_L         g06788(.A(new_n7040), .Y(new_n7045));
  OAI21xp33_ASAP7_75t_L     g06789(.A1(new_n7043), .A2(new_n7044), .B(new_n7045), .Y(new_n7046));
  NOR2xp33_ASAP7_75t_L      g06790(.A(new_n6774), .B(new_n6771), .Y(new_n7047));
  MAJIxp5_ASAP7_75t_L       g06791(.A(new_n6782), .B(new_n6777), .C(new_n7047), .Y(new_n7048));
  AND3x1_ASAP7_75t_L        g06792(.A(new_n7048), .B(new_n7046), .C(new_n7041), .Y(new_n7049));
  AOI21xp33_ASAP7_75t_L     g06793(.A1(new_n7046), .A2(new_n7041), .B(new_n7048), .Y(new_n7050));
  NOR2xp33_ASAP7_75t_L      g06794(.A(new_n7050), .B(new_n7049), .Y(new_n7051));
  AOI22xp33_ASAP7_75t_L     g06795(.A1(new_n444), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n471), .Y(new_n7052));
  OAI221xp5_ASAP7_75t_L     g06796(.A1(new_n468), .A2(new_n5321), .B1(new_n469), .B2(new_n5346), .C(new_n7052), .Y(new_n7053));
  XNOR2x2_ASAP7_75t_L       g06797(.A(\a[8] ), .B(new_n7053), .Y(new_n7054));
  NAND2xp33_ASAP7_75t_L     g06798(.A(new_n7054), .B(new_n7051), .Y(new_n7055));
  NAND3xp33_ASAP7_75t_L     g06799(.A(new_n7048), .B(new_n7046), .C(new_n7041), .Y(new_n7056));
  AO21x2_ASAP7_75t_L        g06800(.A1(new_n7041), .A2(new_n7046), .B(new_n7048), .Y(new_n7057));
  NAND2xp33_ASAP7_75t_L     g06801(.A(new_n7056), .B(new_n7057), .Y(new_n7058));
  INVx1_ASAP7_75t_L         g06802(.A(new_n7054), .Y(new_n7059));
  NAND2xp33_ASAP7_75t_L     g06803(.A(new_n7059), .B(new_n7058), .Y(new_n7060));
  OAI21xp33_ASAP7_75t_L     g06804(.A1(new_n6796), .A2(new_n6802), .B(new_n6799), .Y(new_n7061));
  NAND3xp33_ASAP7_75t_L     g06805(.A(new_n7055), .B(new_n7060), .C(new_n7061), .Y(new_n7062));
  AO21x2_ASAP7_75t_L        g06806(.A1(new_n7060), .A2(new_n7055), .B(new_n7061), .Y(new_n7063));
  NOR2xp33_ASAP7_75t_L      g06807(.A(new_n5829), .B(new_n429), .Y(new_n7064));
  INVx1_ASAP7_75t_L         g06808(.A(new_n7064), .Y(new_n7065));
  INVx1_ASAP7_75t_L         g06809(.A(new_n6329), .Y(new_n7066));
  NAND2xp33_ASAP7_75t_L     g06810(.A(new_n341), .B(new_n7066), .Y(new_n7067));
  AOI22xp33_ASAP7_75t_L     g06811(.A1(new_n344), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n370), .Y(new_n7068));
  AND4x1_ASAP7_75t_L        g06812(.A(new_n7068), .B(new_n7067), .C(new_n7065), .D(\a[5] ), .Y(new_n7069));
  AOI31xp33_ASAP7_75t_L     g06813(.A1(new_n7067), .A2(new_n7065), .A3(new_n7068), .B(\a[5] ), .Y(new_n7070));
  NOR2xp33_ASAP7_75t_L      g06814(.A(new_n7070), .B(new_n7069), .Y(new_n7071));
  AOI21xp33_ASAP7_75t_L     g06815(.A1(new_n7063), .A2(new_n7062), .B(new_n7071), .Y(new_n7072));
  AND3x1_ASAP7_75t_L        g06816(.A(new_n7063), .B(new_n7071), .C(new_n7062), .Y(new_n7073));
  NOR3xp33_ASAP7_75t_L      g06817(.A(new_n6845), .B(new_n7072), .C(new_n7073), .Y(new_n7074));
  INVx1_ASAP7_75t_L         g06818(.A(new_n7072), .Y(new_n7075));
  NAND3xp33_ASAP7_75t_L     g06819(.A(new_n7063), .B(new_n7062), .C(new_n7071), .Y(new_n7076));
  AOI221xp5_ASAP7_75t_L     g06820(.A1(new_n6809), .A2(new_n6584), .B1(new_n7076), .B2(new_n7075), .C(new_n6808), .Y(new_n7077));
  OAI21xp33_ASAP7_75t_L     g06821(.A1(new_n7074), .A2(new_n7077), .B(new_n6840), .Y(new_n7078));
  NOR3xp33_ASAP7_75t_L      g06822(.A(new_n7077), .B(new_n7074), .C(new_n6840), .Y(new_n7079));
  INVx1_ASAP7_75t_L         g06823(.A(new_n7079), .Y(new_n7080));
  NAND2xp33_ASAP7_75t_L     g06824(.A(new_n7078), .B(new_n7080), .Y(new_n7081));
  O2A1O1Ixp33_ASAP7_75t_L   g06825(.A1(new_n6810), .A2(new_n6823), .B(new_n6827), .C(new_n7081), .Y(new_n7082));
  MAJIxp5_ASAP7_75t_L       g06826(.A(new_n6825), .B(new_n6810), .C(new_n6823), .Y(new_n7083));
  AOI21xp33_ASAP7_75t_L     g06827(.A1(new_n7080), .A2(new_n7078), .B(new_n7083), .Y(new_n7084));
  NOR2xp33_ASAP7_75t_L      g06828(.A(new_n7084), .B(new_n7082), .Y(\f[48] ));
  INVx1_ASAP7_75t_L         g06829(.A(new_n7083), .Y(new_n7086));
  NOR3xp33_ASAP7_75t_L      g06830(.A(new_n6997), .B(new_n6998), .C(new_n6995), .Y(new_n7087));
  OAI22xp33_ASAP7_75t_L     g06831(.A1(new_n1829), .A2(new_n2348), .B1(new_n2666), .B2(new_n1696), .Y(new_n7088));
  AOI221xp5_ASAP7_75t_L     g06832(.A1(\b[27] ), .A2(new_n1706), .B1(new_n1695), .B2(new_n4237), .C(new_n7088), .Y(new_n7089));
  XNOR2x2_ASAP7_75t_L       g06833(.A(new_n1689), .B(new_n7089), .Y(new_n7090));
  NAND2xp33_ASAP7_75t_L     g06834(.A(new_n6924), .B(new_n6919), .Y(new_n7091));
  MAJIxp5_ASAP7_75t_L       g06835(.A(new_n6933), .B(new_n6868), .C(new_n7091), .Y(new_n7092));
  AOI22xp33_ASAP7_75t_L     g06836(.A1(new_n4283), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n4512), .Y(new_n7093));
  OAI221xp5_ASAP7_75t_L     g06837(.A1(new_n4277), .A2(new_n760), .B1(new_n4499), .B2(new_n790), .C(new_n7093), .Y(new_n7094));
  XNOR2x2_ASAP7_75t_L       g06838(.A(\a[38] ), .B(new_n7094), .Y(new_n7095));
  NOR3xp33_ASAP7_75t_L      g06839(.A(new_n6650), .B(new_n6878), .C(new_n6870), .Y(new_n7096));
  NAND2xp33_ASAP7_75t_L     g06840(.A(\b[3] ), .B(new_n6380), .Y(new_n7097));
  AOI22xp33_ASAP7_75t_L     g06841(.A1(new_n6376), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n6648), .Y(new_n7098));
  OA21x2_ASAP7_75t_L        g06842(.A1(new_n6636), .A2(new_n330), .B(new_n7098), .Y(new_n7099));
  NAND3xp33_ASAP7_75t_L     g06843(.A(new_n7099), .B(new_n7097), .C(\a[47] ), .Y(new_n7100));
  OAI211xp5_ASAP7_75t_L     g06844(.A1(new_n6636), .A2(new_n330), .B(new_n7097), .C(new_n7098), .Y(new_n7101));
  NAND2xp33_ASAP7_75t_L     g06845(.A(new_n6371), .B(new_n7101), .Y(new_n7102));
  NAND2xp33_ASAP7_75t_L     g06846(.A(\a[50] ), .B(new_n6875), .Y(new_n7103));
  INVx1_ASAP7_75t_L         g06847(.A(\a[49] ), .Y(new_n7104));
  NAND2xp33_ASAP7_75t_L     g06848(.A(\a[50] ), .B(new_n7104), .Y(new_n7105));
  INVx1_ASAP7_75t_L         g06849(.A(\a[50] ), .Y(new_n7106));
  NAND2xp33_ASAP7_75t_L     g06850(.A(\a[49] ), .B(new_n7106), .Y(new_n7107));
  AOI21xp33_ASAP7_75t_L     g06851(.A1(new_n7107), .A2(new_n7105), .B(new_n6874), .Y(new_n7108));
  NAND2xp33_ASAP7_75t_L     g06852(.A(new_n269), .B(new_n7108), .Y(new_n7109));
  NAND2xp33_ASAP7_75t_L     g06853(.A(new_n7107), .B(new_n7105), .Y(new_n7110));
  NOR2xp33_ASAP7_75t_L      g06854(.A(new_n7110), .B(new_n6874), .Y(new_n7111));
  NAND2xp33_ASAP7_75t_L     g06855(.A(\b[1] ), .B(new_n7111), .Y(new_n7112));
  NAND2xp33_ASAP7_75t_L     g06856(.A(new_n6873), .B(new_n6872), .Y(new_n7113));
  XNOR2x2_ASAP7_75t_L       g06857(.A(\a[49] ), .B(\a[48] ), .Y(new_n7114));
  NOR2xp33_ASAP7_75t_L      g06858(.A(new_n7114), .B(new_n7113), .Y(new_n7115));
  NAND2xp33_ASAP7_75t_L     g06859(.A(\b[0] ), .B(new_n7115), .Y(new_n7116));
  NAND3xp33_ASAP7_75t_L     g06860(.A(new_n7109), .B(new_n7112), .C(new_n7116), .Y(new_n7117));
  XOR2x2_ASAP7_75t_L        g06861(.A(new_n7103), .B(new_n7117), .Y(new_n7118));
  NAND3xp33_ASAP7_75t_L     g06862(.A(new_n7100), .B(new_n7102), .C(new_n7118), .Y(new_n7119));
  NOR2xp33_ASAP7_75t_L      g06863(.A(new_n6371), .B(new_n7101), .Y(new_n7120));
  O2A1O1Ixp33_ASAP7_75t_L   g06864(.A1(new_n298), .A2(new_n6646), .B(new_n7099), .C(\a[47] ), .Y(new_n7121));
  XNOR2x2_ASAP7_75t_L       g06865(.A(new_n7103), .B(new_n7117), .Y(new_n7122));
  OAI21xp33_ASAP7_75t_L     g06866(.A1(new_n7120), .A2(new_n7121), .B(new_n7122), .Y(new_n7123));
  OAI211xp5_ASAP7_75t_L     g06867(.A1(new_n7096), .A2(new_n6897), .B(new_n7119), .C(new_n7123), .Y(new_n7124));
  NOR2xp33_ASAP7_75t_L      g06868(.A(new_n6870), .B(new_n6650), .Y(new_n7125));
  NAND2xp33_ASAP7_75t_L     g06869(.A(new_n6886), .B(new_n6883), .Y(new_n7126));
  MAJIxp5_ASAP7_75t_L       g06870(.A(new_n7126), .B(new_n6875), .C(new_n7125), .Y(new_n7127));
  NOR3xp33_ASAP7_75t_L      g06871(.A(new_n7121), .B(new_n7122), .C(new_n7120), .Y(new_n7128));
  AOI21xp33_ASAP7_75t_L     g06872(.A1(new_n7100), .A2(new_n7102), .B(new_n7118), .Y(new_n7129));
  OAI21xp33_ASAP7_75t_L     g06873(.A1(new_n7129), .A2(new_n7128), .B(new_n7127), .Y(new_n7130));
  AOI22xp33_ASAP7_75t_L     g06874(.A1(new_n5624), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n5901), .Y(new_n7131));
  OAI221xp5_ASAP7_75t_L     g06875(.A1(new_n5900), .A2(new_n418), .B1(new_n5892), .B2(new_n425), .C(new_n7131), .Y(new_n7132));
  XNOR2x2_ASAP7_75t_L       g06876(.A(\a[44] ), .B(new_n7132), .Y(new_n7133));
  NAND3xp33_ASAP7_75t_L     g06877(.A(new_n7124), .B(new_n7130), .C(new_n7133), .Y(new_n7134));
  AO21x2_ASAP7_75t_L        g06878(.A1(new_n7130), .A2(new_n7124), .B(new_n7133), .Y(new_n7135));
  NAND2xp33_ASAP7_75t_L     g06879(.A(new_n7134), .B(new_n7135), .Y(new_n7136));
  AOI211xp5_ASAP7_75t_L     g06880(.A1(new_n6895), .A2(new_n6893), .B(new_n6897), .C(new_n6898), .Y(new_n7137));
  INVx1_ASAP7_75t_L         g06881(.A(new_n7137), .Y(new_n7138));
  A2O1A1Ixp33_ASAP7_75t_L   g06882(.A1(new_n6900), .A2(new_n6896), .B(new_n6903), .C(new_n7138), .Y(new_n7139));
  NOR2xp33_ASAP7_75t_L      g06883(.A(new_n7136), .B(new_n7139), .Y(new_n7140));
  A2O1A1O1Ixp25_ASAP7_75t_L g06884(.A1(new_n6658), .A2(new_n6657), .B(new_n6902), .C(new_n6905), .D(new_n7137), .Y(new_n7141));
  AOI21xp33_ASAP7_75t_L     g06885(.A1(new_n7135), .A2(new_n7134), .B(new_n7141), .Y(new_n7142));
  AOI22xp33_ASAP7_75t_L     g06886(.A1(new_n4920), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n5167), .Y(new_n7143));
  OAI221xp5_ASAP7_75t_L     g06887(.A1(new_n5154), .A2(new_n540), .B1(new_n5158), .B2(new_n624), .C(new_n7143), .Y(new_n7144));
  XNOR2x2_ASAP7_75t_L       g06888(.A(\a[41] ), .B(new_n7144), .Y(new_n7145));
  OAI21xp33_ASAP7_75t_L     g06889(.A1(new_n7142), .A2(new_n7140), .B(new_n7145), .Y(new_n7146));
  NAND3xp33_ASAP7_75t_L     g06890(.A(new_n7141), .B(new_n7135), .C(new_n7134), .Y(new_n7147));
  A2O1A1Ixp33_ASAP7_75t_L   g06891(.A1(new_n6905), .A2(new_n6913), .B(new_n7137), .C(new_n7136), .Y(new_n7148));
  INVx1_ASAP7_75t_L         g06892(.A(new_n7145), .Y(new_n7149));
  NAND3xp33_ASAP7_75t_L     g06893(.A(new_n7148), .B(new_n7147), .C(new_n7149), .Y(new_n7150));
  AOI221xp5_ASAP7_75t_L     g06894(.A1(new_n6929), .A2(new_n6918), .B1(new_n7146), .B2(new_n7150), .C(new_n6917), .Y(new_n7151));
  A2O1A1O1Ixp25_ASAP7_75t_L g06895(.A1(new_n6669), .A2(new_n6621), .B(new_n6869), .C(new_n6921), .D(new_n6917), .Y(new_n7152));
  INVx1_ASAP7_75t_L         g06896(.A(new_n7146), .Y(new_n7153));
  NOR3xp33_ASAP7_75t_L      g06897(.A(new_n7140), .B(new_n7142), .C(new_n7145), .Y(new_n7154));
  NOR3xp33_ASAP7_75t_L      g06898(.A(new_n7153), .B(new_n7154), .C(new_n7152), .Y(new_n7155));
  OAI21xp33_ASAP7_75t_L     g06899(.A1(new_n7151), .A2(new_n7155), .B(new_n7095), .Y(new_n7156));
  OR3x1_ASAP7_75t_L         g06900(.A(new_n7155), .B(new_n7095), .C(new_n7151), .Y(new_n7157));
  NAND3xp33_ASAP7_75t_L     g06901(.A(new_n7092), .B(new_n7157), .C(new_n7156), .Y(new_n7158));
  NOR2xp33_ASAP7_75t_L      g06902(.A(new_n6928), .B(new_n6930), .Y(new_n7159));
  MAJIxp5_ASAP7_75t_L       g06903(.A(new_n6865), .B(new_n6926), .C(new_n7159), .Y(new_n7160));
  INVx1_ASAP7_75t_L         g06904(.A(new_n7156), .Y(new_n7161));
  NOR3xp33_ASAP7_75t_L      g06905(.A(new_n7155), .B(new_n7151), .C(new_n7095), .Y(new_n7162));
  OAI21xp33_ASAP7_75t_L     g06906(.A1(new_n7162), .A2(new_n7161), .B(new_n7160), .Y(new_n7163));
  AOI22xp33_ASAP7_75t_L     g06907(.A1(new_n3633), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n3858), .Y(new_n7164));
  OAI221xp5_ASAP7_75t_L     g06908(.A1(new_n3853), .A2(new_n942), .B1(new_n3856), .B2(new_n1035), .C(new_n7164), .Y(new_n7165));
  XNOR2x2_ASAP7_75t_L       g06909(.A(\a[35] ), .B(new_n7165), .Y(new_n7166));
  NAND3xp33_ASAP7_75t_L     g06910(.A(new_n7163), .B(new_n7158), .C(new_n7166), .Y(new_n7167));
  AO21x2_ASAP7_75t_L        g06911(.A1(new_n7158), .A2(new_n7163), .B(new_n7166), .Y(new_n7168));
  NAND3xp33_ASAP7_75t_L     g06912(.A(new_n6167), .B(new_n6172), .C(new_n6174), .Y(new_n7169));
  A2O1A1Ixp33_ASAP7_75t_L   g06913(.A1(new_n6179), .A2(new_n7169), .B(new_n6421), .C(new_n6426), .Y(new_n7170));
  NOR3xp33_ASAP7_75t_L      g06914(.A(new_n6939), .B(new_n6938), .C(new_n6863), .Y(new_n7171));
  A2O1A1O1Ixp25_ASAP7_75t_L g06915(.A1(new_n6693), .A2(new_n7170), .B(new_n6858), .C(new_n6940), .D(new_n7171), .Y(new_n7172));
  NAND3xp33_ASAP7_75t_L     g06916(.A(new_n7172), .B(new_n7168), .C(new_n7167), .Y(new_n7173));
  AO21x2_ASAP7_75t_L        g06917(.A1(new_n7167), .A2(new_n7168), .B(new_n7172), .Y(new_n7174));
  AOI22xp33_ASAP7_75t_L     g06918(.A1(new_n3029), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n3258), .Y(new_n7175));
  OAI221xp5_ASAP7_75t_L     g06919(.A1(new_n3024), .A2(new_n1313), .B1(new_n3256), .B2(new_n1438), .C(new_n7175), .Y(new_n7176));
  XNOR2x2_ASAP7_75t_L       g06920(.A(\a[32] ), .B(new_n7176), .Y(new_n7177));
  NAND3xp33_ASAP7_75t_L     g06921(.A(new_n7174), .B(new_n7173), .C(new_n7177), .Y(new_n7178));
  AND3x1_ASAP7_75t_L        g06922(.A(new_n7172), .B(new_n7168), .C(new_n7167), .Y(new_n7179));
  AOI21xp33_ASAP7_75t_L     g06923(.A1(new_n7168), .A2(new_n7167), .B(new_n7172), .Y(new_n7180));
  INVx1_ASAP7_75t_L         g06924(.A(new_n7177), .Y(new_n7181));
  OAI21xp33_ASAP7_75t_L     g06925(.A1(new_n7180), .A2(new_n7179), .B(new_n7181), .Y(new_n7182));
  NAND2xp33_ASAP7_75t_L     g06926(.A(new_n7178), .B(new_n7182), .Y(new_n7183));
  NOR3xp33_ASAP7_75t_L      g06927(.A(new_n6949), .B(new_n6950), .C(new_n6947), .Y(new_n7184));
  AOI211xp5_ASAP7_75t_L     g06928(.A1(new_n6955), .A2(new_n6953), .B(new_n7184), .C(new_n7183), .Y(new_n7185));
  O2A1O1Ixp33_ASAP7_75t_L   g06929(.A1(new_n6957), .A2(new_n6958), .B(new_n6955), .C(new_n7184), .Y(new_n7186));
  AOI21xp33_ASAP7_75t_L     g06930(.A1(new_n7182), .A2(new_n7178), .B(new_n7186), .Y(new_n7187));
  AOI22xp33_ASAP7_75t_L     g06931(.A1(new_n2552), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n2736), .Y(new_n7188));
  OAI221xp5_ASAP7_75t_L     g06932(.A1(new_n2547), .A2(new_n1655), .B1(new_n2734), .B2(new_n1780), .C(new_n7188), .Y(new_n7189));
  XNOR2x2_ASAP7_75t_L       g06933(.A(\a[29] ), .B(new_n7189), .Y(new_n7190));
  INVx1_ASAP7_75t_L         g06934(.A(new_n7190), .Y(new_n7191));
  NOR3xp33_ASAP7_75t_L      g06935(.A(new_n7185), .B(new_n7187), .C(new_n7191), .Y(new_n7192));
  NAND3xp33_ASAP7_75t_L     g06936(.A(new_n7186), .B(new_n7182), .C(new_n7178), .Y(new_n7193));
  A2O1A1Ixp33_ASAP7_75t_L   g06937(.A1(new_n6953), .A2(new_n6955), .B(new_n7184), .C(new_n7183), .Y(new_n7194));
  AOI21xp33_ASAP7_75t_L     g06938(.A1(new_n7193), .A2(new_n7194), .B(new_n7190), .Y(new_n7195));
  XNOR2x2_ASAP7_75t_L       g06939(.A(new_n6955), .B(new_n6953), .Y(new_n7196));
  MAJIxp5_ASAP7_75t_L       g06940(.A(new_n6976), .B(new_n6965), .C(new_n7196), .Y(new_n7197));
  NOR3xp33_ASAP7_75t_L      g06941(.A(new_n7197), .B(new_n7195), .C(new_n7192), .Y(new_n7198));
  NAND3xp33_ASAP7_75t_L     g06942(.A(new_n7193), .B(new_n7194), .C(new_n7190), .Y(new_n7199));
  OAI21xp33_ASAP7_75t_L     g06943(.A1(new_n7187), .A2(new_n7185), .B(new_n7191), .Y(new_n7200));
  NOR2xp33_ASAP7_75t_L      g06944(.A(new_n6956), .B(new_n6962), .Y(new_n7201));
  MAJIxp5_ASAP7_75t_L       g06945(.A(new_n6972), .B(new_n6966), .C(new_n7201), .Y(new_n7202));
  AOI21xp33_ASAP7_75t_L     g06946(.A1(new_n7200), .A2(new_n7199), .B(new_n7202), .Y(new_n7203));
  OAI22xp33_ASAP7_75t_L     g06947(.A1(new_n2269), .A2(new_n1909), .B1(new_n2067), .B2(new_n2107), .Y(new_n7204));
  AOI221xp5_ASAP7_75t_L     g06948(.A1(new_n2115), .A2(\b[24] ), .B1(new_n2106), .B2(new_n2648), .C(new_n7204), .Y(new_n7205));
  XNOR2x2_ASAP7_75t_L       g06949(.A(\a[26] ), .B(new_n7205), .Y(new_n7206));
  NOR3xp33_ASAP7_75t_L      g06950(.A(new_n7203), .B(new_n7198), .C(new_n7206), .Y(new_n7207));
  NAND2xp33_ASAP7_75t_L     g06951(.A(new_n6966), .B(new_n7201), .Y(new_n7208));
  NAND4xp25_ASAP7_75t_L     g06952(.A(new_n6985), .B(new_n7208), .C(new_n7200), .D(new_n7199), .Y(new_n7209));
  OAI21xp33_ASAP7_75t_L     g06953(.A1(new_n7192), .A2(new_n7195), .B(new_n7197), .Y(new_n7210));
  XNOR2x2_ASAP7_75t_L       g06954(.A(new_n2100), .B(new_n7205), .Y(new_n7211));
  AOI21xp33_ASAP7_75t_L     g06955(.A1(new_n7209), .A2(new_n7210), .B(new_n7211), .Y(new_n7212));
  NOR3xp33_ASAP7_75t_L      g06956(.A(new_n6982), .B(new_n6973), .C(new_n6977), .Y(new_n7213));
  AO31x2_ASAP7_75t_L        g06957(.A1(new_n6987), .A2(new_n6983), .A3(new_n6715), .B(new_n7213), .Y(new_n7214));
  OAI21xp33_ASAP7_75t_L     g06958(.A1(new_n7207), .A2(new_n7212), .B(new_n7214), .Y(new_n7215));
  NAND3xp33_ASAP7_75t_L     g06959(.A(new_n7209), .B(new_n7210), .C(new_n7211), .Y(new_n7216));
  OAI21xp33_ASAP7_75t_L     g06960(.A1(new_n7198), .A2(new_n7203), .B(new_n7206), .Y(new_n7217));
  AOI31xp33_ASAP7_75t_L     g06961(.A1(new_n6987), .A2(new_n6983), .A3(new_n6715), .B(new_n7213), .Y(new_n7218));
  NAND3xp33_ASAP7_75t_L     g06962(.A(new_n7218), .B(new_n7217), .C(new_n7216), .Y(new_n7219));
  AOI21xp33_ASAP7_75t_L     g06963(.A1(new_n7215), .A2(new_n7219), .B(new_n7090), .Y(new_n7220));
  XNOR2x2_ASAP7_75t_L       g06964(.A(\a[23] ), .B(new_n7089), .Y(new_n7221));
  AOI21xp33_ASAP7_75t_L     g06965(.A1(new_n7217), .A2(new_n7216), .B(new_n7218), .Y(new_n7222));
  AND4x1_ASAP7_75t_L        g06966(.A(new_n6988), .B(new_n6986), .C(new_n7217), .D(new_n7216), .Y(new_n7223));
  NOR3xp33_ASAP7_75t_L      g06967(.A(new_n7223), .B(new_n7221), .C(new_n7222), .Y(new_n7224));
  NOR2xp33_ASAP7_75t_L      g06968(.A(new_n7220), .B(new_n7224), .Y(new_n7225));
  A2O1A1Ixp33_ASAP7_75t_L   g06969(.A1(new_n7000), .A2(new_n7009), .B(new_n7087), .C(new_n7225), .Y(new_n7226));
  AOI21xp33_ASAP7_75t_L     g06970(.A1(new_n7009), .A2(new_n7000), .B(new_n7087), .Y(new_n7227));
  OAI21xp33_ASAP7_75t_L     g06971(.A1(new_n7222), .A2(new_n7223), .B(new_n7221), .Y(new_n7228));
  NAND3xp33_ASAP7_75t_L     g06972(.A(new_n7215), .B(new_n7219), .C(new_n7090), .Y(new_n7229));
  NAND2xp33_ASAP7_75t_L     g06973(.A(new_n7229), .B(new_n7228), .Y(new_n7230));
  NAND2xp33_ASAP7_75t_L     g06974(.A(new_n7230), .B(new_n7227), .Y(new_n7231));
  AOI22xp33_ASAP7_75t_L     g06975(.A1(new_n1360), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1581), .Y(new_n7232));
  OAI221xp5_ASAP7_75t_L     g06976(.A1(new_n1373), .A2(new_n2982), .B1(new_n1359), .B2(new_n3187), .C(new_n7232), .Y(new_n7233));
  XNOR2x2_ASAP7_75t_L       g06977(.A(\a[20] ), .B(new_n7233), .Y(new_n7234));
  AOI21xp33_ASAP7_75t_L     g06978(.A1(new_n7226), .A2(new_n7231), .B(new_n7234), .Y(new_n7235));
  NOR2xp33_ASAP7_75t_L      g06979(.A(new_n7230), .B(new_n7227), .Y(new_n7236));
  INVx1_ASAP7_75t_L         g06980(.A(new_n7087), .Y(new_n7237));
  A2O1A1Ixp33_ASAP7_75t_L   g06981(.A1(new_n6996), .A2(new_n6999), .B(new_n7004), .C(new_n7237), .Y(new_n7238));
  NOR2xp33_ASAP7_75t_L      g06982(.A(new_n7238), .B(new_n7225), .Y(new_n7239));
  INVx1_ASAP7_75t_L         g06983(.A(new_n7234), .Y(new_n7240));
  NOR3xp33_ASAP7_75t_L      g06984(.A(new_n7236), .B(new_n7239), .C(new_n7240), .Y(new_n7241));
  OAI221xp5_ASAP7_75t_L     g06985(.A1(new_n7014), .A2(new_n7013), .B1(new_n7235), .B2(new_n7241), .C(new_n7006), .Y(new_n7242));
  AOI21xp33_ASAP7_75t_L     g06986(.A1(new_n7001), .A2(new_n7005), .B(new_n6857), .Y(new_n7243));
  OAI21xp33_ASAP7_75t_L     g06987(.A1(new_n7243), .A2(new_n7013), .B(new_n7006), .Y(new_n7244));
  OAI21xp33_ASAP7_75t_L     g06988(.A1(new_n7239), .A2(new_n7236), .B(new_n7240), .Y(new_n7245));
  NAND3xp33_ASAP7_75t_L     g06989(.A(new_n7226), .B(new_n7231), .C(new_n7234), .Y(new_n7246));
  NAND3xp33_ASAP7_75t_L     g06990(.A(new_n7244), .B(new_n7245), .C(new_n7246), .Y(new_n7247));
  NAND2xp33_ASAP7_75t_L     g06991(.A(\b[33] ), .B(new_n1080), .Y(new_n7248));
  NAND3xp33_ASAP7_75t_L     g06992(.A(new_n3587), .B(new_n1073), .C(new_n3590), .Y(new_n7249));
  AOI22xp33_ASAP7_75t_L     g06993(.A1(new_n1076), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1253), .Y(new_n7250));
  AND4x1_ASAP7_75t_L        g06994(.A(new_n7250), .B(new_n7249), .C(new_n7248), .D(\a[17] ), .Y(new_n7251));
  AOI31xp33_ASAP7_75t_L     g06995(.A1(new_n7249), .A2(new_n7248), .A3(new_n7250), .B(\a[17] ), .Y(new_n7252));
  NOR2xp33_ASAP7_75t_L      g06996(.A(new_n7252), .B(new_n7251), .Y(new_n7253));
  AND3x1_ASAP7_75t_L        g06997(.A(new_n7247), .B(new_n7242), .C(new_n7253), .Y(new_n7254));
  AOI21xp33_ASAP7_75t_L     g06998(.A1(new_n7247), .A2(new_n7242), .B(new_n7253), .Y(new_n7255));
  NOR2xp33_ASAP7_75t_L      g06999(.A(new_n7255), .B(new_n7254), .Y(new_n7256));
  OAI21xp33_ASAP7_75t_L     g07000(.A1(new_n6753), .A2(new_n6752), .B(new_n6749), .Y(new_n7257));
  NOR2xp33_ASAP7_75t_L      g07001(.A(new_n7021), .B(new_n7020), .Y(new_n7258));
  MAJIxp5_ASAP7_75t_L       g07002(.A(new_n7257), .B(new_n7258), .C(new_n7022), .Y(new_n7259));
  NAND2xp33_ASAP7_75t_L     g07003(.A(new_n7256), .B(new_n7259), .Y(new_n7260));
  NAND2xp33_ASAP7_75t_L     g07004(.A(new_n7015), .B(new_n7012), .Y(new_n7261));
  MAJIxp5_ASAP7_75t_L       g07005(.A(new_n6852), .B(new_n7018), .C(new_n7261), .Y(new_n7262));
  OAI21xp33_ASAP7_75t_L     g07006(.A1(new_n7254), .A2(new_n7255), .B(new_n7262), .Y(new_n7263));
  AOI22xp33_ASAP7_75t_L     g07007(.A1(new_n811), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n900), .Y(new_n7264));
  OAI221xp5_ASAP7_75t_L     g07008(.A1(new_n904), .A2(new_n4216), .B1(new_n898), .B2(new_n4431), .C(new_n7264), .Y(new_n7265));
  XNOR2x2_ASAP7_75t_L       g07009(.A(\a[14] ), .B(new_n7265), .Y(new_n7266));
  NAND3xp33_ASAP7_75t_L     g07010(.A(new_n7260), .B(new_n7266), .C(new_n7263), .Y(new_n7267));
  AO21x2_ASAP7_75t_L        g07011(.A1(new_n7263), .A2(new_n7260), .B(new_n7266), .Y(new_n7268));
  A2O1A1O1Ixp25_ASAP7_75t_L g07012(.A1(new_n6770), .A2(new_n6767), .B(new_n7033), .C(new_n7030), .D(new_n7034), .Y(new_n7269));
  NAND3xp33_ASAP7_75t_L     g07013(.A(new_n7269), .B(new_n7268), .C(new_n7267), .Y(new_n7270));
  AO21x2_ASAP7_75t_L        g07014(.A1(new_n7267), .A2(new_n7268), .B(new_n7269), .Y(new_n7271));
  NAND2xp33_ASAP7_75t_L     g07015(.A(new_n578), .B(new_n4876), .Y(new_n7272));
  AOI22xp33_ASAP7_75t_L     g07016(.A1(\b[38] ), .A2(new_n651), .B1(\b[40] ), .B2(new_n581), .Y(new_n7273));
  NAND2xp33_ASAP7_75t_L     g07017(.A(new_n7273), .B(new_n7272), .Y(new_n7274));
  AOI21xp33_ASAP7_75t_L     g07018(.A1(new_n584), .A2(\b[39] ), .B(new_n7274), .Y(new_n7275));
  NAND2xp33_ASAP7_75t_L     g07019(.A(\a[11] ), .B(new_n7275), .Y(new_n7276));
  A2O1A1Ixp33_ASAP7_75t_L   g07020(.A1(\b[39] ), .A2(new_n584), .B(new_n7274), .C(new_n574), .Y(new_n7277));
  NAND4xp25_ASAP7_75t_L     g07021(.A(new_n7271), .B(new_n7276), .C(new_n7277), .D(new_n7270), .Y(new_n7278));
  AND3x1_ASAP7_75t_L        g07022(.A(new_n7269), .B(new_n7268), .C(new_n7267), .Y(new_n7279));
  AOI21xp33_ASAP7_75t_L     g07023(.A1(new_n7268), .A2(new_n7267), .B(new_n7269), .Y(new_n7280));
  NAND2xp33_ASAP7_75t_L     g07024(.A(new_n7277), .B(new_n7276), .Y(new_n7281));
  OAI21xp33_ASAP7_75t_L     g07025(.A1(new_n7280), .A2(new_n7279), .B(new_n7281), .Y(new_n7282));
  NAND3xp33_ASAP7_75t_L     g07026(.A(new_n7037), .B(new_n7032), .C(new_n7045), .Y(new_n7283));
  NAND4xp25_ASAP7_75t_L     g07027(.A(new_n7057), .B(new_n7283), .C(new_n7282), .D(new_n7278), .Y(new_n7284));
  NAND2xp33_ASAP7_75t_L     g07028(.A(new_n7278), .B(new_n7282), .Y(new_n7285));
  A2O1A1Ixp33_ASAP7_75t_L   g07029(.A1(new_n7046), .A2(new_n7041), .B(new_n7048), .C(new_n7283), .Y(new_n7286));
  NAND2xp33_ASAP7_75t_L     g07030(.A(new_n7286), .B(new_n7285), .Y(new_n7287));
  AOI22xp33_ASAP7_75t_L     g07031(.A1(new_n444), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n471), .Y(new_n7288));
  INVx1_ASAP7_75t_L         g07032(.A(new_n7288), .Y(new_n7289));
  AOI221xp5_ASAP7_75t_L     g07033(.A1(\b[42] ), .A2(new_n447), .B1(new_n441), .B2(new_n5812), .C(new_n7289), .Y(new_n7290));
  AND2x2_ASAP7_75t_L        g07034(.A(\a[8] ), .B(new_n7290), .Y(new_n7291));
  NOR2xp33_ASAP7_75t_L      g07035(.A(\a[8] ), .B(new_n7290), .Y(new_n7292));
  NOR2xp33_ASAP7_75t_L      g07036(.A(new_n7292), .B(new_n7291), .Y(new_n7293));
  NAND3xp33_ASAP7_75t_L     g07037(.A(new_n7284), .B(new_n7287), .C(new_n7293), .Y(new_n7294));
  NOR2xp33_ASAP7_75t_L      g07038(.A(new_n7286), .B(new_n7285), .Y(new_n7295));
  AOI22xp33_ASAP7_75t_L     g07039(.A1(new_n7278), .A2(new_n7282), .B1(new_n7283), .B2(new_n7057), .Y(new_n7296));
  INVx1_ASAP7_75t_L         g07040(.A(new_n7293), .Y(new_n7297));
  OAI21xp33_ASAP7_75t_L     g07041(.A1(new_n7295), .A2(new_n7296), .B(new_n7297), .Y(new_n7298));
  MAJIxp5_ASAP7_75t_L       g07042(.A(new_n7061), .B(new_n7051), .C(new_n7059), .Y(new_n7299));
  NAND3xp33_ASAP7_75t_L     g07043(.A(new_n7299), .B(new_n7298), .C(new_n7294), .Y(new_n7300));
  NAND2xp33_ASAP7_75t_L     g07044(.A(new_n7294), .B(new_n7298), .Y(new_n7301));
  A2O1A1O1Ixp25_ASAP7_75t_L g07045(.A1(new_n6554), .A2(new_n6559), .B(new_n6552), .C(new_n6800), .D(new_n6792), .Y(new_n7302));
  MAJIxp5_ASAP7_75t_L       g07046(.A(new_n7302), .B(new_n7058), .C(new_n7054), .Y(new_n7303));
  NAND2xp33_ASAP7_75t_L     g07047(.A(new_n7303), .B(new_n7301), .Y(new_n7304));
  AOI22xp33_ASAP7_75t_L     g07048(.A1(new_n344), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n370), .Y(new_n7305));
  OAI221xp5_ASAP7_75t_L     g07049(.A1(new_n429), .A2(new_n6321), .B1(new_n366), .B2(new_n6573), .C(new_n7305), .Y(new_n7306));
  XNOR2x2_ASAP7_75t_L       g07050(.A(\a[5] ), .B(new_n7306), .Y(new_n7307));
  NAND3xp33_ASAP7_75t_L     g07051(.A(new_n7304), .B(new_n7300), .C(new_n7307), .Y(new_n7308));
  INVx1_ASAP7_75t_L         g07052(.A(new_n7308), .Y(new_n7309));
  AOI21xp33_ASAP7_75t_L     g07053(.A1(new_n7304), .A2(new_n7300), .B(new_n7307), .Y(new_n7310));
  OAI21xp33_ASAP7_75t_L     g07054(.A1(new_n7073), .A2(new_n6845), .B(new_n7075), .Y(new_n7311));
  NOR3xp33_ASAP7_75t_L      g07055(.A(new_n7311), .B(new_n7309), .C(new_n7310), .Y(new_n7312));
  INVx1_ASAP7_75t_L         g07056(.A(new_n7310), .Y(new_n7313));
  A2O1A1O1Ixp25_ASAP7_75t_L g07057(.A1(new_n6844), .A2(new_n6584), .B(new_n6808), .C(new_n7076), .D(new_n7072), .Y(new_n7314));
  AOI21xp33_ASAP7_75t_L     g07058(.A1(new_n7313), .A2(new_n7308), .B(new_n7314), .Y(new_n7315));
  NOR2xp33_ASAP7_75t_L      g07059(.A(\b[48] ), .B(\b[49] ), .Y(new_n7316));
  INVx1_ASAP7_75t_L         g07060(.A(\b[49] ), .Y(new_n7317));
  NOR2xp33_ASAP7_75t_L      g07061(.A(new_n6830), .B(new_n7317), .Y(new_n7318));
  NOR2xp33_ASAP7_75t_L      g07062(.A(new_n7316), .B(new_n7318), .Y(new_n7319));
  A2O1A1Ixp33_ASAP7_75t_L   g07063(.A1(\b[48] ), .A2(\b[47] ), .B(new_n6834), .C(new_n7319), .Y(new_n7320));
  O2A1O1Ixp33_ASAP7_75t_L   g07064(.A1(new_n6813), .A2(new_n6816), .B(new_n6832), .C(new_n6831), .Y(new_n7321));
  OAI21xp33_ASAP7_75t_L     g07065(.A1(new_n7316), .A2(new_n7318), .B(new_n7321), .Y(new_n7322));
  NAND2xp33_ASAP7_75t_L     g07066(.A(new_n7320), .B(new_n7322), .Y(new_n7323));
  AOI22xp33_ASAP7_75t_L     g07067(.A1(\b[47] ), .A2(new_n282), .B1(\b[49] ), .B2(new_n303), .Y(new_n7324));
  OAI221xp5_ASAP7_75t_L     g07068(.A1(new_n291), .A2(new_n6830), .B1(new_n268), .B2(new_n7323), .C(new_n7324), .Y(new_n7325));
  XNOR2x2_ASAP7_75t_L       g07069(.A(\a[2] ), .B(new_n7325), .Y(new_n7326));
  OAI21xp33_ASAP7_75t_L     g07070(.A1(new_n7315), .A2(new_n7312), .B(new_n7326), .Y(new_n7327));
  NOR3xp33_ASAP7_75t_L      g07071(.A(new_n7312), .B(new_n7315), .C(new_n7326), .Y(new_n7328));
  INVx1_ASAP7_75t_L         g07072(.A(new_n7328), .Y(new_n7329));
  NAND2xp33_ASAP7_75t_L     g07073(.A(new_n7327), .B(new_n7329), .Y(new_n7330));
  O2A1O1Ixp33_ASAP7_75t_L   g07074(.A1(new_n7086), .A2(new_n7081), .B(new_n7080), .C(new_n7330), .Y(new_n7331));
  AOI211xp5_ASAP7_75t_L     g07075(.A1(new_n7329), .A2(new_n7327), .B(new_n7079), .C(new_n7082), .Y(new_n7332));
  NOR2xp33_ASAP7_75t_L      g07076(.A(new_n7331), .B(new_n7332), .Y(\f[49] ));
  OAI21xp33_ASAP7_75t_L     g07077(.A1(new_n7310), .A2(new_n7309), .B(new_n7311), .Y(new_n7334));
  AOI22xp33_ASAP7_75t_L     g07078(.A1(new_n344), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n370), .Y(new_n7335));
  OAI221xp5_ASAP7_75t_L     g07079(.A1(new_n429), .A2(new_n6568), .B1(new_n366), .B2(new_n6820), .C(new_n7335), .Y(new_n7336));
  XNOR2x2_ASAP7_75t_L       g07080(.A(\a[5] ), .B(new_n7336), .Y(new_n7337));
  NOR2xp33_ASAP7_75t_L      g07081(.A(new_n7295), .B(new_n7296), .Y(new_n7338));
  MAJIxp5_ASAP7_75t_L       g07082(.A(new_n7303), .B(new_n7338), .C(new_n7297), .Y(new_n7339));
  AO21x2_ASAP7_75t_L        g07083(.A1(new_n7246), .A2(new_n7244), .B(new_n7235), .Y(new_n7340));
  NOR2xp33_ASAP7_75t_L      g07084(.A(new_n3180), .B(new_n1373), .Y(new_n7341));
  INVx1_ASAP7_75t_L         g07085(.A(new_n7341), .Y(new_n7342));
  NAND3xp33_ASAP7_75t_L     g07086(.A(new_n3210), .B(new_n1365), .C(new_n3213), .Y(new_n7343));
  AOI22xp33_ASAP7_75t_L     g07087(.A1(new_n1360), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1581), .Y(new_n7344));
  AND4x1_ASAP7_75t_L        g07088(.A(new_n7344), .B(new_n7343), .C(new_n7342), .D(\a[20] ), .Y(new_n7345));
  AOI31xp33_ASAP7_75t_L     g07089(.A1(new_n7343), .A2(new_n7342), .A3(new_n7344), .B(\a[20] ), .Y(new_n7346));
  NOR2xp33_ASAP7_75t_L      g07090(.A(new_n7346), .B(new_n7345), .Y(new_n7347));
  NOR3xp33_ASAP7_75t_L      g07091(.A(new_n7223), .B(new_n7222), .C(new_n7090), .Y(new_n7348));
  O2A1O1Ixp33_ASAP7_75t_L   g07092(.A1(new_n7220), .A2(new_n7224), .B(new_n7238), .C(new_n7348), .Y(new_n7349));
  AOI22xp33_ASAP7_75t_L     g07093(.A1(new_n1704), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1837), .Y(new_n7350));
  OAI221xp5_ASAP7_75t_L     g07094(.A1(new_n1699), .A2(new_n2666), .B1(new_n1827), .B2(new_n2695), .C(new_n7350), .Y(new_n7351));
  XNOR2x2_ASAP7_75t_L       g07095(.A(new_n1689), .B(new_n7351), .Y(new_n7352));
  NAND2xp33_ASAP7_75t_L     g07096(.A(new_n7210), .B(new_n7209), .Y(new_n7353));
  MAJIxp5_ASAP7_75t_L       g07097(.A(new_n7218), .B(new_n7353), .C(new_n7211), .Y(new_n7354));
  AOI22xp33_ASAP7_75t_L     g07098(.A1(new_n2114), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n2259), .Y(new_n7355));
  OAI221xp5_ASAP7_75t_L     g07099(.A1(new_n2109), .A2(new_n2067), .B1(new_n2257), .B2(new_n2355), .C(new_n7355), .Y(new_n7356));
  XNOR2x2_ASAP7_75t_L       g07100(.A(\a[26] ), .B(new_n7356), .Y(new_n7357));
  NAND2xp33_ASAP7_75t_L     g07101(.A(new_n7199), .B(new_n7200), .Y(new_n7358));
  NAND2xp33_ASAP7_75t_L     g07102(.A(new_n7194), .B(new_n7193), .Y(new_n7359));
  NOR2xp33_ASAP7_75t_L      g07103(.A(new_n7190), .B(new_n7359), .Y(new_n7360));
  INVx1_ASAP7_75t_L         g07104(.A(new_n7184), .Y(new_n7361));
  OAI21xp33_ASAP7_75t_L     g07105(.A1(new_n6959), .A2(new_n6961), .B(new_n7361), .Y(new_n7362));
  NOR3xp33_ASAP7_75t_L      g07106(.A(new_n7179), .B(new_n7180), .C(new_n7177), .Y(new_n7363));
  NAND2xp33_ASAP7_75t_L     g07107(.A(new_n7158), .B(new_n7163), .Y(new_n7364));
  MAJIxp5_ASAP7_75t_L       g07108(.A(new_n7172), .B(new_n7166), .C(new_n7364), .Y(new_n7365));
  AOI22xp33_ASAP7_75t_L     g07109(.A1(new_n3633), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n3858), .Y(new_n7366));
  OAI221xp5_ASAP7_75t_L     g07110(.A1(new_n3853), .A2(new_n1030), .B1(new_n3856), .B2(new_n1209), .C(new_n7366), .Y(new_n7367));
  XNOR2x2_ASAP7_75t_L       g07111(.A(new_n3628), .B(new_n7367), .Y(new_n7368));
  AOI21xp33_ASAP7_75t_L     g07112(.A1(new_n7092), .A2(new_n7156), .B(new_n7162), .Y(new_n7369));
  INVx1_ASAP7_75t_L         g07113(.A(new_n7133), .Y(new_n7370));
  NAND3xp33_ASAP7_75t_L     g07114(.A(new_n7370), .B(new_n7130), .C(new_n7124), .Y(new_n7371));
  A2O1A1Ixp33_ASAP7_75t_L   g07115(.A1(new_n7135), .A2(new_n7134), .B(new_n7141), .C(new_n7371), .Y(new_n7372));
  AOI22xp33_ASAP7_75t_L     g07116(.A1(new_n5624), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n5901), .Y(new_n7373));
  OAI221xp5_ASAP7_75t_L     g07117(.A1(new_n5900), .A2(new_n420), .B1(new_n5892), .B2(new_n494), .C(new_n7373), .Y(new_n7374));
  XNOR2x2_ASAP7_75t_L       g07118(.A(\a[44] ), .B(new_n7374), .Y(new_n7375));
  INVx1_ASAP7_75t_L         g07119(.A(new_n7375), .Y(new_n7376));
  NAND2xp33_ASAP7_75t_L     g07120(.A(new_n6876), .B(new_n6879), .Y(new_n7377));
  A2O1A1O1Ixp25_ASAP7_75t_L g07121(.A1(new_n7126), .A2(new_n7377), .B(new_n7096), .C(new_n7119), .D(new_n7129), .Y(new_n7378));
  NAND2xp33_ASAP7_75t_L     g07122(.A(\b[4] ), .B(new_n6380), .Y(new_n7379));
  INVx1_ASAP7_75t_L         g07123(.A(new_n7379), .Y(new_n7380));
  NOR3xp33_ASAP7_75t_L      g07124(.A(new_n357), .B(new_n358), .C(new_n6636), .Y(new_n7381));
  OAI22xp33_ASAP7_75t_L     g07125(.A1(new_n6638), .A2(new_n298), .B1(new_n354), .B2(new_n6880), .Y(new_n7382));
  NOR4xp25_ASAP7_75t_L      g07126(.A(new_n7381), .B(new_n6371), .C(new_n7382), .D(new_n7380), .Y(new_n7383));
  OAI31xp33_ASAP7_75t_L     g07127(.A1(new_n7381), .A2(new_n7380), .A3(new_n7382), .B(new_n6371), .Y(new_n7384));
  INVx1_ASAP7_75t_L         g07128(.A(new_n7384), .Y(new_n7385));
  NOR2xp33_ASAP7_75t_L      g07129(.A(new_n7383), .B(new_n7385), .Y(new_n7386));
  A2O1A1Ixp33_ASAP7_75t_L   g07130(.A1(\b[0] ), .A2(new_n7113), .B(new_n7117), .C(\a[50] ), .Y(new_n7387));
  NAND2xp33_ASAP7_75t_L     g07131(.A(\b[1] ), .B(new_n7115), .Y(new_n7388));
  NAND3xp33_ASAP7_75t_L     g07132(.A(new_n7113), .B(new_n7105), .C(new_n7107), .Y(new_n7389));
  NOR2xp33_ASAP7_75t_L      g07133(.A(new_n276), .B(new_n7389), .Y(new_n7390));
  AND3x1_ASAP7_75t_L        g07134(.A(new_n6874), .B(new_n7114), .C(new_n7110), .Y(new_n7391));
  AOI221xp5_ASAP7_75t_L     g07135(.A1(\b[0] ), .A2(new_n7391), .B1(new_n7108), .B2(new_n281), .C(new_n7390), .Y(new_n7392));
  NAND3xp33_ASAP7_75t_L     g07136(.A(new_n7387), .B(new_n7388), .C(new_n7392), .Y(new_n7393));
  NAND5xp2_ASAP7_75t_L      g07137(.A(\a[50] ), .B(new_n7109), .C(new_n7112), .D(new_n7116), .E(new_n6878), .Y(new_n7394));
  NAND2xp33_ASAP7_75t_L     g07138(.A(new_n7388), .B(new_n7392), .Y(new_n7395));
  NAND3xp33_ASAP7_75t_L     g07139(.A(new_n7395), .B(new_n7394), .C(\a[50] ), .Y(new_n7396));
  NAND3xp33_ASAP7_75t_L     g07140(.A(new_n7386), .B(new_n7393), .C(new_n7396), .Y(new_n7397));
  INVx1_ASAP7_75t_L         g07141(.A(new_n7383), .Y(new_n7398));
  NAND2xp33_ASAP7_75t_L     g07142(.A(new_n7384), .B(new_n7398), .Y(new_n7399));
  NAND2xp33_ASAP7_75t_L     g07143(.A(new_n7396), .B(new_n7393), .Y(new_n7400));
  NAND2xp33_ASAP7_75t_L     g07144(.A(new_n7399), .B(new_n7400), .Y(new_n7401));
  AOI21xp33_ASAP7_75t_L     g07145(.A1(new_n7401), .A2(new_n7397), .B(new_n7378), .Y(new_n7402));
  OAI21xp33_ASAP7_75t_L     g07146(.A1(new_n7128), .A2(new_n7127), .B(new_n7123), .Y(new_n7403));
  NAND2xp33_ASAP7_75t_L     g07147(.A(new_n7397), .B(new_n7401), .Y(new_n7404));
  NOR2xp33_ASAP7_75t_L      g07148(.A(new_n7403), .B(new_n7404), .Y(new_n7405));
  OAI21xp33_ASAP7_75t_L     g07149(.A1(new_n7402), .A2(new_n7405), .B(new_n7376), .Y(new_n7406));
  NAND2xp33_ASAP7_75t_L     g07150(.A(new_n7403), .B(new_n7404), .Y(new_n7407));
  NAND3xp33_ASAP7_75t_L     g07151(.A(new_n7378), .B(new_n7397), .C(new_n7401), .Y(new_n7408));
  NAND3xp33_ASAP7_75t_L     g07152(.A(new_n7407), .B(new_n7408), .C(new_n7375), .Y(new_n7409));
  AND2x2_ASAP7_75t_L        g07153(.A(new_n7409), .B(new_n7406), .Y(new_n7410));
  NAND2xp33_ASAP7_75t_L     g07154(.A(new_n7372), .B(new_n7410), .Y(new_n7411));
  NAND2xp33_ASAP7_75t_L     g07155(.A(new_n7409), .B(new_n7406), .Y(new_n7412));
  NAND3xp33_ASAP7_75t_L     g07156(.A(new_n7148), .B(new_n7412), .C(new_n7371), .Y(new_n7413));
  AOI22xp33_ASAP7_75t_L     g07157(.A1(new_n4920), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n5167), .Y(new_n7414));
  OAI221xp5_ASAP7_75t_L     g07158(.A1(new_n5154), .A2(new_n617), .B1(new_n5158), .B2(new_n685), .C(new_n7414), .Y(new_n7415));
  XNOR2x2_ASAP7_75t_L       g07159(.A(\a[41] ), .B(new_n7415), .Y(new_n7416));
  NAND3xp33_ASAP7_75t_L     g07160(.A(new_n7411), .B(new_n7413), .C(new_n7416), .Y(new_n7417));
  A2O1A1O1Ixp25_ASAP7_75t_L g07161(.A1(new_n7135), .A2(new_n7134), .B(new_n7141), .C(new_n7371), .D(new_n7412), .Y(new_n7418));
  NOR2xp33_ASAP7_75t_L      g07162(.A(new_n7372), .B(new_n7410), .Y(new_n7419));
  INVx1_ASAP7_75t_L         g07163(.A(new_n7416), .Y(new_n7420));
  OAI21xp33_ASAP7_75t_L     g07164(.A1(new_n7418), .A2(new_n7419), .B(new_n7420), .Y(new_n7421));
  NAND2xp33_ASAP7_75t_L     g07165(.A(new_n7150), .B(new_n7152), .Y(new_n7422));
  NAND4xp25_ASAP7_75t_L     g07166(.A(new_n7422), .B(new_n7421), .C(new_n7417), .D(new_n7146), .Y(new_n7423));
  NOR3xp33_ASAP7_75t_L      g07167(.A(new_n7419), .B(new_n7418), .C(new_n7420), .Y(new_n7424));
  AOI21xp33_ASAP7_75t_L     g07168(.A1(new_n7411), .A2(new_n7413), .B(new_n7416), .Y(new_n7425));
  AOI211xp5_ASAP7_75t_L     g07169(.A1(new_n6929), .A2(new_n6918), .B(new_n7154), .C(new_n6917), .Y(new_n7426));
  OAI22xp33_ASAP7_75t_L     g07170(.A1(new_n7426), .A2(new_n7153), .B1(new_n7424), .B2(new_n7425), .Y(new_n7427));
  AOI22xp33_ASAP7_75t_L     g07171(.A1(new_n4283), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n4512), .Y(new_n7428));
  OAI221xp5_ASAP7_75t_L     g07172(.A1(new_n4277), .A2(new_n784), .B1(new_n4499), .B2(new_n875), .C(new_n7428), .Y(new_n7429));
  XNOR2x2_ASAP7_75t_L       g07173(.A(\a[38] ), .B(new_n7429), .Y(new_n7430));
  NAND3xp33_ASAP7_75t_L     g07174(.A(new_n7427), .B(new_n7423), .C(new_n7430), .Y(new_n7431));
  NOR4xp25_ASAP7_75t_L      g07175(.A(new_n7426), .B(new_n7424), .C(new_n7153), .D(new_n7425), .Y(new_n7432));
  AOI22xp33_ASAP7_75t_L     g07176(.A1(new_n7421), .A2(new_n7417), .B1(new_n7146), .B2(new_n7422), .Y(new_n7433));
  INVx1_ASAP7_75t_L         g07177(.A(new_n7430), .Y(new_n7434));
  OAI21xp33_ASAP7_75t_L     g07178(.A1(new_n7433), .A2(new_n7432), .B(new_n7434), .Y(new_n7435));
  AOI21xp33_ASAP7_75t_L     g07179(.A1(new_n7435), .A2(new_n7431), .B(new_n7369), .Y(new_n7436));
  NAND2xp33_ASAP7_75t_L     g07180(.A(new_n6926), .B(new_n7159), .Y(new_n7437));
  A2O1A1Ixp33_ASAP7_75t_L   g07181(.A1(new_n6932), .A2(new_n7437), .B(new_n7161), .C(new_n7157), .Y(new_n7438));
  NAND2xp33_ASAP7_75t_L     g07182(.A(new_n7431), .B(new_n7435), .Y(new_n7439));
  NOR2xp33_ASAP7_75t_L      g07183(.A(new_n7439), .B(new_n7438), .Y(new_n7440));
  OAI21xp33_ASAP7_75t_L     g07184(.A1(new_n7436), .A2(new_n7440), .B(new_n7368), .Y(new_n7441));
  XNOR2x2_ASAP7_75t_L       g07185(.A(\a[35] ), .B(new_n7367), .Y(new_n7442));
  A2O1A1Ixp33_ASAP7_75t_L   g07186(.A1(new_n7156), .A2(new_n7092), .B(new_n7162), .C(new_n7439), .Y(new_n7443));
  NAND3xp33_ASAP7_75t_L     g07187(.A(new_n7369), .B(new_n7431), .C(new_n7435), .Y(new_n7444));
  NAND3xp33_ASAP7_75t_L     g07188(.A(new_n7443), .B(new_n7444), .C(new_n7442), .Y(new_n7445));
  NAND3xp33_ASAP7_75t_L     g07189(.A(new_n7365), .B(new_n7441), .C(new_n7445), .Y(new_n7446));
  AND3x1_ASAP7_75t_L        g07190(.A(new_n7163), .B(new_n7158), .C(new_n7166), .Y(new_n7447));
  AOI21xp33_ASAP7_75t_L     g07191(.A1(new_n7163), .A2(new_n7158), .B(new_n7166), .Y(new_n7448));
  NOR2xp33_ASAP7_75t_L      g07192(.A(new_n7448), .B(new_n7447), .Y(new_n7449));
  OR2x4_ASAP7_75t_L         g07193(.A(new_n7166), .B(new_n7364), .Y(new_n7450));
  AOI21xp33_ASAP7_75t_L     g07194(.A1(new_n7443), .A2(new_n7444), .B(new_n7442), .Y(new_n7451));
  NOR3xp33_ASAP7_75t_L      g07195(.A(new_n7440), .B(new_n7436), .C(new_n7368), .Y(new_n7452));
  OAI221xp5_ASAP7_75t_L     g07196(.A1(new_n7452), .A2(new_n7451), .B1(new_n7172), .B2(new_n7449), .C(new_n7450), .Y(new_n7453));
  OAI22xp33_ASAP7_75t_L     g07197(.A1(new_n3402), .A2(new_n1313), .B1(new_n1539), .B2(new_n3022), .Y(new_n7454));
  AOI221xp5_ASAP7_75t_L     g07198(.A1(new_n3030), .A2(\b[19] ), .B1(new_n3021), .B2(new_n1886), .C(new_n7454), .Y(new_n7455));
  XNOR2x2_ASAP7_75t_L       g07199(.A(new_n3015), .B(new_n7455), .Y(new_n7456));
  AO21x2_ASAP7_75t_L        g07200(.A1(new_n7453), .A2(new_n7446), .B(new_n7456), .Y(new_n7457));
  NAND3xp33_ASAP7_75t_L     g07201(.A(new_n7446), .B(new_n7453), .C(new_n7456), .Y(new_n7458));
  AOI221xp5_ASAP7_75t_L     g07202(.A1(new_n7457), .A2(new_n7458), .B1(new_n7183), .B2(new_n7362), .C(new_n7363), .Y(new_n7459));
  A2O1A1O1Ixp25_ASAP7_75t_L g07203(.A1(new_n6955), .A2(new_n6953), .B(new_n7184), .C(new_n7183), .D(new_n7363), .Y(new_n7460));
  NAND2xp33_ASAP7_75t_L     g07204(.A(new_n7458), .B(new_n7457), .Y(new_n7461));
  NOR2xp33_ASAP7_75t_L      g07205(.A(new_n7461), .B(new_n7460), .Y(new_n7462));
  AOI22xp33_ASAP7_75t_L     g07206(.A1(new_n2552), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n2736), .Y(new_n7463));
  OAI221xp5_ASAP7_75t_L     g07207(.A1(new_n2547), .A2(new_n1774), .B1(new_n2734), .B2(new_n1915), .C(new_n7463), .Y(new_n7464));
  XNOR2x2_ASAP7_75t_L       g07208(.A(\a[29] ), .B(new_n7464), .Y(new_n7465));
  OAI21xp33_ASAP7_75t_L     g07209(.A1(new_n7459), .A2(new_n7462), .B(new_n7465), .Y(new_n7466));
  NAND2xp33_ASAP7_75t_L     g07210(.A(new_n7461), .B(new_n7460), .Y(new_n7467));
  INVx1_ASAP7_75t_L         g07211(.A(new_n7363), .Y(new_n7468));
  A2O1A1Ixp33_ASAP7_75t_L   g07212(.A1(new_n7182), .A2(new_n7178), .B(new_n7186), .C(new_n7468), .Y(new_n7469));
  NAND3xp33_ASAP7_75t_L     g07213(.A(new_n7469), .B(new_n7457), .C(new_n7458), .Y(new_n7470));
  INVx1_ASAP7_75t_L         g07214(.A(new_n7465), .Y(new_n7471));
  NAND3xp33_ASAP7_75t_L     g07215(.A(new_n7470), .B(new_n7467), .C(new_n7471), .Y(new_n7472));
  AOI221xp5_ASAP7_75t_L     g07216(.A1(new_n7358), .A2(new_n7197), .B1(new_n7466), .B2(new_n7472), .C(new_n7360), .Y(new_n7473));
  NOR2xp33_ASAP7_75t_L      g07217(.A(new_n7187), .B(new_n7185), .Y(new_n7474));
  MAJIxp5_ASAP7_75t_L       g07218(.A(new_n7197), .B(new_n7191), .C(new_n7474), .Y(new_n7475));
  AOI21xp33_ASAP7_75t_L     g07219(.A1(new_n7470), .A2(new_n7467), .B(new_n7471), .Y(new_n7476));
  NOR3xp33_ASAP7_75t_L      g07220(.A(new_n7462), .B(new_n7465), .C(new_n7459), .Y(new_n7477));
  NOR3xp33_ASAP7_75t_L      g07221(.A(new_n7475), .B(new_n7476), .C(new_n7477), .Y(new_n7478));
  OAI21xp33_ASAP7_75t_L     g07222(.A1(new_n7473), .A2(new_n7478), .B(new_n7357), .Y(new_n7479));
  INVx1_ASAP7_75t_L         g07223(.A(new_n7357), .Y(new_n7480));
  OAI21xp33_ASAP7_75t_L     g07224(.A1(new_n7476), .A2(new_n7477), .B(new_n7475), .Y(new_n7481));
  MAJIxp5_ASAP7_75t_L       g07225(.A(new_n7202), .B(new_n7359), .C(new_n7190), .Y(new_n7482));
  NAND3xp33_ASAP7_75t_L     g07226(.A(new_n7482), .B(new_n7466), .C(new_n7472), .Y(new_n7483));
  NAND3xp33_ASAP7_75t_L     g07227(.A(new_n7483), .B(new_n7481), .C(new_n7480), .Y(new_n7484));
  NAND3xp33_ASAP7_75t_L     g07228(.A(new_n7354), .B(new_n7479), .C(new_n7484), .Y(new_n7485));
  NOR2xp33_ASAP7_75t_L      g07229(.A(new_n7212), .B(new_n7207), .Y(new_n7486));
  NOR2xp33_ASAP7_75t_L      g07230(.A(new_n7211), .B(new_n7353), .Y(new_n7487));
  INVx1_ASAP7_75t_L         g07231(.A(new_n7487), .Y(new_n7488));
  AOI21xp33_ASAP7_75t_L     g07232(.A1(new_n7483), .A2(new_n7481), .B(new_n7480), .Y(new_n7489));
  NOR3xp33_ASAP7_75t_L      g07233(.A(new_n7478), .B(new_n7473), .C(new_n7357), .Y(new_n7490));
  OAI221xp5_ASAP7_75t_L     g07234(.A1(new_n7486), .A2(new_n7218), .B1(new_n7490), .B2(new_n7489), .C(new_n7488), .Y(new_n7491));
  AO21x2_ASAP7_75t_L        g07235(.A1(new_n7491), .A2(new_n7485), .B(new_n7352), .Y(new_n7492));
  NAND3xp33_ASAP7_75t_L     g07236(.A(new_n7485), .B(new_n7491), .C(new_n7352), .Y(new_n7493));
  NAND2xp33_ASAP7_75t_L     g07237(.A(new_n7493), .B(new_n7492), .Y(new_n7494));
  NOR2xp33_ASAP7_75t_L      g07238(.A(new_n7349), .B(new_n7494), .Y(new_n7495));
  AOI221xp5_ASAP7_75t_L     g07239(.A1(new_n7238), .A2(new_n7230), .B1(new_n7493), .B2(new_n7492), .C(new_n7348), .Y(new_n7496));
  OAI21xp33_ASAP7_75t_L     g07240(.A1(new_n7496), .A2(new_n7495), .B(new_n7347), .Y(new_n7497));
  INVx1_ASAP7_75t_L         g07241(.A(new_n7347), .Y(new_n7498));
  INVx1_ASAP7_75t_L         g07242(.A(new_n7348), .Y(new_n7499));
  A2O1A1Ixp33_ASAP7_75t_L   g07243(.A1(new_n7228), .A2(new_n7229), .B(new_n7227), .C(new_n7499), .Y(new_n7500));
  NAND3xp33_ASAP7_75t_L     g07244(.A(new_n7500), .B(new_n7492), .C(new_n7493), .Y(new_n7501));
  INVx1_ASAP7_75t_L         g07245(.A(new_n7496), .Y(new_n7502));
  NAND3xp33_ASAP7_75t_L     g07246(.A(new_n7502), .B(new_n7501), .C(new_n7498), .Y(new_n7503));
  NAND3xp33_ASAP7_75t_L     g07247(.A(new_n7340), .B(new_n7497), .C(new_n7503), .Y(new_n7504));
  INVx1_ASAP7_75t_L         g07248(.A(new_n7006), .Y(new_n7505));
  A2O1A1O1Ixp25_ASAP7_75t_L g07249(.A1(new_n7011), .A2(new_n6853), .B(new_n7505), .C(new_n7246), .D(new_n7235), .Y(new_n7506));
  AOI21xp33_ASAP7_75t_L     g07250(.A1(new_n7502), .A2(new_n7501), .B(new_n7498), .Y(new_n7507));
  NOR3xp33_ASAP7_75t_L      g07251(.A(new_n7495), .B(new_n7496), .C(new_n7347), .Y(new_n7508));
  OAI21xp33_ASAP7_75t_L     g07252(.A1(new_n7508), .A2(new_n7507), .B(new_n7506), .Y(new_n7509));
  NOR2xp33_ASAP7_75t_L      g07253(.A(new_n3584), .B(new_n1154), .Y(new_n7510));
  INVx1_ASAP7_75t_L         g07254(.A(new_n7510), .Y(new_n7511));
  NAND2xp33_ASAP7_75t_L     g07255(.A(new_n1073), .B(new_n3811), .Y(new_n7512));
  AOI22xp33_ASAP7_75t_L     g07256(.A1(new_n1076), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1253), .Y(new_n7513));
  AND4x1_ASAP7_75t_L        g07257(.A(new_n7513), .B(new_n7512), .C(new_n7511), .D(\a[17] ), .Y(new_n7514));
  AOI31xp33_ASAP7_75t_L     g07258(.A1(new_n7512), .A2(new_n7511), .A3(new_n7513), .B(\a[17] ), .Y(new_n7515));
  NOR2xp33_ASAP7_75t_L      g07259(.A(new_n7515), .B(new_n7514), .Y(new_n7516));
  NAND3xp33_ASAP7_75t_L     g07260(.A(new_n7504), .B(new_n7516), .C(new_n7509), .Y(new_n7517));
  NOR3xp33_ASAP7_75t_L      g07261(.A(new_n7506), .B(new_n7507), .C(new_n7508), .Y(new_n7518));
  AOI21xp33_ASAP7_75t_L     g07262(.A1(new_n7503), .A2(new_n7497), .B(new_n7340), .Y(new_n7519));
  OAI22xp33_ASAP7_75t_L     g07263(.A1(new_n7519), .A2(new_n7518), .B1(new_n7515), .B2(new_n7514), .Y(new_n7520));
  AND2x2_ASAP7_75t_L        g07264(.A(new_n7517), .B(new_n7520), .Y(new_n7521));
  INVx1_ASAP7_75t_L         g07265(.A(new_n7253), .Y(new_n7522));
  NAND3xp33_ASAP7_75t_L     g07266(.A(new_n7247), .B(new_n7242), .C(new_n7522), .Y(new_n7523));
  INVx1_ASAP7_75t_L         g07267(.A(new_n7523), .Y(new_n7524));
  O2A1O1Ixp33_ASAP7_75t_L   g07268(.A1(new_n7254), .A2(new_n7255), .B(new_n7262), .C(new_n7524), .Y(new_n7525));
  NAND2xp33_ASAP7_75t_L     g07269(.A(new_n7525), .B(new_n7521), .Y(new_n7526));
  NAND2xp33_ASAP7_75t_L     g07270(.A(new_n7517), .B(new_n7520), .Y(new_n7527));
  OAI21xp33_ASAP7_75t_L     g07271(.A1(new_n7256), .A2(new_n7259), .B(new_n7523), .Y(new_n7528));
  NAND2xp33_ASAP7_75t_L     g07272(.A(new_n7527), .B(new_n7528), .Y(new_n7529));
  OAI22xp33_ASAP7_75t_L     g07273(.A1(new_n978), .A2(new_n4216), .B1(new_n4632), .B2(new_n977), .Y(new_n7530));
  AOI221xp5_ASAP7_75t_L     g07274(.A1(\b[37] ), .A2(new_n815), .B1(new_n808), .B2(new_n4640), .C(new_n7530), .Y(new_n7531));
  XNOR2x2_ASAP7_75t_L       g07275(.A(new_n806), .B(new_n7531), .Y(new_n7532));
  NAND3xp33_ASAP7_75t_L     g07276(.A(new_n7526), .B(new_n7532), .C(new_n7529), .Y(new_n7533));
  NOR2xp33_ASAP7_75t_L      g07277(.A(new_n7527), .B(new_n7528), .Y(new_n7534));
  AOI21xp33_ASAP7_75t_L     g07278(.A1(new_n7520), .A2(new_n7517), .B(new_n7525), .Y(new_n7535));
  INVx1_ASAP7_75t_L         g07279(.A(new_n7532), .Y(new_n7536));
  OAI21xp33_ASAP7_75t_L     g07280(.A1(new_n7535), .A2(new_n7534), .B(new_n7536), .Y(new_n7537));
  INVx1_ASAP7_75t_L         g07281(.A(new_n7266), .Y(new_n7538));
  NAND3xp33_ASAP7_75t_L     g07282(.A(new_n7260), .B(new_n7263), .C(new_n7538), .Y(new_n7539));
  NAND4xp25_ASAP7_75t_L     g07283(.A(new_n7271), .B(new_n7539), .C(new_n7537), .D(new_n7533), .Y(new_n7540));
  NOR3xp33_ASAP7_75t_L      g07284(.A(new_n7534), .B(new_n7535), .C(new_n7536), .Y(new_n7541));
  AOI21xp33_ASAP7_75t_L     g07285(.A1(new_n7526), .A2(new_n7529), .B(new_n7532), .Y(new_n7542));
  NAND2xp33_ASAP7_75t_L     g07286(.A(new_n7263), .B(new_n7260), .Y(new_n7543));
  MAJIxp5_ASAP7_75t_L       g07287(.A(new_n7269), .B(new_n7543), .C(new_n7266), .Y(new_n7544));
  OAI21xp33_ASAP7_75t_L     g07288(.A1(new_n7541), .A2(new_n7542), .B(new_n7544), .Y(new_n7545));
  NAND2xp33_ASAP7_75t_L     g07289(.A(\b[40] ), .B(new_n584), .Y(new_n7546));
  NAND3xp33_ASAP7_75t_L     g07290(.A(new_n5326), .B(new_n5324), .C(new_n578), .Y(new_n7547));
  AOI22xp33_ASAP7_75t_L     g07291(.A1(\b[39] ), .A2(new_n651), .B1(\b[41] ), .B2(new_n581), .Y(new_n7548));
  AND4x1_ASAP7_75t_L        g07292(.A(new_n7548), .B(new_n7547), .C(new_n7546), .D(\a[11] ), .Y(new_n7549));
  AOI31xp33_ASAP7_75t_L     g07293(.A1(new_n7547), .A2(new_n7546), .A3(new_n7548), .B(\a[11] ), .Y(new_n7550));
  NOR2xp33_ASAP7_75t_L      g07294(.A(new_n7550), .B(new_n7549), .Y(new_n7551));
  NAND3xp33_ASAP7_75t_L     g07295(.A(new_n7540), .B(new_n7545), .C(new_n7551), .Y(new_n7552));
  NOR3xp33_ASAP7_75t_L      g07296(.A(new_n7544), .B(new_n7542), .C(new_n7541), .Y(new_n7553));
  OA21x2_ASAP7_75t_L        g07297(.A1(new_n7541), .A2(new_n7542), .B(new_n7544), .Y(new_n7554));
  INVx1_ASAP7_75t_L         g07298(.A(new_n7551), .Y(new_n7555));
  OAI21xp33_ASAP7_75t_L     g07299(.A1(new_n7553), .A2(new_n7554), .B(new_n7555), .Y(new_n7556));
  NAND2xp33_ASAP7_75t_L     g07300(.A(new_n7552), .B(new_n7556), .Y(new_n7557));
  AOI211xp5_ASAP7_75t_L     g07301(.A1(new_n7276), .A2(new_n7277), .B(new_n7280), .C(new_n7279), .Y(new_n7558));
  AO21x2_ASAP7_75t_L        g07302(.A1(new_n7286), .A2(new_n7285), .B(new_n7558), .Y(new_n7559));
  NOR2xp33_ASAP7_75t_L      g07303(.A(new_n7557), .B(new_n7559), .Y(new_n7560));
  AND2x2_ASAP7_75t_L        g07304(.A(new_n7552), .B(new_n7556), .Y(new_n7561));
  NOR2xp33_ASAP7_75t_L      g07305(.A(new_n7280), .B(new_n7279), .Y(new_n7562));
  MAJIxp5_ASAP7_75t_L       g07306(.A(new_n7286), .B(new_n7562), .C(new_n7281), .Y(new_n7563));
  NOR2xp33_ASAP7_75t_L      g07307(.A(new_n7563), .B(new_n7561), .Y(new_n7564));
  AOI22xp33_ASAP7_75t_L     g07308(.A1(new_n444), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n471), .Y(new_n7565));
  OAI221xp5_ASAP7_75t_L     g07309(.A1(new_n468), .A2(new_n5805), .B1(new_n469), .B2(new_n5835), .C(new_n7565), .Y(new_n7566));
  XNOR2x2_ASAP7_75t_L       g07310(.A(\a[8] ), .B(new_n7566), .Y(new_n7567));
  NOR3xp33_ASAP7_75t_L      g07311(.A(new_n7564), .B(new_n7560), .C(new_n7567), .Y(new_n7568));
  NAND2xp33_ASAP7_75t_L     g07312(.A(new_n7563), .B(new_n7561), .Y(new_n7569));
  A2O1A1Ixp33_ASAP7_75t_L   g07313(.A1(new_n7285), .A2(new_n7286), .B(new_n7558), .C(new_n7557), .Y(new_n7570));
  INVx1_ASAP7_75t_L         g07314(.A(new_n7567), .Y(new_n7571));
  AOI21xp33_ASAP7_75t_L     g07315(.A1(new_n7569), .A2(new_n7570), .B(new_n7571), .Y(new_n7572));
  OAI21xp33_ASAP7_75t_L     g07316(.A1(new_n7568), .A2(new_n7572), .B(new_n7339), .Y(new_n7573));
  NAND2xp33_ASAP7_75t_L     g07317(.A(new_n7287), .B(new_n7284), .Y(new_n7574));
  MAJIxp5_ASAP7_75t_L       g07318(.A(new_n7299), .B(new_n7574), .C(new_n7293), .Y(new_n7575));
  NAND3xp33_ASAP7_75t_L     g07319(.A(new_n7569), .B(new_n7570), .C(new_n7571), .Y(new_n7576));
  OAI21xp33_ASAP7_75t_L     g07320(.A1(new_n7560), .A2(new_n7564), .B(new_n7567), .Y(new_n7577));
  NAND3xp33_ASAP7_75t_L     g07321(.A(new_n7575), .B(new_n7576), .C(new_n7577), .Y(new_n7578));
  NAND3xp33_ASAP7_75t_L     g07322(.A(new_n7578), .B(new_n7573), .C(new_n7337), .Y(new_n7579));
  INVx1_ASAP7_75t_L         g07323(.A(new_n7337), .Y(new_n7580));
  AOI21xp33_ASAP7_75t_L     g07324(.A1(new_n7577), .A2(new_n7576), .B(new_n7575), .Y(new_n7581));
  NOR3xp33_ASAP7_75t_L      g07325(.A(new_n7339), .B(new_n7568), .C(new_n7572), .Y(new_n7582));
  OAI21xp33_ASAP7_75t_L     g07326(.A1(new_n7581), .A2(new_n7582), .B(new_n7580), .Y(new_n7583));
  NAND2xp33_ASAP7_75t_L     g07327(.A(new_n7300), .B(new_n7304), .Y(new_n7584));
  NOR2xp33_ASAP7_75t_L      g07328(.A(new_n7307), .B(new_n7584), .Y(new_n7585));
  INVx1_ASAP7_75t_L         g07329(.A(new_n7585), .Y(new_n7586));
  NAND4xp25_ASAP7_75t_L     g07330(.A(new_n7334), .B(new_n7586), .C(new_n7583), .D(new_n7579), .Y(new_n7587));
  NAND2xp33_ASAP7_75t_L     g07331(.A(new_n7579), .B(new_n7583), .Y(new_n7588));
  MAJIxp5_ASAP7_75t_L       g07332(.A(new_n7314), .B(new_n7307), .C(new_n7584), .Y(new_n7589));
  NAND2xp33_ASAP7_75t_L     g07333(.A(new_n7589), .B(new_n7588), .Y(new_n7590));
  NAND2xp33_ASAP7_75t_L     g07334(.A(new_n7590), .B(new_n7587), .Y(new_n7591));
  NOR2xp33_ASAP7_75t_L      g07335(.A(\b[49] ), .B(\b[50] ), .Y(new_n7592));
  INVx1_ASAP7_75t_L         g07336(.A(\b[50] ), .Y(new_n7593));
  NOR2xp33_ASAP7_75t_L      g07337(.A(new_n7317), .B(new_n7593), .Y(new_n7594));
  NOR2xp33_ASAP7_75t_L      g07338(.A(new_n7592), .B(new_n7594), .Y(new_n7595));
  INVx1_ASAP7_75t_L         g07339(.A(new_n7595), .Y(new_n7596));
  O2A1O1Ixp33_ASAP7_75t_L   g07340(.A1(new_n6830), .A2(new_n7317), .B(new_n7320), .C(new_n7596), .Y(new_n7597));
  O2A1O1Ixp33_ASAP7_75t_L   g07341(.A1(new_n6831), .A2(new_n6834), .B(new_n7319), .C(new_n7318), .Y(new_n7598));
  NAND2xp33_ASAP7_75t_L     g07342(.A(new_n7596), .B(new_n7598), .Y(new_n7599));
  INVx1_ASAP7_75t_L         g07343(.A(new_n7599), .Y(new_n7600));
  NOR2xp33_ASAP7_75t_L      g07344(.A(new_n7597), .B(new_n7600), .Y(new_n7601));
  INVx1_ASAP7_75t_L         g07345(.A(new_n7601), .Y(new_n7602));
  AOI22xp33_ASAP7_75t_L     g07346(.A1(\b[48] ), .A2(new_n282), .B1(\b[50] ), .B2(new_n303), .Y(new_n7603));
  OAI221xp5_ASAP7_75t_L     g07347(.A1(new_n291), .A2(new_n7317), .B1(new_n268), .B2(new_n7602), .C(new_n7603), .Y(new_n7604));
  XNOR2x2_ASAP7_75t_L       g07348(.A(\a[2] ), .B(new_n7604), .Y(new_n7605));
  INVx1_ASAP7_75t_L         g07349(.A(new_n7605), .Y(new_n7606));
  XNOR2x2_ASAP7_75t_L       g07350(.A(new_n7606), .B(new_n7591), .Y(new_n7607));
  A2O1A1O1Ixp25_ASAP7_75t_L g07351(.A1(new_n7078), .A2(new_n7083), .B(new_n7079), .C(new_n7327), .D(new_n7328), .Y(new_n7608));
  INVx1_ASAP7_75t_L         g07352(.A(new_n7608), .Y(new_n7609));
  AND2x2_ASAP7_75t_L        g07353(.A(new_n7609), .B(new_n7607), .Y(new_n7610));
  NOR2xp33_ASAP7_75t_L      g07354(.A(new_n7609), .B(new_n7607), .Y(new_n7611));
  NOR2xp33_ASAP7_75t_L      g07355(.A(new_n7611), .B(new_n7610), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g07356(.A(new_n7608), .B(new_n7591), .C(new_n7605), .Y(new_n7613));
  INVx1_ASAP7_75t_L         g07357(.A(new_n7594), .Y(new_n7614));
  NOR2xp33_ASAP7_75t_L      g07358(.A(\b[50] ), .B(\b[51] ), .Y(new_n7615));
  INVx1_ASAP7_75t_L         g07359(.A(\b[51] ), .Y(new_n7616));
  NOR2xp33_ASAP7_75t_L      g07360(.A(new_n7593), .B(new_n7616), .Y(new_n7617));
  NOR2xp33_ASAP7_75t_L      g07361(.A(new_n7615), .B(new_n7617), .Y(new_n7618));
  INVx1_ASAP7_75t_L         g07362(.A(new_n7618), .Y(new_n7619));
  O2A1O1Ixp33_ASAP7_75t_L   g07363(.A1(new_n7596), .A2(new_n7598), .B(new_n7614), .C(new_n7619), .Y(new_n7620));
  NOR3xp33_ASAP7_75t_L      g07364(.A(new_n7597), .B(new_n7618), .C(new_n7594), .Y(new_n7621));
  NOR2xp33_ASAP7_75t_L      g07365(.A(new_n7620), .B(new_n7621), .Y(new_n7622));
  INVx1_ASAP7_75t_L         g07366(.A(new_n7622), .Y(new_n7623));
  AOI22xp33_ASAP7_75t_L     g07367(.A1(\b[49] ), .A2(new_n282), .B1(\b[51] ), .B2(new_n303), .Y(new_n7624));
  OAI221xp5_ASAP7_75t_L     g07368(.A1(new_n291), .A2(new_n7593), .B1(new_n268), .B2(new_n7623), .C(new_n7624), .Y(new_n7625));
  XNOR2x2_ASAP7_75t_L       g07369(.A(\a[2] ), .B(new_n7625), .Y(new_n7626));
  NOR3xp33_ASAP7_75t_L      g07370(.A(new_n7582), .B(new_n7581), .C(new_n7337), .Y(new_n7627));
  O2A1O1Ixp33_ASAP7_75t_L   g07371(.A1(new_n7585), .A2(new_n7315), .B(new_n7588), .C(new_n7627), .Y(new_n7628));
  NAND2xp33_ASAP7_75t_L     g07372(.A(\b[47] ), .B(new_n347), .Y(new_n7629));
  INVx1_ASAP7_75t_L         g07373(.A(new_n6837), .Y(new_n7630));
  NAND2xp33_ASAP7_75t_L     g07374(.A(new_n341), .B(new_n7630), .Y(new_n7631));
  AOI22xp33_ASAP7_75t_L     g07375(.A1(new_n344), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n370), .Y(new_n7632));
  AND4x1_ASAP7_75t_L        g07376(.A(new_n7632), .B(new_n7631), .C(new_n7629), .D(\a[5] ), .Y(new_n7633));
  AOI31xp33_ASAP7_75t_L     g07377(.A1(new_n7631), .A2(new_n7629), .A3(new_n7632), .B(\a[5] ), .Y(new_n7634));
  NOR2xp33_ASAP7_75t_L      g07378(.A(new_n7634), .B(new_n7633), .Y(new_n7635));
  O2A1O1Ixp33_ASAP7_75t_L   g07379(.A1(new_n7261), .A2(new_n7018), .B(new_n7024), .C(new_n7256), .Y(new_n7636));
  NOR3xp33_ASAP7_75t_L      g07380(.A(new_n7519), .B(new_n7518), .C(new_n7516), .Y(new_n7637));
  O2A1O1Ixp33_ASAP7_75t_L   g07381(.A1(new_n7524), .A2(new_n7636), .B(new_n7527), .C(new_n7637), .Y(new_n7638));
  OAI22xp33_ASAP7_75t_L     g07382(.A1(new_n1158), .A2(new_n3584), .B1(new_n4216), .B2(new_n1259), .Y(new_n7639));
  AOI221xp5_ASAP7_75t_L     g07383(.A1(\b[35] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n6848), .C(new_n7639), .Y(new_n7640));
  XNOR2x2_ASAP7_75t_L       g07384(.A(new_n1071), .B(new_n7640), .Y(new_n7641));
  INVx1_ASAP7_75t_L         g07385(.A(new_n7641), .Y(new_n7642));
  OAI21xp33_ASAP7_75t_L     g07386(.A1(new_n7507), .A2(new_n7506), .B(new_n7503), .Y(new_n7643));
  AND3x1_ASAP7_75t_L        g07387(.A(new_n7485), .B(new_n7491), .C(new_n7352), .Y(new_n7644));
  A2O1A1O1Ixp25_ASAP7_75t_L g07388(.A1(new_n7230), .A2(new_n7238), .B(new_n7348), .C(new_n7492), .D(new_n7644), .Y(new_n7645));
  AOI22xp33_ASAP7_75t_L     g07389(.A1(new_n1704), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1837), .Y(new_n7646));
  OAI221xp5_ASAP7_75t_L     g07390(.A1(new_n1699), .A2(new_n2688), .B1(new_n1827), .B2(new_n2990), .C(new_n7646), .Y(new_n7647));
  XNOR2x2_ASAP7_75t_L       g07391(.A(\a[23] ), .B(new_n7647), .Y(new_n7648));
  NAND2xp33_ASAP7_75t_L     g07392(.A(new_n7216), .B(new_n7217), .Y(new_n7649));
  A2O1A1O1Ixp25_ASAP7_75t_L g07393(.A1(new_n7214), .A2(new_n7649), .B(new_n7487), .C(new_n7479), .D(new_n7490), .Y(new_n7650));
  NAND2xp33_ASAP7_75t_L     g07394(.A(new_n7445), .B(new_n7441), .Y(new_n7651));
  NOR3xp33_ASAP7_75t_L      g07395(.A(new_n7440), .B(new_n7436), .C(new_n7442), .Y(new_n7652));
  AOI22xp33_ASAP7_75t_L     g07396(.A1(new_n3633), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n3858), .Y(new_n7653));
  OAI221xp5_ASAP7_75t_L     g07397(.A1(new_n3853), .A2(new_n1201), .B1(new_n3856), .B2(new_n1320), .C(new_n7653), .Y(new_n7654));
  XNOR2x2_ASAP7_75t_L       g07398(.A(\a[35] ), .B(new_n7654), .Y(new_n7655));
  NAND2xp33_ASAP7_75t_L     g07399(.A(new_n7423), .B(new_n7427), .Y(new_n7656));
  AOI22xp33_ASAP7_75t_L     g07400(.A1(new_n4283), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n4512), .Y(new_n7657));
  OAI221xp5_ASAP7_75t_L     g07401(.A1(new_n4277), .A2(new_n869), .B1(new_n4499), .B2(new_n950), .C(new_n7657), .Y(new_n7658));
  XNOR2x2_ASAP7_75t_L       g07402(.A(\a[38] ), .B(new_n7658), .Y(new_n7659));
  INVx1_ASAP7_75t_L         g07403(.A(new_n7659), .Y(new_n7660));
  OAI31xp33_ASAP7_75t_L     g07404(.A1(new_n7426), .A2(new_n7424), .A3(new_n7153), .B(new_n7421), .Y(new_n7661));
  AOI22xp33_ASAP7_75t_L     g07405(.A1(new_n4920), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n5167), .Y(new_n7662));
  OAI221xp5_ASAP7_75t_L     g07406(.A1(new_n5154), .A2(new_n679), .B1(new_n5158), .B2(new_n768), .C(new_n7662), .Y(new_n7663));
  XNOR2x2_ASAP7_75t_L       g07407(.A(\a[41] ), .B(new_n7663), .Y(new_n7664));
  NOR3xp33_ASAP7_75t_L      g07408(.A(new_n7405), .B(new_n7402), .C(new_n7375), .Y(new_n7665));
  INVx1_ASAP7_75t_L         g07409(.A(\a[51] ), .Y(new_n7666));
  NAND2xp33_ASAP7_75t_L     g07410(.A(\a[50] ), .B(new_n7666), .Y(new_n7667));
  NAND2xp33_ASAP7_75t_L     g07411(.A(\a[51] ), .B(new_n7106), .Y(new_n7668));
  AND2x2_ASAP7_75t_L        g07412(.A(new_n7667), .B(new_n7668), .Y(new_n7669));
  NOR2xp33_ASAP7_75t_L      g07413(.A(new_n258), .B(new_n7669), .Y(new_n7670));
  OAI21xp33_ASAP7_75t_L     g07414(.A1(new_n7394), .A2(new_n7395), .B(new_n7670), .Y(new_n7671));
  NOR2xp33_ASAP7_75t_L      g07415(.A(new_n7106), .B(new_n6875), .Y(new_n7672));
  AND4x1_ASAP7_75t_L        g07416(.A(new_n7109), .B(new_n7672), .C(new_n7112), .D(new_n7116), .Y(new_n7673));
  INVx1_ASAP7_75t_L         g07417(.A(new_n7670), .Y(new_n7674));
  NAND4xp25_ASAP7_75t_L     g07418(.A(new_n7673), .B(new_n7674), .C(new_n7392), .D(new_n7388), .Y(new_n7675));
  NAND3xp33_ASAP7_75t_L     g07419(.A(new_n6874), .B(new_n7110), .C(new_n7114), .Y(new_n7676));
  OAI22xp33_ASAP7_75t_L     g07420(.A1(new_n7676), .A2(new_n261), .B1(new_n298), .B2(new_n7389), .Y(new_n7677));
  AOI221xp5_ASAP7_75t_L     g07421(.A1(\b[2] ), .A2(new_n7115), .B1(new_n406), .B2(new_n7108), .C(new_n7677), .Y(new_n7678));
  NAND2xp33_ASAP7_75t_L     g07422(.A(\a[50] ), .B(new_n7678), .Y(new_n7679));
  AO21x2_ASAP7_75t_L        g07423(.A1(new_n406), .A2(new_n7108), .B(new_n7677), .Y(new_n7680));
  A2O1A1Ixp33_ASAP7_75t_L   g07424(.A1(\b[2] ), .A2(new_n7115), .B(new_n7680), .C(new_n7106), .Y(new_n7681));
  AO22x1_ASAP7_75t_L        g07425(.A1(new_n7681), .A2(new_n7679), .B1(new_n7675), .B2(new_n7671), .Y(new_n7682));
  NAND4xp25_ASAP7_75t_L     g07426(.A(new_n7671), .B(new_n7681), .C(new_n7679), .D(new_n7675), .Y(new_n7683));
  NOR2xp33_ASAP7_75t_L      g07427(.A(new_n354), .B(new_n6646), .Y(new_n7684));
  INVx1_ASAP7_75t_L         g07428(.A(new_n7684), .Y(new_n7685));
  NAND2xp33_ASAP7_75t_L     g07429(.A(new_n6373), .B(new_n526), .Y(new_n7686));
  AOI22xp33_ASAP7_75t_L     g07430(.A1(new_n6376), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n6648), .Y(new_n7687));
  NAND4xp25_ASAP7_75t_L     g07431(.A(new_n7686), .B(\a[47] ), .C(new_n7685), .D(new_n7687), .Y(new_n7688));
  AOI31xp33_ASAP7_75t_L     g07432(.A1(new_n7686), .A2(new_n7685), .A3(new_n7687), .B(\a[47] ), .Y(new_n7689));
  INVx1_ASAP7_75t_L         g07433(.A(new_n7689), .Y(new_n7690));
  NAND4xp25_ASAP7_75t_L     g07434(.A(new_n7682), .B(new_n7690), .C(new_n7688), .D(new_n7683), .Y(new_n7691));
  AOI22xp33_ASAP7_75t_L     g07435(.A1(new_n7679), .A2(new_n7681), .B1(new_n7675), .B2(new_n7671), .Y(new_n7692));
  AND4x1_ASAP7_75t_L        g07436(.A(new_n7671), .B(new_n7681), .C(new_n7675), .D(new_n7679), .Y(new_n7693));
  INVx1_ASAP7_75t_L         g07437(.A(new_n7688), .Y(new_n7694));
  OAI22xp33_ASAP7_75t_L     g07438(.A1(new_n7693), .A2(new_n7692), .B1(new_n7689), .B2(new_n7694), .Y(new_n7695));
  AND2x2_ASAP7_75t_L        g07439(.A(new_n7691), .B(new_n7695), .Y(new_n7696));
  INVx1_ASAP7_75t_L         g07440(.A(new_n7400), .Y(new_n7697));
  MAJIxp5_ASAP7_75t_L       g07441(.A(new_n7403), .B(new_n7399), .C(new_n7697), .Y(new_n7698));
  NAND2xp33_ASAP7_75t_L     g07442(.A(new_n7698), .B(new_n7696), .Y(new_n7699));
  NAND2xp33_ASAP7_75t_L     g07443(.A(new_n7691), .B(new_n7695), .Y(new_n7700));
  NOR2xp33_ASAP7_75t_L      g07444(.A(new_n7386), .B(new_n7400), .Y(new_n7701));
  A2O1A1Ixp33_ASAP7_75t_L   g07445(.A1(new_n7403), .A2(new_n7404), .B(new_n7701), .C(new_n7700), .Y(new_n7702));
  AOI22xp33_ASAP7_75t_L     g07446(.A1(new_n5624), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n5901), .Y(new_n7703));
  OAI221xp5_ASAP7_75t_L     g07447(.A1(new_n5900), .A2(new_n488), .B1(new_n5892), .B2(new_n548), .C(new_n7703), .Y(new_n7704));
  XNOR2x2_ASAP7_75t_L       g07448(.A(new_n5619), .B(new_n7704), .Y(new_n7705));
  AOI21xp33_ASAP7_75t_L     g07449(.A1(new_n7699), .A2(new_n7702), .B(new_n7705), .Y(new_n7706));
  INVx1_ASAP7_75t_L         g07450(.A(new_n7701), .Y(new_n7707));
  A2O1A1Ixp33_ASAP7_75t_L   g07451(.A1(new_n7397), .A2(new_n7401), .B(new_n7378), .C(new_n7707), .Y(new_n7708));
  NOR2xp33_ASAP7_75t_L      g07452(.A(new_n7700), .B(new_n7708), .Y(new_n7709));
  O2A1O1Ixp33_ASAP7_75t_L   g07453(.A1(new_n7386), .A2(new_n7400), .B(new_n7407), .C(new_n7696), .Y(new_n7710));
  XNOR2x2_ASAP7_75t_L       g07454(.A(\a[44] ), .B(new_n7704), .Y(new_n7711));
  NOR3xp33_ASAP7_75t_L      g07455(.A(new_n7710), .B(new_n7711), .C(new_n7709), .Y(new_n7712));
  NOR2xp33_ASAP7_75t_L      g07456(.A(new_n7706), .B(new_n7712), .Y(new_n7713));
  A2O1A1Ixp33_ASAP7_75t_L   g07457(.A1(new_n7412), .A2(new_n7372), .B(new_n7665), .C(new_n7713), .Y(new_n7714));
  AOI21xp33_ASAP7_75t_L     g07458(.A1(new_n7372), .A2(new_n7412), .B(new_n7665), .Y(new_n7715));
  OAI21xp33_ASAP7_75t_L     g07459(.A1(new_n7709), .A2(new_n7710), .B(new_n7711), .Y(new_n7716));
  NAND3xp33_ASAP7_75t_L     g07460(.A(new_n7705), .B(new_n7699), .C(new_n7702), .Y(new_n7717));
  NAND2xp33_ASAP7_75t_L     g07461(.A(new_n7717), .B(new_n7716), .Y(new_n7718));
  NAND2xp33_ASAP7_75t_L     g07462(.A(new_n7718), .B(new_n7715), .Y(new_n7719));
  AOI21xp33_ASAP7_75t_L     g07463(.A1(new_n7714), .A2(new_n7719), .B(new_n7664), .Y(new_n7720));
  INVx1_ASAP7_75t_L         g07464(.A(new_n7664), .Y(new_n7721));
  NOR2xp33_ASAP7_75t_L      g07465(.A(new_n7718), .B(new_n7715), .Y(new_n7722));
  AOI221xp5_ASAP7_75t_L     g07466(.A1(new_n7372), .A2(new_n7412), .B1(new_n7716), .B2(new_n7717), .C(new_n7665), .Y(new_n7723));
  NOR3xp33_ASAP7_75t_L      g07467(.A(new_n7722), .B(new_n7721), .C(new_n7723), .Y(new_n7724));
  OAI21xp33_ASAP7_75t_L     g07468(.A1(new_n7720), .A2(new_n7724), .B(new_n7661), .Y(new_n7725));
  AOI31xp33_ASAP7_75t_L     g07469(.A1(new_n7422), .A2(new_n7417), .A3(new_n7146), .B(new_n7425), .Y(new_n7726));
  OAI21xp33_ASAP7_75t_L     g07470(.A1(new_n7723), .A2(new_n7722), .B(new_n7721), .Y(new_n7727));
  NAND3xp33_ASAP7_75t_L     g07471(.A(new_n7714), .B(new_n7664), .C(new_n7719), .Y(new_n7728));
  NAND3xp33_ASAP7_75t_L     g07472(.A(new_n7726), .B(new_n7727), .C(new_n7728), .Y(new_n7729));
  NAND3xp33_ASAP7_75t_L     g07473(.A(new_n7725), .B(new_n7660), .C(new_n7729), .Y(new_n7730));
  AOI21xp33_ASAP7_75t_L     g07474(.A1(new_n7728), .A2(new_n7727), .B(new_n7726), .Y(new_n7731));
  NOR3xp33_ASAP7_75t_L      g07475(.A(new_n7661), .B(new_n7720), .C(new_n7724), .Y(new_n7732));
  OAI21xp33_ASAP7_75t_L     g07476(.A1(new_n7731), .A2(new_n7732), .B(new_n7659), .Y(new_n7733));
  NAND2xp33_ASAP7_75t_L     g07477(.A(new_n7730), .B(new_n7733), .Y(new_n7734));
  O2A1O1Ixp33_ASAP7_75t_L   g07478(.A1(new_n7656), .A2(new_n7430), .B(new_n7443), .C(new_n7734), .Y(new_n7735));
  NAND3xp33_ASAP7_75t_L     g07479(.A(new_n7427), .B(new_n7434), .C(new_n7423), .Y(new_n7736));
  A2O1A1Ixp33_ASAP7_75t_L   g07480(.A1(new_n7431), .A2(new_n7435), .B(new_n7369), .C(new_n7736), .Y(new_n7737));
  AOI21xp33_ASAP7_75t_L     g07481(.A1(new_n7733), .A2(new_n7730), .B(new_n7737), .Y(new_n7738));
  NOR3xp33_ASAP7_75t_L      g07482(.A(new_n7735), .B(new_n7738), .C(new_n7655), .Y(new_n7739));
  XNOR2x2_ASAP7_75t_L       g07483(.A(new_n3628), .B(new_n7654), .Y(new_n7740));
  NAND3xp33_ASAP7_75t_L     g07484(.A(new_n7737), .B(new_n7730), .C(new_n7733), .Y(new_n7741));
  NOR2xp33_ASAP7_75t_L      g07485(.A(new_n7430), .B(new_n7656), .Y(new_n7742));
  A2O1A1O1Ixp25_ASAP7_75t_L g07486(.A1(new_n7156), .A2(new_n7092), .B(new_n7162), .C(new_n7439), .D(new_n7742), .Y(new_n7743));
  NAND2xp33_ASAP7_75t_L     g07487(.A(new_n7734), .B(new_n7743), .Y(new_n7744));
  AOI21xp33_ASAP7_75t_L     g07488(.A1(new_n7744), .A2(new_n7741), .B(new_n7740), .Y(new_n7745));
  NOR2xp33_ASAP7_75t_L      g07489(.A(new_n7745), .B(new_n7739), .Y(new_n7746));
  A2O1A1Ixp33_ASAP7_75t_L   g07490(.A1(new_n7651), .A2(new_n7365), .B(new_n7652), .C(new_n7746), .Y(new_n7747));
  O2A1O1Ixp33_ASAP7_75t_L   g07491(.A1(new_n7451), .A2(new_n7452), .B(new_n7365), .C(new_n7652), .Y(new_n7748));
  NAND3xp33_ASAP7_75t_L     g07492(.A(new_n7744), .B(new_n7741), .C(new_n7740), .Y(new_n7749));
  OAI21xp33_ASAP7_75t_L     g07493(.A1(new_n7738), .A2(new_n7735), .B(new_n7655), .Y(new_n7750));
  NAND2xp33_ASAP7_75t_L     g07494(.A(new_n7749), .B(new_n7750), .Y(new_n7751));
  NAND2xp33_ASAP7_75t_L     g07495(.A(new_n7748), .B(new_n7751), .Y(new_n7752));
  AOI22xp33_ASAP7_75t_L     g07496(.A1(new_n3029), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n3258), .Y(new_n7753));
  OAI221xp5_ASAP7_75t_L     g07497(.A1(new_n3024), .A2(new_n1539), .B1(new_n3256), .B2(new_n1662), .C(new_n7753), .Y(new_n7754));
  NOR2xp33_ASAP7_75t_L      g07498(.A(new_n3015), .B(new_n7754), .Y(new_n7755));
  AND2x2_ASAP7_75t_L        g07499(.A(new_n3015), .B(new_n7754), .Y(new_n7756));
  NOR2xp33_ASAP7_75t_L      g07500(.A(new_n7755), .B(new_n7756), .Y(new_n7757));
  NAND3xp33_ASAP7_75t_L     g07501(.A(new_n7747), .B(new_n7752), .C(new_n7757), .Y(new_n7758));
  NOR2xp33_ASAP7_75t_L      g07502(.A(new_n7748), .B(new_n7751), .Y(new_n7759));
  AOI221xp5_ASAP7_75t_L     g07503(.A1(new_n7365), .A2(new_n7651), .B1(new_n7749), .B2(new_n7750), .C(new_n7652), .Y(new_n7760));
  OAI22xp33_ASAP7_75t_L     g07504(.A1(new_n7759), .A2(new_n7760), .B1(new_n7756), .B2(new_n7755), .Y(new_n7761));
  NAND2xp33_ASAP7_75t_L     g07505(.A(new_n7761), .B(new_n7758), .Y(new_n7762));
  A2O1A1Ixp33_ASAP7_75t_L   g07506(.A1(new_n7194), .A2(new_n7468), .B(new_n7461), .C(new_n7457), .Y(new_n7763));
  NOR2xp33_ASAP7_75t_L      g07507(.A(new_n7763), .B(new_n7762), .Y(new_n7764));
  AOI21xp33_ASAP7_75t_L     g07508(.A1(new_n7446), .A2(new_n7453), .B(new_n7456), .Y(new_n7765));
  A2O1A1O1Ixp25_ASAP7_75t_L g07509(.A1(new_n7183), .A2(new_n7362), .B(new_n7363), .C(new_n7458), .D(new_n7765), .Y(new_n7766));
  AOI21xp33_ASAP7_75t_L     g07510(.A1(new_n7761), .A2(new_n7758), .B(new_n7766), .Y(new_n7767));
  AOI22xp33_ASAP7_75t_L     g07511(.A1(new_n2552), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n2736), .Y(new_n7768));
  OAI221xp5_ASAP7_75t_L     g07512(.A1(new_n2547), .A2(new_n1909), .B1(new_n2734), .B2(new_n2477), .C(new_n7768), .Y(new_n7769));
  XNOR2x2_ASAP7_75t_L       g07513(.A(\a[29] ), .B(new_n7769), .Y(new_n7770));
  OAI21xp33_ASAP7_75t_L     g07514(.A1(new_n7767), .A2(new_n7764), .B(new_n7770), .Y(new_n7771));
  NAND3xp33_ASAP7_75t_L     g07515(.A(new_n7766), .B(new_n7761), .C(new_n7758), .Y(new_n7772));
  NAND2xp33_ASAP7_75t_L     g07516(.A(new_n7763), .B(new_n7762), .Y(new_n7773));
  XNOR2x2_ASAP7_75t_L       g07517(.A(new_n2538), .B(new_n7769), .Y(new_n7774));
  NAND3xp33_ASAP7_75t_L     g07518(.A(new_n7773), .B(new_n7772), .C(new_n7774), .Y(new_n7775));
  NAND2xp33_ASAP7_75t_L     g07519(.A(new_n7191), .B(new_n7474), .Y(new_n7776));
  NAND3xp33_ASAP7_75t_L     g07520(.A(new_n7210), .B(new_n7776), .C(new_n7472), .Y(new_n7777));
  NAND4xp25_ASAP7_75t_L     g07521(.A(new_n7777), .B(new_n7771), .C(new_n7775), .D(new_n7466), .Y(new_n7778));
  AOI21xp33_ASAP7_75t_L     g07522(.A1(new_n7773), .A2(new_n7772), .B(new_n7774), .Y(new_n7779));
  NOR3xp33_ASAP7_75t_L      g07523(.A(new_n7764), .B(new_n7767), .C(new_n7770), .Y(new_n7780));
  AOI211xp5_ASAP7_75t_L     g07524(.A1(new_n7358), .A2(new_n7197), .B(new_n7360), .C(new_n7477), .Y(new_n7781));
  OAI22xp33_ASAP7_75t_L     g07525(.A1(new_n7781), .A2(new_n7476), .B1(new_n7779), .B2(new_n7780), .Y(new_n7782));
  AOI22xp33_ASAP7_75t_L     g07526(.A1(new_n2114), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n2259), .Y(new_n7783));
  OAI221xp5_ASAP7_75t_L     g07527(.A1(new_n2109), .A2(new_n2348), .B1(new_n2257), .B2(new_n2505), .C(new_n7783), .Y(new_n7784));
  XNOR2x2_ASAP7_75t_L       g07528(.A(\a[26] ), .B(new_n7784), .Y(new_n7785));
  NAND3xp33_ASAP7_75t_L     g07529(.A(new_n7782), .B(new_n7778), .C(new_n7785), .Y(new_n7786));
  NOR4xp25_ASAP7_75t_L      g07530(.A(new_n7781), .B(new_n7780), .C(new_n7779), .D(new_n7476), .Y(new_n7787));
  AOI22xp33_ASAP7_75t_L     g07531(.A1(new_n7775), .A2(new_n7771), .B1(new_n7466), .B2(new_n7777), .Y(new_n7788));
  INVx1_ASAP7_75t_L         g07532(.A(new_n7785), .Y(new_n7789));
  OAI21xp33_ASAP7_75t_L     g07533(.A1(new_n7788), .A2(new_n7787), .B(new_n7789), .Y(new_n7790));
  AOI21xp33_ASAP7_75t_L     g07534(.A1(new_n7790), .A2(new_n7786), .B(new_n7650), .Y(new_n7791));
  A2O1A1Ixp33_ASAP7_75t_L   g07535(.A1(new_n7215), .A2(new_n7488), .B(new_n7489), .C(new_n7484), .Y(new_n7792));
  NAND2xp33_ASAP7_75t_L     g07536(.A(new_n7786), .B(new_n7790), .Y(new_n7793));
  NOR2xp33_ASAP7_75t_L      g07537(.A(new_n7792), .B(new_n7793), .Y(new_n7794));
  NOR3xp33_ASAP7_75t_L      g07538(.A(new_n7794), .B(new_n7791), .C(new_n7648), .Y(new_n7795));
  INVx1_ASAP7_75t_L         g07539(.A(new_n7648), .Y(new_n7796));
  NAND2xp33_ASAP7_75t_L     g07540(.A(new_n7792), .B(new_n7793), .Y(new_n7797));
  NOR3xp33_ASAP7_75t_L      g07541(.A(new_n7787), .B(new_n7788), .C(new_n7789), .Y(new_n7798));
  AOI21xp33_ASAP7_75t_L     g07542(.A1(new_n7782), .A2(new_n7778), .B(new_n7785), .Y(new_n7799));
  NOR2xp33_ASAP7_75t_L      g07543(.A(new_n7799), .B(new_n7798), .Y(new_n7800));
  NAND2xp33_ASAP7_75t_L     g07544(.A(new_n7650), .B(new_n7800), .Y(new_n7801));
  AOI21xp33_ASAP7_75t_L     g07545(.A1(new_n7801), .A2(new_n7797), .B(new_n7796), .Y(new_n7802));
  NOR3xp33_ASAP7_75t_L      g07546(.A(new_n7645), .B(new_n7802), .C(new_n7795), .Y(new_n7803));
  NAND3xp33_ASAP7_75t_L     g07547(.A(new_n7801), .B(new_n7797), .C(new_n7796), .Y(new_n7804));
  OAI21xp33_ASAP7_75t_L     g07548(.A1(new_n7791), .A2(new_n7794), .B(new_n7648), .Y(new_n7805));
  AOI221xp5_ASAP7_75t_L     g07549(.A1(new_n7500), .A2(new_n7492), .B1(new_n7804), .B2(new_n7805), .C(new_n7644), .Y(new_n7806));
  AOI22xp33_ASAP7_75t_L     g07550(.A1(new_n1360), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1581), .Y(new_n7807));
  OAI221xp5_ASAP7_75t_L     g07551(.A1(new_n1373), .A2(new_n3207), .B1(new_n1359), .B2(new_n3572), .C(new_n7807), .Y(new_n7808));
  NOR2xp33_ASAP7_75t_L      g07552(.A(new_n1356), .B(new_n7808), .Y(new_n7809));
  AND2x2_ASAP7_75t_L        g07553(.A(new_n1356), .B(new_n7808), .Y(new_n7810));
  NOR2xp33_ASAP7_75t_L      g07554(.A(new_n7809), .B(new_n7810), .Y(new_n7811));
  INVx1_ASAP7_75t_L         g07555(.A(new_n7811), .Y(new_n7812));
  NOR3xp33_ASAP7_75t_L      g07556(.A(new_n7812), .B(new_n7806), .C(new_n7803), .Y(new_n7813));
  OR3x1_ASAP7_75t_L         g07557(.A(new_n7645), .B(new_n7795), .C(new_n7802), .Y(new_n7814));
  OAI21xp33_ASAP7_75t_L     g07558(.A1(new_n7795), .A2(new_n7802), .B(new_n7645), .Y(new_n7815));
  AOI21xp33_ASAP7_75t_L     g07559(.A1(new_n7814), .A2(new_n7815), .B(new_n7811), .Y(new_n7816));
  OAI21xp33_ASAP7_75t_L     g07560(.A1(new_n7813), .A2(new_n7816), .B(new_n7643), .Y(new_n7817));
  A2O1A1O1Ixp25_ASAP7_75t_L g07561(.A1(new_n7244), .A2(new_n7246), .B(new_n7235), .C(new_n7497), .D(new_n7508), .Y(new_n7818));
  INVx1_ASAP7_75t_L         g07562(.A(new_n7813), .Y(new_n7819));
  INVx1_ASAP7_75t_L         g07563(.A(new_n7816), .Y(new_n7820));
  NAND3xp33_ASAP7_75t_L     g07564(.A(new_n7820), .B(new_n7819), .C(new_n7818), .Y(new_n7821));
  NAND3xp33_ASAP7_75t_L     g07565(.A(new_n7642), .B(new_n7821), .C(new_n7817), .Y(new_n7822));
  AOI21xp33_ASAP7_75t_L     g07566(.A1(new_n7820), .A2(new_n7819), .B(new_n7818), .Y(new_n7823));
  NOR3xp33_ASAP7_75t_L      g07567(.A(new_n7643), .B(new_n7813), .C(new_n7816), .Y(new_n7824));
  OAI21xp33_ASAP7_75t_L     g07568(.A1(new_n7824), .A2(new_n7823), .B(new_n7641), .Y(new_n7825));
  NAND2xp33_ASAP7_75t_L     g07569(.A(new_n7822), .B(new_n7825), .Y(new_n7826));
  NAND2xp33_ASAP7_75t_L     g07570(.A(new_n7826), .B(new_n7638), .Y(new_n7827));
  NOR3xp33_ASAP7_75t_L      g07571(.A(new_n7823), .B(new_n7824), .C(new_n7641), .Y(new_n7828));
  AOI21xp33_ASAP7_75t_L     g07572(.A1(new_n7821), .A2(new_n7817), .B(new_n7642), .Y(new_n7829));
  NOR2xp33_ASAP7_75t_L      g07573(.A(new_n7829), .B(new_n7828), .Y(new_n7830));
  A2O1A1Ixp33_ASAP7_75t_L   g07574(.A1(new_n7528), .A2(new_n7527), .B(new_n7637), .C(new_n7830), .Y(new_n7831));
  AOI22xp33_ASAP7_75t_L     g07575(.A1(new_n811), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n900), .Y(new_n7832));
  OAI221xp5_ASAP7_75t_L     g07576(.A1(new_n904), .A2(new_n4632), .B1(new_n898), .B2(new_n4858), .C(new_n7832), .Y(new_n7833));
  XNOR2x2_ASAP7_75t_L       g07577(.A(\a[14] ), .B(new_n7833), .Y(new_n7834));
  NAND3xp33_ASAP7_75t_L     g07578(.A(new_n7827), .B(new_n7831), .C(new_n7834), .Y(new_n7835));
  INVx1_ASAP7_75t_L         g07579(.A(new_n7637), .Y(new_n7836));
  A2O1A1Ixp33_ASAP7_75t_L   g07580(.A1(new_n7520), .A2(new_n7517), .B(new_n7525), .C(new_n7836), .Y(new_n7837));
  NOR2xp33_ASAP7_75t_L      g07581(.A(new_n7837), .B(new_n7830), .Y(new_n7838));
  O2A1O1Ixp33_ASAP7_75t_L   g07582(.A1(new_n7521), .A2(new_n7525), .B(new_n7836), .C(new_n7826), .Y(new_n7839));
  INVx1_ASAP7_75t_L         g07583(.A(new_n7834), .Y(new_n7840));
  OAI21xp33_ASAP7_75t_L     g07584(.A1(new_n7838), .A2(new_n7839), .B(new_n7840), .Y(new_n7841));
  NOR2xp33_ASAP7_75t_L      g07585(.A(new_n7535), .B(new_n7534), .Y(new_n7842));
  MAJIxp5_ASAP7_75t_L       g07586(.A(new_n7544), .B(new_n7536), .C(new_n7842), .Y(new_n7843));
  NAND3xp33_ASAP7_75t_L     g07587(.A(new_n7843), .B(new_n7841), .C(new_n7835), .Y(new_n7844));
  NAND2xp33_ASAP7_75t_L     g07588(.A(new_n7536), .B(new_n7842), .Y(new_n7845));
  AO22x1_ASAP7_75t_L        g07589(.A1(new_n7835), .A2(new_n7841), .B1(new_n7845), .B2(new_n7545), .Y(new_n7846));
  NOR2xp33_ASAP7_75t_L      g07590(.A(new_n5321), .B(new_n821), .Y(new_n7847));
  INVx1_ASAP7_75t_L         g07591(.A(new_n7847), .Y(new_n7848));
  NAND3xp33_ASAP7_75t_L     g07592(.A(new_n5343), .B(new_n578), .C(new_n5345), .Y(new_n7849));
  AOI22xp33_ASAP7_75t_L     g07593(.A1(\b[40] ), .A2(new_n651), .B1(\b[42] ), .B2(new_n581), .Y(new_n7850));
  AND4x1_ASAP7_75t_L        g07594(.A(new_n7850), .B(new_n7849), .C(new_n7848), .D(\a[11] ), .Y(new_n7851));
  AOI31xp33_ASAP7_75t_L     g07595(.A1(new_n7849), .A2(new_n7848), .A3(new_n7850), .B(\a[11] ), .Y(new_n7852));
  NOR2xp33_ASAP7_75t_L      g07596(.A(new_n7852), .B(new_n7851), .Y(new_n7853));
  INVx1_ASAP7_75t_L         g07597(.A(new_n7853), .Y(new_n7854));
  AOI21xp33_ASAP7_75t_L     g07598(.A1(new_n7846), .A2(new_n7844), .B(new_n7854), .Y(new_n7855));
  AND4x1_ASAP7_75t_L        g07599(.A(new_n7545), .B(new_n7845), .C(new_n7835), .D(new_n7841), .Y(new_n7856));
  AOI21xp33_ASAP7_75t_L     g07600(.A1(new_n7841), .A2(new_n7835), .B(new_n7843), .Y(new_n7857));
  NOR3xp33_ASAP7_75t_L      g07601(.A(new_n7856), .B(new_n7857), .C(new_n7853), .Y(new_n7858));
  NOR2xp33_ASAP7_75t_L      g07602(.A(new_n7858), .B(new_n7855), .Y(new_n7859));
  NAND2xp33_ASAP7_75t_L     g07603(.A(new_n7545), .B(new_n7540), .Y(new_n7860));
  MAJIxp5_ASAP7_75t_L       g07604(.A(new_n7563), .B(new_n7860), .C(new_n7551), .Y(new_n7861));
  NAND2xp33_ASAP7_75t_L     g07605(.A(new_n7861), .B(new_n7859), .Y(new_n7862));
  NOR2xp33_ASAP7_75t_L      g07606(.A(new_n7551), .B(new_n7860), .Y(new_n7863));
  INVx1_ASAP7_75t_L         g07607(.A(new_n7863), .Y(new_n7864));
  OAI221xp5_ASAP7_75t_L     g07608(.A1(new_n7855), .A2(new_n7858), .B1(new_n7563), .B2(new_n7561), .C(new_n7864), .Y(new_n7865));
  NAND2xp33_ASAP7_75t_L     g07609(.A(\b[44] ), .B(new_n447), .Y(new_n7866));
  NAND2xp33_ASAP7_75t_L     g07610(.A(new_n441), .B(new_n7066), .Y(new_n7867));
  AOI22xp33_ASAP7_75t_L     g07611(.A1(new_n444), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n471), .Y(new_n7868));
  AND4x1_ASAP7_75t_L        g07612(.A(new_n7868), .B(new_n7867), .C(new_n7866), .D(\a[8] ), .Y(new_n7869));
  AOI31xp33_ASAP7_75t_L     g07613(.A1(new_n7867), .A2(new_n7866), .A3(new_n7868), .B(\a[8] ), .Y(new_n7870));
  NOR2xp33_ASAP7_75t_L      g07614(.A(new_n7870), .B(new_n7869), .Y(new_n7871));
  NAND3xp33_ASAP7_75t_L     g07615(.A(new_n7862), .B(new_n7865), .C(new_n7871), .Y(new_n7872));
  OAI21xp33_ASAP7_75t_L     g07616(.A1(new_n7857), .A2(new_n7856), .B(new_n7853), .Y(new_n7873));
  NAND3xp33_ASAP7_75t_L     g07617(.A(new_n7846), .B(new_n7844), .C(new_n7854), .Y(new_n7874));
  NAND2xp33_ASAP7_75t_L     g07618(.A(new_n7873), .B(new_n7874), .Y(new_n7875));
  O2A1O1Ixp33_ASAP7_75t_L   g07619(.A1(new_n7563), .A2(new_n7561), .B(new_n7864), .C(new_n7875), .Y(new_n7876));
  NOR2xp33_ASAP7_75t_L      g07620(.A(new_n7861), .B(new_n7859), .Y(new_n7877));
  INVx1_ASAP7_75t_L         g07621(.A(new_n7871), .Y(new_n7878));
  OAI21xp33_ASAP7_75t_L     g07622(.A1(new_n7877), .A2(new_n7876), .B(new_n7878), .Y(new_n7879));
  NOR2xp33_ASAP7_75t_L      g07623(.A(new_n7293), .B(new_n7574), .Y(new_n7880));
  A2O1A1O1Ixp25_ASAP7_75t_L g07624(.A1(new_n7303), .A2(new_n7301), .B(new_n7880), .C(new_n7577), .D(new_n7568), .Y(new_n7881));
  AOI21xp33_ASAP7_75t_L     g07625(.A1(new_n7879), .A2(new_n7872), .B(new_n7881), .Y(new_n7882));
  NAND2xp33_ASAP7_75t_L     g07626(.A(new_n7872), .B(new_n7879), .Y(new_n7883));
  OAI21xp33_ASAP7_75t_L     g07627(.A1(new_n7572), .A2(new_n7339), .B(new_n7576), .Y(new_n7884));
  NOR2xp33_ASAP7_75t_L      g07628(.A(new_n7884), .B(new_n7883), .Y(new_n7885));
  OAI21xp33_ASAP7_75t_L     g07629(.A1(new_n7882), .A2(new_n7885), .B(new_n7635), .Y(new_n7886));
  INVx1_ASAP7_75t_L         g07630(.A(new_n7886), .Y(new_n7887));
  NOR3xp33_ASAP7_75t_L      g07631(.A(new_n7885), .B(new_n7635), .C(new_n7882), .Y(new_n7888));
  NOR3xp33_ASAP7_75t_L      g07632(.A(new_n7628), .B(new_n7887), .C(new_n7888), .Y(new_n7889));
  INVx1_ASAP7_75t_L         g07633(.A(new_n7888), .Y(new_n7890));
  AOI221xp5_ASAP7_75t_L     g07634(.A1(new_n7588), .A2(new_n7589), .B1(new_n7886), .B2(new_n7890), .C(new_n7627), .Y(new_n7891));
  NOR3xp33_ASAP7_75t_L      g07635(.A(new_n7889), .B(new_n7891), .C(new_n7626), .Y(new_n7892));
  INVx1_ASAP7_75t_L         g07636(.A(new_n7892), .Y(new_n7893));
  OAI21xp33_ASAP7_75t_L     g07637(.A1(new_n7891), .A2(new_n7889), .B(new_n7626), .Y(new_n7894));
  NAND2xp33_ASAP7_75t_L     g07638(.A(new_n7894), .B(new_n7893), .Y(new_n7895));
  XNOR2x2_ASAP7_75t_L       g07639(.A(new_n7613), .B(new_n7895), .Y(\f[51] ));
  INVx1_ASAP7_75t_L         g07640(.A(new_n7591), .Y(new_n7897));
  A2O1A1O1Ixp25_ASAP7_75t_L g07641(.A1(new_n7606), .A2(new_n7897), .B(new_n7610), .C(new_n7894), .D(new_n7892), .Y(new_n7898));
  NOR2xp33_ASAP7_75t_L      g07642(.A(\b[51] ), .B(\b[52] ), .Y(new_n7899));
  INVx1_ASAP7_75t_L         g07643(.A(\b[52] ), .Y(new_n7900));
  NOR2xp33_ASAP7_75t_L      g07644(.A(new_n7616), .B(new_n7900), .Y(new_n7901));
  NOR2xp33_ASAP7_75t_L      g07645(.A(new_n7899), .B(new_n7901), .Y(new_n7902));
  A2O1A1Ixp33_ASAP7_75t_L   g07646(.A1(\b[51] ), .A2(\b[50] ), .B(new_n7620), .C(new_n7902), .Y(new_n7903));
  O2A1O1Ixp33_ASAP7_75t_L   g07647(.A1(new_n7594), .A2(new_n7597), .B(new_n7618), .C(new_n7617), .Y(new_n7904));
  OAI21xp33_ASAP7_75t_L     g07648(.A1(new_n7899), .A2(new_n7901), .B(new_n7904), .Y(new_n7905));
  NAND2xp33_ASAP7_75t_L     g07649(.A(new_n7903), .B(new_n7905), .Y(new_n7906));
  AOI22xp33_ASAP7_75t_L     g07650(.A1(\b[50] ), .A2(new_n282), .B1(\b[52] ), .B2(new_n303), .Y(new_n7907));
  OAI221xp5_ASAP7_75t_L     g07651(.A1(new_n291), .A2(new_n7616), .B1(new_n268), .B2(new_n7906), .C(new_n7907), .Y(new_n7908));
  XNOR2x2_ASAP7_75t_L       g07652(.A(\a[2] ), .B(new_n7908), .Y(new_n7909));
  A2O1A1O1Ixp25_ASAP7_75t_L g07653(.A1(new_n7589), .A2(new_n7588), .B(new_n7627), .C(new_n7886), .D(new_n7888), .Y(new_n7910));
  NOR3xp33_ASAP7_75t_L      g07654(.A(new_n7876), .B(new_n7877), .C(new_n7878), .Y(new_n7911));
  AOI21xp33_ASAP7_75t_L     g07655(.A1(new_n7862), .A2(new_n7865), .B(new_n7871), .Y(new_n7912));
  NOR2xp33_ASAP7_75t_L      g07656(.A(new_n7912), .B(new_n7911), .Y(new_n7913));
  NAND2xp33_ASAP7_75t_L     g07657(.A(new_n7865), .B(new_n7862), .Y(new_n7914));
  NOR2xp33_ASAP7_75t_L      g07658(.A(new_n7871), .B(new_n7914), .Y(new_n7915));
  INVx1_ASAP7_75t_L         g07659(.A(new_n7915), .Y(new_n7916));
  NOR2xp33_ASAP7_75t_L      g07660(.A(new_n6321), .B(new_n468), .Y(new_n7917));
  INVx1_ASAP7_75t_L         g07661(.A(new_n7917), .Y(new_n7918));
  INVx1_ASAP7_75t_L         g07662(.A(new_n6573), .Y(new_n7919));
  NAND2xp33_ASAP7_75t_L     g07663(.A(new_n441), .B(new_n7919), .Y(new_n7920));
  AOI22xp33_ASAP7_75t_L     g07664(.A1(new_n444), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n471), .Y(new_n7921));
  AND4x1_ASAP7_75t_L        g07665(.A(new_n7921), .B(new_n7920), .C(new_n7918), .D(\a[8] ), .Y(new_n7922));
  AOI31xp33_ASAP7_75t_L     g07666(.A1(new_n7920), .A2(new_n7918), .A3(new_n7921), .B(\a[8] ), .Y(new_n7923));
  NOR2xp33_ASAP7_75t_L      g07667(.A(new_n7923), .B(new_n7922), .Y(new_n7924));
  NAND3xp33_ASAP7_75t_L     g07668(.A(new_n7782), .B(new_n7778), .C(new_n7789), .Y(new_n7925));
  AOI22xp33_ASAP7_75t_L     g07669(.A1(new_n2114), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n2259), .Y(new_n7926));
  OAI221xp5_ASAP7_75t_L     g07670(.A1(new_n2109), .A2(new_n2497), .B1(new_n2257), .B2(new_n2672), .C(new_n7926), .Y(new_n7927));
  XNOR2x2_ASAP7_75t_L       g07671(.A(\a[26] ), .B(new_n7927), .Y(new_n7928));
  AOI31xp33_ASAP7_75t_L     g07672(.A1(new_n7777), .A2(new_n7771), .A3(new_n7466), .B(new_n7780), .Y(new_n7929));
  XNOR2x2_ASAP7_75t_L       g07673(.A(new_n7748), .B(new_n7751), .Y(new_n7930));
  NOR2xp33_ASAP7_75t_L      g07674(.A(new_n7757), .B(new_n7930), .Y(new_n7931));
  INVx1_ASAP7_75t_L         g07675(.A(new_n7931), .Y(new_n7932));
  AOI22xp33_ASAP7_75t_L     g07676(.A1(new_n3029), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n3258), .Y(new_n7933));
  OAI221xp5_ASAP7_75t_L     g07677(.A1(new_n3024), .A2(new_n1655), .B1(new_n3256), .B2(new_n1780), .C(new_n7933), .Y(new_n7934));
  NOR2xp33_ASAP7_75t_L      g07678(.A(new_n3015), .B(new_n7934), .Y(new_n7935));
  AND2x2_ASAP7_75t_L        g07679(.A(new_n3015), .B(new_n7934), .Y(new_n7936));
  A2O1A1O1Ixp25_ASAP7_75t_L g07680(.A1(new_n7365), .A2(new_n7651), .B(new_n7652), .C(new_n7750), .D(new_n7739), .Y(new_n7937));
  NAND2xp33_ASAP7_75t_L     g07681(.A(new_n7719), .B(new_n7714), .Y(new_n7938));
  MAJIxp5_ASAP7_75t_L       g07682(.A(new_n7726), .B(new_n7664), .C(new_n7938), .Y(new_n7939));
  AOI22xp33_ASAP7_75t_L     g07683(.A1(new_n4920), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n5167), .Y(new_n7940));
  OAI221xp5_ASAP7_75t_L     g07684(.A1(new_n5154), .A2(new_n760), .B1(new_n5158), .B2(new_n790), .C(new_n7940), .Y(new_n7941));
  XNOR2x2_ASAP7_75t_L       g07685(.A(\a[41] ), .B(new_n7941), .Y(new_n7942));
  NOR3xp33_ASAP7_75t_L      g07686(.A(new_n7395), .B(new_n7674), .C(new_n7394), .Y(new_n7943));
  NAND2xp33_ASAP7_75t_L     g07687(.A(\b[3] ), .B(new_n7115), .Y(new_n7944));
  NAND2xp33_ASAP7_75t_L     g07688(.A(new_n7108), .B(new_n329), .Y(new_n7945));
  AOI22xp33_ASAP7_75t_L     g07689(.A1(new_n7111), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n7391), .Y(new_n7946));
  NAND4xp25_ASAP7_75t_L     g07690(.A(new_n7945), .B(\a[50] ), .C(new_n7944), .D(new_n7946), .Y(new_n7947));
  AOI31xp33_ASAP7_75t_L     g07691(.A1(new_n7945), .A2(new_n7944), .A3(new_n7946), .B(\a[50] ), .Y(new_n7948));
  INVx1_ASAP7_75t_L         g07692(.A(new_n7948), .Y(new_n7949));
  NAND2xp33_ASAP7_75t_L     g07693(.A(\a[53] ), .B(new_n7670), .Y(new_n7950));
  NAND2xp33_ASAP7_75t_L     g07694(.A(new_n7668), .B(new_n7667), .Y(new_n7951));
  INVx1_ASAP7_75t_L         g07695(.A(\a[52] ), .Y(new_n7952));
  NAND2xp33_ASAP7_75t_L     g07696(.A(\a[53] ), .B(new_n7952), .Y(new_n7953));
  INVx1_ASAP7_75t_L         g07697(.A(\a[53] ), .Y(new_n7954));
  NAND2xp33_ASAP7_75t_L     g07698(.A(\a[52] ), .B(new_n7954), .Y(new_n7955));
  NAND2xp33_ASAP7_75t_L     g07699(.A(new_n7955), .B(new_n7953), .Y(new_n7956));
  NAND2xp33_ASAP7_75t_L     g07700(.A(new_n7956), .B(new_n7951), .Y(new_n7957));
  INVx1_ASAP7_75t_L         g07701(.A(new_n7957), .Y(new_n7958));
  NAND2xp33_ASAP7_75t_L     g07702(.A(new_n269), .B(new_n7958), .Y(new_n7959));
  NOR2xp33_ASAP7_75t_L      g07703(.A(new_n7956), .B(new_n7669), .Y(new_n7960));
  NAND2xp33_ASAP7_75t_L     g07704(.A(\b[1] ), .B(new_n7960), .Y(new_n7961));
  XNOR2x2_ASAP7_75t_L       g07705(.A(\a[52] ), .B(\a[51] ), .Y(new_n7962));
  NOR2xp33_ASAP7_75t_L      g07706(.A(new_n7962), .B(new_n7951), .Y(new_n7963));
  NAND2xp33_ASAP7_75t_L     g07707(.A(\b[0] ), .B(new_n7963), .Y(new_n7964));
  NAND3xp33_ASAP7_75t_L     g07708(.A(new_n7959), .B(new_n7961), .C(new_n7964), .Y(new_n7965));
  XOR2x2_ASAP7_75t_L        g07709(.A(new_n7950), .B(new_n7965), .Y(new_n7966));
  NAND3xp33_ASAP7_75t_L     g07710(.A(new_n7966), .B(new_n7949), .C(new_n7947), .Y(new_n7967));
  INVx1_ASAP7_75t_L         g07711(.A(new_n7947), .Y(new_n7968));
  XNOR2x2_ASAP7_75t_L       g07712(.A(new_n7950), .B(new_n7965), .Y(new_n7969));
  OAI21xp33_ASAP7_75t_L     g07713(.A1(new_n7948), .A2(new_n7968), .B(new_n7969), .Y(new_n7970));
  OAI211xp5_ASAP7_75t_L     g07714(.A1(new_n7943), .A2(new_n7692), .B(new_n7967), .C(new_n7970), .Y(new_n7971));
  NOR2xp33_ASAP7_75t_L      g07715(.A(new_n7394), .B(new_n7395), .Y(new_n7972));
  NAND2xp33_ASAP7_75t_L     g07716(.A(new_n7679), .B(new_n7681), .Y(new_n7973));
  MAJIxp5_ASAP7_75t_L       g07717(.A(new_n7973), .B(new_n7670), .C(new_n7972), .Y(new_n7974));
  NOR3xp33_ASAP7_75t_L      g07718(.A(new_n7969), .B(new_n7948), .C(new_n7968), .Y(new_n7975));
  AOI21xp33_ASAP7_75t_L     g07719(.A1(new_n7949), .A2(new_n7947), .B(new_n7966), .Y(new_n7976));
  OAI21xp33_ASAP7_75t_L     g07720(.A1(new_n7975), .A2(new_n7976), .B(new_n7974), .Y(new_n7977));
  AOI22xp33_ASAP7_75t_L     g07721(.A1(new_n6376), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n6648), .Y(new_n7978));
  OAI221xp5_ASAP7_75t_L     g07722(.A1(new_n6646), .A2(new_n418), .B1(new_n6636), .B2(new_n425), .C(new_n7978), .Y(new_n7979));
  XNOR2x2_ASAP7_75t_L       g07723(.A(\a[47] ), .B(new_n7979), .Y(new_n7980));
  NAND3xp33_ASAP7_75t_L     g07724(.A(new_n7977), .B(new_n7971), .C(new_n7980), .Y(new_n7981));
  NOR3xp33_ASAP7_75t_L      g07725(.A(new_n7974), .B(new_n7975), .C(new_n7976), .Y(new_n7982));
  AOI211xp5_ASAP7_75t_L     g07726(.A1(new_n7967), .A2(new_n7970), .B(new_n7943), .C(new_n7692), .Y(new_n7983));
  XNOR2x2_ASAP7_75t_L       g07727(.A(new_n6371), .B(new_n7979), .Y(new_n7984));
  OAI21xp33_ASAP7_75t_L     g07728(.A1(new_n7983), .A2(new_n7982), .B(new_n7984), .Y(new_n7985));
  AOI211xp5_ASAP7_75t_L     g07729(.A1(new_n7690), .A2(new_n7688), .B(new_n7692), .C(new_n7693), .Y(new_n7986));
  A2O1A1O1Ixp25_ASAP7_75t_L g07730(.A1(new_n7404), .A2(new_n7403), .B(new_n7701), .C(new_n7700), .D(new_n7986), .Y(new_n7987));
  NAND3xp33_ASAP7_75t_L     g07731(.A(new_n7987), .B(new_n7985), .C(new_n7981), .Y(new_n7988));
  NAND2xp33_ASAP7_75t_L     g07732(.A(new_n7981), .B(new_n7985), .Y(new_n7989));
  INVx1_ASAP7_75t_L         g07733(.A(new_n7986), .Y(new_n7990));
  A2O1A1Ixp33_ASAP7_75t_L   g07734(.A1(new_n7695), .A2(new_n7691), .B(new_n7698), .C(new_n7990), .Y(new_n7991));
  NAND2xp33_ASAP7_75t_L     g07735(.A(new_n7989), .B(new_n7991), .Y(new_n7992));
  AOI22xp33_ASAP7_75t_L     g07736(.A1(new_n5624), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n5901), .Y(new_n7993));
  OAI221xp5_ASAP7_75t_L     g07737(.A1(new_n5900), .A2(new_n540), .B1(new_n5892), .B2(new_n624), .C(new_n7993), .Y(new_n7994));
  XNOR2x2_ASAP7_75t_L       g07738(.A(\a[44] ), .B(new_n7994), .Y(new_n7995));
  INVx1_ASAP7_75t_L         g07739(.A(new_n7995), .Y(new_n7996));
  AOI21xp33_ASAP7_75t_L     g07740(.A1(new_n7992), .A2(new_n7988), .B(new_n7996), .Y(new_n7997));
  NOR2xp33_ASAP7_75t_L      g07741(.A(new_n7989), .B(new_n7991), .Y(new_n7998));
  AOI21xp33_ASAP7_75t_L     g07742(.A1(new_n7985), .A2(new_n7981), .B(new_n7987), .Y(new_n7999));
  NOR3xp33_ASAP7_75t_L      g07743(.A(new_n7998), .B(new_n7999), .C(new_n7995), .Y(new_n8000));
  NOR2xp33_ASAP7_75t_L      g07744(.A(new_n7997), .B(new_n8000), .Y(new_n8001));
  NOR3xp33_ASAP7_75t_L      g07745(.A(new_n7722), .B(new_n8001), .C(new_n7712), .Y(new_n8002));
  OAI21xp33_ASAP7_75t_L     g07746(.A1(new_n7999), .A2(new_n7998), .B(new_n7995), .Y(new_n8003));
  NAND3xp33_ASAP7_75t_L     g07747(.A(new_n7996), .B(new_n7992), .C(new_n7988), .Y(new_n8004));
  NAND2xp33_ASAP7_75t_L     g07748(.A(new_n8004), .B(new_n8003), .Y(new_n8005));
  O2A1O1Ixp33_ASAP7_75t_L   g07749(.A1(new_n7715), .A2(new_n7706), .B(new_n7717), .C(new_n8005), .Y(new_n8006));
  OAI21xp33_ASAP7_75t_L     g07750(.A1(new_n8006), .A2(new_n8002), .B(new_n7942), .Y(new_n8007));
  INVx1_ASAP7_75t_L         g07751(.A(new_n7942), .Y(new_n8008));
  A2O1A1O1Ixp25_ASAP7_75t_L g07752(.A1(new_n7412), .A2(new_n7372), .B(new_n7665), .C(new_n7716), .D(new_n7712), .Y(new_n8009));
  NAND2xp33_ASAP7_75t_L     g07753(.A(new_n8009), .B(new_n8005), .Y(new_n8010));
  NOR2xp33_ASAP7_75t_L      g07754(.A(new_n7709), .B(new_n7710), .Y(new_n8011));
  A2O1A1Ixp33_ASAP7_75t_L   g07755(.A1(new_n7705), .A2(new_n8011), .B(new_n7722), .C(new_n8001), .Y(new_n8012));
  NAND3xp33_ASAP7_75t_L     g07756(.A(new_n8012), .B(new_n8010), .C(new_n8008), .Y(new_n8013));
  NAND3xp33_ASAP7_75t_L     g07757(.A(new_n7939), .B(new_n8007), .C(new_n8013), .Y(new_n8014));
  NOR2xp33_ASAP7_75t_L      g07758(.A(new_n7723), .B(new_n7722), .Y(new_n8015));
  NAND2xp33_ASAP7_75t_L     g07759(.A(new_n7721), .B(new_n8015), .Y(new_n8016));
  AOI21xp33_ASAP7_75t_L     g07760(.A1(new_n8012), .A2(new_n8010), .B(new_n8008), .Y(new_n8017));
  NOR3xp33_ASAP7_75t_L      g07761(.A(new_n8002), .B(new_n8006), .C(new_n7942), .Y(new_n8018));
  OAI211xp5_ASAP7_75t_L     g07762(.A1(new_n8017), .A2(new_n8018), .B(new_n7725), .C(new_n8016), .Y(new_n8019));
  AOI22xp33_ASAP7_75t_L     g07763(.A1(new_n4283), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n4512), .Y(new_n8020));
  OAI221xp5_ASAP7_75t_L     g07764(.A1(new_n4277), .A2(new_n942), .B1(new_n4499), .B2(new_n1035), .C(new_n8020), .Y(new_n8021));
  XNOR2x2_ASAP7_75t_L       g07765(.A(\a[38] ), .B(new_n8021), .Y(new_n8022));
  NAND3xp33_ASAP7_75t_L     g07766(.A(new_n8019), .B(new_n8014), .C(new_n8022), .Y(new_n8023));
  AO21x2_ASAP7_75t_L        g07767(.A1(new_n8014), .A2(new_n8019), .B(new_n8022), .Y(new_n8024));
  NOR3xp33_ASAP7_75t_L      g07768(.A(new_n7732), .B(new_n7731), .C(new_n7659), .Y(new_n8025));
  A2O1A1O1Ixp25_ASAP7_75t_L g07769(.A1(new_n7439), .A2(new_n7438), .B(new_n7742), .C(new_n7733), .D(new_n8025), .Y(new_n8026));
  NAND3xp33_ASAP7_75t_L     g07770(.A(new_n8026), .B(new_n8024), .C(new_n8023), .Y(new_n8027));
  AO21x2_ASAP7_75t_L        g07771(.A1(new_n8023), .A2(new_n8024), .B(new_n8026), .Y(new_n8028));
  AOI22xp33_ASAP7_75t_L     g07772(.A1(new_n3633), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n3858), .Y(new_n8029));
  OAI221xp5_ASAP7_75t_L     g07773(.A1(new_n3853), .A2(new_n1313), .B1(new_n3856), .B2(new_n1438), .C(new_n8029), .Y(new_n8030));
  XNOR2x2_ASAP7_75t_L       g07774(.A(new_n3628), .B(new_n8030), .Y(new_n8031));
  AOI21xp33_ASAP7_75t_L     g07775(.A1(new_n8028), .A2(new_n8027), .B(new_n8031), .Y(new_n8032));
  AND3x1_ASAP7_75t_L        g07776(.A(new_n8028), .B(new_n8031), .C(new_n8027), .Y(new_n8033));
  OAI21xp33_ASAP7_75t_L     g07777(.A1(new_n8032), .A2(new_n8033), .B(new_n7937), .Y(new_n8034));
  OAI21xp33_ASAP7_75t_L     g07778(.A1(new_n7745), .A2(new_n7748), .B(new_n7749), .Y(new_n8035));
  INVx1_ASAP7_75t_L         g07779(.A(new_n8032), .Y(new_n8036));
  NAND3xp33_ASAP7_75t_L     g07780(.A(new_n8028), .B(new_n8027), .C(new_n8031), .Y(new_n8037));
  NAND3xp33_ASAP7_75t_L     g07781(.A(new_n8035), .B(new_n8036), .C(new_n8037), .Y(new_n8038));
  OAI211xp5_ASAP7_75t_L     g07782(.A1(new_n7935), .A2(new_n7936), .B(new_n8038), .C(new_n8034), .Y(new_n8039));
  NOR2xp33_ASAP7_75t_L      g07783(.A(new_n7935), .B(new_n7936), .Y(new_n8040));
  OA21x2_ASAP7_75t_L        g07784(.A1(new_n8032), .A2(new_n8033), .B(new_n7937), .Y(new_n8041));
  NOR3xp33_ASAP7_75t_L      g07785(.A(new_n7937), .B(new_n8032), .C(new_n8033), .Y(new_n8042));
  OAI21xp33_ASAP7_75t_L     g07786(.A1(new_n8042), .A2(new_n8041), .B(new_n8040), .Y(new_n8043));
  NAND2xp33_ASAP7_75t_L     g07787(.A(new_n8043), .B(new_n8039), .Y(new_n8044));
  NAND3xp33_ASAP7_75t_L     g07788(.A(new_n7773), .B(new_n7932), .C(new_n8044), .Y(new_n8045));
  NOR3xp33_ASAP7_75t_L      g07789(.A(new_n8041), .B(new_n8042), .C(new_n8040), .Y(new_n8046));
  OA21x2_ASAP7_75t_L        g07790(.A1(new_n8042), .A2(new_n8041), .B(new_n8040), .Y(new_n8047));
  NOR2xp33_ASAP7_75t_L      g07791(.A(new_n8046), .B(new_n8047), .Y(new_n8048));
  A2O1A1Ixp33_ASAP7_75t_L   g07792(.A1(new_n7763), .A2(new_n7762), .B(new_n7931), .C(new_n8048), .Y(new_n8049));
  AOI22xp33_ASAP7_75t_L     g07793(.A1(new_n2552), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n2736), .Y(new_n8050));
  OAI221xp5_ASAP7_75t_L     g07794(.A1(new_n2547), .A2(new_n1929), .B1(new_n2734), .B2(new_n2075), .C(new_n8050), .Y(new_n8051));
  XNOR2x2_ASAP7_75t_L       g07795(.A(\a[29] ), .B(new_n8051), .Y(new_n8052));
  NAND3xp33_ASAP7_75t_L     g07796(.A(new_n8049), .B(new_n8045), .C(new_n8052), .Y(new_n8053));
  MAJIxp5_ASAP7_75t_L       g07797(.A(new_n7766), .B(new_n7930), .C(new_n7757), .Y(new_n8054));
  NOR2xp33_ASAP7_75t_L      g07798(.A(new_n8054), .B(new_n8048), .Y(new_n8055));
  AND2x2_ASAP7_75t_L        g07799(.A(new_n7761), .B(new_n7758), .Y(new_n8056));
  O2A1O1Ixp33_ASAP7_75t_L   g07800(.A1(new_n8056), .A2(new_n7766), .B(new_n7932), .C(new_n8044), .Y(new_n8057));
  INVx1_ASAP7_75t_L         g07801(.A(new_n8052), .Y(new_n8058));
  OAI21xp33_ASAP7_75t_L     g07802(.A1(new_n8055), .A2(new_n8057), .B(new_n8058), .Y(new_n8059));
  AOI21xp33_ASAP7_75t_L     g07803(.A1(new_n8059), .A2(new_n8053), .B(new_n7929), .Y(new_n8060));
  OAI31xp33_ASAP7_75t_L     g07804(.A1(new_n7781), .A2(new_n7779), .A3(new_n7476), .B(new_n7775), .Y(new_n8061));
  NOR3xp33_ASAP7_75t_L      g07805(.A(new_n8058), .B(new_n8057), .C(new_n8055), .Y(new_n8062));
  AOI21xp33_ASAP7_75t_L     g07806(.A1(new_n8049), .A2(new_n8045), .B(new_n8052), .Y(new_n8063));
  NOR3xp33_ASAP7_75t_L      g07807(.A(new_n8061), .B(new_n8062), .C(new_n8063), .Y(new_n8064));
  NOR3xp33_ASAP7_75t_L      g07808(.A(new_n8064), .B(new_n8060), .C(new_n7928), .Y(new_n8065));
  INVx1_ASAP7_75t_L         g07809(.A(new_n7928), .Y(new_n8066));
  OAI21xp33_ASAP7_75t_L     g07810(.A1(new_n8062), .A2(new_n8063), .B(new_n8061), .Y(new_n8067));
  NAND3xp33_ASAP7_75t_L     g07811(.A(new_n7929), .B(new_n8053), .C(new_n8059), .Y(new_n8068));
  AOI21xp33_ASAP7_75t_L     g07812(.A1(new_n8068), .A2(new_n8067), .B(new_n8066), .Y(new_n8069));
  OAI221xp5_ASAP7_75t_L     g07813(.A1(new_n7800), .A2(new_n7650), .B1(new_n8069), .B2(new_n8065), .C(new_n7925), .Y(new_n8070));
  A2O1A1Ixp33_ASAP7_75t_L   g07814(.A1(new_n7786), .A2(new_n7790), .B(new_n7650), .C(new_n7925), .Y(new_n8071));
  NAND3xp33_ASAP7_75t_L     g07815(.A(new_n8068), .B(new_n8067), .C(new_n8066), .Y(new_n8072));
  OAI21xp33_ASAP7_75t_L     g07816(.A1(new_n8060), .A2(new_n8064), .B(new_n7928), .Y(new_n8073));
  NAND3xp33_ASAP7_75t_L     g07817(.A(new_n8071), .B(new_n8072), .C(new_n8073), .Y(new_n8074));
  AOI22xp33_ASAP7_75t_L     g07818(.A1(new_n1704), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1837), .Y(new_n8075));
  OAI221xp5_ASAP7_75t_L     g07819(.A1(new_n1699), .A2(new_n2982), .B1(new_n1827), .B2(new_n3187), .C(new_n8075), .Y(new_n8076));
  XNOR2x2_ASAP7_75t_L       g07820(.A(\a[23] ), .B(new_n8076), .Y(new_n8077));
  NAND3xp33_ASAP7_75t_L     g07821(.A(new_n8074), .B(new_n8070), .C(new_n8077), .Y(new_n8078));
  AO21x2_ASAP7_75t_L        g07822(.A1(new_n8070), .A2(new_n8074), .B(new_n8077), .Y(new_n8079));
  A2O1A1O1Ixp25_ASAP7_75t_L g07823(.A1(new_n7492), .A2(new_n7500), .B(new_n7644), .C(new_n7805), .D(new_n7795), .Y(new_n8080));
  NAND3xp33_ASAP7_75t_L     g07824(.A(new_n8080), .B(new_n8079), .C(new_n8078), .Y(new_n8081));
  AND3x1_ASAP7_75t_L        g07825(.A(new_n8074), .B(new_n8070), .C(new_n8077), .Y(new_n8082));
  AOI21xp33_ASAP7_75t_L     g07826(.A1(new_n8074), .A2(new_n8070), .B(new_n8077), .Y(new_n8083));
  OAI21xp33_ASAP7_75t_L     g07827(.A1(new_n7802), .A2(new_n7645), .B(new_n7804), .Y(new_n8084));
  OAI21xp33_ASAP7_75t_L     g07828(.A1(new_n8082), .A2(new_n8083), .B(new_n8084), .Y(new_n8085));
  AOI22xp33_ASAP7_75t_L     g07829(.A1(new_n1360), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1581), .Y(new_n8086));
  OAI221xp5_ASAP7_75t_L     g07830(.A1(new_n1373), .A2(new_n3565), .B1(new_n1359), .B2(new_n3591), .C(new_n8086), .Y(new_n8087));
  XNOR2x2_ASAP7_75t_L       g07831(.A(\a[20] ), .B(new_n8087), .Y(new_n8088));
  NAND3xp33_ASAP7_75t_L     g07832(.A(new_n8081), .B(new_n8085), .C(new_n8088), .Y(new_n8089));
  NAND2xp33_ASAP7_75t_L     g07833(.A(new_n8078), .B(new_n8079), .Y(new_n8090));
  NOR2xp33_ASAP7_75t_L      g07834(.A(new_n8084), .B(new_n8090), .Y(new_n8091));
  AOI21xp33_ASAP7_75t_L     g07835(.A1(new_n8079), .A2(new_n8078), .B(new_n8080), .Y(new_n8092));
  INVx1_ASAP7_75t_L         g07836(.A(new_n8088), .Y(new_n8093));
  OAI21xp33_ASAP7_75t_L     g07837(.A1(new_n8092), .A2(new_n8091), .B(new_n8093), .Y(new_n8094));
  NOR2xp33_ASAP7_75t_L      g07838(.A(new_n7803), .B(new_n7806), .Y(new_n8095));
  NAND2xp33_ASAP7_75t_L     g07839(.A(new_n7812), .B(new_n8095), .Y(new_n8096));
  NAND4xp25_ASAP7_75t_L     g07840(.A(new_n7817), .B(new_n8096), .C(new_n8094), .D(new_n8089), .Y(new_n8097));
  NOR3xp33_ASAP7_75t_L      g07841(.A(new_n8091), .B(new_n8092), .C(new_n8093), .Y(new_n8098));
  AOI21xp33_ASAP7_75t_L     g07842(.A1(new_n8081), .A2(new_n8085), .B(new_n8088), .Y(new_n8099));
  NAND2xp33_ASAP7_75t_L     g07843(.A(new_n7815), .B(new_n7814), .Y(new_n8100));
  MAJIxp5_ASAP7_75t_L       g07844(.A(new_n7818), .B(new_n7811), .C(new_n8100), .Y(new_n8101));
  OAI21xp33_ASAP7_75t_L     g07845(.A1(new_n8098), .A2(new_n8099), .B(new_n8101), .Y(new_n8102));
  AOI22xp33_ASAP7_75t_L     g07846(.A1(new_n1076), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1253), .Y(new_n8103));
  OAI221xp5_ASAP7_75t_L     g07847(.A1(new_n1154), .A2(new_n4216), .B1(new_n1156), .B2(new_n4431), .C(new_n8103), .Y(new_n8104));
  XNOR2x2_ASAP7_75t_L       g07848(.A(\a[17] ), .B(new_n8104), .Y(new_n8105));
  NAND3xp33_ASAP7_75t_L     g07849(.A(new_n8097), .B(new_n8102), .C(new_n8105), .Y(new_n8106));
  NOR3xp33_ASAP7_75t_L      g07850(.A(new_n8101), .B(new_n8099), .C(new_n8098), .Y(new_n8107));
  MAJIxp5_ASAP7_75t_L       g07851(.A(new_n7643), .B(new_n8095), .C(new_n7812), .Y(new_n8108));
  AOI21xp33_ASAP7_75t_L     g07852(.A1(new_n8094), .A2(new_n8089), .B(new_n8108), .Y(new_n8109));
  INVx1_ASAP7_75t_L         g07853(.A(new_n8105), .Y(new_n8110));
  OAI21xp33_ASAP7_75t_L     g07854(.A1(new_n8107), .A2(new_n8109), .B(new_n8110), .Y(new_n8111));
  A2O1A1O1Ixp25_ASAP7_75t_L g07855(.A1(new_n7527), .A2(new_n7528), .B(new_n7637), .C(new_n7825), .D(new_n7828), .Y(new_n8112));
  NAND3xp33_ASAP7_75t_L     g07856(.A(new_n8112), .B(new_n8111), .C(new_n8106), .Y(new_n8113));
  NAND2xp33_ASAP7_75t_L     g07857(.A(new_n8106), .B(new_n8111), .Y(new_n8114));
  A2O1A1Ixp33_ASAP7_75t_L   g07858(.A1(new_n7830), .A2(new_n7837), .B(new_n7828), .C(new_n8114), .Y(new_n8115));
  NOR2xp33_ASAP7_75t_L      g07859(.A(new_n4848), .B(new_n904), .Y(new_n8116));
  INVx1_ASAP7_75t_L         g07860(.A(new_n8116), .Y(new_n8117));
  NAND2xp33_ASAP7_75t_L     g07861(.A(new_n808), .B(new_n4876), .Y(new_n8118));
  AOI22xp33_ASAP7_75t_L     g07862(.A1(new_n811), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n900), .Y(new_n8119));
  AND4x1_ASAP7_75t_L        g07863(.A(new_n8119), .B(new_n8118), .C(new_n8117), .D(\a[14] ), .Y(new_n8120));
  AOI31xp33_ASAP7_75t_L     g07864(.A1(new_n8118), .A2(new_n8117), .A3(new_n8119), .B(\a[14] ), .Y(new_n8121));
  NOR2xp33_ASAP7_75t_L      g07865(.A(new_n8121), .B(new_n8120), .Y(new_n8122));
  NAND3xp33_ASAP7_75t_L     g07866(.A(new_n8115), .B(new_n8122), .C(new_n8113), .Y(new_n8123));
  AND3x1_ASAP7_75t_L        g07867(.A(new_n8112), .B(new_n8111), .C(new_n8106), .Y(new_n8124));
  AOI21xp33_ASAP7_75t_L     g07868(.A1(new_n8111), .A2(new_n8106), .B(new_n8112), .Y(new_n8125));
  INVx1_ASAP7_75t_L         g07869(.A(new_n8122), .Y(new_n8126));
  OAI21xp33_ASAP7_75t_L     g07870(.A1(new_n8125), .A2(new_n8124), .B(new_n8126), .Y(new_n8127));
  NAND3xp33_ASAP7_75t_L     g07871(.A(new_n7827), .B(new_n7831), .C(new_n7840), .Y(new_n8128));
  NAND4xp25_ASAP7_75t_L     g07872(.A(new_n7846), .B(new_n8128), .C(new_n8127), .D(new_n8123), .Y(new_n8129));
  NAND2xp33_ASAP7_75t_L     g07873(.A(new_n8123), .B(new_n8127), .Y(new_n8130));
  A2O1A1Ixp33_ASAP7_75t_L   g07874(.A1(new_n7841), .A2(new_n7835), .B(new_n7843), .C(new_n8128), .Y(new_n8131));
  NAND2xp33_ASAP7_75t_L     g07875(.A(new_n8131), .B(new_n8130), .Y(new_n8132));
  AOI22xp33_ASAP7_75t_L     g07876(.A1(\b[41] ), .A2(new_n651), .B1(\b[43] ), .B2(new_n581), .Y(new_n8133));
  INVx1_ASAP7_75t_L         g07877(.A(new_n8133), .Y(new_n8134));
  AOI221xp5_ASAP7_75t_L     g07878(.A1(\b[42] ), .A2(new_n584), .B1(new_n578), .B2(new_n5812), .C(new_n8134), .Y(new_n8135));
  XNOR2x2_ASAP7_75t_L       g07879(.A(\a[11] ), .B(new_n8135), .Y(new_n8136));
  AO21x2_ASAP7_75t_L        g07880(.A1(new_n8132), .A2(new_n8129), .B(new_n8136), .Y(new_n8137));
  NAND3xp33_ASAP7_75t_L     g07881(.A(new_n8129), .B(new_n8132), .C(new_n8136), .Y(new_n8138));
  AOI221xp5_ASAP7_75t_L     g07882(.A1(new_n7861), .A2(new_n7873), .B1(new_n8138), .B2(new_n8137), .C(new_n7858), .Y(new_n8139));
  A2O1A1O1Ixp25_ASAP7_75t_L g07883(.A1(new_n7557), .A2(new_n7559), .B(new_n7863), .C(new_n7873), .D(new_n7858), .Y(new_n8140));
  XOR2x2_ASAP7_75t_L        g07884(.A(new_n8131), .B(new_n8130), .Y(new_n8141));
  NOR2xp33_ASAP7_75t_L      g07885(.A(new_n8136), .B(new_n8141), .Y(new_n8142));
  INVx1_ASAP7_75t_L         g07886(.A(new_n8138), .Y(new_n8143));
  NOR3xp33_ASAP7_75t_L      g07887(.A(new_n8142), .B(new_n8143), .C(new_n8140), .Y(new_n8144));
  NOR3xp33_ASAP7_75t_L      g07888(.A(new_n8144), .B(new_n8139), .C(new_n7924), .Y(new_n8145));
  OA21x2_ASAP7_75t_L        g07889(.A1(new_n8139), .A2(new_n8144), .B(new_n7924), .Y(new_n8146));
  OAI221xp5_ASAP7_75t_L     g07890(.A1(new_n7913), .A2(new_n7881), .B1(new_n8145), .B2(new_n8146), .C(new_n7916), .Y(new_n8147));
  MAJIxp5_ASAP7_75t_L       g07891(.A(new_n7881), .B(new_n7914), .C(new_n7871), .Y(new_n8148));
  OR3x1_ASAP7_75t_L         g07892(.A(new_n8144), .B(new_n7924), .C(new_n8139), .Y(new_n8149));
  OAI21xp33_ASAP7_75t_L     g07893(.A1(new_n8139), .A2(new_n8144), .B(new_n7924), .Y(new_n8150));
  NAND3xp33_ASAP7_75t_L     g07894(.A(new_n8148), .B(new_n8149), .C(new_n8150), .Y(new_n8151));
  AOI22xp33_ASAP7_75t_L     g07895(.A1(new_n344), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n370), .Y(new_n8152));
  OAI221xp5_ASAP7_75t_L     g07896(.A1(new_n429), .A2(new_n6830), .B1(new_n366), .B2(new_n7323), .C(new_n8152), .Y(new_n8153));
  XNOR2x2_ASAP7_75t_L       g07897(.A(\a[5] ), .B(new_n8153), .Y(new_n8154));
  NAND3xp33_ASAP7_75t_L     g07898(.A(new_n8151), .B(new_n8147), .C(new_n8154), .Y(new_n8155));
  AO21x2_ASAP7_75t_L        g07899(.A1(new_n8147), .A2(new_n8151), .B(new_n8154), .Y(new_n8156));
  AOI21xp33_ASAP7_75t_L     g07900(.A1(new_n8156), .A2(new_n8155), .B(new_n7910), .Y(new_n8157));
  AND3x1_ASAP7_75t_L        g07901(.A(new_n7910), .B(new_n8156), .C(new_n8155), .Y(new_n8158));
  NOR3xp33_ASAP7_75t_L      g07902(.A(new_n8158), .B(new_n8157), .C(new_n7909), .Y(new_n8159));
  INVx1_ASAP7_75t_L         g07903(.A(new_n8159), .Y(new_n8160));
  OAI21xp33_ASAP7_75t_L     g07904(.A1(new_n8157), .A2(new_n8158), .B(new_n7909), .Y(new_n8161));
  NAND2xp33_ASAP7_75t_L     g07905(.A(new_n8161), .B(new_n8160), .Y(new_n8162));
  XOR2x2_ASAP7_75t_L        g07906(.A(new_n8162), .B(new_n7898), .Y(\f[52] ));
  NOR2xp33_ASAP7_75t_L      g07907(.A(\b[52] ), .B(\b[53] ), .Y(new_n8164));
  INVx1_ASAP7_75t_L         g07908(.A(\b[53] ), .Y(new_n8165));
  NOR2xp33_ASAP7_75t_L      g07909(.A(new_n7900), .B(new_n8165), .Y(new_n8166));
  NOR2xp33_ASAP7_75t_L      g07910(.A(new_n8164), .B(new_n8166), .Y(new_n8167));
  INVx1_ASAP7_75t_L         g07911(.A(new_n8167), .Y(new_n8168));
  O2A1O1Ixp33_ASAP7_75t_L   g07912(.A1(new_n7616), .A2(new_n7900), .B(new_n7903), .C(new_n8168), .Y(new_n8169));
  INVx1_ASAP7_75t_L         g07913(.A(new_n8169), .Y(new_n8170));
  O2A1O1Ixp33_ASAP7_75t_L   g07914(.A1(new_n7617), .A2(new_n7620), .B(new_n7902), .C(new_n7901), .Y(new_n8171));
  NAND2xp33_ASAP7_75t_L     g07915(.A(new_n8168), .B(new_n8171), .Y(new_n8172));
  AND2x2_ASAP7_75t_L        g07916(.A(new_n8172), .B(new_n8170), .Y(new_n8173));
  INVx1_ASAP7_75t_L         g07917(.A(new_n8173), .Y(new_n8174));
  AOI22xp33_ASAP7_75t_L     g07918(.A1(\b[51] ), .A2(new_n282), .B1(\b[53] ), .B2(new_n303), .Y(new_n8175));
  OAI221xp5_ASAP7_75t_L     g07919(.A1(new_n291), .A2(new_n7900), .B1(new_n268), .B2(new_n8174), .C(new_n8175), .Y(new_n8176));
  XNOR2x2_ASAP7_75t_L       g07920(.A(\a[2] ), .B(new_n8176), .Y(new_n8177));
  AND3x1_ASAP7_75t_L        g07921(.A(new_n8151), .B(new_n8147), .C(new_n8154), .Y(new_n8178));
  AOI21xp33_ASAP7_75t_L     g07922(.A1(new_n8151), .A2(new_n8147), .B(new_n8154), .Y(new_n8179));
  NOR2xp33_ASAP7_75t_L      g07923(.A(new_n8179), .B(new_n8178), .Y(new_n8180));
  NAND2xp33_ASAP7_75t_L     g07924(.A(new_n8147), .B(new_n8151), .Y(new_n8181));
  INVx1_ASAP7_75t_L         g07925(.A(new_n8181), .Y(new_n8182));
  INVx1_ASAP7_75t_L         g07926(.A(new_n8154), .Y(new_n8183));
  NAND2xp33_ASAP7_75t_L     g07927(.A(new_n8183), .B(new_n8182), .Y(new_n8184));
  NAND2xp33_ASAP7_75t_L     g07928(.A(\b[46] ), .B(new_n447), .Y(new_n8185));
  INVx1_ASAP7_75t_L         g07929(.A(new_n6820), .Y(new_n8186));
  NAND2xp33_ASAP7_75t_L     g07930(.A(new_n441), .B(new_n8186), .Y(new_n8187));
  AOI22xp33_ASAP7_75t_L     g07931(.A1(new_n444), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n471), .Y(new_n8188));
  AND4x1_ASAP7_75t_L        g07932(.A(new_n8188), .B(new_n8187), .C(new_n8185), .D(\a[8] ), .Y(new_n8189));
  AOI31xp33_ASAP7_75t_L     g07933(.A1(new_n8187), .A2(new_n8185), .A3(new_n8188), .B(\a[8] ), .Y(new_n8190));
  NOR2xp33_ASAP7_75t_L      g07934(.A(new_n8190), .B(new_n8189), .Y(new_n8191));
  NAND2xp33_ASAP7_75t_L     g07935(.A(new_n8070), .B(new_n8074), .Y(new_n8192));
  MAJIxp5_ASAP7_75t_L       g07936(.A(new_n8080), .B(new_n8192), .C(new_n8077), .Y(new_n8193));
  NOR2xp33_ASAP7_75t_L      g07937(.A(new_n3180), .B(new_n1699), .Y(new_n8194));
  INVx1_ASAP7_75t_L         g07938(.A(new_n8194), .Y(new_n8195));
  NAND3xp33_ASAP7_75t_L     g07939(.A(new_n3210), .B(new_n1695), .C(new_n3213), .Y(new_n8196));
  AOI22xp33_ASAP7_75t_L     g07940(.A1(new_n1704), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1837), .Y(new_n8197));
  NAND4xp25_ASAP7_75t_L     g07941(.A(new_n8196), .B(\a[23] ), .C(new_n8195), .D(new_n8197), .Y(new_n8198));
  AOI31xp33_ASAP7_75t_L     g07942(.A1(new_n8196), .A2(new_n8195), .A3(new_n8197), .B(\a[23] ), .Y(new_n8199));
  INVx1_ASAP7_75t_L         g07943(.A(new_n8199), .Y(new_n8200));
  NAND2xp33_ASAP7_75t_L     g07944(.A(new_n8198), .B(new_n8200), .Y(new_n8201));
  INVx1_ASAP7_75t_L         g07945(.A(new_n8201), .Y(new_n8202));
  NOR3xp33_ASAP7_75t_L      g07946(.A(new_n7787), .B(new_n7788), .C(new_n7785), .Y(new_n8203));
  A2O1A1O1Ixp25_ASAP7_75t_L g07947(.A1(new_n7792), .A2(new_n7793), .B(new_n8203), .C(new_n8073), .D(new_n8065), .Y(new_n8204));
  AOI22xp33_ASAP7_75t_L     g07948(.A1(new_n2114), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n2259), .Y(new_n8205));
  OAI221xp5_ASAP7_75t_L     g07949(.A1(new_n2109), .A2(new_n2666), .B1(new_n2257), .B2(new_n2695), .C(new_n8205), .Y(new_n8206));
  XNOR2x2_ASAP7_75t_L       g07950(.A(\a[26] ), .B(new_n8206), .Y(new_n8207));
  INVx1_ASAP7_75t_L         g07951(.A(new_n8207), .Y(new_n8208));
  NAND2xp33_ASAP7_75t_L     g07952(.A(new_n8045), .B(new_n8049), .Y(new_n8209));
  MAJIxp5_ASAP7_75t_L       g07953(.A(new_n7929), .B(new_n8052), .C(new_n8209), .Y(new_n8210));
  AOI22xp33_ASAP7_75t_L     g07954(.A1(new_n2552), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n2736), .Y(new_n8211));
  OAI221xp5_ASAP7_75t_L     g07955(.A1(new_n2547), .A2(new_n2067), .B1(new_n2734), .B2(new_n2355), .C(new_n8211), .Y(new_n8212));
  XNOR2x2_ASAP7_75t_L       g07956(.A(\a[29] ), .B(new_n8212), .Y(new_n8213));
  O2A1O1Ixp33_ASAP7_75t_L   g07957(.A1(new_n7765), .A2(new_n7462), .B(new_n7762), .C(new_n7931), .Y(new_n8214));
  AOI22xp33_ASAP7_75t_L     g07958(.A1(new_n3029), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n3258), .Y(new_n8215));
  OAI221xp5_ASAP7_75t_L     g07959(.A1(new_n3024), .A2(new_n1774), .B1(new_n3256), .B2(new_n1915), .C(new_n8215), .Y(new_n8216));
  XNOR2x2_ASAP7_75t_L       g07960(.A(new_n3015), .B(new_n8216), .Y(new_n8217));
  INVx1_ASAP7_75t_L         g07961(.A(new_n8217), .Y(new_n8218));
  INVx1_ASAP7_75t_L         g07962(.A(new_n8022), .Y(new_n8219));
  NAND3xp33_ASAP7_75t_L     g07963(.A(new_n8019), .B(new_n8014), .C(new_n8219), .Y(new_n8220));
  A2O1A1Ixp33_ASAP7_75t_L   g07964(.A1(new_n8024), .A2(new_n8023), .B(new_n8026), .C(new_n8220), .Y(new_n8221));
  AOI22xp33_ASAP7_75t_L     g07965(.A1(new_n4283), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n4512), .Y(new_n8222));
  OAI221xp5_ASAP7_75t_L     g07966(.A1(new_n4277), .A2(new_n1030), .B1(new_n4499), .B2(new_n1209), .C(new_n8222), .Y(new_n8223));
  XNOR2x2_ASAP7_75t_L       g07967(.A(\a[38] ), .B(new_n8223), .Y(new_n8224));
  INVx1_ASAP7_75t_L         g07968(.A(new_n8224), .Y(new_n8225));
  NAND2xp33_ASAP7_75t_L     g07969(.A(new_n7727), .B(new_n7728), .Y(new_n8226));
  NOR2xp33_ASAP7_75t_L      g07970(.A(new_n7664), .B(new_n7938), .Y(new_n8227));
  A2O1A1O1Ixp25_ASAP7_75t_L g07971(.A1(new_n7661), .A2(new_n8226), .B(new_n8227), .C(new_n8007), .D(new_n8018), .Y(new_n8228));
  AOI22xp33_ASAP7_75t_L     g07972(.A1(new_n5624), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n5901), .Y(new_n8229));
  OAI221xp5_ASAP7_75t_L     g07973(.A1(new_n5900), .A2(new_n617), .B1(new_n5892), .B2(new_n685), .C(new_n8229), .Y(new_n8230));
  XNOR2x2_ASAP7_75t_L       g07974(.A(\a[44] ), .B(new_n8230), .Y(new_n8231));
  NAND3xp33_ASAP7_75t_L     g07975(.A(new_n7977), .B(new_n7971), .C(new_n7984), .Y(new_n8232));
  AOI22xp33_ASAP7_75t_L     g07976(.A1(new_n6376), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n6648), .Y(new_n8233));
  OAI221xp5_ASAP7_75t_L     g07977(.A1(new_n6646), .A2(new_n420), .B1(new_n6636), .B2(new_n494), .C(new_n8233), .Y(new_n8234));
  XNOR2x2_ASAP7_75t_L       g07978(.A(new_n6371), .B(new_n8234), .Y(new_n8235));
  O2A1O1Ixp33_ASAP7_75t_L   g07979(.A1(new_n7943), .A2(new_n7692), .B(new_n7967), .C(new_n7976), .Y(new_n8236));
  INVx1_ASAP7_75t_L         g07980(.A(new_n7108), .Y(new_n8237));
  NAND2xp33_ASAP7_75t_L     g07981(.A(\b[4] ), .B(new_n7115), .Y(new_n8238));
  AOI22xp33_ASAP7_75t_L     g07982(.A1(new_n7111), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n7391), .Y(new_n8239));
  OAI311xp33_ASAP7_75t_L    g07983(.A1(new_n357), .A2(new_n8237), .A3(new_n358), .B1(new_n8238), .C1(new_n8239), .Y(new_n8240));
  NOR2xp33_ASAP7_75t_L      g07984(.A(new_n7106), .B(new_n8240), .Y(new_n8241));
  AND2x2_ASAP7_75t_L        g07985(.A(new_n7106), .B(new_n8240), .Y(new_n8242));
  NAND3xp33_ASAP7_75t_L     g07986(.A(new_n7951), .B(new_n7953), .C(new_n7955), .Y(new_n8243));
  OAI21xp33_ASAP7_75t_L     g07987(.A1(new_n261), .A2(new_n8243), .B(new_n7964), .Y(new_n8244));
  AOI21xp33_ASAP7_75t_L     g07988(.A1(new_n7958), .A2(new_n269), .B(new_n8244), .Y(new_n8245));
  NAND2xp33_ASAP7_75t_L     g07989(.A(\b[2] ), .B(new_n7960), .Y(new_n8246));
  NAND3xp33_ASAP7_75t_L     g07990(.A(new_n7669), .B(new_n7956), .C(new_n7962), .Y(new_n8247));
  OAI221xp5_ASAP7_75t_L     g07991(.A1(new_n258), .A2(new_n8247), .B1(new_n280), .B2(new_n7957), .C(new_n8246), .Y(new_n8248));
  AOI21xp33_ASAP7_75t_L     g07992(.A1(new_n7963), .A2(\b[1] ), .B(new_n8248), .Y(new_n8249));
  A2O1A1Ixp33_ASAP7_75t_L   g07993(.A1(new_n7674), .A2(new_n8245), .B(new_n7954), .C(new_n8249), .Y(new_n8250));
  O2A1O1Ixp33_ASAP7_75t_L   g07994(.A1(new_n258), .A2(new_n7669), .B(new_n8245), .C(new_n7954), .Y(new_n8251));
  A2O1A1Ixp33_ASAP7_75t_L   g07995(.A1(\b[1] ), .A2(new_n7963), .B(new_n8248), .C(new_n8251), .Y(new_n8252));
  AOI211xp5_ASAP7_75t_L     g07996(.A1(new_n8252), .A2(new_n8250), .B(new_n8241), .C(new_n8242), .Y(new_n8253));
  OAI211xp5_ASAP7_75t_L     g07997(.A1(new_n8241), .A2(new_n8242), .B(new_n8252), .C(new_n8250), .Y(new_n8254));
  INVx1_ASAP7_75t_L         g07998(.A(new_n8254), .Y(new_n8255));
  OAI21xp33_ASAP7_75t_L     g07999(.A1(new_n8253), .A2(new_n8255), .B(new_n8236), .Y(new_n8256));
  INVx1_ASAP7_75t_L         g08000(.A(new_n7943), .Y(new_n8257));
  A2O1A1Ixp33_ASAP7_75t_L   g08001(.A1(new_n7682), .A2(new_n8257), .B(new_n7975), .C(new_n7970), .Y(new_n8258));
  NOR2xp33_ASAP7_75t_L      g08002(.A(new_n8241), .B(new_n8242), .Y(new_n8259));
  NAND2xp33_ASAP7_75t_L     g08003(.A(new_n8250), .B(new_n8252), .Y(new_n8260));
  NAND2xp33_ASAP7_75t_L     g08004(.A(new_n8259), .B(new_n8260), .Y(new_n8261));
  NAND3xp33_ASAP7_75t_L     g08005(.A(new_n8258), .B(new_n8261), .C(new_n8254), .Y(new_n8262));
  AO21x2_ASAP7_75t_L        g08006(.A1(new_n8256), .A2(new_n8262), .B(new_n8235), .Y(new_n8263));
  NAND3xp33_ASAP7_75t_L     g08007(.A(new_n8262), .B(new_n8256), .C(new_n8235), .Y(new_n8264));
  NAND2xp33_ASAP7_75t_L     g08008(.A(new_n8264), .B(new_n8263), .Y(new_n8265));
  A2O1A1O1Ixp25_ASAP7_75t_L g08009(.A1(new_n7985), .A2(new_n7981), .B(new_n7987), .C(new_n8232), .D(new_n8265), .Y(new_n8266));
  A2O1A1Ixp33_ASAP7_75t_L   g08010(.A1(new_n7985), .A2(new_n7981), .B(new_n7987), .C(new_n8232), .Y(new_n8267));
  AOI21xp33_ASAP7_75t_L     g08011(.A1(new_n8264), .A2(new_n8263), .B(new_n8267), .Y(new_n8268));
  OAI21xp33_ASAP7_75t_L     g08012(.A1(new_n8268), .A2(new_n8266), .B(new_n8231), .Y(new_n8269));
  INVx1_ASAP7_75t_L         g08013(.A(new_n8231), .Y(new_n8270));
  INVx1_ASAP7_75t_L         g08014(.A(new_n8232), .Y(new_n8271));
  AND2x2_ASAP7_75t_L        g08015(.A(new_n8264), .B(new_n8263), .Y(new_n8272));
  A2O1A1Ixp33_ASAP7_75t_L   g08016(.A1(new_n7991), .A2(new_n7989), .B(new_n8271), .C(new_n8272), .Y(new_n8273));
  A2O1A1O1Ixp25_ASAP7_75t_L g08017(.A1(new_n7708), .A2(new_n7700), .B(new_n7986), .C(new_n7989), .D(new_n8271), .Y(new_n8274));
  NAND2xp33_ASAP7_75t_L     g08018(.A(new_n8265), .B(new_n8274), .Y(new_n8275));
  NAND3xp33_ASAP7_75t_L     g08019(.A(new_n8273), .B(new_n8270), .C(new_n8275), .Y(new_n8276));
  OAI211xp5_ASAP7_75t_L     g08020(.A1(new_n7718), .A2(new_n7715), .B(new_n7717), .C(new_n8004), .Y(new_n8277));
  NAND4xp25_ASAP7_75t_L     g08021(.A(new_n8276), .B(new_n8277), .C(new_n8003), .D(new_n8269), .Y(new_n8278));
  AO22x1_ASAP7_75t_L        g08022(.A1(new_n8003), .A2(new_n8277), .B1(new_n8269), .B2(new_n8276), .Y(new_n8279));
  AOI22xp33_ASAP7_75t_L     g08023(.A1(new_n4920), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n5167), .Y(new_n8280));
  OAI221xp5_ASAP7_75t_L     g08024(.A1(new_n5154), .A2(new_n784), .B1(new_n5158), .B2(new_n875), .C(new_n8280), .Y(new_n8281));
  XNOR2x2_ASAP7_75t_L       g08025(.A(\a[41] ), .B(new_n8281), .Y(new_n8282));
  NAND3xp33_ASAP7_75t_L     g08026(.A(new_n8279), .B(new_n8278), .C(new_n8282), .Y(new_n8283));
  AND4x1_ASAP7_75t_L        g08027(.A(new_n8277), .B(new_n8276), .C(new_n8269), .D(new_n8003), .Y(new_n8284));
  AOI22xp33_ASAP7_75t_L     g08028(.A1(new_n8277), .A2(new_n8003), .B1(new_n8269), .B2(new_n8276), .Y(new_n8285));
  INVx1_ASAP7_75t_L         g08029(.A(new_n8282), .Y(new_n8286));
  OAI21xp33_ASAP7_75t_L     g08030(.A1(new_n8285), .A2(new_n8284), .B(new_n8286), .Y(new_n8287));
  AOI21xp33_ASAP7_75t_L     g08031(.A1(new_n8287), .A2(new_n8283), .B(new_n8228), .Y(new_n8288));
  A2O1A1Ixp33_ASAP7_75t_L   g08032(.A1(new_n7725), .A2(new_n8016), .B(new_n8017), .C(new_n8013), .Y(new_n8289));
  NAND2xp33_ASAP7_75t_L     g08033(.A(new_n8287), .B(new_n8283), .Y(new_n8290));
  NOR2xp33_ASAP7_75t_L      g08034(.A(new_n8290), .B(new_n8289), .Y(new_n8291));
  OAI21xp33_ASAP7_75t_L     g08035(.A1(new_n8288), .A2(new_n8291), .B(new_n8225), .Y(new_n8292));
  A2O1A1Ixp33_ASAP7_75t_L   g08036(.A1(new_n8007), .A2(new_n7939), .B(new_n8018), .C(new_n8290), .Y(new_n8293));
  AND2x2_ASAP7_75t_L        g08037(.A(new_n8287), .B(new_n8283), .Y(new_n8294));
  NAND2xp33_ASAP7_75t_L     g08038(.A(new_n8228), .B(new_n8294), .Y(new_n8295));
  NAND3xp33_ASAP7_75t_L     g08039(.A(new_n8295), .B(new_n8293), .C(new_n8224), .Y(new_n8296));
  NAND3xp33_ASAP7_75t_L     g08040(.A(new_n8221), .B(new_n8292), .C(new_n8296), .Y(new_n8297));
  AND3x1_ASAP7_75t_L        g08041(.A(new_n8019), .B(new_n8014), .C(new_n8022), .Y(new_n8298));
  AOI21xp33_ASAP7_75t_L     g08042(.A1(new_n8019), .A2(new_n8014), .B(new_n8022), .Y(new_n8299));
  NOR2xp33_ASAP7_75t_L      g08043(.A(new_n8299), .B(new_n8298), .Y(new_n8300));
  AOI21xp33_ASAP7_75t_L     g08044(.A1(new_n8295), .A2(new_n8293), .B(new_n8224), .Y(new_n8301));
  NOR3xp33_ASAP7_75t_L      g08045(.A(new_n8225), .B(new_n8291), .C(new_n8288), .Y(new_n8302));
  OAI221xp5_ASAP7_75t_L     g08046(.A1(new_n8300), .A2(new_n8026), .B1(new_n8302), .B2(new_n8301), .C(new_n8220), .Y(new_n8303));
  AOI22xp33_ASAP7_75t_L     g08047(.A1(new_n3633), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n3858), .Y(new_n8304));
  OAI221xp5_ASAP7_75t_L     g08048(.A1(new_n3853), .A2(new_n1432), .B1(new_n3856), .B2(new_n1547), .C(new_n8304), .Y(new_n8305));
  XNOR2x2_ASAP7_75t_L       g08049(.A(\a[35] ), .B(new_n8305), .Y(new_n8306));
  AO21x2_ASAP7_75t_L        g08050(.A1(new_n8303), .A2(new_n8297), .B(new_n8306), .Y(new_n8307));
  NAND3xp33_ASAP7_75t_L     g08051(.A(new_n8297), .B(new_n8303), .C(new_n8306), .Y(new_n8308));
  OAI211xp5_ASAP7_75t_L     g08052(.A1(new_n7748), .A2(new_n7745), .B(new_n8037), .C(new_n7749), .Y(new_n8309));
  NAND4xp25_ASAP7_75t_L     g08053(.A(new_n8307), .B(new_n8309), .C(new_n8036), .D(new_n8308), .Y(new_n8310));
  AO22x1_ASAP7_75t_L        g08054(.A1(new_n8036), .A2(new_n8309), .B1(new_n8307), .B2(new_n8308), .Y(new_n8311));
  AOI21xp33_ASAP7_75t_L     g08055(.A1(new_n8311), .A2(new_n8310), .B(new_n8218), .Y(new_n8312));
  AND4x1_ASAP7_75t_L        g08056(.A(new_n8307), .B(new_n8036), .C(new_n8309), .D(new_n8308), .Y(new_n8313));
  AOI22xp33_ASAP7_75t_L     g08057(.A1(new_n8309), .A2(new_n8036), .B1(new_n8307), .B2(new_n8308), .Y(new_n8314));
  NOR3xp33_ASAP7_75t_L      g08058(.A(new_n8313), .B(new_n8314), .C(new_n8217), .Y(new_n8315));
  NOR2xp33_ASAP7_75t_L      g08059(.A(new_n8315), .B(new_n8312), .Y(new_n8316));
  O2A1O1Ixp33_ASAP7_75t_L   g08060(.A1(new_n8047), .A2(new_n8214), .B(new_n8039), .C(new_n8316), .Y(new_n8317));
  OAI21xp33_ASAP7_75t_L     g08061(.A1(new_n8314), .A2(new_n8313), .B(new_n8217), .Y(new_n8318));
  NAND3xp33_ASAP7_75t_L     g08062(.A(new_n8311), .B(new_n8218), .C(new_n8310), .Y(new_n8319));
  NAND2xp33_ASAP7_75t_L     g08063(.A(new_n8319), .B(new_n8318), .Y(new_n8320));
  AOI211xp5_ASAP7_75t_L     g08064(.A1(new_n8048), .A2(new_n8054), .B(new_n8046), .C(new_n8320), .Y(new_n8321));
  OAI21xp33_ASAP7_75t_L     g08065(.A1(new_n8317), .A2(new_n8321), .B(new_n8213), .Y(new_n8322));
  INVx1_ASAP7_75t_L         g08066(.A(new_n8213), .Y(new_n8323));
  A2O1A1Ixp33_ASAP7_75t_L   g08067(.A1(new_n8048), .A2(new_n8054), .B(new_n8046), .C(new_n8320), .Y(new_n8324));
  A2O1A1O1Ixp25_ASAP7_75t_L g08068(.A1(new_n7763), .A2(new_n7762), .B(new_n7931), .C(new_n8043), .D(new_n8046), .Y(new_n8325));
  NAND2xp33_ASAP7_75t_L     g08069(.A(new_n8316), .B(new_n8325), .Y(new_n8326));
  NAND3xp33_ASAP7_75t_L     g08070(.A(new_n8326), .B(new_n8324), .C(new_n8323), .Y(new_n8327));
  NAND3xp33_ASAP7_75t_L     g08071(.A(new_n8210), .B(new_n8322), .C(new_n8327), .Y(new_n8328));
  XNOR2x2_ASAP7_75t_L       g08072(.A(new_n8054), .B(new_n8044), .Y(new_n8329));
  MAJIxp5_ASAP7_75t_L       g08073(.A(new_n8061), .B(new_n8329), .C(new_n8058), .Y(new_n8330));
  NAND2xp33_ASAP7_75t_L     g08074(.A(new_n8327), .B(new_n8322), .Y(new_n8331));
  NAND2xp33_ASAP7_75t_L     g08075(.A(new_n8330), .B(new_n8331), .Y(new_n8332));
  AOI21xp33_ASAP7_75t_L     g08076(.A1(new_n8332), .A2(new_n8328), .B(new_n8208), .Y(new_n8333));
  NOR2xp33_ASAP7_75t_L      g08077(.A(new_n8330), .B(new_n8331), .Y(new_n8334));
  AOI21xp33_ASAP7_75t_L     g08078(.A1(new_n8327), .A2(new_n8322), .B(new_n8210), .Y(new_n8335));
  NOR3xp33_ASAP7_75t_L      g08079(.A(new_n8334), .B(new_n8335), .C(new_n8207), .Y(new_n8336));
  NOR3xp33_ASAP7_75t_L      g08080(.A(new_n8204), .B(new_n8333), .C(new_n8336), .Y(new_n8337));
  OAI21xp33_ASAP7_75t_L     g08081(.A1(new_n8335), .A2(new_n8334), .B(new_n8207), .Y(new_n8338));
  NAND3xp33_ASAP7_75t_L     g08082(.A(new_n8332), .B(new_n8328), .C(new_n8208), .Y(new_n8339));
  AOI221xp5_ASAP7_75t_L     g08083(.A1(new_n8073), .A2(new_n8071), .B1(new_n8339), .B2(new_n8338), .C(new_n8065), .Y(new_n8340));
  OAI21xp33_ASAP7_75t_L     g08084(.A1(new_n8340), .A2(new_n8337), .B(new_n8202), .Y(new_n8341));
  AO21x2_ASAP7_75t_L        g08085(.A1(new_n8073), .A2(new_n8071), .B(new_n8065), .Y(new_n8342));
  NAND3xp33_ASAP7_75t_L     g08086(.A(new_n8342), .B(new_n8338), .C(new_n8339), .Y(new_n8343));
  OAI21xp33_ASAP7_75t_L     g08087(.A1(new_n8333), .A2(new_n8336), .B(new_n8204), .Y(new_n8344));
  NAND3xp33_ASAP7_75t_L     g08088(.A(new_n8343), .B(new_n8201), .C(new_n8344), .Y(new_n8345));
  NAND3xp33_ASAP7_75t_L     g08089(.A(new_n8193), .B(new_n8341), .C(new_n8345), .Y(new_n8346));
  INVx1_ASAP7_75t_L         g08090(.A(new_n8077), .Y(new_n8347));
  AND3x1_ASAP7_75t_L        g08091(.A(new_n8074), .B(new_n8070), .C(new_n8347), .Y(new_n8348));
  O2A1O1Ixp33_ASAP7_75t_L   g08092(.A1(new_n8083), .A2(new_n8082), .B(new_n8084), .C(new_n8348), .Y(new_n8349));
  AOI21xp33_ASAP7_75t_L     g08093(.A1(new_n8343), .A2(new_n8344), .B(new_n8201), .Y(new_n8350));
  NOR3xp33_ASAP7_75t_L      g08094(.A(new_n8337), .B(new_n8340), .C(new_n8202), .Y(new_n8351));
  OAI21xp33_ASAP7_75t_L     g08095(.A1(new_n8350), .A2(new_n8351), .B(new_n8349), .Y(new_n8352));
  NOR2xp33_ASAP7_75t_L      g08096(.A(new_n3584), .B(new_n1373), .Y(new_n8353));
  INVx1_ASAP7_75t_L         g08097(.A(new_n8353), .Y(new_n8354));
  NAND2xp33_ASAP7_75t_L     g08098(.A(new_n1365), .B(new_n3811), .Y(new_n8355));
  AOI22xp33_ASAP7_75t_L     g08099(.A1(new_n1360), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1581), .Y(new_n8356));
  AND4x1_ASAP7_75t_L        g08100(.A(new_n8356), .B(new_n8355), .C(new_n8354), .D(\a[20] ), .Y(new_n8357));
  AOI31xp33_ASAP7_75t_L     g08101(.A1(new_n8355), .A2(new_n8354), .A3(new_n8356), .B(\a[20] ), .Y(new_n8358));
  NOR2xp33_ASAP7_75t_L      g08102(.A(new_n8358), .B(new_n8357), .Y(new_n8359));
  NAND3xp33_ASAP7_75t_L     g08103(.A(new_n8346), .B(new_n8352), .C(new_n8359), .Y(new_n8360));
  NOR3xp33_ASAP7_75t_L      g08104(.A(new_n8349), .B(new_n8350), .C(new_n8351), .Y(new_n8361));
  AOI221xp5_ASAP7_75t_L     g08105(.A1(new_n8090), .A2(new_n8084), .B1(new_n8341), .B2(new_n8345), .C(new_n8348), .Y(new_n8362));
  INVx1_ASAP7_75t_L         g08106(.A(new_n8359), .Y(new_n8363));
  OAI21xp33_ASAP7_75t_L     g08107(.A1(new_n8362), .A2(new_n8361), .B(new_n8363), .Y(new_n8364));
  NAND2xp33_ASAP7_75t_L     g08108(.A(new_n8085), .B(new_n8081), .Y(new_n8365));
  NOR2xp33_ASAP7_75t_L      g08109(.A(new_n8088), .B(new_n8365), .Y(new_n8366));
  O2A1O1Ixp33_ASAP7_75t_L   g08110(.A1(new_n8098), .A2(new_n8099), .B(new_n8101), .C(new_n8366), .Y(new_n8367));
  NAND3xp33_ASAP7_75t_L     g08111(.A(new_n8367), .B(new_n8364), .C(new_n8360), .Y(new_n8368));
  INVx1_ASAP7_75t_L         g08112(.A(new_n8365), .Y(new_n8369));
  NAND2xp33_ASAP7_75t_L     g08113(.A(new_n8364), .B(new_n8360), .Y(new_n8370));
  A2O1A1Ixp33_ASAP7_75t_L   g08114(.A1(new_n8093), .A2(new_n8369), .B(new_n8109), .C(new_n8370), .Y(new_n8371));
  NAND2xp33_ASAP7_75t_L     g08115(.A(\b[37] ), .B(new_n1080), .Y(new_n8372));
  NAND2xp33_ASAP7_75t_L     g08116(.A(new_n1073), .B(new_n4640), .Y(new_n8373));
  AOI22xp33_ASAP7_75t_L     g08117(.A1(new_n1076), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1253), .Y(new_n8374));
  NAND4xp25_ASAP7_75t_L     g08118(.A(new_n8373), .B(\a[17] ), .C(new_n8372), .D(new_n8374), .Y(new_n8375));
  NAND2xp33_ASAP7_75t_L     g08119(.A(new_n8374), .B(new_n8373), .Y(new_n8376));
  A2O1A1Ixp33_ASAP7_75t_L   g08120(.A1(\b[37] ), .A2(new_n1080), .B(new_n8376), .C(new_n1071), .Y(new_n8377));
  NAND2xp33_ASAP7_75t_L     g08121(.A(new_n8375), .B(new_n8377), .Y(new_n8378));
  INVx1_ASAP7_75t_L         g08122(.A(new_n8378), .Y(new_n8379));
  NAND3xp33_ASAP7_75t_L     g08123(.A(new_n8371), .B(new_n8368), .C(new_n8379), .Y(new_n8380));
  MAJIxp5_ASAP7_75t_L       g08124(.A(new_n8108), .B(new_n8365), .C(new_n8088), .Y(new_n8381));
  NOR2xp33_ASAP7_75t_L      g08125(.A(new_n8370), .B(new_n8381), .Y(new_n8382));
  AOI21xp33_ASAP7_75t_L     g08126(.A1(new_n8364), .A2(new_n8360), .B(new_n8367), .Y(new_n8383));
  OAI21xp33_ASAP7_75t_L     g08127(.A1(new_n8383), .A2(new_n8382), .B(new_n8378), .Y(new_n8384));
  NAND3xp33_ASAP7_75t_L     g08128(.A(new_n8097), .B(new_n8102), .C(new_n8110), .Y(new_n8385));
  NAND4xp25_ASAP7_75t_L     g08129(.A(new_n8115), .B(new_n8385), .C(new_n8384), .D(new_n8380), .Y(new_n8386));
  NAND2xp33_ASAP7_75t_L     g08130(.A(new_n8384), .B(new_n8380), .Y(new_n8387));
  A2O1A1Ixp33_ASAP7_75t_L   g08131(.A1(new_n8111), .A2(new_n8106), .B(new_n8112), .C(new_n8385), .Y(new_n8388));
  NAND2xp33_ASAP7_75t_L     g08132(.A(new_n8388), .B(new_n8387), .Y(new_n8389));
  NAND2xp33_ASAP7_75t_L     g08133(.A(\b[40] ), .B(new_n815), .Y(new_n8390));
  NAND3xp33_ASAP7_75t_L     g08134(.A(new_n5326), .B(new_n5324), .C(new_n808), .Y(new_n8391));
  AOI22xp33_ASAP7_75t_L     g08135(.A1(new_n811), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n900), .Y(new_n8392));
  AND4x1_ASAP7_75t_L        g08136(.A(new_n8392), .B(new_n8391), .C(new_n8390), .D(\a[14] ), .Y(new_n8393));
  AOI31xp33_ASAP7_75t_L     g08137(.A1(new_n8391), .A2(new_n8390), .A3(new_n8392), .B(\a[14] ), .Y(new_n8394));
  NOR2xp33_ASAP7_75t_L      g08138(.A(new_n8394), .B(new_n8393), .Y(new_n8395));
  NAND3xp33_ASAP7_75t_L     g08139(.A(new_n8386), .B(new_n8389), .C(new_n8395), .Y(new_n8396));
  NOR2xp33_ASAP7_75t_L      g08140(.A(new_n8388), .B(new_n8387), .Y(new_n8397));
  NOR3xp33_ASAP7_75t_L      g08141(.A(new_n8382), .B(new_n8383), .C(new_n8378), .Y(new_n8398));
  AOI21xp33_ASAP7_75t_L     g08142(.A1(new_n8371), .A2(new_n8368), .B(new_n8379), .Y(new_n8399));
  OA21x2_ASAP7_75t_L        g08143(.A1(new_n8398), .A2(new_n8399), .B(new_n8388), .Y(new_n8400));
  INVx1_ASAP7_75t_L         g08144(.A(new_n8395), .Y(new_n8401));
  OAI21xp33_ASAP7_75t_L     g08145(.A1(new_n8397), .A2(new_n8400), .B(new_n8401), .Y(new_n8402));
  NOR3xp33_ASAP7_75t_L      g08146(.A(new_n8124), .B(new_n8125), .C(new_n8122), .Y(new_n8403));
  AOI21xp33_ASAP7_75t_L     g08147(.A1(new_n8130), .A2(new_n8131), .B(new_n8403), .Y(new_n8404));
  NAND3xp33_ASAP7_75t_L     g08148(.A(new_n8404), .B(new_n8402), .C(new_n8396), .Y(new_n8405));
  NAND2xp33_ASAP7_75t_L     g08149(.A(new_n8396), .B(new_n8402), .Y(new_n8406));
  A2O1A1Ixp33_ASAP7_75t_L   g08150(.A1(new_n8130), .A2(new_n8131), .B(new_n8403), .C(new_n8406), .Y(new_n8407));
  AOI22xp33_ASAP7_75t_L     g08151(.A1(\b[42] ), .A2(new_n651), .B1(\b[44] ), .B2(new_n581), .Y(new_n8408));
  OAI221xp5_ASAP7_75t_L     g08152(.A1(new_n821), .A2(new_n5805), .B1(new_n577), .B2(new_n5835), .C(new_n8408), .Y(new_n8409));
  XNOR2x2_ASAP7_75t_L       g08153(.A(\a[11] ), .B(new_n8409), .Y(new_n8410));
  INVx1_ASAP7_75t_L         g08154(.A(new_n8410), .Y(new_n8411));
  NAND3xp33_ASAP7_75t_L     g08155(.A(new_n8407), .B(new_n8405), .C(new_n8411), .Y(new_n8412));
  AO21x2_ASAP7_75t_L        g08156(.A1(new_n8131), .A2(new_n8130), .B(new_n8403), .Y(new_n8413));
  NOR2xp33_ASAP7_75t_L      g08157(.A(new_n8406), .B(new_n8413), .Y(new_n8414));
  AOI21xp33_ASAP7_75t_L     g08158(.A1(new_n8402), .A2(new_n8396), .B(new_n8404), .Y(new_n8415));
  OAI21xp33_ASAP7_75t_L     g08159(.A1(new_n8415), .A2(new_n8414), .B(new_n8410), .Y(new_n8416));
  A2O1A1O1Ixp25_ASAP7_75t_L g08160(.A1(new_n7286), .A2(new_n7285), .B(new_n7558), .C(new_n7557), .D(new_n7863), .Y(new_n8417));
  OAI211xp5_ASAP7_75t_L     g08161(.A1(new_n7875), .A2(new_n8417), .B(new_n7874), .C(new_n8138), .Y(new_n8418));
  NAND4xp25_ASAP7_75t_L     g08162(.A(new_n8418), .B(new_n8137), .C(new_n8416), .D(new_n8412), .Y(new_n8419));
  NOR3xp33_ASAP7_75t_L      g08163(.A(new_n8414), .B(new_n8415), .C(new_n8410), .Y(new_n8420));
  AOI21xp33_ASAP7_75t_L     g08164(.A1(new_n8407), .A2(new_n8405), .B(new_n8411), .Y(new_n8421));
  AOI221xp5_ASAP7_75t_L     g08165(.A1(new_n8141), .A2(new_n8136), .B1(new_n7873), .B2(new_n7861), .C(new_n7858), .Y(new_n8422));
  OAI22xp33_ASAP7_75t_L     g08166(.A1(new_n8422), .A2(new_n8142), .B1(new_n8421), .B2(new_n8420), .Y(new_n8423));
  NAND3xp33_ASAP7_75t_L     g08167(.A(new_n8423), .B(new_n8419), .C(new_n8191), .Y(new_n8424));
  OR2x4_ASAP7_75t_L         g08168(.A(new_n8190), .B(new_n8189), .Y(new_n8425));
  NOR4xp25_ASAP7_75t_L      g08169(.A(new_n8422), .B(new_n8420), .C(new_n8421), .D(new_n8142), .Y(new_n8426));
  AOI22xp33_ASAP7_75t_L     g08170(.A1(new_n8416), .A2(new_n8412), .B1(new_n8137), .B2(new_n8418), .Y(new_n8427));
  OAI21xp33_ASAP7_75t_L     g08171(.A1(new_n8427), .A2(new_n8426), .B(new_n8425), .Y(new_n8428));
  A2O1A1O1Ixp25_ASAP7_75t_L g08172(.A1(new_n7884), .A2(new_n7883), .B(new_n7915), .C(new_n8150), .D(new_n8145), .Y(new_n8429));
  NAND3xp33_ASAP7_75t_L     g08173(.A(new_n8429), .B(new_n8428), .C(new_n8424), .Y(new_n8430));
  INVx1_ASAP7_75t_L         g08174(.A(new_n8430), .Y(new_n8431));
  AOI21xp33_ASAP7_75t_L     g08175(.A1(new_n8428), .A2(new_n8424), .B(new_n8429), .Y(new_n8432));
  NAND2xp33_ASAP7_75t_L     g08176(.A(\b[49] ), .B(new_n347), .Y(new_n8433));
  NAND2xp33_ASAP7_75t_L     g08177(.A(new_n341), .B(new_n7601), .Y(new_n8434));
  AOI22xp33_ASAP7_75t_L     g08178(.A1(new_n344), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n370), .Y(new_n8435));
  AND4x1_ASAP7_75t_L        g08179(.A(new_n8435), .B(new_n8434), .C(new_n8433), .D(\a[5] ), .Y(new_n8436));
  AOI31xp33_ASAP7_75t_L     g08180(.A1(new_n8434), .A2(new_n8433), .A3(new_n8435), .B(\a[5] ), .Y(new_n8437));
  NOR2xp33_ASAP7_75t_L      g08181(.A(new_n8437), .B(new_n8436), .Y(new_n8438));
  NOR3xp33_ASAP7_75t_L      g08182(.A(new_n8431), .B(new_n8432), .C(new_n8438), .Y(new_n8439));
  NAND2xp33_ASAP7_75t_L     g08183(.A(new_n8424), .B(new_n8428), .Y(new_n8440));
  A2O1A1Ixp33_ASAP7_75t_L   g08184(.A1(new_n8150), .A2(new_n8148), .B(new_n8145), .C(new_n8440), .Y(new_n8441));
  INVx1_ASAP7_75t_L         g08185(.A(new_n8438), .Y(new_n8442));
  AOI21xp33_ASAP7_75t_L     g08186(.A1(new_n8441), .A2(new_n8430), .B(new_n8442), .Y(new_n8443));
  OAI221xp5_ASAP7_75t_L     g08187(.A1(new_n8180), .A2(new_n7910), .B1(new_n8443), .B2(new_n8439), .C(new_n8184), .Y(new_n8444));
  MAJIxp5_ASAP7_75t_L       g08188(.A(new_n7910), .B(new_n8181), .C(new_n8154), .Y(new_n8445));
  NAND3xp33_ASAP7_75t_L     g08189(.A(new_n8441), .B(new_n8430), .C(new_n8442), .Y(new_n8446));
  INVx1_ASAP7_75t_L         g08190(.A(new_n8443), .Y(new_n8447));
  NAND3xp33_ASAP7_75t_L     g08191(.A(new_n8445), .B(new_n8447), .C(new_n8446), .Y(new_n8448));
  NAND2xp33_ASAP7_75t_L     g08192(.A(new_n8448), .B(new_n8444), .Y(new_n8449));
  XNOR2x2_ASAP7_75t_L       g08193(.A(new_n8177), .B(new_n8449), .Y(new_n8450));
  O2A1O1Ixp33_ASAP7_75t_L   g08194(.A1(new_n8162), .A2(new_n7898), .B(new_n8160), .C(new_n8450), .Y(new_n8451));
  A2O1A1O1Ixp25_ASAP7_75t_L g08195(.A1(new_n7894), .A2(new_n7613), .B(new_n7892), .C(new_n8161), .D(new_n8159), .Y(new_n8452));
  AND2x2_ASAP7_75t_L        g08196(.A(new_n8452), .B(new_n8450), .Y(new_n8453));
  NOR2xp33_ASAP7_75t_L      g08197(.A(new_n8451), .B(new_n8453), .Y(\f[53] ));
  MAJIxp5_ASAP7_75t_L       g08198(.A(new_n8452), .B(new_n8177), .C(new_n8449), .Y(new_n8455));
  INVx1_ASAP7_75t_L         g08199(.A(new_n8166), .Y(new_n8456));
  NOR2xp33_ASAP7_75t_L      g08200(.A(\b[53] ), .B(\b[54] ), .Y(new_n8457));
  INVx1_ASAP7_75t_L         g08201(.A(\b[54] ), .Y(new_n8458));
  NOR2xp33_ASAP7_75t_L      g08202(.A(new_n8165), .B(new_n8458), .Y(new_n8459));
  NOR2xp33_ASAP7_75t_L      g08203(.A(new_n8457), .B(new_n8459), .Y(new_n8460));
  INVx1_ASAP7_75t_L         g08204(.A(new_n8460), .Y(new_n8461));
  O2A1O1Ixp33_ASAP7_75t_L   g08205(.A1(new_n8168), .A2(new_n8171), .B(new_n8456), .C(new_n8461), .Y(new_n8462));
  NOR3xp33_ASAP7_75t_L      g08206(.A(new_n8169), .B(new_n8460), .C(new_n8166), .Y(new_n8463));
  NOR2xp33_ASAP7_75t_L      g08207(.A(new_n8462), .B(new_n8463), .Y(new_n8464));
  INVx1_ASAP7_75t_L         g08208(.A(new_n8464), .Y(new_n8465));
  AOI22xp33_ASAP7_75t_L     g08209(.A1(\b[52] ), .A2(new_n282), .B1(\b[54] ), .B2(new_n303), .Y(new_n8466));
  OAI221xp5_ASAP7_75t_L     g08210(.A1(new_n291), .A2(new_n8165), .B1(new_n268), .B2(new_n8465), .C(new_n8466), .Y(new_n8467));
  XNOR2x2_ASAP7_75t_L       g08211(.A(\a[2] ), .B(new_n8467), .Y(new_n8468));
  AOI22xp33_ASAP7_75t_L     g08212(.A1(new_n444), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n471), .Y(new_n8469));
  OAI21xp33_ASAP7_75t_L     g08213(.A1(new_n469), .A2(new_n6837), .B(new_n8469), .Y(new_n8470));
  AOI211xp5_ASAP7_75t_L     g08214(.A1(\b[47] ), .A2(new_n447), .B(new_n435), .C(new_n8470), .Y(new_n8471));
  NOR2xp33_ASAP7_75t_L      g08215(.A(new_n6812), .B(new_n468), .Y(new_n8472));
  OA21x2_ASAP7_75t_L        g08216(.A1(new_n8472), .A2(new_n8470), .B(new_n435), .Y(new_n8473));
  NOR2xp33_ASAP7_75t_L      g08217(.A(new_n8471), .B(new_n8473), .Y(new_n8474));
  NOR2xp33_ASAP7_75t_L      g08218(.A(new_n5829), .B(new_n821), .Y(new_n8475));
  INVx1_ASAP7_75t_L         g08219(.A(new_n8475), .Y(new_n8476));
  NAND2xp33_ASAP7_75t_L     g08220(.A(new_n578), .B(new_n7066), .Y(new_n8477));
  AOI22xp33_ASAP7_75t_L     g08221(.A1(\b[43] ), .A2(new_n651), .B1(\b[45] ), .B2(new_n581), .Y(new_n8478));
  AND4x1_ASAP7_75t_L        g08222(.A(new_n8478), .B(new_n8477), .C(new_n8476), .D(\a[11] ), .Y(new_n8479));
  AOI31xp33_ASAP7_75t_L     g08223(.A1(new_n8477), .A2(new_n8476), .A3(new_n8478), .B(\a[11] ), .Y(new_n8480));
  NOR2xp33_ASAP7_75t_L      g08224(.A(new_n8480), .B(new_n8479), .Y(new_n8481));
  NAND3xp33_ASAP7_75t_L     g08225(.A(new_n8386), .B(new_n8389), .C(new_n8401), .Y(new_n8482));
  INVx1_ASAP7_75t_L         g08226(.A(new_n8482), .Y(new_n8483));
  NAND2xp33_ASAP7_75t_L     g08227(.A(new_n8352), .B(new_n8346), .Y(new_n8484));
  NOR2xp33_ASAP7_75t_L      g08228(.A(new_n8359), .B(new_n8484), .Y(new_n8485));
  O2A1O1Ixp33_ASAP7_75t_L   g08229(.A1(new_n8366), .A2(new_n8109), .B(new_n8370), .C(new_n8485), .Y(new_n8486));
  AOI22xp33_ASAP7_75t_L     g08230(.A1(new_n1360), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n1581), .Y(new_n8487));
  OAI221xp5_ASAP7_75t_L     g08231(.A1(new_n1373), .A2(new_n3804), .B1(new_n1359), .B2(new_n4223), .C(new_n8487), .Y(new_n8488));
  XNOR2x2_ASAP7_75t_L       g08232(.A(\a[20] ), .B(new_n8488), .Y(new_n8489));
  INVx1_ASAP7_75t_L         g08233(.A(new_n8489), .Y(new_n8490));
  OAI21xp33_ASAP7_75t_L     g08234(.A1(new_n8333), .A2(new_n8204), .B(new_n8339), .Y(new_n8491));
  AOI22xp33_ASAP7_75t_L     g08235(.A1(new_n2114), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n2259), .Y(new_n8492));
  OAI221xp5_ASAP7_75t_L     g08236(.A1(new_n2109), .A2(new_n2688), .B1(new_n2257), .B2(new_n2990), .C(new_n8492), .Y(new_n8493));
  XNOR2x2_ASAP7_75t_L       g08237(.A(\a[26] ), .B(new_n8493), .Y(new_n8494));
  INVx1_ASAP7_75t_L         g08238(.A(new_n8494), .Y(new_n8495));
  INVx1_ASAP7_75t_L         g08239(.A(new_n8327), .Y(new_n8496));
  AOI22xp33_ASAP7_75t_L     g08240(.A1(new_n2552), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n2736), .Y(new_n8497));
  OAI221xp5_ASAP7_75t_L     g08241(.A1(new_n2547), .A2(new_n2348), .B1(new_n2734), .B2(new_n2505), .C(new_n8497), .Y(new_n8498));
  XNOR2x2_ASAP7_75t_L       g08242(.A(\a[29] ), .B(new_n8498), .Y(new_n8499));
  NAND2xp33_ASAP7_75t_L     g08243(.A(new_n8310), .B(new_n8311), .Y(new_n8500));
  AOI22xp33_ASAP7_75t_L     g08244(.A1(new_n3029), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n3258), .Y(new_n8501));
  INVx1_ASAP7_75t_L         g08245(.A(new_n8501), .Y(new_n8502));
  AOI221xp5_ASAP7_75t_L     g08246(.A1(new_n3030), .A2(\b[23] ), .B1(new_n3021), .B2(new_n1935), .C(new_n8502), .Y(new_n8503));
  XNOR2x2_ASAP7_75t_L       g08247(.A(\a[32] ), .B(new_n8503), .Y(new_n8504));
  AOI21xp33_ASAP7_75t_L     g08248(.A1(new_n8297), .A2(new_n8303), .B(new_n8306), .Y(new_n8505));
  AOI31xp33_ASAP7_75t_L     g08249(.A1(new_n8309), .A2(new_n8036), .A3(new_n8308), .B(new_n8505), .Y(new_n8506));
  AOI22xp33_ASAP7_75t_L     g08250(.A1(new_n3633), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n3858), .Y(new_n8507));
  OAI221xp5_ASAP7_75t_L     g08251(.A1(new_n3853), .A2(new_n1539), .B1(new_n3856), .B2(new_n1662), .C(new_n8507), .Y(new_n8508));
  XNOR2x2_ASAP7_75t_L       g08252(.A(\a[35] ), .B(new_n8508), .Y(new_n8509));
  NOR3xp33_ASAP7_75t_L      g08253(.A(new_n8291), .B(new_n8288), .C(new_n8224), .Y(new_n8510));
  O2A1O1Ixp33_ASAP7_75t_L   g08254(.A1(new_n8301), .A2(new_n8302), .B(new_n8221), .C(new_n8510), .Y(new_n8511));
  AOI22xp33_ASAP7_75t_L     g08255(.A1(new_n4283), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n4512), .Y(new_n8512));
  OAI221xp5_ASAP7_75t_L     g08256(.A1(new_n4277), .A2(new_n1201), .B1(new_n4499), .B2(new_n1320), .C(new_n8512), .Y(new_n8513));
  XNOR2x2_ASAP7_75t_L       g08257(.A(new_n4268), .B(new_n8513), .Y(new_n8514));
  NOR3xp33_ASAP7_75t_L      g08258(.A(new_n8284), .B(new_n8285), .C(new_n8282), .Y(new_n8515));
  INVx1_ASAP7_75t_L         g08259(.A(new_n8515), .Y(new_n8516));
  AOI22xp33_ASAP7_75t_L     g08260(.A1(new_n4920), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n5167), .Y(new_n8517));
  OAI221xp5_ASAP7_75t_L     g08261(.A1(new_n5154), .A2(new_n869), .B1(new_n5158), .B2(new_n950), .C(new_n8517), .Y(new_n8518));
  XNOR2x2_ASAP7_75t_L       g08262(.A(\a[41] ), .B(new_n8518), .Y(new_n8519));
  INVx1_ASAP7_75t_L         g08263(.A(new_n8519), .Y(new_n8520));
  NOR3xp33_ASAP7_75t_L      g08264(.A(new_n8266), .B(new_n8268), .C(new_n8231), .Y(new_n8521));
  AO31x2_ASAP7_75t_L        g08265(.A1(new_n8277), .A2(new_n8269), .A3(new_n8003), .B(new_n8521), .Y(new_n8522));
  AOI22xp33_ASAP7_75t_L     g08266(.A1(new_n5624), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n5901), .Y(new_n8523));
  INVx1_ASAP7_75t_L         g08267(.A(new_n8523), .Y(new_n8524));
  AOI221xp5_ASAP7_75t_L     g08268(.A1(new_n5628), .A2(\b[11] ), .B1(new_n5621), .B2(new_n1232), .C(new_n8524), .Y(new_n8525));
  XNOR2x2_ASAP7_75t_L       g08269(.A(\a[44] ), .B(new_n8525), .Y(new_n8526));
  AND3x1_ASAP7_75t_L        g08270(.A(new_n8262), .B(new_n8256), .C(new_n8235), .Y(new_n8527));
  A2O1A1O1Ixp25_ASAP7_75t_L g08271(.A1(new_n7989), .A2(new_n7991), .B(new_n8271), .C(new_n8263), .D(new_n8527), .Y(new_n8528));
  AOI22xp33_ASAP7_75t_L     g08272(.A1(new_n6376), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n6648), .Y(new_n8529));
  OAI221xp5_ASAP7_75t_L     g08273(.A1(new_n6646), .A2(new_n488), .B1(new_n6636), .B2(new_n548), .C(new_n8529), .Y(new_n8530));
  NOR2xp33_ASAP7_75t_L      g08274(.A(new_n6371), .B(new_n8530), .Y(new_n8531));
  NAND2xp33_ASAP7_75t_L     g08275(.A(new_n6371), .B(new_n8530), .Y(new_n8532));
  INVx1_ASAP7_75t_L         g08276(.A(new_n8532), .Y(new_n8533));
  NAND5xp2_ASAP7_75t_L      g08277(.A(\a[53] ), .B(new_n7959), .C(new_n7961), .D(new_n7964), .E(new_n7674), .Y(new_n8534));
  NAND2xp33_ASAP7_75t_L     g08278(.A(\b[1] ), .B(new_n7963), .Y(new_n8535));
  NOR2xp33_ASAP7_75t_L      g08279(.A(new_n280), .B(new_n7957), .Y(new_n8536));
  AND3x1_ASAP7_75t_L        g08280(.A(new_n7669), .B(new_n7962), .C(new_n7956), .Y(new_n8537));
  AOI221xp5_ASAP7_75t_L     g08281(.A1(new_n7960), .A2(\b[2] ), .B1(new_n8537), .B2(\b[0] ), .C(new_n8536), .Y(new_n8538));
  NAND2xp33_ASAP7_75t_L     g08282(.A(new_n8535), .B(new_n8538), .Y(new_n8539));
  INVx1_ASAP7_75t_L         g08283(.A(\a[54] ), .Y(new_n8540));
  NAND2xp33_ASAP7_75t_L     g08284(.A(\a[53] ), .B(new_n8540), .Y(new_n8541));
  NAND2xp33_ASAP7_75t_L     g08285(.A(\a[54] ), .B(new_n7954), .Y(new_n8542));
  AND2x2_ASAP7_75t_L        g08286(.A(new_n8541), .B(new_n8542), .Y(new_n8543));
  NOR2xp33_ASAP7_75t_L      g08287(.A(new_n258), .B(new_n8543), .Y(new_n8544));
  OAI21xp33_ASAP7_75t_L     g08288(.A1(new_n8534), .A2(new_n8539), .B(new_n8544), .Y(new_n8545));
  A2O1A1Ixp33_ASAP7_75t_L   g08289(.A1(new_n7667), .A2(new_n7668), .B(new_n258), .C(\a[53] ), .Y(new_n8546));
  AOI211xp5_ASAP7_75t_L     g08290(.A1(new_n7958), .A2(new_n269), .B(new_n8546), .C(new_n8244), .Y(new_n8547));
  INVx1_ASAP7_75t_L         g08291(.A(new_n8544), .Y(new_n8548));
  NAND4xp25_ASAP7_75t_L     g08292(.A(new_n8547), .B(new_n8548), .C(new_n8538), .D(new_n8535), .Y(new_n8549));
  OAI22xp33_ASAP7_75t_L     g08293(.A1(new_n8247), .A2(new_n261), .B1(new_n298), .B2(new_n8243), .Y(new_n8550));
  AOI221xp5_ASAP7_75t_L     g08294(.A1(\b[2] ), .A2(new_n7963), .B1(new_n406), .B2(new_n7958), .C(new_n8550), .Y(new_n8551));
  NAND2xp33_ASAP7_75t_L     g08295(.A(\a[53] ), .B(new_n8551), .Y(new_n8552));
  AO21x2_ASAP7_75t_L        g08296(.A1(new_n406), .A2(new_n7958), .B(new_n8550), .Y(new_n8553));
  A2O1A1Ixp33_ASAP7_75t_L   g08297(.A1(\b[2] ), .A2(new_n7963), .B(new_n8553), .C(new_n7954), .Y(new_n8554));
  AO22x1_ASAP7_75t_L        g08298(.A1(new_n8554), .A2(new_n8552), .B1(new_n8549), .B2(new_n8545), .Y(new_n8555));
  XNOR2x2_ASAP7_75t_L       g08299(.A(new_n7954), .B(new_n8551), .Y(new_n8556));
  NAND3xp33_ASAP7_75t_L     g08300(.A(new_n8556), .B(new_n8549), .C(new_n8545), .Y(new_n8557));
  INVx1_ASAP7_75t_L         g08301(.A(new_n7115), .Y(new_n8558));
  NOR2xp33_ASAP7_75t_L      g08302(.A(new_n354), .B(new_n8558), .Y(new_n8559));
  INVx1_ASAP7_75t_L         g08303(.A(new_n8559), .Y(new_n8560));
  NAND2xp33_ASAP7_75t_L     g08304(.A(new_n7108), .B(new_n526), .Y(new_n8561));
  AOI22xp33_ASAP7_75t_L     g08305(.A1(new_n7111), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n7391), .Y(new_n8562));
  NAND4xp25_ASAP7_75t_L     g08306(.A(new_n8561), .B(\a[50] ), .C(new_n8560), .D(new_n8562), .Y(new_n8563));
  AOI31xp33_ASAP7_75t_L     g08307(.A1(new_n8561), .A2(new_n8560), .A3(new_n8562), .B(\a[50] ), .Y(new_n8564));
  INVx1_ASAP7_75t_L         g08308(.A(new_n8564), .Y(new_n8565));
  NAND4xp25_ASAP7_75t_L     g08309(.A(new_n8557), .B(new_n8565), .C(new_n8555), .D(new_n8563), .Y(new_n8566));
  AOI21xp33_ASAP7_75t_L     g08310(.A1(new_n8549), .A2(new_n8545), .B(new_n8556), .Y(new_n8567));
  AND4x1_ASAP7_75t_L        g08311(.A(new_n8545), .B(new_n8554), .C(new_n8549), .D(new_n8552), .Y(new_n8568));
  INVx1_ASAP7_75t_L         g08312(.A(new_n8563), .Y(new_n8569));
  OAI22xp33_ASAP7_75t_L     g08313(.A1(new_n8567), .A2(new_n8568), .B1(new_n8564), .B2(new_n8569), .Y(new_n8570));
  AOI221xp5_ASAP7_75t_L     g08314(.A1(new_n8236), .A2(new_n8254), .B1(new_n8566), .B2(new_n8570), .C(new_n8253), .Y(new_n8571));
  NAND2xp33_ASAP7_75t_L     g08315(.A(new_n8566), .B(new_n8570), .Y(new_n8572));
  O2A1O1Ixp33_ASAP7_75t_L   g08316(.A1(new_n8258), .A2(new_n8255), .B(new_n8261), .C(new_n8572), .Y(new_n8573));
  OAI22xp33_ASAP7_75t_L     g08317(.A1(new_n8573), .A2(new_n8571), .B1(new_n8533), .B2(new_n8531), .Y(new_n8574));
  INVx1_ASAP7_75t_L         g08318(.A(new_n8531), .Y(new_n8575));
  NOR4xp25_ASAP7_75t_L      g08319(.A(new_n8567), .B(new_n8569), .C(new_n8568), .D(new_n8564), .Y(new_n8576));
  AOI22xp33_ASAP7_75t_L     g08320(.A1(new_n8563), .A2(new_n8565), .B1(new_n8555), .B2(new_n8557), .Y(new_n8577));
  OAI211xp5_ASAP7_75t_L     g08321(.A1(new_n7975), .A2(new_n7974), .B(new_n7970), .C(new_n8254), .Y(new_n8578));
  OAI211xp5_ASAP7_75t_L     g08322(.A1(new_n8576), .A2(new_n8577), .B(new_n8578), .C(new_n8261), .Y(new_n8579));
  NOR2xp33_ASAP7_75t_L      g08323(.A(new_n8577), .B(new_n8576), .Y(new_n8580));
  A2O1A1Ixp33_ASAP7_75t_L   g08324(.A1(new_n8254), .A2(new_n8236), .B(new_n8253), .C(new_n8580), .Y(new_n8581));
  NAND4xp25_ASAP7_75t_L     g08325(.A(new_n8581), .B(new_n8575), .C(new_n8532), .D(new_n8579), .Y(new_n8582));
  AOI21xp33_ASAP7_75t_L     g08326(.A1(new_n8582), .A2(new_n8574), .B(new_n8528), .Y(new_n8583));
  AND3x1_ASAP7_75t_L        g08327(.A(new_n8528), .B(new_n8582), .C(new_n8574), .Y(new_n8584));
  OAI21xp33_ASAP7_75t_L     g08328(.A1(new_n8583), .A2(new_n8584), .B(new_n8526), .Y(new_n8585));
  XNOR2x2_ASAP7_75t_L       g08329(.A(new_n5619), .B(new_n8525), .Y(new_n8586));
  NAND2xp33_ASAP7_75t_L     g08330(.A(new_n8582), .B(new_n8574), .Y(new_n8587));
  A2O1A1Ixp33_ASAP7_75t_L   g08331(.A1(new_n8272), .A2(new_n8267), .B(new_n8527), .C(new_n8587), .Y(new_n8588));
  NAND3xp33_ASAP7_75t_L     g08332(.A(new_n8528), .B(new_n8574), .C(new_n8582), .Y(new_n8589));
  NAND3xp33_ASAP7_75t_L     g08333(.A(new_n8588), .B(new_n8586), .C(new_n8589), .Y(new_n8590));
  NAND2xp33_ASAP7_75t_L     g08334(.A(new_n8590), .B(new_n8585), .Y(new_n8591));
  NAND2xp33_ASAP7_75t_L     g08335(.A(new_n8522), .B(new_n8591), .Y(new_n8592));
  AOI31xp33_ASAP7_75t_L     g08336(.A1(new_n8277), .A2(new_n8269), .A3(new_n8003), .B(new_n8521), .Y(new_n8593));
  NAND3xp33_ASAP7_75t_L     g08337(.A(new_n8593), .B(new_n8585), .C(new_n8590), .Y(new_n8594));
  NAND3xp33_ASAP7_75t_L     g08338(.A(new_n8592), .B(new_n8594), .C(new_n8520), .Y(new_n8595));
  AOI21xp33_ASAP7_75t_L     g08339(.A1(new_n8590), .A2(new_n8585), .B(new_n8593), .Y(new_n8596));
  NOR2xp33_ASAP7_75t_L      g08340(.A(new_n8522), .B(new_n8591), .Y(new_n8597));
  OAI21xp33_ASAP7_75t_L     g08341(.A1(new_n8596), .A2(new_n8597), .B(new_n8519), .Y(new_n8598));
  NAND2xp33_ASAP7_75t_L     g08342(.A(new_n8595), .B(new_n8598), .Y(new_n8599));
  O2A1O1Ixp33_ASAP7_75t_L   g08343(.A1(new_n8228), .A2(new_n8294), .B(new_n8516), .C(new_n8599), .Y(new_n8600));
  AOI221xp5_ASAP7_75t_L     g08344(.A1(new_n8598), .A2(new_n8595), .B1(new_n8289), .B2(new_n8290), .C(new_n8515), .Y(new_n8601));
  OAI21xp33_ASAP7_75t_L     g08345(.A1(new_n8601), .A2(new_n8600), .B(new_n8514), .Y(new_n8602));
  XNOR2x2_ASAP7_75t_L       g08346(.A(\a[38] ), .B(new_n8513), .Y(new_n8603));
  A2O1A1Ixp33_ASAP7_75t_L   g08347(.A1(new_n8283), .A2(new_n8287), .B(new_n8228), .C(new_n8516), .Y(new_n8604));
  NAND3xp33_ASAP7_75t_L     g08348(.A(new_n8604), .B(new_n8595), .C(new_n8598), .Y(new_n8605));
  AO221x2_ASAP7_75t_L       g08349(.A1(new_n8598), .A2(new_n8595), .B1(new_n8289), .B2(new_n8290), .C(new_n8515), .Y(new_n8606));
  NAND3xp33_ASAP7_75t_L     g08350(.A(new_n8605), .B(new_n8606), .C(new_n8603), .Y(new_n8607));
  AOI21xp33_ASAP7_75t_L     g08351(.A1(new_n8607), .A2(new_n8602), .B(new_n8511), .Y(new_n8608));
  INVx1_ASAP7_75t_L         g08352(.A(new_n8510), .Y(new_n8609));
  OAI21xp33_ASAP7_75t_L     g08353(.A1(new_n8301), .A2(new_n8302), .B(new_n8221), .Y(new_n8610));
  AND4x1_ASAP7_75t_L        g08354(.A(new_n8610), .B(new_n8609), .C(new_n8607), .D(new_n8602), .Y(new_n8611));
  NOR3xp33_ASAP7_75t_L      g08355(.A(new_n8611), .B(new_n8608), .C(new_n8509), .Y(new_n8612));
  INVx1_ASAP7_75t_L         g08356(.A(new_n8509), .Y(new_n8613));
  NAND2xp33_ASAP7_75t_L     g08357(.A(new_n8292), .B(new_n8296), .Y(new_n8614));
  NAND2xp33_ASAP7_75t_L     g08358(.A(new_n8607), .B(new_n8602), .Y(new_n8615));
  A2O1A1Ixp33_ASAP7_75t_L   g08359(.A1(new_n8614), .A2(new_n8221), .B(new_n8510), .C(new_n8615), .Y(new_n8616));
  AOI21xp33_ASAP7_75t_L     g08360(.A1(new_n8605), .A2(new_n8606), .B(new_n8603), .Y(new_n8617));
  NOR3xp33_ASAP7_75t_L      g08361(.A(new_n8600), .B(new_n8601), .C(new_n8514), .Y(new_n8618));
  NOR2xp33_ASAP7_75t_L      g08362(.A(new_n8617), .B(new_n8618), .Y(new_n8619));
  NAND2xp33_ASAP7_75t_L     g08363(.A(new_n8511), .B(new_n8619), .Y(new_n8620));
  AOI21xp33_ASAP7_75t_L     g08364(.A1(new_n8616), .A2(new_n8620), .B(new_n8613), .Y(new_n8621));
  OR3x1_ASAP7_75t_L         g08365(.A(new_n8506), .B(new_n8612), .C(new_n8621), .Y(new_n8622));
  OAI21xp33_ASAP7_75t_L     g08366(.A1(new_n8612), .A2(new_n8621), .B(new_n8506), .Y(new_n8623));
  NAND3xp33_ASAP7_75t_L     g08367(.A(new_n8622), .B(new_n8504), .C(new_n8623), .Y(new_n8624));
  XNOR2x2_ASAP7_75t_L       g08368(.A(new_n3015), .B(new_n8503), .Y(new_n8625));
  NOR3xp33_ASAP7_75t_L      g08369(.A(new_n8506), .B(new_n8621), .C(new_n8612), .Y(new_n8626));
  NAND3xp33_ASAP7_75t_L     g08370(.A(new_n8616), .B(new_n8620), .C(new_n8613), .Y(new_n8627));
  OAI21xp33_ASAP7_75t_L     g08371(.A1(new_n8608), .A2(new_n8611), .B(new_n8509), .Y(new_n8628));
  AOI211xp5_ASAP7_75t_L     g08372(.A1(new_n8628), .A2(new_n8627), .B(new_n8505), .C(new_n8313), .Y(new_n8629));
  OAI21xp33_ASAP7_75t_L     g08373(.A1(new_n8626), .A2(new_n8629), .B(new_n8625), .Y(new_n8630));
  NAND2xp33_ASAP7_75t_L     g08374(.A(new_n8630), .B(new_n8624), .Y(new_n8631));
  O2A1O1Ixp33_ASAP7_75t_L   g08375(.A1(new_n8218), .A2(new_n8500), .B(new_n8324), .C(new_n8631), .Y(new_n8632));
  NOR2xp33_ASAP7_75t_L      g08376(.A(new_n8314), .B(new_n8313), .Y(new_n8633));
  NAND2xp33_ASAP7_75t_L     g08377(.A(new_n8217), .B(new_n8633), .Y(new_n8634));
  OAI21xp33_ASAP7_75t_L     g08378(.A1(new_n8316), .A2(new_n8325), .B(new_n8634), .Y(new_n8635));
  NOR3xp33_ASAP7_75t_L      g08379(.A(new_n8629), .B(new_n8626), .C(new_n8625), .Y(new_n8636));
  AOI21xp33_ASAP7_75t_L     g08380(.A1(new_n8622), .A2(new_n8623), .B(new_n8504), .Y(new_n8637));
  NOR2xp33_ASAP7_75t_L      g08381(.A(new_n8636), .B(new_n8637), .Y(new_n8638));
  NOR2xp33_ASAP7_75t_L      g08382(.A(new_n8635), .B(new_n8638), .Y(new_n8639));
  NOR3xp33_ASAP7_75t_L      g08383(.A(new_n8632), .B(new_n8639), .C(new_n8499), .Y(new_n8640));
  INVx1_ASAP7_75t_L         g08384(.A(new_n8499), .Y(new_n8641));
  A2O1A1Ixp33_ASAP7_75t_L   g08385(.A1(new_n8633), .A2(new_n8217), .B(new_n8317), .C(new_n8638), .Y(new_n8642));
  NOR2xp33_ASAP7_75t_L      g08386(.A(new_n8218), .B(new_n8500), .Y(new_n8643));
  A2O1A1O1Ixp25_ASAP7_75t_L g08387(.A1(new_n8054), .A2(new_n8048), .B(new_n8046), .C(new_n8320), .D(new_n8643), .Y(new_n8644));
  NAND2xp33_ASAP7_75t_L     g08388(.A(new_n8631), .B(new_n8644), .Y(new_n8645));
  AOI21xp33_ASAP7_75t_L     g08389(.A1(new_n8642), .A2(new_n8645), .B(new_n8641), .Y(new_n8646));
  NOR2xp33_ASAP7_75t_L      g08390(.A(new_n8640), .B(new_n8646), .Y(new_n8647));
  OAI21xp33_ASAP7_75t_L     g08391(.A1(new_n8496), .A2(new_n8334), .B(new_n8647), .Y(new_n8648));
  NAND2xp33_ASAP7_75t_L     g08392(.A(new_n8059), .B(new_n8053), .Y(new_n8649));
  NOR2xp33_ASAP7_75t_L      g08393(.A(new_n8052), .B(new_n8209), .Y(new_n8650));
  A2O1A1O1Ixp25_ASAP7_75t_L g08394(.A1(new_n8061), .A2(new_n8649), .B(new_n8650), .C(new_n8322), .D(new_n8496), .Y(new_n8651));
  OAI21xp33_ASAP7_75t_L     g08395(.A1(new_n8640), .A2(new_n8646), .B(new_n8651), .Y(new_n8652));
  NAND3xp33_ASAP7_75t_L     g08396(.A(new_n8648), .B(new_n8495), .C(new_n8652), .Y(new_n8653));
  NOR3xp33_ASAP7_75t_L      g08397(.A(new_n8651), .B(new_n8640), .C(new_n8646), .Y(new_n8654));
  NAND3xp33_ASAP7_75t_L     g08398(.A(new_n8642), .B(new_n8645), .C(new_n8641), .Y(new_n8655));
  OAI21xp33_ASAP7_75t_L     g08399(.A1(new_n8639), .A2(new_n8632), .B(new_n8499), .Y(new_n8656));
  AOI221xp5_ASAP7_75t_L     g08400(.A1(new_n8210), .A2(new_n8322), .B1(new_n8656), .B2(new_n8655), .C(new_n8496), .Y(new_n8657));
  OAI21xp33_ASAP7_75t_L     g08401(.A1(new_n8657), .A2(new_n8654), .B(new_n8494), .Y(new_n8658));
  NAND3xp33_ASAP7_75t_L     g08402(.A(new_n8491), .B(new_n8653), .C(new_n8658), .Y(new_n8659));
  A2O1A1O1Ixp25_ASAP7_75t_L g08403(.A1(new_n8071), .A2(new_n8073), .B(new_n8065), .C(new_n8338), .D(new_n8336), .Y(new_n8660));
  NOR3xp33_ASAP7_75t_L      g08404(.A(new_n8654), .B(new_n8657), .C(new_n8494), .Y(new_n8661));
  AOI21xp33_ASAP7_75t_L     g08405(.A1(new_n8648), .A2(new_n8652), .B(new_n8495), .Y(new_n8662));
  OAI21xp33_ASAP7_75t_L     g08406(.A1(new_n8661), .A2(new_n8662), .B(new_n8660), .Y(new_n8663));
  AOI22xp33_ASAP7_75t_L     g08407(.A1(new_n1704), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1837), .Y(new_n8664));
  INVx1_ASAP7_75t_L         g08408(.A(new_n8664), .Y(new_n8665));
  AOI221xp5_ASAP7_75t_L     g08409(.A1(\b[32] ), .A2(new_n1706), .B1(new_n1695), .B2(new_n4821), .C(new_n8665), .Y(new_n8666));
  XNOR2x2_ASAP7_75t_L       g08410(.A(new_n1689), .B(new_n8666), .Y(new_n8667));
  NAND3xp33_ASAP7_75t_L     g08411(.A(new_n8659), .B(new_n8663), .C(new_n8667), .Y(new_n8668));
  NOR3xp33_ASAP7_75t_L      g08412(.A(new_n8660), .B(new_n8662), .C(new_n8661), .Y(new_n8669));
  AOI21xp33_ASAP7_75t_L     g08413(.A1(new_n8658), .A2(new_n8653), .B(new_n8491), .Y(new_n8670));
  INVx1_ASAP7_75t_L         g08414(.A(new_n8667), .Y(new_n8671));
  OAI21xp33_ASAP7_75t_L     g08415(.A1(new_n8670), .A2(new_n8669), .B(new_n8671), .Y(new_n8672));
  NAND2xp33_ASAP7_75t_L     g08416(.A(new_n8668), .B(new_n8672), .Y(new_n8673));
  A2O1A1Ixp33_ASAP7_75t_L   g08417(.A1(new_n8341), .A2(new_n8193), .B(new_n8351), .C(new_n8673), .Y(new_n8674));
  A2O1A1O1Ixp25_ASAP7_75t_L g08418(.A1(new_n8084), .A2(new_n8090), .B(new_n8348), .C(new_n8341), .D(new_n8351), .Y(new_n8675));
  NAND3xp33_ASAP7_75t_L     g08419(.A(new_n8675), .B(new_n8668), .C(new_n8672), .Y(new_n8676));
  NAND3xp33_ASAP7_75t_L     g08420(.A(new_n8674), .B(new_n8490), .C(new_n8676), .Y(new_n8677));
  AOI21xp33_ASAP7_75t_L     g08421(.A1(new_n8672), .A2(new_n8668), .B(new_n8675), .Y(new_n8678));
  INVx1_ASAP7_75t_L         g08422(.A(new_n8348), .Y(new_n8679));
  A2O1A1Ixp33_ASAP7_75t_L   g08423(.A1(new_n8085), .A2(new_n8679), .B(new_n8350), .C(new_n8345), .Y(new_n8680));
  NOR2xp33_ASAP7_75t_L      g08424(.A(new_n8680), .B(new_n8673), .Y(new_n8681));
  OAI21xp33_ASAP7_75t_L     g08425(.A1(new_n8678), .A2(new_n8681), .B(new_n8489), .Y(new_n8682));
  NAND2xp33_ASAP7_75t_L     g08426(.A(new_n8682), .B(new_n8677), .Y(new_n8683));
  NAND2xp33_ASAP7_75t_L     g08427(.A(new_n8683), .B(new_n8486), .Y(new_n8684));
  OAI211xp5_ASAP7_75t_L     g08428(.A1(new_n8485), .A2(new_n8383), .B(new_n8677), .C(new_n8682), .Y(new_n8685));
  AOI22xp33_ASAP7_75t_L     g08429(.A1(new_n1076), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1253), .Y(new_n8686));
  OAI221xp5_ASAP7_75t_L     g08430(.A1(new_n1154), .A2(new_n4632), .B1(new_n1156), .B2(new_n4858), .C(new_n8686), .Y(new_n8687));
  XNOR2x2_ASAP7_75t_L       g08431(.A(\a[17] ), .B(new_n8687), .Y(new_n8688));
  NAND3xp33_ASAP7_75t_L     g08432(.A(new_n8685), .B(new_n8684), .C(new_n8688), .Y(new_n8689));
  AOI211xp5_ASAP7_75t_L     g08433(.A1(new_n8677), .A2(new_n8682), .B(new_n8485), .C(new_n8383), .Y(new_n8690));
  O2A1O1Ixp33_ASAP7_75t_L   g08434(.A1(new_n8484), .A2(new_n8359), .B(new_n8371), .C(new_n8683), .Y(new_n8691));
  INVx1_ASAP7_75t_L         g08435(.A(new_n8688), .Y(new_n8692));
  OAI21xp33_ASAP7_75t_L     g08436(.A1(new_n8690), .A2(new_n8691), .B(new_n8692), .Y(new_n8693));
  NOR3xp33_ASAP7_75t_L      g08437(.A(new_n8382), .B(new_n8383), .C(new_n8379), .Y(new_n8694));
  O2A1O1Ixp33_ASAP7_75t_L   g08438(.A1(new_n8398), .A2(new_n8399), .B(new_n8388), .C(new_n8694), .Y(new_n8695));
  NAND3xp33_ASAP7_75t_L     g08439(.A(new_n8695), .B(new_n8693), .C(new_n8689), .Y(new_n8696));
  NAND2xp33_ASAP7_75t_L     g08440(.A(new_n8689), .B(new_n8693), .Y(new_n8697));
  OAI21xp33_ASAP7_75t_L     g08441(.A1(new_n8694), .A2(new_n8400), .B(new_n8697), .Y(new_n8698));
  NAND2xp33_ASAP7_75t_L     g08442(.A(\b[40] ), .B(new_n900), .Y(new_n8699));
  OAI221xp5_ASAP7_75t_L     g08443(.A1(new_n977), .A2(new_n5338), .B1(new_n898), .B2(new_n5346), .C(new_n8699), .Y(new_n8700));
  AOI21xp33_ASAP7_75t_L     g08444(.A1(new_n815), .A2(\b[41] ), .B(new_n8700), .Y(new_n8701));
  NAND2xp33_ASAP7_75t_L     g08445(.A(\a[14] ), .B(new_n8701), .Y(new_n8702));
  A2O1A1Ixp33_ASAP7_75t_L   g08446(.A1(\b[41] ), .A2(new_n815), .B(new_n8700), .C(new_n806), .Y(new_n8703));
  NAND2xp33_ASAP7_75t_L     g08447(.A(new_n8703), .B(new_n8702), .Y(new_n8704));
  AOI21xp33_ASAP7_75t_L     g08448(.A1(new_n8698), .A2(new_n8696), .B(new_n8704), .Y(new_n8705));
  AND3x1_ASAP7_75t_L        g08449(.A(new_n8695), .B(new_n8693), .C(new_n8689), .Y(new_n8706));
  AOI21xp33_ASAP7_75t_L     g08450(.A1(new_n8693), .A2(new_n8689), .B(new_n8695), .Y(new_n8707));
  INVx1_ASAP7_75t_L         g08451(.A(new_n8704), .Y(new_n8708));
  NOR3xp33_ASAP7_75t_L      g08452(.A(new_n8706), .B(new_n8708), .C(new_n8707), .Y(new_n8709));
  NOR2xp33_ASAP7_75t_L      g08453(.A(new_n8705), .B(new_n8709), .Y(new_n8710));
  A2O1A1Ixp33_ASAP7_75t_L   g08454(.A1(new_n8413), .A2(new_n8406), .B(new_n8483), .C(new_n8710), .Y(new_n8711));
  A2O1A1O1Ixp25_ASAP7_75t_L g08455(.A1(new_n8131), .A2(new_n8130), .B(new_n8403), .C(new_n8406), .D(new_n8483), .Y(new_n8712));
  OAI21xp33_ASAP7_75t_L     g08456(.A1(new_n8707), .A2(new_n8706), .B(new_n8708), .Y(new_n8713));
  NAND3xp33_ASAP7_75t_L     g08457(.A(new_n8698), .B(new_n8696), .C(new_n8704), .Y(new_n8714));
  NAND2xp33_ASAP7_75t_L     g08458(.A(new_n8714), .B(new_n8713), .Y(new_n8715));
  NAND2xp33_ASAP7_75t_L     g08459(.A(new_n8715), .B(new_n8712), .Y(new_n8716));
  AOI21xp33_ASAP7_75t_L     g08460(.A1(new_n8711), .A2(new_n8716), .B(new_n8481), .Y(new_n8717));
  INVx1_ASAP7_75t_L         g08461(.A(new_n8481), .Y(new_n8718));
  NOR2xp33_ASAP7_75t_L      g08462(.A(new_n8715), .B(new_n8712), .Y(new_n8719));
  A2O1A1Ixp33_ASAP7_75t_L   g08463(.A1(new_n8402), .A2(new_n8396), .B(new_n8404), .C(new_n8482), .Y(new_n8720));
  NOR2xp33_ASAP7_75t_L      g08464(.A(new_n8720), .B(new_n8710), .Y(new_n8721));
  NOR3xp33_ASAP7_75t_L      g08465(.A(new_n8721), .B(new_n8719), .C(new_n8718), .Y(new_n8722));
  OAI31xp33_ASAP7_75t_L     g08466(.A1(new_n8422), .A2(new_n8142), .A3(new_n8421), .B(new_n8412), .Y(new_n8723));
  OAI21xp33_ASAP7_75t_L     g08467(.A1(new_n8722), .A2(new_n8717), .B(new_n8723), .Y(new_n8724));
  OAI21xp33_ASAP7_75t_L     g08468(.A1(new_n8719), .A2(new_n8721), .B(new_n8718), .Y(new_n8725));
  NAND3xp33_ASAP7_75t_L     g08469(.A(new_n8711), .B(new_n8481), .C(new_n8716), .Y(new_n8726));
  AOI31xp33_ASAP7_75t_L     g08470(.A1(new_n8418), .A2(new_n8137), .A3(new_n8416), .B(new_n8420), .Y(new_n8727));
  NAND3xp33_ASAP7_75t_L     g08471(.A(new_n8727), .B(new_n8726), .C(new_n8725), .Y(new_n8728));
  NAND3xp33_ASAP7_75t_L     g08472(.A(new_n8728), .B(new_n8724), .C(new_n8474), .Y(new_n8729));
  INVx1_ASAP7_75t_L         g08473(.A(new_n8474), .Y(new_n8730));
  AOI21xp33_ASAP7_75t_L     g08474(.A1(new_n8726), .A2(new_n8725), .B(new_n8727), .Y(new_n8731));
  NOR3xp33_ASAP7_75t_L      g08475(.A(new_n8723), .B(new_n8722), .C(new_n8717), .Y(new_n8732));
  OAI21xp33_ASAP7_75t_L     g08476(.A1(new_n8731), .A2(new_n8732), .B(new_n8730), .Y(new_n8733));
  NAND2xp33_ASAP7_75t_L     g08477(.A(new_n8729), .B(new_n8733), .Y(new_n8734));
  NAND3xp33_ASAP7_75t_L     g08478(.A(new_n8425), .B(new_n8423), .C(new_n8419), .Y(new_n8735));
  A2O1A1Ixp33_ASAP7_75t_L   g08479(.A1(new_n8428), .A2(new_n8424), .B(new_n8429), .C(new_n8735), .Y(new_n8736));
  NOR2xp33_ASAP7_75t_L      g08480(.A(new_n8736), .B(new_n8734), .Y(new_n8737));
  NOR3xp33_ASAP7_75t_L      g08481(.A(new_n8732), .B(new_n8731), .C(new_n8730), .Y(new_n8738));
  AOI21xp33_ASAP7_75t_L     g08482(.A1(new_n8728), .A2(new_n8724), .B(new_n8474), .Y(new_n8739));
  NOR2xp33_ASAP7_75t_L      g08483(.A(new_n8739), .B(new_n8738), .Y(new_n8740));
  AOI21xp33_ASAP7_75t_L     g08484(.A1(new_n8441), .A2(new_n8735), .B(new_n8740), .Y(new_n8741));
  NOR2xp33_ASAP7_75t_L      g08485(.A(new_n7593), .B(new_n429), .Y(new_n8742));
  INVx1_ASAP7_75t_L         g08486(.A(new_n8742), .Y(new_n8743));
  NAND2xp33_ASAP7_75t_L     g08487(.A(new_n341), .B(new_n7622), .Y(new_n8744));
  AOI22xp33_ASAP7_75t_L     g08488(.A1(new_n344), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n370), .Y(new_n8745));
  AND4x1_ASAP7_75t_L        g08489(.A(new_n8745), .B(new_n8744), .C(new_n8743), .D(\a[5] ), .Y(new_n8746));
  AOI31xp33_ASAP7_75t_L     g08490(.A1(new_n8744), .A2(new_n8743), .A3(new_n8745), .B(\a[5] ), .Y(new_n8747));
  NOR2xp33_ASAP7_75t_L      g08491(.A(new_n8747), .B(new_n8746), .Y(new_n8748));
  OAI21xp33_ASAP7_75t_L     g08492(.A1(new_n8737), .A2(new_n8741), .B(new_n8748), .Y(new_n8749));
  INVx1_ASAP7_75t_L         g08493(.A(new_n8749), .Y(new_n8750));
  NOR3xp33_ASAP7_75t_L      g08494(.A(new_n8741), .B(new_n8737), .C(new_n8748), .Y(new_n8751));
  A2O1A1O1Ixp25_ASAP7_75t_L g08495(.A1(new_n8183), .A2(new_n8182), .B(new_n8157), .C(new_n8447), .D(new_n8439), .Y(new_n8752));
  NOR3xp33_ASAP7_75t_L      g08496(.A(new_n8752), .B(new_n8750), .C(new_n8751), .Y(new_n8753));
  OA21x2_ASAP7_75t_L        g08497(.A1(new_n8751), .A2(new_n8750), .B(new_n8752), .Y(new_n8754));
  NOR3xp33_ASAP7_75t_L      g08498(.A(new_n8754), .B(new_n8753), .C(new_n8468), .Y(new_n8755));
  INVx1_ASAP7_75t_L         g08499(.A(new_n8755), .Y(new_n8756));
  OAI21xp33_ASAP7_75t_L     g08500(.A1(new_n8753), .A2(new_n8754), .B(new_n8468), .Y(new_n8757));
  NAND2xp33_ASAP7_75t_L     g08501(.A(new_n8757), .B(new_n8756), .Y(new_n8758));
  XNOR2x2_ASAP7_75t_L       g08502(.A(new_n8455), .B(new_n8758), .Y(\f[54] ));
  INVx1_ASAP7_75t_L         g08503(.A(new_n8455), .Y(new_n8760));
  NOR2xp33_ASAP7_75t_L      g08504(.A(\b[54] ), .B(\b[55] ), .Y(new_n8761));
  INVx1_ASAP7_75t_L         g08505(.A(\b[55] ), .Y(new_n8762));
  NOR2xp33_ASAP7_75t_L      g08506(.A(new_n8458), .B(new_n8762), .Y(new_n8763));
  NOR2xp33_ASAP7_75t_L      g08507(.A(new_n8761), .B(new_n8763), .Y(new_n8764));
  A2O1A1Ixp33_ASAP7_75t_L   g08508(.A1(\b[54] ), .A2(\b[53] ), .B(new_n8462), .C(new_n8764), .Y(new_n8765));
  O2A1O1Ixp33_ASAP7_75t_L   g08509(.A1(new_n8166), .A2(new_n8169), .B(new_n8460), .C(new_n8459), .Y(new_n8766));
  OAI21xp33_ASAP7_75t_L     g08510(.A1(new_n8761), .A2(new_n8763), .B(new_n8766), .Y(new_n8767));
  NAND2xp33_ASAP7_75t_L     g08511(.A(new_n8765), .B(new_n8767), .Y(new_n8768));
  AOI22xp33_ASAP7_75t_L     g08512(.A1(\b[53] ), .A2(new_n282), .B1(\b[55] ), .B2(new_n303), .Y(new_n8769));
  OAI221xp5_ASAP7_75t_L     g08513(.A1(new_n291), .A2(new_n8458), .B1(new_n268), .B2(new_n8768), .C(new_n8769), .Y(new_n8770));
  XNOR2x2_ASAP7_75t_L       g08514(.A(\a[2] ), .B(new_n8770), .Y(new_n8771));
  A2O1A1O1Ixp25_ASAP7_75t_L g08515(.A1(new_n8445), .A2(new_n8447), .B(new_n8439), .C(new_n8749), .D(new_n8751), .Y(new_n8772));
  NOR3xp33_ASAP7_75t_L      g08516(.A(new_n8732), .B(new_n8731), .C(new_n8474), .Y(new_n8773));
  INVx1_ASAP7_75t_L         g08517(.A(new_n8773), .Y(new_n8774));
  A2O1A1Ixp33_ASAP7_75t_L   g08518(.A1(new_n8441), .A2(new_n8735), .B(new_n8740), .C(new_n8774), .Y(new_n8775));
  AOI22xp33_ASAP7_75t_L     g08519(.A1(new_n444), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n471), .Y(new_n8776));
  OAI221xp5_ASAP7_75t_L     g08520(.A1(new_n468), .A2(new_n6830), .B1(new_n469), .B2(new_n7323), .C(new_n8776), .Y(new_n8777));
  XNOR2x2_ASAP7_75t_L       g08521(.A(\a[8] ), .B(new_n8777), .Y(new_n8778));
  NOR2xp33_ASAP7_75t_L      g08522(.A(new_n8719), .B(new_n8721), .Y(new_n8779));
  MAJIxp5_ASAP7_75t_L       g08523(.A(new_n8723), .B(new_n8718), .C(new_n8779), .Y(new_n8780));
  NAND2xp33_ASAP7_75t_L     g08524(.A(\b[45] ), .B(new_n584), .Y(new_n8781));
  NAND2xp33_ASAP7_75t_L     g08525(.A(new_n578), .B(new_n7919), .Y(new_n8782));
  AOI22xp33_ASAP7_75t_L     g08526(.A1(\b[44] ), .A2(new_n651), .B1(\b[46] ), .B2(new_n581), .Y(new_n8783));
  NAND4xp25_ASAP7_75t_L     g08527(.A(new_n8782), .B(\a[11] ), .C(new_n8781), .D(new_n8783), .Y(new_n8784));
  NAND2xp33_ASAP7_75t_L     g08528(.A(new_n8783), .B(new_n8782), .Y(new_n8785));
  A2O1A1Ixp33_ASAP7_75t_L   g08529(.A1(\b[45] ), .A2(new_n584), .B(new_n8785), .C(new_n574), .Y(new_n8786));
  AND2x2_ASAP7_75t_L        g08530(.A(new_n8784), .B(new_n8786), .Y(new_n8787));
  A2O1A1O1Ixp25_ASAP7_75t_L g08531(.A1(new_n8406), .A2(new_n8413), .B(new_n8483), .C(new_n8713), .D(new_n8709), .Y(new_n8788));
  OAI21xp33_ASAP7_75t_L     g08532(.A1(new_n8621), .A2(new_n8506), .B(new_n8627), .Y(new_n8789));
  AOI22xp33_ASAP7_75t_L     g08533(.A1(new_n3633), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n3858), .Y(new_n8790));
  OAI221xp5_ASAP7_75t_L     g08534(.A1(new_n3853), .A2(new_n1655), .B1(new_n3856), .B2(new_n1780), .C(new_n8790), .Y(new_n8791));
  XNOR2x2_ASAP7_75t_L       g08535(.A(\a[35] ), .B(new_n8791), .Y(new_n8792));
  INVx1_ASAP7_75t_L         g08536(.A(new_n8792), .Y(new_n8793));
  NAND3xp33_ASAP7_75t_L     g08537(.A(new_n8605), .B(new_n8606), .C(new_n8514), .Y(new_n8794));
  NAND3xp33_ASAP7_75t_L     g08538(.A(new_n8588), .B(new_n8526), .C(new_n8589), .Y(new_n8795));
  A2O1A1Ixp33_ASAP7_75t_L   g08539(.A1(new_n8585), .A2(new_n8590), .B(new_n8593), .C(new_n8795), .Y(new_n8796));
  AOI22xp33_ASAP7_75t_L     g08540(.A1(new_n5624), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n5901), .Y(new_n8797));
  OAI221xp5_ASAP7_75t_L     g08541(.A1(new_n5900), .A2(new_n760), .B1(new_n5892), .B2(new_n790), .C(new_n8797), .Y(new_n8798));
  XNOR2x2_ASAP7_75t_L       g08542(.A(\a[44] ), .B(new_n8798), .Y(new_n8799));
  INVx1_ASAP7_75t_L         g08543(.A(new_n8799), .Y(new_n8800));
  AOI211xp5_ASAP7_75t_L     g08544(.A1(new_n8575), .A2(new_n8532), .B(new_n8571), .C(new_n8573), .Y(new_n8801));
  INVx1_ASAP7_75t_L         g08545(.A(new_n8801), .Y(new_n8802));
  A2O1A1Ixp33_ASAP7_75t_L   g08546(.A1(new_n8574), .A2(new_n8582), .B(new_n8528), .C(new_n8802), .Y(new_n8803));
  AOI22xp33_ASAP7_75t_L     g08547(.A1(new_n6376), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n6648), .Y(new_n8804));
  OAI221xp5_ASAP7_75t_L     g08548(.A1(new_n6646), .A2(new_n540), .B1(new_n6636), .B2(new_n624), .C(new_n8804), .Y(new_n8805));
  XNOR2x2_ASAP7_75t_L       g08549(.A(new_n6371), .B(new_n8805), .Y(new_n8806));
  INVx1_ASAP7_75t_L         g08550(.A(new_n8806), .Y(new_n8807));
  AOI211xp5_ASAP7_75t_L     g08551(.A1(new_n8563), .A2(new_n8565), .B(new_n8568), .C(new_n8567), .Y(new_n8808));
  INVx1_ASAP7_75t_L         g08552(.A(new_n8808), .Y(new_n8809));
  AOI22xp33_ASAP7_75t_L     g08553(.A1(new_n7111), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n7391), .Y(new_n8810));
  OAI221xp5_ASAP7_75t_L     g08554(.A1(new_n8558), .A2(new_n418), .B1(new_n8237), .B2(new_n425), .C(new_n8810), .Y(new_n8811));
  XNOR2x2_ASAP7_75t_L       g08555(.A(\a[50] ), .B(new_n8811), .Y(new_n8812));
  INVx1_ASAP7_75t_L         g08556(.A(new_n8812), .Y(new_n8813));
  NOR3xp33_ASAP7_75t_L      g08557(.A(new_n8539), .B(new_n8548), .C(new_n8534), .Y(new_n8814));
  INVx1_ASAP7_75t_L         g08558(.A(new_n8814), .Y(new_n8815));
  A2O1A1Ixp33_ASAP7_75t_L   g08559(.A1(new_n8549), .A2(new_n8545), .B(new_n8556), .C(new_n8815), .Y(new_n8816));
  INVx1_ASAP7_75t_L         g08560(.A(new_n7963), .Y(new_n8817));
  OAI22xp33_ASAP7_75t_L     g08561(.A1(new_n8247), .A2(new_n276), .B1(new_n324), .B2(new_n8243), .Y(new_n8818));
  AOI21xp33_ASAP7_75t_L     g08562(.A1(new_n329), .A2(new_n7958), .B(new_n8818), .Y(new_n8819));
  OAI211xp5_ASAP7_75t_L     g08563(.A1(new_n298), .A2(new_n8817), .B(new_n8819), .C(\a[53] ), .Y(new_n8820));
  O2A1O1Ixp33_ASAP7_75t_L   g08564(.A1(new_n298), .A2(new_n8817), .B(new_n8819), .C(\a[53] ), .Y(new_n8821));
  INVx1_ASAP7_75t_L         g08565(.A(new_n8821), .Y(new_n8822));
  NAND2xp33_ASAP7_75t_L     g08566(.A(\a[56] ), .B(new_n8544), .Y(new_n8823));
  INVx1_ASAP7_75t_L         g08567(.A(\a[55] ), .Y(new_n8824));
  NAND2xp33_ASAP7_75t_L     g08568(.A(\a[56] ), .B(new_n8824), .Y(new_n8825));
  INVx1_ASAP7_75t_L         g08569(.A(\a[56] ), .Y(new_n8826));
  NAND2xp33_ASAP7_75t_L     g08570(.A(\a[55] ), .B(new_n8826), .Y(new_n8827));
  AOI21xp33_ASAP7_75t_L     g08571(.A1(new_n8827), .A2(new_n8825), .B(new_n8543), .Y(new_n8828));
  NAND2xp33_ASAP7_75t_L     g08572(.A(new_n269), .B(new_n8828), .Y(new_n8829));
  NAND2xp33_ASAP7_75t_L     g08573(.A(new_n8827), .B(new_n8825), .Y(new_n8830));
  NOR2xp33_ASAP7_75t_L      g08574(.A(new_n8830), .B(new_n8543), .Y(new_n8831));
  NAND2xp33_ASAP7_75t_L     g08575(.A(\b[1] ), .B(new_n8831), .Y(new_n8832));
  NAND2xp33_ASAP7_75t_L     g08576(.A(new_n8542), .B(new_n8541), .Y(new_n8833));
  XNOR2x2_ASAP7_75t_L       g08577(.A(\a[55] ), .B(\a[54] ), .Y(new_n8834));
  NOR2xp33_ASAP7_75t_L      g08578(.A(new_n8834), .B(new_n8833), .Y(new_n8835));
  NAND2xp33_ASAP7_75t_L     g08579(.A(\b[0] ), .B(new_n8835), .Y(new_n8836));
  NAND3xp33_ASAP7_75t_L     g08580(.A(new_n8829), .B(new_n8832), .C(new_n8836), .Y(new_n8837));
  XOR2x2_ASAP7_75t_L        g08581(.A(new_n8823), .B(new_n8837), .Y(new_n8838));
  NAND3xp33_ASAP7_75t_L     g08582(.A(new_n8822), .B(new_n8820), .C(new_n8838), .Y(new_n8839));
  INVx1_ASAP7_75t_L         g08583(.A(new_n8820), .Y(new_n8840));
  XNOR2x2_ASAP7_75t_L       g08584(.A(new_n8823), .B(new_n8837), .Y(new_n8841));
  OAI21xp33_ASAP7_75t_L     g08585(.A1(new_n8821), .A2(new_n8840), .B(new_n8841), .Y(new_n8842));
  NAND3xp33_ASAP7_75t_L     g08586(.A(new_n8816), .B(new_n8839), .C(new_n8842), .Y(new_n8843));
  NOR2xp33_ASAP7_75t_L      g08587(.A(new_n8534), .B(new_n8539), .Y(new_n8844));
  NAND2xp33_ASAP7_75t_L     g08588(.A(new_n8552), .B(new_n8554), .Y(new_n8845));
  MAJIxp5_ASAP7_75t_L       g08589(.A(new_n8845), .B(new_n8544), .C(new_n8844), .Y(new_n8846));
  NOR3xp33_ASAP7_75t_L      g08590(.A(new_n8840), .B(new_n8821), .C(new_n8841), .Y(new_n8847));
  AOI21xp33_ASAP7_75t_L     g08591(.A1(new_n8822), .A2(new_n8820), .B(new_n8838), .Y(new_n8848));
  OAI21xp33_ASAP7_75t_L     g08592(.A1(new_n8847), .A2(new_n8848), .B(new_n8846), .Y(new_n8849));
  AOI21xp33_ASAP7_75t_L     g08593(.A1(new_n8849), .A2(new_n8843), .B(new_n8813), .Y(new_n8850));
  NOR3xp33_ASAP7_75t_L      g08594(.A(new_n8846), .B(new_n8847), .C(new_n8848), .Y(new_n8851));
  AOI21xp33_ASAP7_75t_L     g08595(.A1(new_n8842), .A2(new_n8839), .B(new_n8816), .Y(new_n8852));
  NOR3xp33_ASAP7_75t_L      g08596(.A(new_n8851), .B(new_n8852), .C(new_n8812), .Y(new_n8853));
  AOI211xp5_ASAP7_75t_L     g08597(.A1(new_n8579), .A2(new_n8809), .B(new_n8850), .C(new_n8853), .Y(new_n8854));
  OAI21xp33_ASAP7_75t_L     g08598(.A1(new_n8852), .A2(new_n8851), .B(new_n8812), .Y(new_n8855));
  NAND3xp33_ASAP7_75t_L     g08599(.A(new_n8813), .B(new_n8843), .C(new_n8849), .Y(new_n8856));
  AOI211xp5_ASAP7_75t_L     g08600(.A1(new_n8856), .A2(new_n8855), .B(new_n8571), .C(new_n8808), .Y(new_n8857));
  OAI21xp33_ASAP7_75t_L     g08601(.A1(new_n8854), .A2(new_n8857), .B(new_n8807), .Y(new_n8858));
  OAI211xp5_ASAP7_75t_L     g08602(.A1(new_n8571), .A2(new_n8808), .B(new_n8856), .C(new_n8855), .Y(new_n8859));
  AOI21xp33_ASAP7_75t_L     g08603(.A1(new_n8236), .A2(new_n8254), .B(new_n8253), .Y(new_n8860));
  O2A1O1Ixp33_ASAP7_75t_L   g08604(.A1(new_n8576), .A2(new_n8577), .B(new_n8860), .C(new_n8808), .Y(new_n8861));
  OAI21xp33_ASAP7_75t_L     g08605(.A1(new_n8850), .A2(new_n8853), .B(new_n8861), .Y(new_n8862));
  NAND3xp33_ASAP7_75t_L     g08606(.A(new_n8862), .B(new_n8859), .C(new_n8806), .Y(new_n8863));
  NAND3xp33_ASAP7_75t_L     g08607(.A(new_n8803), .B(new_n8858), .C(new_n8863), .Y(new_n8864));
  NAND2xp33_ASAP7_75t_L     g08608(.A(new_n8863), .B(new_n8858), .Y(new_n8865));
  NAND3xp33_ASAP7_75t_L     g08609(.A(new_n8588), .B(new_n8802), .C(new_n8865), .Y(new_n8866));
  AOI21xp33_ASAP7_75t_L     g08610(.A1(new_n8866), .A2(new_n8864), .B(new_n8800), .Y(new_n8867));
  INVx1_ASAP7_75t_L         g08611(.A(new_n8587), .Y(new_n8868));
  O2A1O1Ixp33_ASAP7_75t_L   g08612(.A1(new_n8528), .A2(new_n8868), .B(new_n8802), .C(new_n8865), .Y(new_n8869));
  AOI21xp33_ASAP7_75t_L     g08613(.A1(new_n8863), .A2(new_n8858), .B(new_n8803), .Y(new_n8870));
  NOR3xp33_ASAP7_75t_L      g08614(.A(new_n8869), .B(new_n8870), .C(new_n8799), .Y(new_n8871));
  NOR2xp33_ASAP7_75t_L      g08615(.A(new_n8871), .B(new_n8867), .Y(new_n8872));
  NAND2xp33_ASAP7_75t_L     g08616(.A(new_n8796), .B(new_n8872), .Y(new_n8873));
  INVx1_ASAP7_75t_L         g08617(.A(new_n8795), .Y(new_n8874));
  OAI21xp33_ASAP7_75t_L     g08618(.A1(new_n8870), .A2(new_n8869), .B(new_n8799), .Y(new_n8875));
  NAND3xp33_ASAP7_75t_L     g08619(.A(new_n8866), .B(new_n8864), .C(new_n8800), .Y(new_n8876));
  AO221x2_ASAP7_75t_L       g08620(.A1(new_n8591), .A2(new_n8522), .B1(new_n8875), .B2(new_n8876), .C(new_n8874), .Y(new_n8877));
  AOI22xp33_ASAP7_75t_L     g08621(.A1(new_n4920), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n5167), .Y(new_n8878));
  OAI221xp5_ASAP7_75t_L     g08622(.A1(new_n5154), .A2(new_n942), .B1(new_n5158), .B2(new_n1035), .C(new_n8878), .Y(new_n8879));
  XNOR2x2_ASAP7_75t_L       g08623(.A(\a[41] ), .B(new_n8879), .Y(new_n8880));
  NAND3xp33_ASAP7_75t_L     g08624(.A(new_n8873), .B(new_n8877), .C(new_n8880), .Y(new_n8881));
  NAND2xp33_ASAP7_75t_L     g08625(.A(new_n8589), .B(new_n8588), .Y(new_n8882));
  NAND2xp33_ASAP7_75t_L     g08626(.A(new_n8876), .B(new_n8875), .Y(new_n8883));
  O2A1O1Ixp33_ASAP7_75t_L   g08627(.A1(new_n8586), .A2(new_n8882), .B(new_n8592), .C(new_n8883), .Y(new_n8884));
  NOR2xp33_ASAP7_75t_L      g08628(.A(new_n8796), .B(new_n8872), .Y(new_n8885));
  INVx1_ASAP7_75t_L         g08629(.A(new_n8880), .Y(new_n8886));
  OAI21xp33_ASAP7_75t_L     g08630(.A1(new_n8885), .A2(new_n8884), .B(new_n8886), .Y(new_n8887));
  NOR3xp33_ASAP7_75t_L      g08631(.A(new_n8597), .B(new_n8596), .C(new_n8519), .Y(new_n8888));
  A2O1A1O1Ixp25_ASAP7_75t_L g08632(.A1(new_n8290), .A2(new_n8289), .B(new_n8515), .C(new_n8598), .D(new_n8888), .Y(new_n8889));
  AND3x1_ASAP7_75t_L        g08633(.A(new_n8889), .B(new_n8887), .C(new_n8881), .Y(new_n8890));
  AOI21xp33_ASAP7_75t_L     g08634(.A1(new_n8887), .A2(new_n8881), .B(new_n8889), .Y(new_n8891));
  AOI22xp33_ASAP7_75t_L     g08635(.A1(new_n4283), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n4512), .Y(new_n8892));
  OAI221xp5_ASAP7_75t_L     g08636(.A1(new_n4277), .A2(new_n1313), .B1(new_n4499), .B2(new_n1438), .C(new_n8892), .Y(new_n8893));
  XNOR2x2_ASAP7_75t_L       g08637(.A(\a[38] ), .B(new_n8893), .Y(new_n8894));
  OAI21xp33_ASAP7_75t_L     g08638(.A1(new_n8891), .A2(new_n8890), .B(new_n8894), .Y(new_n8895));
  NAND3xp33_ASAP7_75t_L     g08639(.A(new_n8889), .B(new_n8887), .C(new_n8881), .Y(new_n8896));
  NAND2xp33_ASAP7_75t_L     g08640(.A(new_n8881), .B(new_n8887), .Y(new_n8897));
  A2O1A1Ixp33_ASAP7_75t_L   g08641(.A1(new_n8598), .A2(new_n8604), .B(new_n8888), .C(new_n8897), .Y(new_n8898));
  INVx1_ASAP7_75t_L         g08642(.A(new_n8894), .Y(new_n8899));
  NAND3xp33_ASAP7_75t_L     g08643(.A(new_n8898), .B(new_n8896), .C(new_n8899), .Y(new_n8900));
  NAND2xp33_ASAP7_75t_L     g08644(.A(new_n8895), .B(new_n8900), .Y(new_n8901));
  NAND3xp33_ASAP7_75t_L     g08645(.A(new_n8616), .B(new_n8901), .C(new_n8794), .Y(new_n8902));
  A2O1A1Ixp33_ASAP7_75t_L   g08646(.A1(new_n8602), .A2(new_n8607), .B(new_n8511), .C(new_n8794), .Y(new_n8903));
  AOI21xp33_ASAP7_75t_L     g08647(.A1(new_n8898), .A2(new_n8896), .B(new_n8899), .Y(new_n8904));
  NOR3xp33_ASAP7_75t_L      g08648(.A(new_n8890), .B(new_n8891), .C(new_n8894), .Y(new_n8905));
  NOR2xp33_ASAP7_75t_L      g08649(.A(new_n8905), .B(new_n8904), .Y(new_n8906));
  NAND2xp33_ASAP7_75t_L     g08650(.A(new_n8903), .B(new_n8906), .Y(new_n8907));
  NAND3xp33_ASAP7_75t_L     g08651(.A(new_n8902), .B(new_n8907), .C(new_n8793), .Y(new_n8908));
  NOR2xp33_ASAP7_75t_L      g08652(.A(new_n8903), .B(new_n8906), .Y(new_n8909));
  O2A1O1Ixp33_ASAP7_75t_L   g08653(.A1(new_n8511), .A2(new_n8619), .B(new_n8794), .C(new_n8901), .Y(new_n8910));
  OAI21xp33_ASAP7_75t_L     g08654(.A1(new_n8909), .A2(new_n8910), .B(new_n8792), .Y(new_n8911));
  AOI21xp33_ASAP7_75t_L     g08655(.A1(new_n8911), .A2(new_n8908), .B(new_n8789), .Y(new_n8912));
  AOI21xp33_ASAP7_75t_L     g08656(.A1(new_n7937), .A2(new_n8037), .B(new_n8032), .Y(new_n8913));
  A2O1A1O1Ixp25_ASAP7_75t_L g08657(.A1(new_n8308), .A2(new_n8913), .B(new_n8505), .C(new_n8628), .D(new_n8612), .Y(new_n8914));
  NOR3xp33_ASAP7_75t_L      g08658(.A(new_n8910), .B(new_n8909), .C(new_n8792), .Y(new_n8915));
  AOI21xp33_ASAP7_75t_L     g08659(.A1(new_n8902), .A2(new_n8907), .B(new_n8793), .Y(new_n8916));
  NOR3xp33_ASAP7_75t_L      g08660(.A(new_n8914), .B(new_n8915), .C(new_n8916), .Y(new_n8917));
  OAI22xp33_ASAP7_75t_L     g08661(.A1(new_n3402), .A2(new_n1909), .B1(new_n2067), .B2(new_n3022), .Y(new_n8918));
  AOI221xp5_ASAP7_75t_L     g08662(.A1(new_n3030), .A2(\b[24] ), .B1(new_n3021), .B2(new_n2648), .C(new_n8918), .Y(new_n8919));
  XNOR2x2_ASAP7_75t_L       g08663(.A(\a[32] ), .B(new_n8919), .Y(new_n8920));
  NOR3xp33_ASAP7_75t_L      g08664(.A(new_n8917), .B(new_n8912), .C(new_n8920), .Y(new_n8921));
  OAI21xp33_ASAP7_75t_L     g08665(.A1(new_n8916), .A2(new_n8915), .B(new_n8914), .Y(new_n8922));
  NAND3xp33_ASAP7_75t_L     g08666(.A(new_n8789), .B(new_n8911), .C(new_n8908), .Y(new_n8923));
  XNOR2x2_ASAP7_75t_L       g08667(.A(new_n3015), .B(new_n8919), .Y(new_n8924));
  AOI21xp33_ASAP7_75t_L     g08668(.A1(new_n8922), .A2(new_n8923), .B(new_n8924), .Y(new_n8925));
  NOR2xp33_ASAP7_75t_L      g08669(.A(new_n8925), .B(new_n8921), .Y(new_n8926));
  AO21x2_ASAP7_75t_L        g08670(.A1(new_n8043), .A2(new_n8054), .B(new_n8046), .Y(new_n8927));
  A2O1A1O1Ixp25_ASAP7_75t_L g08671(.A1(new_n8320), .A2(new_n8927), .B(new_n8643), .C(new_n8630), .D(new_n8636), .Y(new_n8928));
  NAND2xp33_ASAP7_75t_L     g08672(.A(new_n8926), .B(new_n8928), .Y(new_n8929));
  NAND3xp33_ASAP7_75t_L     g08673(.A(new_n8922), .B(new_n8923), .C(new_n8924), .Y(new_n8930));
  OAI21xp33_ASAP7_75t_L     g08674(.A1(new_n8912), .A2(new_n8917), .B(new_n8920), .Y(new_n8931));
  NAND2xp33_ASAP7_75t_L     g08675(.A(new_n8930), .B(new_n8931), .Y(new_n8932));
  A2O1A1Ixp33_ASAP7_75t_L   g08676(.A1(new_n8638), .A2(new_n8635), .B(new_n8636), .C(new_n8932), .Y(new_n8933));
  AOI22xp33_ASAP7_75t_L     g08677(.A1(new_n2552), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n2736), .Y(new_n8934));
  OAI221xp5_ASAP7_75t_L     g08678(.A1(new_n2547), .A2(new_n2497), .B1(new_n2734), .B2(new_n2672), .C(new_n8934), .Y(new_n8935));
  XNOR2x2_ASAP7_75t_L       g08679(.A(\a[29] ), .B(new_n8935), .Y(new_n8936));
  NAND3xp33_ASAP7_75t_L     g08680(.A(new_n8929), .B(new_n8933), .C(new_n8936), .Y(new_n8937));
  AOI211xp5_ASAP7_75t_L     g08681(.A1(new_n8638), .A2(new_n8635), .B(new_n8636), .C(new_n8932), .Y(new_n8938));
  O2A1O1Ixp33_ASAP7_75t_L   g08682(.A1(new_n8644), .A2(new_n8637), .B(new_n8624), .C(new_n8926), .Y(new_n8939));
  INVx1_ASAP7_75t_L         g08683(.A(new_n8936), .Y(new_n8940));
  OAI21xp33_ASAP7_75t_L     g08684(.A1(new_n8939), .A2(new_n8938), .B(new_n8940), .Y(new_n8941));
  NAND2xp33_ASAP7_75t_L     g08685(.A(new_n8937), .B(new_n8941), .Y(new_n8942));
  OAI21xp33_ASAP7_75t_L     g08686(.A1(new_n8646), .A2(new_n8651), .B(new_n8655), .Y(new_n8943));
  NOR2xp33_ASAP7_75t_L      g08687(.A(new_n8942), .B(new_n8943), .Y(new_n8944));
  A2O1A1O1Ixp25_ASAP7_75t_L g08688(.A1(new_n8322), .A2(new_n8210), .B(new_n8496), .C(new_n8656), .D(new_n8640), .Y(new_n8945));
  AOI21xp33_ASAP7_75t_L     g08689(.A1(new_n8941), .A2(new_n8937), .B(new_n8945), .Y(new_n8946));
  AOI22xp33_ASAP7_75t_L     g08690(.A1(new_n2114), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n2259), .Y(new_n8947));
  OAI221xp5_ASAP7_75t_L     g08691(.A1(new_n2109), .A2(new_n2982), .B1(new_n2257), .B2(new_n3187), .C(new_n8947), .Y(new_n8948));
  XNOR2x2_ASAP7_75t_L       g08692(.A(\a[26] ), .B(new_n8948), .Y(new_n8949));
  INVx1_ASAP7_75t_L         g08693(.A(new_n8949), .Y(new_n8950));
  NOR3xp33_ASAP7_75t_L      g08694(.A(new_n8944), .B(new_n8946), .C(new_n8950), .Y(new_n8951));
  NAND3xp33_ASAP7_75t_L     g08695(.A(new_n8945), .B(new_n8941), .C(new_n8937), .Y(new_n8952));
  NAND2xp33_ASAP7_75t_L     g08696(.A(new_n8942), .B(new_n8943), .Y(new_n8953));
  AOI21xp33_ASAP7_75t_L     g08697(.A1(new_n8953), .A2(new_n8952), .B(new_n8949), .Y(new_n8954));
  NOR2xp33_ASAP7_75t_L      g08698(.A(new_n8954), .B(new_n8951), .Y(new_n8955));
  A2O1A1O1Ixp25_ASAP7_75t_L g08699(.A1(new_n8338), .A2(new_n8342), .B(new_n8336), .C(new_n8658), .D(new_n8661), .Y(new_n8956));
  NAND2xp33_ASAP7_75t_L     g08700(.A(new_n8956), .B(new_n8955), .Y(new_n8957));
  NAND3xp33_ASAP7_75t_L     g08701(.A(new_n8953), .B(new_n8952), .C(new_n8949), .Y(new_n8958));
  OAI21xp33_ASAP7_75t_L     g08702(.A1(new_n8946), .A2(new_n8944), .B(new_n8950), .Y(new_n8959));
  NAND2xp33_ASAP7_75t_L     g08703(.A(new_n8958), .B(new_n8959), .Y(new_n8960));
  A2O1A1Ixp33_ASAP7_75t_L   g08704(.A1(new_n8658), .A2(new_n8491), .B(new_n8661), .C(new_n8960), .Y(new_n8961));
  AOI22xp33_ASAP7_75t_L     g08705(.A1(new_n1704), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1837), .Y(new_n8962));
  OAI221xp5_ASAP7_75t_L     g08706(.A1(new_n1699), .A2(new_n3565), .B1(new_n1827), .B2(new_n3591), .C(new_n8962), .Y(new_n8963));
  XNOR2x2_ASAP7_75t_L       g08707(.A(\a[23] ), .B(new_n8963), .Y(new_n8964));
  NAND3xp33_ASAP7_75t_L     g08708(.A(new_n8961), .B(new_n8957), .C(new_n8964), .Y(new_n8965));
  OAI21xp33_ASAP7_75t_L     g08709(.A1(new_n8662), .A2(new_n8660), .B(new_n8653), .Y(new_n8966));
  NOR2xp33_ASAP7_75t_L      g08710(.A(new_n8966), .B(new_n8960), .Y(new_n8967));
  O2A1O1Ixp33_ASAP7_75t_L   g08711(.A1(new_n8660), .A2(new_n8662), .B(new_n8653), .C(new_n8955), .Y(new_n8968));
  INVx1_ASAP7_75t_L         g08712(.A(new_n8964), .Y(new_n8969));
  OAI21xp33_ASAP7_75t_L     g08713(.A1(new_n8967), .A2(new_n8968), .B(new_n8969), .Y(new_n8970));
  NOR2xp33_ASAP7_75t_L      g08714(.A(new_n8670), .B(new_n8669), .Y(new_n8971));
  MAJIxp5_ASAP7_75t_L       g08715(.A(new_n8680), .B(new_n8971), .C(new_n8671), .Y(new_n8972));
  NAND3xp33_ASAP7_75t_L     g08716(.A(new_n8972), .B(new_n8970), .C(new_n8965), .Y(new_n8973));
  NOR3xp33_ASAP7_75t_L      g08717(.A(new_n8968), .B(new_n8967), .C(new_n8969), .Y(new_n8974));
  AOI21xp33_ASAP7_75t_L     g08718(.A1(new_n8961), .A2(new_n8957), .B(new_n8964), .Y(new_n8975));
  NAND2xp33_ASAP7_75t_L     g08719(.A(new_n8671), .B(new_n8971), .Y(new_n8976));
  A2O1A1Ixp33_ASAP7_75t_L   g08720(.A1(new_n8668), .A2(new_n8672), .B(new_n8675), .C(new_n8976), .Y(new_n8977));
  OAI21xp33_ASAP7_75t_L     g08721(.A1(new_n8975), .A2(new_n8974), .B(new_n8977), .Y(new_n8978));
  AOI22xp33_ASAP7_75t_L     g08722(.A1(new_n1360), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1581), .Y(new_n8979));
  OAI221xp5_ASAP7_75t_L     g08723(.A1(new_n1373), .A2(new_n4216), .B1(new_n1359), .B2(new_n4431), .C(new_n8979), .Y(new_n8980));
  XNOR2x2_ASAP7_75t_L       g08724(.A(\a[20] ), .B(new_n8980), .Y(new_n8981));
  NAND3xp33_ASAP7_75t_L     g08725(.A(new_n8973), .B(new_n8978), .C(new_n8981), .Y(new_n8982));
  AO21x2_ASAP7_75t_L        g08726(.A1(new_n8978), .A2(new_n8973), .B(new_n8981), .Y(new_n8983));
  NOR3xp33_ASAP7_75t_L      g08727(.A(new_n8681), .B(new_n8678), .C(new_n8489), .Y(new_n8984));
  A2O1A1O1Ixp25_ASAP7_75t_L g08728(.A1(new_n8370), .A2(new_n8381), .B(new_n8485), .C(new_n8682), .D(new_n8984), .Y(new_n8985));
  NAND3xp33_ASAP7_75t_L     g08729(.A(new_n8985), .B(new_n8983), .C(new_n8982), .Y(new_n8986));
  AO21x2_ASAP7_75t_L        g08730(.A1(new_n8982), .A2(new_n8983), .B(new_n8985), .Y(new_n8987));
  NAND2xp33_ASAP7_75t_L     g08731(.A(\b[39] ), .B(new_n1080), .Y(new_n8988));
  NAND2xp33_ASAP7_75t_L     g08732(.A(new_n1073), .B(new_n4876), .Y(new_n8989));
  AOI22xp33_ASAP7_75t_L     g08733(.A1(new_n1076), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n1253), .Y(new_n8990));
  AND4x1_ASAP7_75t_L        g08734(.A(new_n8990), .B(new_n8989), .C(new_n8988), .D(\a[17] ), .Y(new_n8991));
  AOI31xp33_ASAP7_75t_L     g08735(.A1(new_n8989), .A2(new_n8988), .A3(new_n8990), .B(\a[17] ), .Y(new_n8992));
  NOR2xp33_ASAP7_75t_L      g08736(.A(new_n8992), .B(new_n8991), .Y(new_n8993));
  NAND3xp33_ASAP7_75t_L     g08737(.A(new_n8987), .B(new_n8986), .C(new_n8993), .Y(new_n8994));
  AND3x1_ASAP7_75t_L        g08738(.A(new_n8985), .B(new_n8983), .C(new_n8982), .Y(new_n8995));
  AOI21xp33_ASAP7_75t_L     g08739(.A1(new_n8983), .A2(new_n8982), .B(new_n8985), .Y(new_n8996));
  OAI22xp33_ASAP7_75t_L     g08740(.A1(new_n8995), .A2(new_n8996), .B1(new_n8992), .B2(new_n8991), .Y(new_n8997));
  NAND2xp33_ASAP7_75t_L     g08741(.A(new_n8994), .B(new_n8997), .Y(new_n8998));
  NAND3xp33_ASAP7_75t_L     g08742(.A(new_n8685), .B(new_n8684), .C(new_n8692), .Y(new_n8999));
  A2O1A1Ixp33_ASAP7_75t_L   g08743(.A1(new_n8693), .A2(new_n8689), .B(new_n8695), .C(new_n8999), .Y(new_n9000));
  XOR2x2_ASAP7_75t_L        g08744(.A(new_n8998), .B(new_n9000), .Y(new_n9001));
  AOI22xp33_ASAP7_75t_L     g08745(.A1(new_n811), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n900), .Y(new_n9002));
  OAI221xp5_ASAP7_75t_L     g08746(.A1(new_n904), .A2(new_n5338), .B1(new_n898), .B2(new_n6338), .C(new_n9002), .Y(new_n9003));
  XNOR2x2_ASAP7_75t_L       g08747(.A(\a[14] ), .B(new_n9003), .Y(new_n9004));
  INVx1_ASAP7_75t_L         g08748(.A(new_n9004), .Y(new_n9005));
  NOR2xp33_ASAP7_75t_L      g08749(.A(new_n9005), .B(new_n9001), .Y(new_n9006));
  NOR2xp33_ASAP7_75t_L      g08750(.A(new_n8998), .B(new_n9000), .Y(new_n9007));
  AOI22xp33_ASAP7_75t_L     g08751(.A1(new_n8994), .A2(new_n8997), .B1(new_n8999), .B2(new_n8698), .Y(new_n9008));
  NOR3xp33_ASAP7_75t_L      g08752(.A(new_n9008), .B(new_n9004), .C(new_n9007), .Y(new_n9009));
  OA21x2_ASAP7_75t_L        g08753(.A1(new_n9009), .A2(new_n9006), .B(new_n8788), .Y(new_n9010));
  NOR3xp33_ASAP7_75t_L      g08754(.A(new_n9006), .B(new_n8788), .C(new_n9009), .Y(new_n9011));
  OA21x2_ASAP7_75t_L        g08755(.A1(new_n9011), .A2(new_n9010), .B(new_n8787), .Y(new_n9012));
  NOR3xp33_ASAP7_75t_L      g08756(.A(new_n9010), .B(new_n9011), .C(new_n8787), .Y(new_n9013));
  NOR3xp33_ASAP7_75t_L      g08757(.A(new_n8780), .B(new_n9012), .C(new_n9013), .Y(new_n9014));
  NAND2xp33_ASAP7_75t_L     g08758(.A(new_n8716), .B(new_n8711), .Y(new_n9015));
  MAJIxp5_ASAP7_75t_L       g08759(.A(new_n8727), .B(new_n8481), .C(new_n9015), .Y(new_n9016));
  OAI21xp33_ASAP7_75t_L     g08760(.A1(new_n9011), .A2(new_n9010), .B(new_n8787), .Y(new_n9017));
  OR3x1_ASAP7_75t_L         g08761(.A(new_n9010), .B(new_n8787), .C(new_n9011), .Y(new_n9018));
  AOI21xp33_ASAP7_75t_L     g08762(.A1(new_n9018), .A2(new_n9017), .B(new_n9016), .Y(new_n9019));
  OAI21xp33_ASAP7_75t_L     g08763(.A1(new_n9019), .A2(new_n9014), .B(new_n8778), .Y(new_n9020));
  INVx1_ASAP7_75t_L         g08764(.A(new_n8778), .Y(new_n9021));
  NAND3xp33_ASAP7_75t_L     g08765(.A(new_n9016), .B(new_n9018), .C(new_n9017), .Y(new_n9022));
  OAI21xp33_ASAP7_75t_L     g08766(.A1(new_n9013), .A2(new_n9012), .B(new_n8780), .Y(new_n9023));
  NAND3xp33_ASAP7_75t_L     g08767(.A(new_n9022), .B(new_n9023), .C(new_n9021), .Y(new_n9024));
  NAND3xp33_ASAP7_75t_L     g08768(.A(new_n8775), .B(new_n9020), .C(new_n9024), .Y(new_n9025));
  O2A1O1Ixp33_ASAP7_75t_L   g08769(.A1(new_n8738), .A2(new_n8739), .B(new_n8736), .C(new_n8773), .Y(new_n9026));
  NAND2xp33_ASAP7_75t_L     g08770(.A(new_n9024), .B(new_n9020), .Y(new_n9027));
  NAND2xp33_ASAP7_75t_L     g08771(.A(new_n9026), .B(new_n9027), .Y(new_n9028));
  AOI22xp33_ASAP7_75t_L     g08772(.A1(new_n344), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n370), .Y(new_n9029));
  OAI221xp5_ASAP7_75t_L     g08773(.A1(new_n429), .A2(new_n7616), .B1(new_n366), .B2(new_n7906), .C(new_n9029), .Y(new_n9030));
  XNOR2x2_ASAP7_75t_L       g08774(.A(\a[5] ), .B(new_n9030), .Y(new_n9031));
  NAND3xp33_ASAP7_75t_L     g08775(.A(new_n9025), .B(new_n9028), .C(new_n9031), .Y(new_n9032));
  NOR2xp33_ASAP7_75t_L      g08776(.A(new_n9026), .B(new_n9027), .Y(new_n9033));
  AOI221xp5_ASAP7_75t_L     g08777(.A1(new_n8734), .A2(new_n8736), .B1(new_n9024), .B2(new_n9020), .C(new_n8773), .Y(new_n9034));
  INVx1_ASAP7_75t_L         g08778(.A(new_n9031), .Y(new_n9035));
  OAI21xp33_ASAP7_75t_L     g08779(.A1(new_n9034), .A2(new_n9033), .B(new_n9035), .Y(new_n9036));
  AOI21xp33_ASAP7_75t_L     g08780(.A1(new_n9036), .A2(new_n9032), .B(new_n8772), .Y(new_n9037));
  AND3x1_ASAP7_75t_L        g08781(.A(new_n8772), .B(new_n9036), .C(new_n9032), .Y(new_n9038));
  NOR3xp33_ASAP7_75t_L      g08782(.A(new_n9038), .B(new_n9037), .C(new_n8771), .Y(new_n9039));
  INVx1_ASAP7_75t_L         g08783(.A(new_n9039), .Y(new_n9040));
  OAI21xp33_ASAP7_75t_L     g08784(.A1(new_n9037), .A2(new_n9038), .B(new_n8771), .Y(new_n9041));
  NAND2xp33_ASAP7_75t_L     g08785(.A(new_n9041), .B(new_n9040), .Y(new_n9042));
  O2A1O1Ixp33_ASAP7_75t_L   g08786(.A1(new_n8760), .A2(new_n8758), .B(new_n8756), .C(new_n9042), .Y(new_n9043));
  AOI221xp5_ASAP7_75t_L     g08787(.A1(new_n8757), .A2(new_n8455), .B1(new_n9041), .B2(new_n9040), .C(new_n8755), .Y(new_n9044));
  NOR2xp33_ASAP7_75t_L      g08788(.A(new_n9044), .B(new_n9043), .Y(\f[55] ));
  XNOR2x2_ASAP7_75t_L       g08789(.A(new_n9026), .B(new_n9027), .Y(new_n9046));
  MAJIxp5_ASAP7_75t_L       g08790(.A(new_n8772), .B(new_n9031), .C(new_n9046), .Y(new_n9047));
  NAND2xp33_ASAP7_75t_L     g08791(.A(\b[52] ), .B(new_n347), .Y(new_n9048));
  NAND2xp33_ASAP7_75t_L     g08792(.A(new_n341), .B(new_n8173), .Y(new_n9049));
  AOI22xp33_ASAP7_75t_L     g08793(.A1(new_n344), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n370), .Y(new_n9050));
  AND4x1_ASAP7_75t_L        g08794(.A(new_n9050), .B(new_n9049), .C(new_n9048), .D(\a[5] ), .Y(new_n9051));
  AOI31xp33_ASAP7_75t_L     g08795(.A1(new_n9049), .A2(new_n9048), .A3(new_n9050), .B(\a[5] ), .Y(new_n9052));
  NOR2xp33_ASAP7_75t_L      g08796(.A(new_n9052), .B(new_n9051), .Y(new_n9053));
  NOR3xp33_ASAP7_75t_L      g08797(.A(new_n9014), .B(new_n9019), .C(new_n8778), .Y(new_n9054));
  A2O1A1O1Ixp25_ASAP7_75t_L g08798(.A1(new_n8736), .A2(new_n8734), .B(new_n8773), .C(new_n9020), .D(new_n9054), .Y(new_n9055));
  NAND2xp33_ASAP7_75t_L     g08799(.A(\b[48] ), .B(new_n471), .Y(new_n9056));
  OAI221xp5_ASAP7_75t_L     g08800(.A1(new_n515), .A2(new_n7593), .B1(new_n469), .B2(new_n7602), .C(new_n9056), .Y(new_n9057));
  AOI21xp33_ASAP7_75t_L     g08801(.A1(new_n447), .A2(\b[49] ), .B(new_n9057), .Y(new_n9058));
  NAND2xp33_ASAP7_75t_L     g08802(.A(\a[8] ), .B(new_n9058), .Y(new_n9059));
  A2O1A1Ixp33_ASAP7_75t_L   g08803(.A1(\b[49] ), .A2(new_n447), .B(new_n9057), .C(new_n435), .Y(new_n9060));
  AND2x2_ASAP7_75t_L        g08804(.A(new_n9060), .B(new_n9059), .Y(new_n9061));
  NAND2xp33_ASAP7_75t_L     g08805(.A(new_n8718), .B(new_n8779), .Y(new_n9062));
  A2O1A1Ixp33_ASAP7_75t_L   g08806(.A1(new_n8724), .A2(new_n9062), .B(new_n9012), .C(new_n9018), .Y(new_n9063));
  AOI22xp33_ASAP7_75t_L     g08807(.A1(\b[45] ), .A2(new_n651), .B1(\b[47] ), .B2(new_n581), .Y(new_n9064));
  OAI221xp5_ASAP7_75t_L     g08808(.A1(new_n821), .A2(new_n6568), .B1(new_n577), .B2(new_n6820), .C(new_n9064), .Y(new_n9065));
  XNOR2x2_ASAP7_75t_L       g08809(.A(\a[11] ), .B(new_n9065), .Y(new_n9066));
  NAND2xp33_ASAP7_75t_L     g08810(.A(new_n8952), .B(new_n8953), .Y(new_n9067));
  MAJIxp5_ASAP7_75t_L       g08811(.A(new_n8956), .B(new_n8949), .C(new_n9067), .Y(new_n9068));
  NOR2xp33_ASAP7_75t_L      g08812(.A(new_n3180), .B(new_n2109), .Y(new_n9069));
  INVx1_ASAP7_75t_L         g08813(.A(new_n9069), .Y(new_n9070));
  NAND3xp33_ASAP7_75t_L     g08814(.A(new_n3210), .B(new_n2106), .C(new_n3213), .Y(new_n9071));
  AOI22xp33_ASAP7_75t_L     g08815(.A1(new_n2114), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n2259), .Y(new_n9072));
  AND4x1_ASAP7_75t_L        g08816(.A(new_n9072), .B(new_n9071), .C(new_n9070), .D(\a[26] ), .Y(new_n9073));
  AOI31xp33_ASAP7_75t_L     g08817(.A1(new_n9071), .A2(new_n9070), .A3(new_n9072), .B(\a[26] ), .Y(new_n9074));
  NOR2xp33_ASAP7_75t_L      g08818(.A(new_n9074), .B(new_n9073), .Y(new_n9075));
  NAND2xp33_ASAP7_75t_L     g08819(.A(new_n8933), .B(new_n8929), .Y(new_n9076));
  AOI22xp33_ASAP7_75t_L     g08820(.A1(new_n2552), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n2736), .Y(new_n9077));
  OAI221xp5_ASAP7_75t_L     g08821(.A1(new_n2547), .A2(new_n2666), .B1(new_n2734), .B2(new_n2695), .C(new_n9077), .Y(new_n9078));
  NOR2xp33_ASAP7_75t_L      g08822(.A(new_n2538), .B(new_n9078), .Y(new_n9079));
  AND2x2_ASAP7_75t_L        g08823(.A(new_n2538), .B(new_n9078), .Y(new_n9080));
  NOR2xp33_ASAP7_75t_L      g08824(.A(new_n9079), .B(new_n9080), .Y(new_n9081));
  NAND3xp33_ASAP7_75t_L     g08825(.A(new_n8923), .B(new_n8922), .C(new_n8920), .Y(new_n9082));
  A2O1A1Ixp33_ASAP7_75t_L   g08826(.A1(new_n8931), .A2(new_n8930), .B(new_n8928), .C(new_n9082), .Y(new_n9083));
  AOI21xp33_ASAP7_75t_L     g08827(.A1(new_n8789), .A2(new_n8911), .B(new_n8915), .Y(new_n9084));
  AOI22xp33_ASAP7_75t_L     g08828(.A1(new_n3633), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n3858), .Y(new_n9085));
  OAI221xp5_ASAP7_75t_L     g08829(.A1(new_n3853), .A2(new_n1774), .B1(new_n3856), .B2(new_n1915), .C(new_n9085), .Y(new_n9086));
  XNOR2x2_ASAP7_75t_L       g08830(.A(\a[35] ), .B(new_n9086), .Y(new_n9087));
  NAND3xp33_ASAP7_75t_L     g08831(.A(new_n8873), .B(new_n8877), .C(new_n8886), .Y(new_n9088));
  AOI22xp33_ASAP7_75t_L     g08832(.A1(new_n4920), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n5167), .Y(new_n9089));
  OAI221xp5_ASAP7_75t_L     g08833(.A1(new_n5154), .A2(new_n1030), .B1(new_n5158), .B2(new_n1209), .C(new_n9089), .Y(new_n9090));
  XNOR2x2_ASAP7_75t_L       g08834(.A(\a[41] ), .B(new_n9090), .Y(new_n9091));
  INVx1_ASAP7_75t_L         g08835(.A(new_n9091), .Y(new_n9092));
  A2O1A1O1Ixp25_ASAP7_75t_L g08836(.A1(new_n8522), .A2(new_n8591), .B(new_n8874), .C(new_n8875), .D(new_n8871), .Y(new_n9093));
  INVx1_ASAP7_75t_L         g08837(.A(new_n8863), .Y(new_n9094));
  AOI22xp33_ASAP7_75t_L     g08838(.A1(new_n6376), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n6648), .Y(new_n9095));
  OAI221xp5_ASAP7_75t_L     g08839(.A1(new_n6646), .A2(new_n617), .B1(new_n6636), .B2(new_n685), .C(new_n9095), .Y(new_n9096));
  XNOR2x2_ASAP7_75t_L       g08840(.A(\a[47] ), .B(new_n9096), .Y(new_n9097));
  A2O1A1O1Ixp25_ASAP7_75t_L g08841(.A1(new_n8860), .A2(new_n8572), .B(new_n8808), .C(new_n8855), .D(new_n8853), .Y(new_n9098));
  AOI22xp33_ASAP7_75t_L     g08842(.A1(new_n7111), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n7391), .Y(new_n9099));
  OAI221xp5_ASAP7_75t_L     g08843(.A1(new_n8558), .A2(new_n420), .B1(new_n8237), .B2(new_n494), .C(new_n9099), .Y(new_n9100));
  XNOR2x2_ASAP7_75t_L       g08844(.A(new_n7106), .B(new_n9100), .Y(new_n9101));
  NAND2xp33_ASAP7_75t_L     g08845(.A(new_n8549), .B(new_n8545), .Y(new_n9102));
  A2O1A1O1Ixp25_ASAP7_75t_L g08846(.A1(new_n8845), .A2(new_n9102), .B(new_n8814), .C(new_n8839), .D(new_n8848), .Y(new_n9103));
  NAND2xp33_ASAP7_75t_L     g08847(.A(\b[4] ), .B(new_n7963), .Y(new_n9104));
  INVx1_ASAP7_75t_L         g08848(.A(new_n9104), .Y(new_n9105));
  NOR3xp33_ASAP7_75t_L      g08849(.A(new_n357), .B(new_n358), .C(new_n7957), .Y(new_n9106));
  OAI22xp33_ASAP7_75t_L     g08850(.A1(new_n8247), .A2(new_n298), .B1(new_n354), .B2(new_n8243), .Y(new_n9107));
  NOR3xp33_ASAP7_75t_L      g08851(.A(new_n9106), .B(new_n9107), .C(new_n9105), .Y(new_n9108));
  NAND2xp33_ASAP7_75t_L     g08852(.A(\a[53] ), .B(new_n9108), .Y(new_n9109));
  INVx1_ASAP7_75t_L         g08853(.A(new_n9109), .Y(new_n9110));
  NOR2xp33_ASAP7_75t_L      g08854(.A(\a[53] ), .B(new_n9108), .Y(new_n9111));
  NAND2xp33_ASAP7_75t_L     g08855(.A(\b[1] ), .B(new_n8835), .Y(new_n9112));
  NAND3xp33_ASAP7_75t_L     g08856(.A(new_n8833), .B(new_n8825), .C(new_n8827), .Y(new_n9113));
  NOR2xp33_ASAP7_75t_L      g08857(.A(new_n276), .B(new_n9113), .Y(new_n9114));
  AND3x1_ASAP7_75t_L        g08858(.A(new_n8543), .B(new_n8834), .C(new_n8830), .Y(new_n9115));
  AOI221xp5_ASAP7_75t_L     g08859(.A1(\b[0] ), .A2(new_n9115), .B1(new_n8828), .B2(new_n281), .C(new_n9114), .Y(new_n9116));
  NAND2xp33_ASAP7_75t_L     g08860(.A(new_n9112), .B(new_n9116), .Y(new_n9117));
  O2A1O1Ixp33_ASAP7_75t_L   g08861(.A1(new_n8544), .A2(new_n8837), .B(\a[56] ), .C(new_n9117), .Y(new_n9118));
  INVx1_ASAP7_75t_L         g08862(.A(new_n9118), .Y(new_n9119));
  NAND5xp2_ASAP7_75t_L      g08863(.A(\a[56] ), .B(new_n8829), .C(new_n8832), .D(new_n8836), .E(new_n8548), .Y(new_n9120));
  NAND3xp33_ASAP7_75t_L     g08864(.A(new_n9117), .B(new_n9120), .C(\a[56] ), .Y(new_n9121));
  AOI211xp5_ASAP7_75t_L     g08865(.A1(new_n9119), .A2(new_n9121), .B(new_n9111), .C(new_n9110), .Y(new_n9122));
  INVx1_ASAP7_75t_L         g08866(.A(new_n9111), .Y(new_n9123));
  INVx1_ASAP7_75t_L         g08867(.A(new_n9121), .Y(new_n9124));
  AOI211xp5_ASAP7_75t_L     g08868(.A1(new_n9123), .A2(new_n9109), .B(new_n9118), .C(new_n9124), .Y(new_n9125));
  OAI21xp33_ASAP7_75t_L     g08869(.A1(new_n9122), .A2(new_n9125), .B(new_n9103), .Y(new_n9126));
  A2O1A1Ixp33_ASAP7_75t_L   g08870(.A1(new_n8555), .A2(new_n8815), .B(new_n8847), .C(new_n8842), .Y(new_n9127));
  INVx1_ASAP7_75t_L         g08871(.A(new_n9122), .Y(new_n9128));
  OAI211xp5_ASAP7_75t_L     g08872(.A1(new_n9111), .A2(new_n9110), .B(new_n9119), .C(new_n9121), .Y(new_n9129));
  NAND3xp33_ASAP7_75t_L     g08873(.A(new_n9128), .B(new_n9127), .C(new_n9129), .Y(new_n9130));
  AOI21xp33_ASAP7_75t_L     g08874(.A1(new_n9130), .A2(new_n9126), .B(new_n9101), .Y(new_n9131));
  AND3x1_ASAP7_75t_L        g08875(.A(new_n9130), .B(new_n9126), .C(new_n9101), .Y(new_n9132));
  NOR3xp33_ASAP7_75t_L      g08876(.A(new_n9098), .B(new_n9132), .C(new_n9131), .Y(new_n9133));
  A2O1A1Ixp33_ASAP7_75t_L   g08877(.A1(new_n8579), .A2(new_n8809), .B(new_n8850), .C(new_n8856), .Y(new_n9134));
  AO21x2_ASAP7_75t_L        g08878(.A1(new_n9126), .A2(new_n9130), .B(new_n9101), .Y(new_n9135));
  NAND3xp33_ASAP7_75t_L     g08879(.A(new_n9130), .B(new_n9126), .C(new_n9101), .Y(new_n9136));
  AOI21xp33_ASAP7_75t_L     g08880(.A1(new_n9136), .A2(new_n9135), .B(new_n9134), .Y(new_n9137));
  OAI21xp33_ASAP7_75t_L     g08881(.A1(new_n9133), .A2(new_n9137), .B(new_n9097), .Y(new_n9138));
  XNOR2x2_ASAP7_75t_L       g08882(.A(new_n6371), .B(new_n9096), .Y(new_n9139));
  NAND3xp33_ASAP7_75t_L     g08883(.A(new_n9134), .B(new_n9135), .C(new_n9136), .Y(new_n9140));
  OAI21xp33_ASAP7_75t_L     g08884(.A1(new_n9131), .A2(new_n9132), .B(new_n9098), .Y(new_n9141));
  NAND3xp33_ASAP7_75t_L     g08885(.A(new_n9140), .B(new_n9139), .C(new_n9141), .Y(new_n9142));
  AND2x2_ASAP7_75t_L        g08886(.A(new_n9142), .B(new_n9138), .Y(new_n9143));
  A2O1A1Ixp33_ASAP7_75t_L   g08887(.A1(new_n8858), .A2(new_n8803), .B(new_n9094), .C(new_n9143), .Y(new_n9144));
  O2A1O1Ixp33_ASAP7_75t_L   g08888(.A1(new_n8801), .A2(new_n8583), .B(new_n8858), .C(new_n9094), .Y(new_n9145));
  NAND2xp33_ASAP7_75t_L     g08889(.A(new_n9142), .B(new_n9138), .Y(new_n9146));
  NAND2xp33_ASAP7_75t_L     g08890(.A(new_n9146), .B(new_n9145), .Y(new_n9147));
  AOI22xp33_ASAP7_75t_L     g08891(.A1(new_n5624), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n5901), .Y(new_n9148));
  OAI221xp5_ASAP7_75t_L     g08892(.A1(new_n5900), .A2(new_n784), .B1(new_n5892), .B2(new_n875), .C(new_n9148), .Y(new_n9149));
  XNOR2x2_ASAP7_75t_L       g08893(.A(\a[44] ), .B(new_n9149), .Y(new_n9150));
  NAND3xp33_ASAP7_75t_L     g08894(.A(new_n9144), .B(new_n9147), .C(new_n9150), .Y(new_n9151));
  A2O1A1O1Ixp25_ASAP7_75t_L g08895(.A1(new_n8267), .A2(new_n8272), .B(new_n8527), .C(new_n8587), .D(new_n8801), .Y(new_n9152));
  O2A1O1Ixp33_ASAP7_75t_L   g08896(.A1(new_n9152), .A2(new_n8865), .B(new_n8863), .C(new_n9146), .Y(new_n9153));
  AO21x2_ASAP7_75t_L        g08897(.A1(new_n8858), .A2(new_n8803), .B(new_n9094), .Y(new_n9154));
  NOR2xp33_ASAP7_75t_L      g08898(.A(new_n9143), .B(new_n9154), .Y(new_n9155));
  INVx1_ASAP7_75t_L         g08899(.A(new_n9150), .Y(new_n9156));
  OAI21xp33_ASAP7_75t_L     g08900(.A1(new_n9153), .A2(new_n9155), .B(new_n9156), .Y(new_n9157));
  AOI21xp33_ASAP7_75t_L     g08901(.A1(new_n9157), .A2(new_n9151), .B(new_n9093), .Y(new_n9158));
  AND3x1_ASAP7_75t_L        g08902(.A(new_n9093), .B(new_n9157), .C(new_n9151), .Y(new_n9159));
  OAI21xp33_ASAP7_75t_L     g08903(.A1(new_n9158), .A2(new_n9159), .B(new_n9092), .Y(new_n9160));
  AO21x2_ASAP7_75t_L        g08904(.A1(new_n9157), .A2(new_n9151), .B(new_n9093), .Y(new_n9161));
  NAND3xp33_ASAP7_75t_L     g08905(.A(new_n9093), .B(new_n9151), .C(new_n9157), .Y(new_n9162));
  NAND3xp33_ASAP7_75t_L     g08906(.A(new_n9161), .B(new_n9091), .C(new_n9162), .Y(new_n9163));
  NAND2xp33_ASAP7_75t_L     g08907(.A(new_n9163), .B(new_n9160), .Y(new_n9164));
  A2O1A1O1Ixp25_ASAP7_75t_L g08908(.A1(new_n8887), .A2(new_n8881), .B(new_n8889), .C(new_n9088), .D(new_n9164), .Y(new_n9165));
  A2O1A1Ixp33_ASAP7_75t_L   g08909(.A1(new_n8887), .A2(new_n8881), .B(new_n8889), .C(new_n9088), .Y(new_n9166));
  AOI21xp33_ASAP7_75t_L     g08910(.A1(new_n9163), .A2(new_n9160), .B(new_n9166), .Y(new_n9167));
  AOI22xp33_ASAP7_75t_L     g08911(.A1(new_n4283), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n4512), .Y(new_n9168));
  OAI221xp5_ASAP7_75t_L     g08912(.A1(new_n4277), .A2(new_n1432), .B1(new_n4499), .B2(new_n1547), .C(new_n9168), .Y(new_n9169));
  XNOR2x2_ASAP7_75t_L       g08913(.A(\a[38] ), .B(new_n9169), .Y(new_n9170));
  INVx1_ASAP7_75t_L         g08914(.A(new_n9170), .Y(new_n9171));
  OAI21xp33_ASAP7_75t_L     g08915(.A1(new_n9167), .A2(new_n9165), .B(new_n9171), .Y(new_n9172));
  NAND3xp33_ASAP7_75t_L     g08916(.A(new_n9166), .B(new_n9160), .C(new_n9163), .Y(new_n9173));
  NAND3xp33_ASAP7_75t_L     g08917(.A(new_n8898), .B(new_n9164), .C(new_n9088), .Y(new_n9174));
  NAND3xp33_ASAP7_75t_L     g08918(.A(new_n9174), .B(new_n9173), .C(new_n9170), .Y(new_n9175));
  OAI211xp5_ASAP7_75t_L     g08919(.A1(new_n8511), .A2(new_n8619), .B(new_n8794), .C(new_n8900), .Y(new_n9176));
  AND4x1_ASAP7_75t_L        g08920(.A(new_n9176), .B(new_n9175), .C(new_n9172), .D(new_n8895), .Y(new_n9177));
  AOI22xp33_ASAP7_75t_L     g08921(.A1(new_n9172), .A2(new_n9175), .B1(new_n8895), .B2(new_n9176), .Y(new_n9178));
  NOR3xp33_ASAP7_75t_L      g08922(.A(new_n9177), .B(new_n9178), .C(new_n9087), .Y(new_n9179));
  INVx1_ASAP7_75t_L         g08923(.A(new_n9087), .Y(new_n9180));
  NAND4xp25_ASAP7_75t_L     g08924(.A(new_n9176), .B(new_n9172), .C(new_n8895), .D(new_n9175), .Y(new_n9181));
  INVx1_ASAP7_75t_L         g08925(.A(new_n9178), .Y(new_n9182));
  AOI21xp33_ASAP7_75t_L     g08926(.A1(new_n9182), .A2(new_n9181), .B(new_n9180), .Y(new_n9183));
  OAI21xp33_ASAP7_75t_L     g08927(.A1(new_n9179), .A2(new_n9183), .B(new_n9084), .Y(new_n9184));
  OAI21xp33_ASAP7_75t_L     g08928(.A1(new_n8916), .A2(new_n8914), .B(new_n8908), .Y(new_n9185));
  NAND3xp33_ASAP7_75t_L     g08929(.A(new_n9182), .B(new_n9181), .C(new_n9180), .Y(new_n9186));
  OAI21xp33_ASAP7_75t_L     g08930(.A1(new_n9178), .A2(new_n9177), .B(new_n9087), .Y(new_n9187));
  NAND3xp33_ASAP7_75t_L     g08931(.A(new_n9185), .B(new_n9186), .C(new_n9187), .Y(new_n9188));
  AOI22xp33_ASAP7_75t_L     g08932(.A1(new_n3029), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n3258), .Y(new_n9189));
  OAI221xp5_ASAP7_75t_L     g08933(.A1(new_n3024), .A2(new_n2067), .B1(new_n3256), .B2(new_n2355), .C(new_n9189), .Y(new_n9190));
  XNOR2x2_ASAP7_75t_L       g08934(.A(\a[32] ), .B(new_n9190), .Y(new_n9191));
  INVx1_ASAP7_75t_L         g08935(.A(new_n9191), .Y(new_n9192));
  AOI21xp33_ASAP7_75t_L     g08936(.A1(new_n9188), .A2(new_n9184), .B(new_n9192), .Y(new_n9193));
  AOI21xp33_ASAP7_75t_L     g08937(.A1(new_n9186), .A2(new_n9187), .B(new_n9185), .Y(new_n9194));
  NOR3xp33_ASAP7_75t_L      g08938(.A(new_n9084), .B(new_n9183), .C(new_n9179), .Y(new_n9195));
  NOR3xp33_ASAP7_75t_L      g08939(.A(new_n9195), .B(new_n9194), .C(new_n9191), .Y(new_n9196));
  NOR2xp33_ASAP7_75t_L      g08940(.A(new_n9193), .B(new_n9196), .Y(new_n9197));
  NOR2xp33_ASAP7_75t_L      g08941(.A(new_n9197), .B(new_n9083), .Y(new_n9198));
  OAI21xp33_ASAP7_75t_L     g08942(.A1(new_n9194), .A2(new_n9195), .B(new_n9191), .Y(new_n9199));
  NAND3xp33_ASAP7_75t_L     g08943(.A(new_n9188), .B(new_n9184), .C(new_n9192), .Y(new_n9200));
  NAND2xp33_ASAP7_75t_L     g08944(.A(new_n9200), .B(new_n9199), .Y(new_n9201));
  O2A1O1Ixp33_ASAP7_75t_L   g08945(.A1(new_n8926), .A2(new_n8928), .B(new_n9082), .C(new_n9201), .Y(new_n9202));
  OAI21xp33_ASAP7_75t_L     g08946(.A1(new_n9202), .A2(new_n9198), .B(new_n9081), .Y(new_n9203));
  INVx1_ASAP7_75t_L         g08947(.A(new_n9082), .Y(new_n9204));
  A2O1A1O1Ixp25_ASAP7_75t_L g08948(.A1(new_n8635), .A2(new_n8638), .B(new_n8636), .C(new_n8932), .D(new_n9204), .Y(new_n9205));
  NAND2xp33_ASAP7_75t_L     g08949(.A(new_n9201), .B(new_n9205), .Y(new_n9206));
  INVx1_ASAP7_75t_L         g08950(.A(new_n8928), .Y(new_n9207));
  A2O1A1Ixp33_ASAP7_75t_L   g08951(.A1(new_n9207), .A2(new_n8932), .B(new_n9204), .C(new_n9197), .Y(new_n9208));
  OAI211xp5_ASAP7_75t_L     g08952(.A1(new_n9079), .A2(new_n9080), .B(new_n9208), .C(new_n9206), .Y(new_n9209));
  NAND2xp33_ASAP7_75t_L     g08953(.A(new_n9209), .B(new_n9203), .Y(new_n9210));
  O2A1O1Ixp33_ASAP7_75t_L   g08954(.A1(new_n9076), .A2(new_n8936), .B(new_n8953), .C(new_n9210), .Y(new_n9211));
  NAND3xp33_ASAP7_75t_L     g08955(.A(new_n8929), .B(new_n8933), .C(new_n8940), .Y(new_n9212));
  A2O1A1Ixp33_ASAP7_75t_L   g08956(.A1(new_n8941), .A2(new_n8937), .B(new_n8945), .C(new_n9212), .Y(new_n9213));
  AOI21xp33_ASAP7_75t_L     g08957(.A1(new_n9209), .A2(new_n9203), .B(new_n9213), .Y(new_n9214));
  OAI21xp33_ASAP7_75t_L     g08958(.A1(new_n9214), .A2(new_n9211), .B(new_n9075), .Y(new_n9215));
  INVx1_ASAP7_75t_L         g08959(.A(new_n9075), .Y(new_n9216));
  AND2x2_ASAP7_75t_L        g08960(.A(new_n9209), .B(new_n9203), .Y(new_n9217));
  NAND2xp33_ASAP7_75t_L     g08961(.A(new_n9213), .B(new_n9217), .Y(new_n9218));
  NAND3xp33_ASAP7_75t_L     g08962(.A(new_n9210), .B(new_n9212), .C(new_n8953), .Y(new_n9219));
  NAND3xp33_ASAP7_75t_L     g08963(.A(new_n9218), .B(new_n9219), .C(new_n9216), .Y(new_n9220));
  NAND3xp33_ASAP7_75t_L     g08964(.A(new_n9068), .B(new_n9215), .C(new_n9220), .Y(new_n9221));
  NOR2xp33_ASAP7_75t_L      g08965(.A(new_n8946), .B(new_n8944), .Y(new_n9222));
  MAJIxp5_ASAP7_75t_L       g08966(.A(new_n8966), .B(new_n8950), .C(new_n9222), .Y(new_n9223));
  AOI21xp33_ASAP7_75t_L     g08967(.A1(new_n9218), .A2(new_n9219), .B(new_n9216), .Y(new_n9224));
  NOR3xp33_ASAP7_75t_L      g08968(.A(new_n9211), .B(new_n9214), .C(new_n9075), .Y(new_n9225));
  OAI21xp33_ASAP7_75t_L     g08969(.A1(new_n9225), .A2(new_n9224), .B(new_n9223), .Y(new_n9226));
  NOR2xp33_ASAP7_75t_L      g08970(.A(new_n3584), .B(new_n1699), .Y(new_n9227));
  INVx1_ASAP7_75t_L         g08971(.A(new_n9227), .Y(new_n9228));
  NAND2xp33_ASAP7_75t_L     g08972(.A(new_n1695), .B(new_n3811), .Y(new_n9229));
  AOI22xp33_ASAP7_75t_L     g08973(.A1(new_n1704), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1837), .Y(new_n9230));
  AND4x1_ASAP7_75t_L        g08974(.A(new_n9230), .B(new_n9229), .C(new_n9228), .D(\a[23] ), .Y(new_n9231));
  AOI31xp33_ASAP7_75t_L     g08975(.A1(new_n9229), .A2(new_n9228), .A3(new_n9230), .B(\a[23] ), .Y(new_n9232));
  NOR2xp33_ASAP7_75t_L      g08976(.A(new_n9232), .B(new_n9231), .Y(new_n9233));
  NAND3xp33_ASAP7_75t_L     g08977(.A(new_n9221), .B(new_n9226), .C(new_n9233), .Y(new_n9234));
  NOR3xp33_ASAP7_75t_L      g08978(.A(new_n9223), .B(new_n9224), .C(new_n9225), .Y(new_n9235));
  AOI21xp33_ASAP7_75t_L     g08979(.A1(new_n9220), .A2(new_n9215), .B(new_n9068), .Y(new_n9236));
  INVx1_ASAP7_75t_L         g08980(.A(new_n9233), .Y(new_n9237));
  OAI21xp33_ASAP7_75t_L     g08981(.A1(new_n9236), .A2(new_n9235), .B(new_n9237), .Y(new_n9238));
  NAND2xp33_ASAP7_75t_L     g08982(.A(new_n9234), .B(new_n9238), .Y(new_n9239));
  NAND2xp33_ASAP7_75t_L     g08983(.A(new_n8957), .B(new_n8961), .Y(new_n9240));
  MAJIxp5_ASAP7_75t_L       g08984(.A(new_n8972), .B(new_n8964), .C(new_n9240), .Y(new_n9241));
  NOR2xp33_ASAP7_75t_L      g08985(.A(new_n9241), .B(new_n9239), .Y(new_n9242));
  NOR2xp33_ASAP7_75t_L      g08986(.A(new_n8967), .B(new_n8968), .Y(new_n9243));
  MAJIxp5_ASAP7_75t_L       g08987(.A(new_n8977), .B(new_n8969), .C(new_n9243), .Y(new_n9244));
  AOI21xp33_ASAP7_75t_L     g08988(.A1(new_n9238), .A2(new_n9234), .B(new_n9244), .Y(new_n9245));
  AOI22xp33_ASAP7_75t_L     g08989(.A1(new_n1360), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1581), .Y(new_n9246));
  OAI221xp5_ASAP7_75t_L     g08990(.A1(new_n1373), .A2(new_n4424), .B1(new_n1359), .B2(new_n4641), .C(new_n9246), .Y(new_n9247));
  XNOR2x2_ASAP7_75t_L       g08991(.A(\a[20] ), .B(new_n9247), .Y(new_n9248));
  INVx1_ASAP7_75t_L         g08992(.A(new_n9248), .Y(new_n9249));
  NOR3xp33_ASAP7_75t_L      g08993(.A(new_n9245), .B(new_n9242), .C(new_n9249), .Y(new_n9250));
  NAND3xp33_ASAP7_75t_L     g08994(.A(new_n9244), .B(new_n9238), .C(new_n9234), .Y(new_n9251));
  NAND2xp33_ASAP7_75t_L     g08995(.A(new_n9241), .B(new_n9239), .Y(new_n9252));
  AOI21xp33_ASAP7_75t_L     g08996(.A1(new_n9251), .A2(new_n9252), .B(new_n9248), .Y(new_n9253));
  NAND2xp33_ASAP7_75t_L     g08997(.A(new_n8978), .B(new_n8973), .Y(new_n9254));
  MAJIxp5_ASAP7_75t_L       g08998(.A(new_n8985), .B(new_n9254), .C(new_n8981), .Y(new_n9255));
  NOR3xp33_ASAP7_75t_L      g08999(.A(new_n9255), .B(new_n9253), .C(new_n9250), .Y(new_n9256));
  OA21x2_ASAP7_75t_L        g09000(.A1(new_n9250), .A2(new_n9253), .B(new_n9255), .Y(new_n9257));
  NOR2xp33_ASAP7_75t_L      g09001(.A(new_n4869), .B(new_n1154), .Y(new_n9258));
  NAND3xp33_ASAP7_75t_L     g09002(.A(new_n5326), .B(new_n5324), .C(new_n1073), .Y(new_n9259));
  AOI22xp33_ASAP7_75t_L     g09003(.A1(new_n1076), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1253), .Y(new_n9260));
  NAND2xp33_ASAP7_75t_L     g09004(.A(new_n9260), .B(new_n9259), .Y(new_n9261));
  OR3x1_ASAP7_75t_L         g09005(.A(new_n9261), .B(new_n1071), .C(new_n9258), .Y(new_n9262));
  A2O1A1Ixp33_ASAP7_75t_L   g09006(.A1(\b[40] ), .A2(new_n1080), .B(new_n9261), .C(new_n1071), .Y(new_n9263));
  NAND2xp33_ASAP7_75t_L     g09007(.A(new_n9263), .B(new_n9262), .Y(new_n9264));
  NOR3xp33_ASAP7_75t_L      g09008(.A(new_n9257), .B(new_n9264), .C(new_n9256), .Y(new_n9265));
  NAND3xp33_ASAP7_75t_L     g09009(.A(new_n9251), .B(new_n9252), .C(new_n9248), .Y(new_n9266));
  OAI21xp33_ASAP7_75t_L     g09010(.A1(new_n9242), .A2(new_n9245), .B(new_n9249), .Y(new_n9267));
  INVx1_ASAP7_75t_L         g09011(.A(new_n8981), .Y(new_n9268));
  NAND3xp33_ASAP7_75t_L     g09012(.A(new_n8973), .B(new_n8978), .C(new_n9268), .Y(new_n9269));
  NAND4xp25_ASAP7_75t_L     g09013(.A(new_n8987), .B(new_n9267), .C(new_n9269), .D(new_n9266), .Y(new_n9270));
  OAI21xp33_ASAP7_75t_L     g09014(.A1(new_n9250), .A2(new_n9253), .B(new_n9255), .Y(new_n9271));
  INVx1_ASAP7_75t_L         g09015(.A(new_n9264), .Y(new_n9272));
  AOI21xp33_ASAP7_75t_L     g09016(.A1(new_n9270), .A2(new_n9271), .B(new_n9272), .Y(new_n9273));
  NOR2xp33_ASAP7_75t_L      g09017(.A(new_n9273), .B(new_n9265), .Y(new_n9274));
  NOR3xp33_ASAP7_75t_L      g09018(.A(new_n8995), .B(new_n8996), .C(new_n8993), .Y(new_n9275));
  AOI21xp33_ASAP7_75t_L     g09019(.A1(new_n9000), .A2(new_n8998), .B(new_n9275), .Y(new_n9276));
  NAND2xp33_ASAP7_75t_L     g09020(.A(new_n9274), .B(new_n9276), .Y(new_n9277));
  NAND3xp33_ASAP7_75t_L     g09021(.A(new_n9270), .B(new_n9272), .C(new_n9271), .Y(new_n9278));
  OAI21xp33_ASAP7_75t_L     g09022(.A1(new_n9256), .A2(new_n9257), .B(new_n9264), .Y(new_n9279));
  NAND2xp33_ASAP7_75t_L     g09023(.A(new_n9278), .B(new_n9279), .Y(new_n9280));
  A2O1A1Ixp33_ASAP7_75t_L   g09024(.A1(new_n8998), .A2(new_n9000), .B(new_n9275), .C(new_n9280), .Y(new_n9281));
  AOI22xp33_ASAP7_75t_L     g09025(.A1(new_n811), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n900), .Y(new_n9282));
  OAI221xp5_ASAP7_75t_L     g09026(.A1(new_n904), .A2(new_n5805), .B1(new_n898), .B2(new_n5835), .C(new_n9282), .Y(new_n9283));
  XNOR2x2_ASAP7_75t_L       g09027(.A(\a[14] ), .B(new_n9283), .Y(new_n9284));
  INVx1_ASAP7_75t_L         g09028(.A(new_n9284), .Y(new_n9285));
  AOI21xp33_ASAP7_75t_L     g09029(.A1(new_n9277), .A2(new_n9281), .B(new_n9285), .Y(new_n9286));
  INVx1_ASAP7_75t_L         g09030(.A(new_n9286), .Y(new_n9287));
  NAND3xp33_ASAP7_75t_L     g09031(.A(new_n9277), .B(new_n9281), .C(new_n9285), .Y(new_n9288));
  AOI211xp5_ASAP7_75t_L     g09032(.A1(new_n8720), .A2(new_n8713), .B(new_n8709), .C(new_n9009), .Y(new_n9289));
  OAI211xp5_ASAP7_75t_L     g09033(.A1(new_n9289), .A2(new_n9006), .B(new_n9287), .C(new_n9288), .Y(new_n9290));
  INVx1_ASAP7_75t_L         g09034(.A(new_n9288), .Y(new_n9291));
  NAND2xp33_ASAP7_75t_L     g09035(.A(new_n9005), .B(new_n9001), .Y(new_n9292));
  NAND2xp33_ASAP7_75t_L     g09036(.A(new_n8788), .B(new_n9292), .Y(new_n9293));
  OAI221xp5_ASAP7_75t_L     g09037(.A1(new_n9001), .A2(new_n9005), .B1(new_n9286), .B2(new_n9291), .C(new_n9293), .Y(new_n9294));
  AOI21xp33_ASAP7_75t_L     g09038(.A1(new_n9294), .A2(new_n9290), .B(new_n9066), .Y(new_n9295));
  INVx1_ASAP7_75t_L         g09039(.A(new_n9295), .Y(new_n9296));
  NAND3xp33_ASAP7_75t_L     g09040(.A(new_n9294), .B(new_n9290), .C(new_n9066), .Y(new_n9297));
  NAND3xp33_ASAP7_75t_L     g09041(.A(new_n9296), .B(new_n9063), .C(new_n9297), .Y(new_n9298));
  NOR2xp33_ASAP7_75t_L      g09042(.A(new_n8481), .B(new_n9015), .Y(new_n9299));
  O2A1O1Ixp33_ASAP7_75t_L   g09043(.A1(new_n9299), .A2(new_n8731), .B(new_n9017), .C(new_n9013), .Y(new_n9300));
  AND3x1_ASAP7_75t_L        g09044(.A(new_n9294), .B(new_n9290), .C(new_n9066), .Y(new_n9301));
  OAI21xp33_ASAP7_75t_L     g09045(.A1(new_n9295), .A2(new_n9301), .B(new_n9300), .Y(new_n9302));
  AO21x2_ASAP7_75t_L        g09046(.A1(new_n9302), .A2(new_n9298), .B(new_n9061), .Y(new_n9303));
  NAND3xp33_ASAP7_75t_L     g09047(.A(new_n9061), .B(new_n9298), .C(new_n9302), .Y(new_n9304));
  AOI21xp33_ASAP7_75t_L     g09048(.A1(new_n9303), .A2(new_n9304), .B(new_n9055), .Y(new_n9305));
  AND3x1_ASAP7_75t_L        g09049(.A(new_n9303), .B(new_n9055), .C(new_n9304), .Y(new_n9306));
  OAI21xp33_ASAP7_75t_L     g09050(.A1(new_n9305), .A2(new_n9306), .B(new_n9053), .Y(new_n9307));
  INVx1_ASAP7_75t_L         g09051(.A(new_n9053), .Y(new_n9308));
  AO21x2_ASAP7_75t_L        g09052(.A1(new_n9304), .A2(new_n9303), .B(new_n9055), .Y(new_n9309));
  NAND3xp33_ASAP7_75t_L     g09053(.A(new_n9303), .B(new_n9055), .C(new_n9304), .Y(new_n9310));
  NAND3xp33_ASAP7_75t_L     g09054(.A(new_n9309), .B(new_n9308), .C(new_n9310), .Y(new_n9311));
  NAND3xp33_ASAP7_75t_L     g09055(.A(new_n9047), .B(new_n9307), .C(new_n9311), .Y(new_n9312));
  NOR3xp33_ASAP7_75t_L      g09056(.A(new_n9033), .B(new_n9034), .C(new_n9035), .Y(new_n9313));
  AOI21xp33_ASAP7_75t_L     g09057(.A1(new_n9025), .A2(new_n9028), .B(new_n9031), .Y(new_n9314));
  NOR2xp33_ASAP7_75t_L      g09058(.A(new_n9313), .B(new_n9314), .Y(new_n9315));
  NOR2xp33_ASAP7_75t_L      g09059(.A(new_n9034), .B(new_n9033), .Y(new_n9316));
  NAND2xp33_ASAP7_75t_L     g09060(.A(new_n9035), .B(new_n9316), .Y(new_n9317));
  AOI21xp33_ASAP7_75t_L     g09061(.A1(new_n9309), .A2(new_n9310), .B(new_n9308), .Y(new_n9318));
  NOR3xp33_ASAP7_75t_L      g09062(.A(new_n9306), .B(new_n9053), .C(new_n9305), .Y(new_n9319));
  OAI221xp5_ASAP7_75t_L     g09063(.A1(new_n9319), .A2(new_n9318), .B1(new_n8772), .B2(new_n9315), .C(new_n9317), .Y(new_n9320));
  NAND2xp33_ASAP7_75t_L     g09064(.A(new_n9320), .B(new_n9312), .Y(new_n9321));
  NOR2xp33_ASAP7_75t_L      g09065(.A(\b[55] ), .B(\b[56] ), .Y(new_n9322));
  INVx1_ASAP7_75t_L         g09066(.A(\b[56] ), .Y(new_n9323));
  NOR2xp33_ASAP7_75t_L      g09067(.A(new_n8762), .B(new_n9323), .Y(new_n9324));
  NOR2xp33_ASAP7_75t_L      g09068(.A(new_n9322), .B(new_n9324), .Y(new_n9325));
  INVx1_ASAP7_75t_L         g09069(.A(new_n9325), .Y(new_n9326));
  O2A1O1Ixp33_ASAP7_75t_L   g09070(.A1(new_n8458), .A2(new_n8762), .B(new_n8765), .C(new_n9326), .Y(new_n9327));
  INVx1_ASAP7_75t_L         g09071(.A(new_n9327), .Y(new_n9328));
  O2A1O1Ixp33_ASAP7_75t_L   g09072(.A1(new_n8459), .A2(new_n8462), .B(new_n8764), .C(new_n8763), .Y(new_n9329));
  NAND2xp33_ASAP7_75t_L     g09073(.A(new_n9326), .B(new_n9329), .Y(new_n9330));
  NAND2xp33_ASAP7_75t_L     g09074(.A(new_n9330), .B(new_n9328), .Y(new_n9331));
  INVx1_ASAP7_75t_L         g09075(.A(new_n9331), .Y(new_n9332));
  OAI22xp33_ASAP7_75t_L     g09076(.A1(new_n271), .A2(new_n9323), .B1(new_n8458), .B2(new_n283), .Y(new_n9333));
  AOI221xp5_ASAP7_75t_L     g09077(.A1(\b[55] ), .A2(new_n272), .B1(new_n267), .B2(new_n9332), .C(new_n9333), .Y(new_n9334));
  XNOR2x2_ASAP7_75t_L       g09078(.A(new_n262), .B(new_n9334), .Y(new_n9335));
  XNOR2x2_ASAP7_75t_L       g09079(.A(new_n9335), .B(new_n9321), .Y(new_n9336));
  A2O1A1O1Ixp25_ASAP7_75t_L g09080(.A1(new_n8455), .A2(new_n8757), .B(new_n8755), .C(new_n9041), .D(new_n9039), .Y(new_n9337));
  XOR2x2_ASAP7_75t_L        g09081(.A(new_n9337), .B(new_n9336), .Y(\f[56] ));
  MAJIxp5_ASAP7_75t_L       g09082(.A(new_n9337), .B(new_n9335), .C(new_n9321), .Y(new_n9339));
  AO21x2_ASAP7_75t_L        g09083(.A1(new_n9307), .A2(new_n9047), .B(new_n9319), .Y(new_n9340));
  AOI22xp33_ASAP7_75t_L     g09084(.A1(new_n344), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n370), .Y(new_n9341));
  OAI221xp5_ASAP7_75t_L     g09085(.A1(new_n429), .A2(new_n8165), .B1(new_n366), .B2(new_n8465), .C(new_n9341), .Y(new_n9342));
  NOR2xp33_ASAP7_75t_L      g09086(.A(new_n338), .B(new_n9342), .Y(new_n9343));
  AND2x2_ASAP7_75t_L        g09087(.A(new_n338), .B(new_n9342), .Y(new_n9344));
  NOR2xp33_ASAP7_75t_L      g09088(.A(new_n9343), .B(new_n9344), .Y(new_n9345));
  INVx1_ASAP7_75t_L         g09089(.A(new_n9345), .Y(new_n9346));
  NAND2xp33_ASAP7_75t_L     g09090(.A(new_n9302), .B(new_n9298), .Y(new_n9347));
  MAJIxp5_ASAP7_75t_L       g09091(.A(new_n9055), .B(new_n9061), .C(new_n9347), .Y(new_n9348));
  OAI22xp33_ASAP7_75t_L     g09092(.A1(new_n516), .A2(new_n7317), .B1(new_n7616), .B2(new_n515), .Y(new_n9349));
  AOI221xp5_ASAP7_75t_L     g09093(.A1(\b[50] ), .A2(new_n447), .B1(new_n441), .B2(new_n7622), .C(new_n9349), .Y(new_n9350));
  XNOR2x2_ASAP7_75t_L       g09094(.A(new_n435), .B(new_n9350), .Y(new_n9351));
  NOR2xp33_ASAP7_75t_L      g09095(.A(new_n6812), .B(new_n821), .Y(new_n9352));
  INVx1_ASAP7_75t_L         g09096(.A(new_n9352), .Y(new_n9353));
  NAND2xp33_ASAP7_75t_L     g09097(.A(new_n578), .B(new_n7630), .Y(new_n9354));
  AOI22xp33_ASAP7_75t_L     g09098(.A1(\b[46] ), .A2(new_n651), .B1(\b[48] ), .B2(new_n581), .Y(new_n9355));
  NAND4xp25_ASAP7_75t_L     g09099(.A(new_n9354), .B(\a[11] ), .C(new_n9353), .D(new_n9355), .Y(new_n9356));
  AOI31xp33_ASAP7_75t_L     g09100(.A1(new_n9354), .A2(new_n9353), .A3(new_n9355), .B(\a[11] ), .Y(new_n9357));
  INVx1_ASAP7_75t_L         g09101(.A(new_n9357), .Y(new_n9358));
  NAND2xp33_ASAP7_75t_L     g09102(.A(new_n9356), .B(new_n9358), .Y(new_n9359));
  NOR2xp33_ASAP7_75t_L      g09103(.A(new_n5829), .B(new_n904), .Y(new_n9360));
  INVx1_ASAP7_75t_L         g09104(.A(new_n9360), .Y(new_n9361));
  NAND2xp33_ASAP7_75t_L     g09105(.A(new_n808), .B(new_n7066), .Y(new_n9362));
  AOI22xp33_ASAP7_75t_L     g09106(.A1(new_n811), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n900), .Y(new_n9363));
  AND4x1_ASAP7_75t_L        g09107(.A(new_n9363), .B(new_n9362), .C(new_n9361), .D(\a[14] ), .Y(new_n9364));
  AOI31xp33_ASAP7_75t_L     g09108(.A1(new_n9362), .A2(new_n9361), .A3(new_n9363), .B(\a[14] ), .Y(new_n9365));
  NOR2xp33_ASAP7_75t_L      g09109(.A(new_n9365), .B(new_n9364), .Y(new_n9366));
  NOR3xp33_ASAP7_75t_L      g09110(.A(new_n9257), .B(new_n9272), .C(new_n9256), .Y(new_n9367));
  INVx1_ASAP7_75t_L         g09111(.A(new_n9367), .Y(new_n9368));
  OAI21xp33_ASAP7_75t_L     g09112(.A1(new_n9274), .A2(new_n9276), .B(new_n9368), .Y(new_n9369));
  NOR3xp33_ASAP7_75t_L      g09113(.A(new_n9235), .B(new_n9236), .C(new_n9233), .Y(new_n9370));
  INVx1_ASAP7_75t_L         g09114(.A(new_n9370), .Y(new_n9371));
  AOI22xp33_ASAP7_75t_L     g09115(.A1(new_n1704), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n1837), .Y(new_n9372));
  OAI221xp5_ASAP7_75t_L     g09116(.A1(new_n1699), .A2(new_n3804), .B1(new_n1827), .B2(new_n4223), .C(new_n9372), .Y(new_n9373));
  XNOR2x2_ASAP7_75t_L       g09117(.A(\a[23] ), .B(new_n9373), .Y(new_n9374));
  INVx1_ASAP7_75t_L         g09118(.A(new_n9374), .Y(new_n9375));
  NOR3xp33_ASAP7_75t_L      g09119(.A(new_n9198), .B(new_n9202), .C(new_n9081), .Y(new_n9376));
  NOR2xp33_ASAP7_75t_L      g09120(.A(new_n2688), .B(new_n2547), .Y(new_n9377));
  INVx1_ASAP7_75t_L         g09121(.A(new_n9377), .Y(new_n9378));
  NAND2xp33_ASAP7_75t_L     g09122(.A(new_n2544), .B(new_n2989), .Y(new_n9379));
  AOI22xp33_ASAP7_75t_L     g09123(.A1(new_n2552), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n2736), .Y(new_n9380));
  AND4x1_ASAP7_75t_L        g09124(.A(new_n9380), .B(new_n9379), .C(new_n9378), .D(\a[29] ), .Y(new_n9381));
  AOI31xp33_ASAP7_75t_L     g09125(.A1(new_n9379), .A2(new_n9378), .A3(new_n9380), .B(\a[29] ), .Y(new_n9382));
  NOR2xp33_ASAP7_75t_L      g09126(.A(new_n9382), .B(new_n9381), .Y(new_n9383));
  AOI21xp33_ASAP7_75t_L     g09127(.A1(new_n9174), .A2(new_n9173), .B(new_n9170), .Y(new_n9384));
  AO31x2_ASAP7_75t_L        g09128(.A1(new_n9176), .A2(new_n8895), .A3(new_n9175), .B(new_n9384), .Y(new_n9385));
  AOI22xp33_ASAP7_75t_L     g09129(.A1(new_n4283), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n4512), .Y(new_n9386));
  OAI221xp5_ASAP7_75t_L     g09130(.A1(new_n4277), .A2(new_n1539), .B1(new_n4499), .B2(new_n1662), .C(new_n9386), .Y(new_n9387));
  XNOR2x2_ASAP7_75t_L       g09131(.A(\a[38] ), .B(new_n9387), .Y(new_n9388));
  INVx1_ASAP7_75t_L         g09132(.A(new_n9388), .Y(new_n9389));
  NOR3xp33_ASAP7_75t_L      g09133(.A(new_n9159), .B(new_n9158), .C(new_n9091), .Y(new_n9390));
  AOI22xp33_ASAP7_75t_L     g09134(.A1(new_n4920), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n5167), .Y(new_n9391));
  OAI221xp5_ASAP7_75t_L     g09135(.A1(new_n5154), .A2(new_n1201), .B1(new_n5158), .B2(new_n1320), .C(new_n9391), .Y(new_n9392));
  XNOR2x2_ASAP7_75t_L       g09136(.A(new_n4915), .B(new_n9392), .Y(new_n9393));
  AND2x2_ASAP7_75t_L        g09137(.A(new_n9151), .B(new_n9157), .Y(new_n9394));
  NAND3xp33_ASAP7_75t_L     g09138(.A(new_n9144), .B(new_n9147), .C(new_n9156), .Y(new_n9395));
  AOI22xp33_ASAP7_75t_L     g09139(.A1(new_n5624), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n5901), .Y(new_n9396));
  OAI221xp5_ASAP7_75t_L     g09140(.A1(new_n5900), .A2(new_n869), .B1(new_n5892), .B2(new_n950), .C(new_n9396), .Y(new_n9397));
  XNOR2x2_ASAP7_75t_L       g09141(.A(\a[44] ), .B(new_n9397), .Y(new_n9398));
  INVx1_ASAP7_75t_L         g09142(.A(new_n9398), .Y(new_n9399));
  NOR3xp33_ASAP7_75t_L      g09143(.A(new_n9137), .B(new_n9133), .C(new_n9097), .Y(new_n9400));
  A2O1A1O1Ixp25_ASAP7_75t_L g09144(.A1(new_n8858), .A2(new_n8803), .B(new_n9094), .C(new_n9138), .D(new_n9400), .Y(new_n9401));
  NOR2xp33_ASAP7_75t_L      g09145(.A(new_n679), .B(new_n6646), .Y(new_n9402));
  NAND2xp33_ASAP7_75t_L     g09146(.A(\b[10] ), .B(new_n6648), .Y(new_n9403));
  OAI221xp5_ASAP7_75t_L     g09147(.A1(new_n6880), .A2(new_n760), .B1(new_n6636), .B2(new_n768), .C(new_n9403), .Y(new_n9404));
  OR3x1_ASAP7_75t_L         g09148(.A(new_n9404), .B(new_n6371), .C(new_n9402), .Y(new_n9405));
  A2O1A1Ixp33_ASAP7_75t_L   g09149(.A1(\b[11] ), .A2(new_n6380), .B(new_n9404), .C(new_n6371), .Y(new_n9406));
  NAND2xp33_ASAP7_75t_L     g09150(.A(new_n9406), .B(new_n9405), .Y(new_n9407));
  A2O1A1Ixp33_ASAP7_75t_L   g09151(.A1(new_n8859), .A2(new_n8856), .B(new_n9131), .C(new_n9136), .Y(new_n9408));
  INVx1_ASAP7_75t_L         g09152(.A(\a[57] ), .Y(new_n9409));
  NAND2xp33_ASAP7_75t_L     g09153(.A(\a[56] ), .B(new_n9409), .Y(new_n9410));
  NAND2xp33_ASAP7_75t_L     g09154(.A(\a[57] ), .B(new_n8826), .Y(new_n9411));
  AND2x2_ASAP7_75t_L        g09155(.A(new_n9410), .B(new_n9411), .Y(new_n9412));
  NOR2xp33_ASAP7_75t_L      g09156(.A(new_n258), .B(new_n9412), .Y(new_n9413));
  OAI21xp33_ASAP7_75t_L     g09157(.A1(new_n9120), .A2(new_n9117), .B(new_n9413), .Y(new_n9414));
  INVx1_ASAP7_75t_L         g09158(.A(new_n9120), .Y(new_n9415));
  INVx1_ASAP7_75t_L         g09159(.A(new_n9413), .Y(new_n9416));
  NAND4xp25_ASAP7_75t_L     g09160(.A(new_n9415), .B(new_n9416), .C(new_n9116), .D(new_n9112), .Y(new_n9417));
  NAND3xp33_ASAP7_75t_L     g09161(.A(new_n8543), .B(new_n8830), .C(new_n8834), .Y(new_n9418));
  OAI22xp33_ASAP7_75t_L     g09162(.A1(new_n9418), .A2(new_n261), .B1(new_n298), .B2(new_n9113), .Y(new_n9419));
  AOI221xp5_ASAP7_75t_L     g09163(.A1(\b[2] ), .A2(new_n8835), .B1(new_n406), .B2(new_n8828), .C(new_n9419), .Y(new_n9420));
  NAND2xp33_ASAP7_75t_L     g09164(.A(\a[56] ), .B(new_n9420), .Y(new_n9421));
  AO21x2_ASAP7_75t_L        g09165(.A1(new_n406), .A2(new_n8828), .B(new_n9419), .Y(new_n9422));
  A2O1A1Ixp33_ASAP7_75t_L   g09166(.A1(\b[2] ), .A2(new_n8835), .B(new_n9422), .C(new_n8826), .Y(new_n9423));
  AO22x1_ASAP7_75t_L        g09167(.A1(new_n9423), .A2(new_n9421), .B1(new_n9414), .B2(new_n9417), .Y(new_n9424));
  XNOR2x2_ASAP7_75t_L       g09168(.A(new_n8826), .B(new_n9420), .Y(new_n9425));
  NAND3xp33_ASAP7_75t_L     g09169(.A(new_n9425), .B(new_n9417), .C(new_n9414), .Y(new_n9426));
  NOR2xp33_ASAP7_75t_L      g09170(.A(new_n354), .B(new_n8817), .Y(new_n9427));
  INVx1_ASAP7_75t_L         g09171(.A(new_n9427), .Y(new_n9428));
  NAND2xp33_ASAP7_75t_L     g09172(.A(new_n7958), .B(new_n526), .Y(new_n9429));
  AOI22xp33_ASAP7_75t_L     g09173(.A1(new_n7960), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n8537), .Y(new_n9430));
  NAND4xp25_ASAP7_75t_L     g09174(.A(new_n9429), .B(\a[53] ), .C(new_n9428), .D(new_n9430), .Y(new_n9431));
  AOI31xp33_ASAP7_75t_L     g09175(.A1(new_n9429), .A2(new_n9428), .A3(new_n9430), .B(\a[53] ), .Y(new_n9432));
  INVx1_ASAP7_75t_L         g09176(.A(new_n9432), .Y(new_n9433));
  NAND4xp25_ASAP7_75t_L     g09177(.A(new_n9424), .B(new_n9426), .C(new_n9433), .D(new_n9431), .Y(new_n9434));
  AOI21xp33_ASAP7_75t_L     g09178(.A1(new_n9417), .A2(new_n9414), .B(new_n9425), .Y(new_n9435));
  AND4x1_ASAP7_75t_L        g09179(.A(new_n9417), .B(new_n9414), .C(new_n9423), .D(new_n9421), .Y(new_n9436));
  INVx1_ASAP7_75t_L         g09180(.A(new_n9431), .Y(new_n9437));
  OAI22xp33_ASAP7_75t_L     g09181(.A1(new_n9435), .A2(new_n9436), .B1(new_n9432), .B2(new_n9437), .Y(new_n9438));
  OAI211xp5_ASAP7_75t_L     g09182(.A1(new_n8846), .A2(new_n8847), .B(new_n9129), .C(new_n8842), .Y(new_n9439));
  AND4x1_ASAP7_75t_L        g09183(.A(new_n9439), .B(new_n9438), .C(new_n9434), .D(new_n9128), .Y(new_n9440));
  AOI21xp33_ASAP7_75t_L     g09184(.A1(new_n9103), .A2(new_n9129), .B(new_n9122), .Y(new_n9441));
  AOI21xp33_ASAP7_75t_L     g09185(.A1(new_n9438), .A2(new_n9434), .B(new_n9441), .Y(new_n9442));
  AOI22xp33_ASAP7_75t_L     g09186(.A1(new_n7111), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n7391), .Y(new_n9443));
  OAI221xp5_ASAP7_75t_L     g09187(.A1(new_n8558), .A2(new_n488), .B1(new_n8237), .B2(new_n548), .C(new_n9443), .Y(new_n9444));
  NOR2xp33_ASAP7_75t_L      g09188(.A(new_n7106), .B(new_n9444), .Y(new_n9445));
  NAND2xp33_ASAP7_75t_L     g09189(.A(new_n7106), .B(new_n9444), .Y(new_n9446));
  INVx1_ASAP7_75t_L         g09190(.A(new_n9446), .Y(new_n9447));
  OAI22xp33_ASAP7_75t_L     g09191(.A1(new_n9442), .A2(new_n9440), .B1(new_n9445), .B2(new_n9447), .Y(new_n9448));
  NAND4xp25_ASAP7_75t_L     g09192(.A(new_n9439), .B(new_n9128), .C(new_n9434), .D(new_n9438), .Y(new_n9449));
  NAND2xp33_ASAP7_75t_L     g09193(.A(new_n9438), .B(new_n9434), .Y(new_n9450));
  A2O1A1Ixp33_ASAP7_75t_L   g09194(.A1(new_n9129), .A2(new_n9103), .B(new_n9122), .C(new_n9450), .Y(new_n9451));
  INVx1_ASAP7_75t_L         g09195(.A(new_n9445), .Y(new_n9452));
  NAND4xp25_ASAP7_75t_L     g09196(.A(new_n9451), .B(new_n9452), .C(new_n9446), .D(new_n9449), .Y(new_n9453));
  NAND3xp33_ASAP7_75t_L     g09197(.A(new_n9408), .B(new_n9448), .C(new_n9453), .Y(new_n9454));
  NAND2xp33_ASAP7_75t_L     g09198(.A(new_n8809), .B(new_n8579), .Y(new_n9455));
  A2O1A1O1Ixp25_ASAP7_75t_L g09199(.A1(new_n8855), .A2(new_n9455), .B(new_n8853), .C(new_n9135), .D(new_n9132), .Y(new_n9456));
  NAND2xp33_ASAP7_75t_L     g09200(.A(new_n9453), .B(new_n9448), .Y(new_n9457));
  NAND2xp33_ASAP7_75t_L     g09201(.A(new_n9457), .B(new_n9456), .Y(new_n9458));
  AOI21xp33_ASAP7_75t_L     g09202(.A1(new_n9458), .A2(new_n9454), .B(new_n9407), .Y(new_n9459));
  NOR2xp33_ASAP7_75t_L      g09203(.A(new_n9457), .B(new_n9456), .Y(new_n9460));
  AOI21xp33_ASAP7_75t_L     g09204(.A1(new_n9453), .A2(new_n9448), .B(new_n9408), .Y(new_n9461));
  AOI211xp5_ASAP7_75t_L     g09205(.A1(new_n9405), .A2(new_n9406), .B(new_n9460), .C(new_n9461), .Y(new_n9462));
  OR3x1_ASAP7_75t_L         g09206(.A(new_n9401), .B(new_n9459), .C(new_n9462), .Y(new_n9463));
  OAI21xp33_ASAP7_75t_L     g09207(.A1(new_n9459), .A2(new_n9462), .B(new_n9401), .Y(new_n9464));
  NAND3xp33_ASAP7_75t_L     g09208(.A(new_n9463), .B(new_n9399), .C(new_n9464), .Y(new_n9465));
  NOR3xp33_ASAP7_75t_L      g09209(.A(new_n9401), .B(new_n9459), .C(new_n9462), .Y(new_n9466));
  OA21x2_ASAP7_75t_L        g09210(.A1(new_n9459), .A2(new_n9462), .B(new_n9401), .Y(new_n9467));
  OAI21xp33_ASAP7_75t_L     g09211(.A1(new_n9466), .A2(new_n9467), .B(new_n9398), .Y(new_n9468));
  NAND2xp33_ASAP7_75t_L     g09212(.A(new_n9468), .B(new_n9465), .Y(new_n9469));
  O2A1O1Ixp33_ASAP7_75t_L   g09213(.A1(new_n9093), .A2(new_n9394), .B(new_n9395), .C(new_n9469), .Y(new_n9470));
  A2O1A1Ixp33_ASAP7_75t_L   g09214(.A1(new_n9151), .A2(new_n9157), .B(new_n9093), .C(new_n9395), .Y(new_n9471));
  AOI21xp33_ASAP7_75t_L     g09215(.A1(new_n9468), .A2(new_n9465), .B(new_n9471), .Y(new_n9472));
  OAI21xp33_ASAP7_75t_L     g09216(.A1(new_n9472), .A2(new_n9470), .B(new_n9393), .Y(new_n9473));
  XNOR2x2_ASAP7_75t_L       g09217(.A(\a[41] ), .B(new_n9392), .Y(new_n9474));
  NAND3xp33_ASAP7_75t_L     g09218(.A(new_n9471), .B(new_n9465), .C(new_n9468), .Y(new_n9475));
  NAND3xp33_ASAP7_75t_L     g09219(.A(new_n9161), .B(new_n9469), .C(new_n9395), .Y(new_n9476));
  NAND3xp33_ASAP7_75t_L     g09220(.A(new_n9476), .B(new_n9475), .C(new_n9474), .Y(new_n9477));
  NAND2xp33_ASAP7_75t_L     g09221(.A(new_n9477), .B(new_n9473), .Y(new_n9478));
  A2O1A1Ixp33_ASAP7_75t_L   g09222(.A1(new_n9164), .A2(new_n9166), .B(new_n9390), .C(new_n9478), .Y(new_n9479));
  AOI21xp33_ASAP7_75t_L     g09223(.A1(new_n9164), .A2(new_n9166), .B(new_n9390), .Y(new_n9480));
  AOI21xp33_ASAP7_75t_L     g09224(.A1(new_n9476), .A2(new_n9475), .B(new_n9474), .Y(new_n9481));
  NOR3xp33_ASAP7_75t_L      g09225(.A(new_n9470), .B(new_n9393), .C(new_n9472), .Y(new_n9482));
  NOR2xp33_ASAP7_75t_L      g09226(.A(new_n9481), .B(new_n9482), .Y(new_n9483));
  NAND2xp33_ASAP7_75t_L     g09227(.A(new_n9480), .B(new_n9483), .Y(new_n9484));
  NAND3xp33_ASAP7_75t_L     g09228(.A(new_n9479), .B(new_n9484), .C(new_n9389), .Y(new_n9485));
  NOR2xp33_ASAP7_75t_L      g09229(.A(new_n9480), .B(new_n9483), .Y(new_n9486));
  AO21x2_ASAP7_75t_L        g09230(.A1(new_n9166), .A2(new_n9164), .B(new_n9390), .Y(new_n9487));
  NOR2xp33_ASAP7_75t_L      g09231(.A(new_n9478), .B(new_n9487), .Y(new_n9488));
  OAI21xp33_ASAP7_75t_L     g09232(.A1(new_n9486), .A2(new_n9488), .B(new_n9388), .Y(new_n9489));
  NAND3xp33_ASAP7_75t_L     g09233(.A(new_n9385), .B(new_n9485), .C(new_n9489), .Y(new_n9490));
  NOR3xp33_ASAP7_75t_L      g09234(.A(new_n9488), .B(new_n9486), .C(new_n9388), .Y(new_n9491));
  AOI21xp33_ASAP7_75t_L     g09235(.A1(new_n9479), .A2(new_n9484), .B(new_n9389), .Y(new_n9492));
  OAI211xp5_ASAP7_75t_L     g09236(.A1(new_n9491), .A2(new_n9492), .B(new_n9181), .C(new_n9172), .Y(new_n9493));
  AOI22xp33_ASAP7_75t_L     g09237(.A1(new_n3633), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n3858), .Y(new_n9494));
  OAI221xp5_ASAP7_75t_L     g09238(.A1(new_n3853), .A2(new_n1909), .B1(new_n3856), .B2(new_n2477), .C(new_n9494), .Y(new_n9495));
  XNOR2x2_ASAP7_75t_L       g09239(.A(\a[35] ), .B(new_n9495), .Y(new_n9496));
  NAND3xp33_ASAP7_75t_L     g09240(.A(new_n9496), .B(new_n9490), .C(new_n9493), .Y(new_n9497));
  AO21x2_ASAP7_75t_L        g09241(.A1(new_n9493), .A2(new_n9490), .B(new_n9496), .Y(new_n9498));
  A2O1A1O1Ixp25_ASAP7_75t_L g09242(.A1(new_n8789), .A2(new_n8911), .B(new_n8915), .C(new_n9187), .D(new_n9179), .Y(new_n9499));
  NAND3xp33_ASAP7_75t_L     g09243(.A(new_n9498), .B(new_n9499), .C(new_n9497), .Y(new_n9500));
  INVx1_ASAP7_75t_L         g09244(.A(new_n9500), .Y(new_n9501));
  AOI21xp33_ASAP7_75t_L     g09245(.A1(new_n9498), .A2(new_n9497), .B(new_n9499), .Y(new_n9502));
  AOI22xp33_ASAP7_75t_L     g09246(.A1(new_n3029), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n3258), .Y(new_n9503));
  OAI221xp5_ASAP7_75t_L     g09247(.A1(new_n3024), .A2(new_n2348), .B1(new_n3256), .B2(new_n2505), .C(new_n9503), .Y(new_n9504));
  XNOR2x2_ASAP7_75t_L       g09248(.A(\a[32] ), .B(new_n9504), .Y(new_n9505));
  OAI21xp33_ASAP7_75t_L     g09249(.A1(new_n9502), .A2(new_n9501), .B(new_n9505), .Y(new_n9506));
  AO21x2_ASAP7_75t_L        g09250(.A1(new_n9497), .A2(new_n9498), .B(new_n9499), .Y(new_n9507));
  INVx1_ASAP7_75t_L         g09251(.A(new_n9505), .Y(new_n9508));
  NAND3xp33_ASAP7_75t_L     g09252(.A(new_n9507), .B(new_n9508), .C(new_n9500), .Y(new_n9509));
  OAI211xp5_ASAP7_75t_L     g09253(.A1(new_n8926), .A2(new_n8928), .B(new_n9082), .C(new_n9200), .Y(new_n9510));
  AND4x1_ASAP7_75t_L        g09254(.A(new_n9510), .B(new_n9509), .C(new_n9506), .D(new_n9199), .Y(new_n9511));
  AOI22xp33_ASAP7_75t_L     g09255(.A1(new_n9506), .A2(new_n9509), .B1(new_n9510), .B2(new_n9199), .Y(new_n9512));
  NOR3xp33_ASAP7_75t_L      g09256(.A(new_n9511), .B(new_n9512), .C(new_n9383), .Y(new_n9513));
  INVx1_ASAP7_75t_L         g09257(.A(new_n9383), .Y(new_n9514));
  NAND4xp25_ASAP7_75t_L     g09258(.A(new_n9510), .B(new_n9506), .C(new_n9199), .D(new_n9509), .Y(new_n9515));
  AO22x1_ASAP7_75t_L        g09259(.A1(new_n9509), .A2(new_n9506), .B1(new_n9510), .B2(new_n9199), .Y(new_n9516));
  AOI21xp33_ASAP7_75t_L     g09260(.A1(new_n9516), .A2(new_n9515), .B(new_n9514), .Y(new_n9517));
  NOR2xp33_ASAP7_75t_L      g09261(.A(new_n9513), .B(new_n9517), .Y(new_n9518));
  A2O1A1Ixp33_ASAP7_75t_L   g09262(.A1(new_n9217), .A2(new_n9213), .B(new_n9376), .C(new_n9518), .Y(new_n9519));
  NOR2xp33_ASAP7_75t_L      g09263(.A(new_n8936), .B(new_n9076), .Y(new_n9520));
  A2O1A1O1Ixp25_ASAP7_75t_L g09264(.A1(new_n8942), .A2(new_n8943), .B(new_n9520), .C(new_n9203), .D(new_n9376), .Y(new_n9521));
  NAND3xp33_ASAP7_75t_L     g09265(.A(new_n9516), .B(new_n9514), .C(new_n9515), .Y(new_n9522));
  OAI21xp33_ASAP7_75t_L     g09266(.A1(new_n9512), .A2(new_n9511), .B(new_n9383), .Y(new_n9523));
  NAND2xp33_ASAP7_75t_L     g09267(.A(new_n9522), .B(new_n9523), .Y(new_n9524));
  NAND2xp33_ASAP7_75t_L     g09268(.A(new_n9521), .B(new_n9524), .Y(new_n9525));
  AOI22xp33_ASAP7_75t_L     g09269(.A1(new_n2114), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n2259), .Y(new_n9526));
  OAI221xp5_ASAP7_75t_L     g09270(.A1(new_n2109), .A2(new_n3207), .B1(new_n2257), .B2(new_n3572), .C(new_n9526), .Y(new_n9527));
  XNOR2x2_ASAP7_75t_L       g09271(.A(\a[26] ), .B(new_n9527), .Y(new_n9528));
  NAND3xp33_ASAP7_75t_L     g09272(.A(new_n9519), .B(new_n9528), .C(new_n9525), .Y(new_n9529));
  INVx1_ASAP7_75t_L         g09273(.A(new_n9213), .Y(new_n9530));
  O2A1O1Ixp33_ASAP7_75t_L   g09274(.A1(new_n9530), .A2(new_n9210), .B(new_n9209), .C(new_n9524), .Y(new_n9531));
  AOI221xp5_ASAP7_75t_L     g09275(.A1(new_n9213), .A2(new_n9203), .B1(new_n9522), .B2(new_n9523), .C(new_n9376), .Y(new_n9532));
  INVx1_ASAP7_75t_L         g09276(.A(new_n9528), .Y(new_n9533));
  OAI21xp33_ASAP7_75t_L     g09277(.A1(new_n9532), .A2(new_n9531), .B(new_n9533), .Y(new_n9534));
  NAND2xp33_ASAP7_75t_L     g09278(.A(new_n9534), .B(new_n9529), .Y(new_n9535));
  A2O1A1Ixp33_ASAP7_75t_L   g09279(.A1(new_n9215), .A2(new_n9068), .B(new_n9225), .C(new_n9535), .Y(new_n9536));
  NOR2xp33_ASAP7_75t_L      g09280(.A(new_n8949), .B(new_n9067), .Y(new_n9537));
  A2O1A1O1Ixp25_ASAP7_75t_L g09281(.A1(new_n8966), .A2(new_n8960), .B(new_n9537), .C(new_n9215), .D(new_n9225), .Y(new_n9538));
  NAND3xp33_ASAP7_75t_L     g09282(.A(new_n9538), .B(new_n9529), .C(new_n9534), .Y(new_n9539));
  NAND3xp33_ASAP7_75t_L     g09283(.A(new_n9536), .B(new_n9375), .C(new_n9539), .Y(new_n9540));
  AOI21xp33_ASAP7_75t_L     g09284(.A1(new_n9534), .A2(new_n9529), .B(new_n9538), .Y(new_n9541));
  AND3x1_ASAP7_75t_L        g09285(.A(new_n9538), .B(new_n9534), .C(new_n9529), .Y(new_n9542));
  OAI21xp33_ASAP7_75t_L     g09286(.A1(new_n9541), .A2(new_n9542), .B(new_n9374), .Y(new_n9543));
  NAND2xp33_ASAP7_75t_L     g09287(.A(new_n9543), .B(new_n9540), .Y(new_n9544));
  NAND3xp33_ASAP7_75t_L     g09288(.A(new_n9544), .B(new_n9371), .C(new_n9252), .Y(new_n9545));
  A2O1A1Ixp33_ASAP7_75t_L   g09289(.A1(new_n9238), .A2(new_n9234), .B(new_n9244), .C(new_n9371), .Y(new_n9546));
  NAND3xp33_ASAP7_75t_L     g09290(.A(new_n9546), .B(new_n9540), .C(new_n9543), .Y(new_n9547));
  AOI22xp33_ASAP7_75t_L     g09291(.A1(new_n1360), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1581), .Y(new_n9548));
  OAI221xp5_ASAP7_75t_L     g09292(.A1(new_n1373), .A2(new_n4632), .B1(new_n1359), .B2(new_n4858), .C(new_n9548), .Y(new_n9549));
  XNOR2x2_ASAP7_75t_L       g09293(.A(\a[20] ), .B(new_n9549), .Y(new_n9550));
  NAND3xp33_ASAP7_75t_L     g09294(.A(new_n9545), .B(new_n9547), .C(new_n9550), .Y(new_n9551));
  AOI21xp33_ASAP7_75t_L     g09295(.A1(new_n9543), .A2(new_n9540), .B(new_n9546), .Y(new_n9552));
  AOI21xp33_ASAP7_75t_L     g09296(.A1(new_n9371), .A2(new_n9252), .B(new_n9544), .Y(new_n9553));
  INVx1_ASAP7_75t_L         g09297(.A(new_n9550), .Y(new_n9554));
  OAI21xp33_ASAP7_75t_L     g09298(.A1(new_n9552), .A2(new_n9553), .B(new_n9554), .Y(new_n9555));
  NOR2xp33_ASAP7_75t_L      g09299(.A(new_n9242), .B(new_n9245), .Y(new_n9556));
  MAJIxp5_ASAP7_75t_L       g09300(.A(new_n9255), .B(new_n9249), .C(new_n9556), .Y(new_n9557));
  NAND3xp33_ASAP7_75t_L     g09301(.A(new_n9557), .B(new_n9555), .C(new_n9551), .Y(new_n9558));
  AO21x2_ASAP7_75t_L        g09302(.A1(new_n9551), .A2(new_n9555), .B(new_n9557), .Y(new_n9559));
  NAND2xp33_ASAP7_75t_L     g09303(.A(\b[41] ), .B(new_n1080), .Y(new_n9560));
  NAND3xp33_ASAP7_75t_L     g09304(.A(new_n5343), .B(new_n1073), .C(new_n5345), .Y(new_n9561));
  AOI22xp33_ASAP7_75t_L     g09305(.A1(new_n1076), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n1253), .Y(new_n9562));
  AND4x1_ASAP7_75t_L        g09306(.A(new_n9562), .B(new_n9561), .C(new_n9560), .D(\a[17] ), .Y(new_n9563));
  AOI31xp33_ASAP7_75t_L     g09307(.A1(new_n9561), .A2(new_n9560), .A3(new_n9562), .B(\a[17] ), .Y(new_n9564));
  NOR2xp33_ASAP7_75t_L      g09308(.A(new_n9564), .B(new_n9563), .Y(new_n9565));
  INVx1_ASAP7_75t_L         g09309(.A(new_n9565), .Y(new_n9566));
  AOI21xp33_ASAP7_75t_L     g09310(.A1(new_n9559), .A2(new_n9558), .B(new_n9566), .Y(new_n9567));
  NAND2xp33_ASAP7_75t_L     g09311(.A(new_n9249), .B(new_n9556), .Y(new_n9568));
  AND4x1_ASAP7_75t_L        g09312(.A(new_n9271), .B(new_n9568), .C(new_n9551), .D(new_n9555), .Y(new_n9569));
  AOI21xp33_ASAP7_75t_L     g09313(.A1(new_n9555), .A2(new_n9551), .B(new_n9557), .Y(new_n9570));
  NOR3xp33_ASAP7_75t_L      g09314(.A(new_n9569), .B(new_n9570), .C(new_n9565), .Y(new_n9571));
  NOR2xp33_ASAP7_75t_L      g09315(.A(new_n9571), .B(new_n9567), .Y(new_n9572));
  NAND2xp33_ASAP7_75t_L     g09316(.A(new_n9572), .B(new_n9369), .Y(new_n9573));
  OAI221xp5_ASAP7_75t_L     g09317(.A1(new_n9276), .A2(new_n9274), .B1(new_n9567), .B2(new_n9571), .C(new_n9368), .Y(new_n9574));
  AOI21xp33_ASAP7_75t_L     g09318(.A1(new_n9573), .A2(new_n9574), .B(new_n9366), .Y(new_n9575));
  INVx1_ASAP7_75t_L         g09319(.A(new_n9366), .Y(new_n9576));
  A2O1A1O1Ixp25_ASAP7_75t_L g09320(.A1(new_n9000), .A2(new_n8998), .B(new_n9275), .C(new_n9280), .D(new_n9367), .Y(new_n9577));
  OAI21xp33_ASAP7_75t_L     g09321(.A1(new_n9570), .A2(new_n9569), .B(new_n9565), .Y(new_n9578));
  NAND3xp33_ASAP7_75t_L     g09322(.A(new_n9559), .B(new_n9558), .C(new_n9566), .Y(new_n9579));
  NAND2xp33_ASAP7_75t_L     g09323(.A(new_n9578), .B(new_n9579), .Y(new_n9580));
  NOR2xp33_ASAP7_75t_L      g09324(.A(new_n9580), .B(new_n9577), .Y(new_n9581));
  AO21x2_ASAP7_75t_L        g09325(.A1(new_n8998), .A2(new_n9000), .B(new_n9275), .Y(new_n9582));
  AOI221xp5_ASAP7_75t_L     g09326(.A1(new_n9579), .A2(new_n9578), .B1(new_n9280), .B2(new_n9582), .C(new_n9367), .Y(new_n9583));
  NOR3xp33_ASAP7_75t_L      g09327(.A(new_n9581), .B(new_n9583), .C(new_n9576), .Y(new_n9584));
  A2O1A1O1Ixp25_ASAP7_75t_L g09328(.A1(new_n8788), .A2(new_n9292), .B(new_n9006), .C(new_n9288), .D(new_n9286), .Y(new_n9585));
  OA21x2_ASAP7_75t_L        g09329(.A1(new_n9575), .A2(new_n9584), .B(new_n9585), .Y(new_n9586));
  NOR3xp33_ASAP7_75t_L      g09330(.A(new_n9585), .B(new_n9584), .C(new_n9575), .Y(new_n9587));
  OAI21xp33_ASAP7_75t_L     g09331(.A1(new_n9587), .A2(new_n9586), .B(new_n9359), .Y(new_n9588));
  INVx1_ASAP7_75t_L         g09332(.A(new_n9356), .Y(new_n9589));
  NOR2xp33_ASAP7_75t_L      g09333(.A(new_n9357), .B(new_n9589), .Y(new_n9590));
  OAI21xp33_ASAP7_75t_L     g09334(.A1(new_n9575), .A2(new_n9584), .B(new_n9585), .Y(new_n9591));
  OR3x1_ASAP7_75t_L         g09335(.A(new_n9585), .B(new_n9584), .C(new_n9575), .Y(new_n9592));
  NAND3xp33_ASAP7_75t_L     g09336(.A(new_n9592), .B(new_n9591), .C(new_n9590), .Y(new_n9593));
  NAND2xp33_ASAP7_75t_L     g09337(.A(new_n9588), .B(new_n9593), .Y(new_n9594));
  A2O1A1Ixp33_ASAP7_75t_L   g09338(.A1(new_n9297), .A2(new_n9063), .B(new_n9295), .C(new_n9594), .Y(new_n9595));
  A2O1A1O1Ixp25_ASAP7_75t_L g09339(.A1(new_n9017), .A2(new_n9016), .B(new_n9013), .C(new_n9297), .D(new_n9295), .Y(new_n9596));
  NAND3xp33_ASAP7_75t_L     g09340(.A(new_n9596), .B(new_n9588), .C(new_n9593), .Y(new_n9597));
  AOI21xp33_ASAP7_75t_L     g09341(.A1(new_n9595), .A2(new_n9597), .B(new_n9351), .Y(new_n9598));
  INVx1_ASAP7_75t_L         g09342(.A(new_n9351), .Y(new_n9599));
  AOI21xp33_ASAP7_75t_L     g09343(.A1(new_n9593), .A2(new_n9588), .B(new_n9596), .Y(new_n9600));
  OAI21xp33_ASAP7_75t_L     g09344(.A1(new_n9301), .A2(new_n9300), .B(new_n9296), .Y(new_n9601));
  NOR2xp33_ASAP7_75t_L      g09345(.A(new_n9594), .B(new_n9601), .Y(new_n9602));
  NOR3xp33_ASAP7_75t_L      g09346(.A(new_n9602), .B(new_n9599), .C(new_n9600), .Y(new_n9603));
  OA21x2_ASAP7_75t_L        g09347(.A1(new_n9598), .A2(new_n9603), .B(new_n9348), .Y(new_n9604));
  OAI21xp33_ASAP7_75t_L     g09348(.A1(new_n9600), .A2(new_n9602), .B(new_n9599), .Y(new_n9605));
  NAND3xp33_ASAP7_75t_L     g09349(.A(new_n9595), .B(new_n9351), .C(new_n9597), .Y(new_n9606));
  NAND2xp33_ASAP7_75t_L     g09350(.A(new_n9606), .B(new_n9605), .Y(new_n9607));
  NOR2xp33_ASAP7_75t_L      g09351(.A(new_n9348), .B(new_n9607), .Y(new_n9608));
  OAI21xp33_ASAP7_75t_L     g09352(.A1(new_n9604), .A2(new_n9608), .B(new_n9346), .Y(new_n9609));
  NAND2xp33_ASAP7_75t_L     g09353(.A(new_n9348), .B(new_n9607), .Y(new_n9610));
  OR3x1_ASAP7_75t_L         g09354(.A(new_n9348), .B(new_n9598), .C(new_n9603), .Y(new_n9611));
  NAND3xp33_ASAP7_75t_L     g09355(.A(new_n9611), .B(new_n9610), .C(new_n9345), .Y(new_n9612));
  NAND3xp33_ASAP7_75t_L     g09356(.A(new_n9340), .B(new_n9609), .C(new_n9612), .Y(new_n9613));
  A2O1A1O1Ixp25_ASAP7_75t_L g09357(.A1(new_n9035), .A2(new_n9316), .B(new_n9037), .C(new_n9307), .D(new_n9319), .Y(new_n9614));
  INVx1_ASAP7_75t_L         g09358(.A(new_n9609), .Y(new_n9615));
  NOR3xp33_ASAP7_75t_L      g09359(.A(new_n9608), .B(new_n9604), .C(new_n9346), .Y(new_n9616));
  OAI21xp33_ASAP7_75t_L     g09360(.A1(new_n9616), .A2(new_n9615), .B(new_n9614), .Y(new_n9617));
  INVx1_ASAP7_75t_L         g09361(.A(new_n9324), .Y(new_n9618));
  NOR2xp33_ASAP7_75t_L      g09362(.A(\b[56] ), .B(\b[57] ), .Y(new_n9619));
  INVx1_ASAP7_75t_L         g09363(.A(\b[57] ), .Y(new_n9620));
  NOR2xp33_ASAP7_75t_L      g09364(.A(new_n9323), .B(new_n9620), .Y(new_n9621));
  NOR2xp33_ASAP7_75t_L      g09365(.A(new_n9619), .B(new_n9621), .Y(new_n9622));
  INVx1_ASAP7_75t_L         g09366(.A(new_n9622), .Y(new_n9623));
  O2A1O1Ixp33_ASAP7_75t_L   g09367(.A1(new_n9326), .A2(new_n9329), .B(new_n9618), .C(new_n9623), .Y(new_n9624));
  INVx1_ASAP7_75t_L         g09368(.A(new_n9624), .Y(new_n9625));
  NAND3xp33_ASAP7_75t_L     g09369(.A(new_n9328), .B(new_n9618), .C(new_n9623), .Y(new_n9626));
  NAND2xp33_ASAP7_75t_L     g09370(.A(new_n9625), .B(new_n9626), .Y(new_n9627));
  AOI22xp33_ASAP7_75t_L     g09371(.A1(\b[55] ), .A2(new_n282), .B1(\b[57] ), .B2(new_n303), .Y(new_n9628));
  OAI221xp5_ASAP7_75t_L     g09372(.A1(new_n291), .A2(new_n9323), .B1(new_n268), .B2(new_n9627), .C(new_n9628), .Y(new_n9629));
  XNOR2x2_ASAP7_75t_L       g09373(.A(\a[2] ), .B(new_n9629), .Y(new_n9630));
  AOI21xp33_ASAP7_75t_L     g09374(.A1(new_n9617), .A2(new_n9613), .B(new_n9630), .Y(new_n9631));
  INVx1_ASAP7_75t_L         g09375(.A(new_n9631), .Y(new_n9632));
  NAND3xp33_ASAP7_75t_L     g09376(.A(new_n9617), .B(new_n9613), .C(new_n9630), .Y(new_n9633));
  AND3x1_ASAP7_75t_L        g09377(.A(new_n9632), .B(new_n9633), .C(new_n9339), .Y(new_n9634));
  AOI21xp33_ASAP7_75t_L     g09378(.A1(new_n9632), .A2(new_n9633), .B(new_n9339), .Y(new_n9635));
  NOR2xp33_ASAP7_75t_L      g09379(.A(new_n9635), .B(new_n9634), .Y(\f[57] ));
  NAND2xp33_ASAP7_75t_L     g09380(.A(new_n9610), .B(new_n9611), .Y(new_n9637));
  MAJIxp5_ASAP7_75t_L       g09381(.A(new_n9614), .B(new_n9345), .C(new_n9637), .Y(new_n9638));
  AOI22xp33_ASAP7_75t_L     g09382(.A1(new_n344), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n370), .Y(new_n9639));
  OAI221xp5_ASAP7_75t_L     g09383(.A1(new_n429), .A2(new_n8458), .B1(new_n366), .B2(new_n8768), .C(new_n9639), .Y(new_n9640));
  XNOR2x2_ASAP7_75t_L       g09384(.A(\a[5] ), .B(new_n9640), .Y(new_n9641));
  NOR3xp33_ASAP7_75t_L      g09385(.A(new_n9602), .B(new_n9600), .C(new_n9351), .Y(new_n9642));
  O2A1O1Ixp33_ASAP7_75t_L   g09386(.A1(new_n9598), .A2(new_n9603), .B(new_n9348), .C(new_n9642), .Y(new_n9643));
  AOI22xp33_ASAP7_75t_L     g09387(.A1(new_n444), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n471), .Y(new_n9644));
  OAI221xp5_ASAP7_75t_L     g09388(.A1(new_n468), .A2(new_n7616), .B1(new_n469), .B2(new_n7906), .C(new_n9644), .Y(new_n9645));
  XNOR2x2_ASAP7_75t_L       g09389(.A(new_n435), .B(new_n9645), .Y(new_n9646));
  NAND2xp33_ASAP7_75t_L     g09390(.A(new_n9591), .B(new_n9592), .Y(new_n9647));
  MAJIxp5_ASAP7_75t_L       g09391(.A(new_n9596), .B(new_n9590), .C(new_n9647), .Y(new_n9648));
  AOI22xp33_ASAP7_75t_L     g09392(.A1(\b[47] ), .A2(new_n651), .B1(\b[49] ), .B2(new_n581), .Y(new_n9649));
  OAI221xp5_ASAP7_75t_L     g09393(.A1(new_n821), .A2(new_n6830), .B1(new_n577), .B2(new_n7323), .C(new_n9649), .Y(new_n9650));
  XNOR2x2_ASAP7_75t_L       g09394(.A(\a[11] ), .B(new_n9650), .Y(new_n9651));
  NOR3xp33_ASAP7_75t_L      g09395(.A(new_n9581), .B(new_n9583), .C(new_n9366), .Y(new_n9652));
  O2A1O1Ixp33_ASAP7_75t_L   g09396(.A1(new_n9575), .A2(new_n9584), .B(new_n9585), .C(new_n9652), .Y(new_n9653));
  AOI22xp33_ASAP7_75t_L     g09397(.A1(new_n811), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n900), .Y(new_n9654));
  OAI221xp5_ASAP7_75t_L     g09398(.A1(new_n904), .A2(new_n6321), .B1(new_n898), .B2(new_n6573), .C(new_n9654), .Y(new_n9655));
  XNOR2x2_ASAP7_75t_L       g09399(.A(\a[14] ), .B(new_n9655), .Y(new_n9656));
  A2O1A1O1Ixp25_ASAP7_75t_L g09400(.A1(new_n9280), .A2(new_n9582), .B(new_n9367), .C(new_n9578), .D(new_n9571), .Y(new_n9657));
  A2O1A1O1Ixp25_ASAP7_75t_L g09401(.A1(new_n9203), .A2(new_n9213), .B(new_n9376), .C(new_n9523), .D(new_n9513), .Y(new_n9658));
  NOR3xp33_ASAP7_75t_L      g09402(.A(new_n9501), .B(new_n9502), .C(new_n9505), .Y(new_n9659));
  AO31x2_ASAP7_75t_L        g09403(.A1(new_n9510), .A2(new_n9506), .A3(new_n9199), .B(new_n9659), .Y(new_n9660));
  A2O1A1Ixp33_ASAP7_75t_L   g09404(.A1(new_n9181), .A2(new_n9172), .B(new_n9492), .C(new_n9485), .Y(new_n9661));
  AOI22xp33_ASAP7_75t_L     g09405(.A1(new_n4283), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n4512), .Y(new_n9662));
  OAI221xp5_ASAP7_75t_L     g09406(.A1(new_n4277), .A2(new_n1655), .B1(new_n4499), .B2(new_n1780), .C(new_n9662), .Y(new_n9663));
  XNOR2x2_ASAP7_75t_L       g09407(.A(\a[38] ), .B(new_n9663), .Y(new_n9664));
  INVx1_ASAP7_75t_L         g09408(.A(new_n9664), .Y(new_n9665));
  NOR3xp33_ASAP7_75t_L      g09409(.A(new_n9470), .B(new_n9472), .C(new_n9474), .Y(new_n9666));
  INVx1_ASAP7_75t_L         g09410(.A(new_n9666), .Y(new_n9667));
  NOR3xp33_ASAP7_75t_L      g09411(.A(new_n9467), .B(new_n9466), .C(new_n9398), .Y(new_n9668));
  AOI22xp33_ASAP7_75t_L     g09412(.A1(new_n5624), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n5901), .Y(new_n9669));
  OAI221xp5_ASAP7_75t_L     g09413(.A1(new_n5900), .A2(new_n942), .B1(new_n5892), .B2(new_n1035), .C(new_n9669), .Y(new_n9670));
  XNOR2x2_ASAP7_75t_L       g09414(.A(\a[44] ), .B(new_n9670), .Y(new_n9671));
  INVx1_ASAP7_75t_L         g09415(.A(new_n9671), .Y(new_n9672));
  OAI211xp5_ASAP7_75t_L     g09416(.A1(new_n9460), .A2(new_n9461), .B(new_n9406), .C(new_n9405), .Y(new_n9673));
  A2O1A1O1Ixp25_ASAP7_75t_L g09417(.A1(new_n9143), .A2(new_n9154), .B(new_n9400), .C(new_n9673), .D(new_n9462), .Y(new_n9674));
  AOI211xp5_ASAP7_75t_L     g09418(.A1(new_n9431), .A2(new_n9433), .B(new_n9436), .C(new_n9435), .Y(new_n9675));
  AOI221xp5_ASAP7_75t_L     g09419(.A1(new_n9129), .A2(new_n9103), .B1(new_n9438), .B2(new_n9434), .C(new_n9122), .Y(new_n9676));
  AOI22xp33_ASAP7_75t_L     g09420(.A1(new_n7960), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n8537), .Y(new_n9677));
  OAI221xp5_ASAP7_75t_L     g09421(.A1(new_n8817), .A2(new_n418), .B1(new_n7957), .B2(new_n425), .C(new_n9677), .Y(new_n9678));
  XNOR2x2_ASAP7_75t_L       g09422(.A(\a[53] ), .B(new_n9678), .Y(new_n9679));
  NOR2xp33_ASAP7_75t_L      g09423(.A(new_n9120), .B(new_n9117), .Y(new_n9680));
  NAND2xp33_ASAP7_75t_L     g09424(.A(new_n9421), .B(new_n9423), .Y(new_n9681));
  MAJIxp5_ASAP7_75t_L       g09425(.A(new_n9681), .B(new_n9413), .C(new_n9680), .Y(new_n9682));
  NAND2xp33_ASAP7_75t_L     g09426(.A(\b[3] ), .B(new_n8835), .Y(new_n9683));
  NAND2xp33_ASAP7_75t_L     g09427(.A(new_n8828), .B(new_n329), .Y(new_n9684));
  AOI22xp33_ASAP7_75t_L     g09428(.A1(new_n8831), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n9115), .Y(new_n9685));
  NAND4xp25_ASAP7_75t_L     g09429(.A(new_n9684), .B(\a[56] ), .C(new_n9683), .D(new_n9685), .Y(new_n9686));
  INVx1_ASAP7_75t_L         g09430(.A(new_n9686), .Y(new_n9687));
  AOI31xp33_ASAP7_75t_L     g09431(.A1(new_n9684), .A2(new_n9683), .A3(new_n9685), .B(\a[56] ), .Y(new_n9688));
  NAND2xp33_ASAP7_75t_L     g09432(.A(\a[59] ), .B(new_n9413), .Y(new_n9689));
  NAND2xp33_ASAP7_75t_L     g09433(.A(new_n9411), .B(new_n9410), .Y(new_n9690));
  INVx1_ASAP7_75t_L         g09434(.A(\a[58] ), .Y(new_n9691));
  NAND2xp33_ASAP7_75t_L     g09435(.A(\a[59] ), .B(new_n9691), .Y(new_n9692));
  INVx1_ASAP7_75t_L         g09436(.A(\a[59] ), .Y(new_n9693));
  NAND2xp33_ASAP7_75t_L     g09437(.A(\a[58] ), .B(new_n9693), .Y(new_n9694));
  NAND2xp33_ASAP7_75t_L     g09438(.A(new_n9694), .B(new_n9692), .Y(new_n9695));
  NAND2xp33_ASAP7_75t_L     g09439(.A(new_n9695), .B(new_n9690), .Y(new_n9696));
  INVx1_ASAP7_75t_L         g09440(.A(new_n9696), .Y(new_n9697));
  NAND2xp33_ASAP7_75t_L     g09441(.A(new_n269), .B(new_n9697), .Y(new_n9698));
  NAND3xp33_ASAP7_75t_L     g09442(.A(new_n9690), .B(new_n9692), .C(new_n9694), .Y(new_n9699));
  INVx1_ASAP7_75t_L         g09443(.A(new_n9699), .Y(new_n9700));
  NAND2xp33_ASAP7_75t_L     g09444(.A(\b[1] ), .B(new_n9700), .Y(new_n9701));
  XNOR2x2_ASAP7_75t_L       g09445(.A(\a[58] ), .B(\a[57] ), .Y(new_n9702));
  NOR2xp33_ASAP7_75t_L      g09446(.A(new_n9702), .B(new_n9690), .Y(new_n9703));
  NAND2xp33_ASAP7_75t_L     g09447(.A(\b[0] ), .B(new_n9703), .Y(new_n9704));
  NAND3xp33_ASAP7_75t_L     g09448(.A(new_n9701), .B(new_n9698), .C(new_n9704), .Y(new_n9705));
  XNOR2x2_ASAP7_75t_L       g09449(.A(new_n9689), .B(new_n9705), .Y(new_n9706));
  NOR3xp33_ASAP7_75t_L      g09450(.A(new_n9706), .B(new_n9688), .C(new_n9687), .Y(new_n9707));
  INVx1_ASAP7_75t_L         g09451(.A(new_n9688), .Y(new_n9708));
  XOR2x2_ASAP7_75t_L        g09452(.A(new_n9689), .B(new_n9705), .Y(new_n9709));
  AOI21xp33_ASAP7_75t_L     g09453(.A1(new_n9708), .A2(new_n9686), .B(new_n9709), .Y(new_n9710));
  NOR3xp33_ASAP7_75t_L      g09454(.A(new_n9682), .B(new_n9707), .C(new_n9710), .Y(new_n9711));
  NAND2xp33_ASAP7_75t_L     g09455(.A(new_n9413), .B(new_n9680), .Y(new_n9712));
  A2O1A1Ixp33_ASAP7_75t_L   g09456(.A1(new_n9417), .A2(new_n9414), .B(new_n9425), .C(new_n9712), .Y(new_n9713));
  NAND3xp33_ASAP7_75t_L     g09457(.A(new_n9709), .B(new_n9708), .C(new_n9686), .Y(new_n9714));
  OAI21xp33_ASAP7_75t_L     g09458(.A1(new_n9688), .A2(new_n9687), .B(new_n9706), .Y(new_n9715));
  AOI21xp33_ASAP7_75t_L     g09459(.A1(new_n9715), .A2(new_n9714), .B(new_n9713), .Y(new_n9716));
  OAI21xp33_ASAP7_75t_L     g09460(.A1(new_n9716), .A2(new_n9711), .B(new_n9679), .Y(new_n9717));
  INVx1_ASAP7_75t_L         g09461(.A(new_n9679), .Y(new_n9718));
  NAND3xp33_ASAP7_75t_L     g09462(.A(new_n9713), .B(new_n9714), .C(new_n9715), .Y(new_n9719));
  OAI21xp33_ASAP7_75t_L     g09463(.A1(new_n9707), .A2(new_n9710), .B(new_n9682), .Y(new_n9720));
  NAND3xp33_ASAP7_75t_L     g09464(.A(new_n9718), .B(new_n9719), .C(new_n9720), .Y(new_n9721));
  OAI211xp5_ASAP7_75t_L     g09465(.A1(new_n9675), .A2(new_n9676), .B(new_n9721), .C(new_n9717), .Y(new_n9722));
  NOR4xp25_ASAP7_75t_L      g09466(.A(new_n9435), .B(new_n9436), .C(new_n9432), .D(new_n9437), .Y(new_n9723));
  AOI22xp33_ASAP7_75t_L     g09467(.A1(new_n9431), .A2(new_n9433), .B1(new_n9426), .B2(new_n9424), .Y(new_n9724));
  O2A1O1Ixp33_ASAP7_75t_L   g09468(.A1(new_n9723), .A2(new_n9724), .B(new_n9441), .C(new_n9675), .Y(new_n9725));
  AOI21xp33_ASAP7_75t_L     g09469(.A1(new_n9720), .A2(new_n9719), .B(new_n9718), .Y(new_n9726));
  NOR3xp33_ASAP7_75t_L      g09470(.A(new_n9711), .B(new_n9716), .C(new_n9679), .Y(new_n9727));
  OAI21xp33_ASAP7_75t_L     g09471(.A1(new_n9726), .A2(new_n9727), .B(new_n9725), .Y(new_n9728));
  AOI22xp33_ASAP7_75t_L     g09472(.A1(new_n7111), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n7391), .Y(new_n9729));
  OAI221xp5_ASAP7_75t_L     g09473(.A1(new_n8558), .A2(new_n540), .B1(new_n8237), .B2(new_n624), .C(new_n9729), .Y(new_n9730));
  XNOR2x2_ASAP7_75t_L       g09474(.A(\a[50] ), .B(new_n9730), .Y(new_n9731));
  NAND3xp33_ASAP7_75t_L     g09475(.A(new_n9728), .B(new_n9722), .C(new_n9731), .Y(new_n9732));
  AO21x2_ASAP7_75t_L        g09476(.A1(new_n9722), .A2(new_n9728), .B(new_n9731), .Y(new_n9733));
  AOI22xp33_ASAP7_75t_L     g09477(.A1(new_n9452), .A2(new_n9446), .B1(new_n9449), .B2(new_n9451), .Y(new_n9734));
  A2O1A1O1Ixp25_ASAP7_75t_L g09478(.A1(new_n9135), .A2(new_n9134), .B(new_n9132), .C(new_n9453), .D(new_n9734), .Y(new_n9735));
  AND3x1_ASAP7_75t_L        g09479(.A(new_n9735), .B(new_n9733), .C(new_n9732), .Y(new_n9736));
  AOI21xp33_ASAP7_75t_L     g09480(.A1(new_n9733), .A2(new_n9732), .B(new_n9735), .Y(new_n9737));
  AOI22xp33_ASAP7_75t_L     g09481(.A1(new_n6376), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n6648), .Y(new_n9738));
  OAI221xp5_ASAP7_75t_L     g09482(.A1(new_n6646), .A2(new_n760), .B1(new_n6636), .B2(new_n790), .C(new_n9738), .Y(new_n9739));
  XNOR2x2_ASAP7_75t_L       g09483(.A(\a[47] ), .B(new_n9739), .Y(new_n9740));
  OAI21xp33_ASAP7_75t_L     g09484(.A1(new_n9737), .A2(new_n9736), .B(new_n9740), .Y(new_n9741));
  NAND3xp33_ASAP7_75t_L     g09485(.A(new_n9735), .B(new_n9733), .C(new_n9732), .Y(new_n9742));
  AO21x2_ASAP7_75t_L        g09486(.A1(new_n9732), .A2(new_n9733), .B(new_n9735), .Y(new_n9743));
  INVx1_ASAP7_75t_L         g09487(.A(new_n9740), .Y(new_n9744));
  NAND3xp33_ASAP7_75t_L     g09488(.A(new_n9744), .B(new_n9743), .C(new_n9742), .Y(new_n9745));
  NAND2xp33_ASAP7_75t_L     g09489(.A(new_n9741), .B(new_n9745), .Y(new_n9746));
  NAND2xp33_ASAP7_75t_L     g09490(.A(new_n9746), .B(new_n9674), .Y(new_n9747));
  NAND3xp33_ASAP7_75t_L     g09491(.A(new_n9407), .B(new_n9454), .C(new_n9458), .Y(new_n9748));
  OAI21xp33_ASAP7_75t_L     g09492(.A1(new_n9459), .A2(new_n9401), .B(new_n9748), .Y(new_n9749));
  NAND3xp33_ASAP7_75t_L     g09493(.A(new_n9749), .B(new_n9741), .C(new_n9745), .Y(new_n9750));
  NAND3xp33_ASAP7_75t_L     g09494(.A(new_n9747), .B(new_n9672), .C(new_n9750), .Y(new_n9751));
  AOI21xp33_ASAP7_75t_L     g09495(.A1(new_n9745), .A2(new_n9741), .B(new_n9749), .Y(new_n9752));
  O2A1O1Ixp33_ASAP7_75t_L   g09496(.A1(new_n9401), .A2(new_n9459), .B(new_n9748), .C(new_n9746), .Y(new_n9753));
  OAI21xp33_ASAP7_75t_L     g09497(.A1(new_n9752), .A2(new_n9753), .B(new_n9671), .Y(new_n9754));
  AOI221xp5_ASAP7_75t_L     g09498(.A1(new_n9471), .A2(new_n9468), .B1(new_n9751), .B2(new_n9754), .C(new_n9668), .Y(new_n9755));
  NAND2xp33_ASAP7_75t_L     g09499(.A(new_n9751), .B(new_n9754), .Y(new_n9756));
  A2O1A1O1Ixp25_ASAP7_75t_L g09500(.A1(new_n9395), .A2(new_n9161), .B(new_n9469), .C(new_n9465), .D(new_n9756), .Y(new_n9757));
  AOI22xp33_ASAP7_75t_L     g09501(.A1(new_n4920), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n5167), .Y(new_n9758));
  OAI221xp5_ASAP7_75t_L     g09502(.A1(new_n5154), .A2(new_n1313), .B1(new_n5158), .B2(new_n1438), .C(new_n9758), .Y(new_n9759));
  XNOR2x2_ASAP7_75t_L       g09503(.A(\a[41] ), .B(new_n9759), .Y(new_n9760));
  OAI21xp33_ASAP7_75t_L     g09504(.A1(new_n9755), .A2(new_n9757), .B(new_n9760), .Y(new_n9761));
  INVx1_ASAP7_75t_L         g09505(.A(new_n9755), .Y(new_n9762));
  AO21x2_ASAP7_75t_L        g09506(.A1(new_n9468), .A2(new_n9471), .B(new_n9668), .Y(new_n9763));
  AND2x2_ASAP7_75t_L        g09507(.A(new_n9751), .B(new_n9754), .Y(new_n9764));
  NAND2xp33_ASAP7_75t_L     g09508(.A(new_n9763), .B(new_n9764), .Y(new_n9765));
  INVx1_ASAP7_75t_L         g09509(.A(new_n9760), .Y(new_n9766));
  NAND3xp33_ASAP7_75t_L     g09510(.A(new_n9765), .B(new_n9762), .C(new_n9766), .Y(new_n9767));
  NAND2xp33_ASAP7_75t_L     g09511(.A(new_n9761), .B(new_n9767), .Y(new_n9768));
  NAND3xp33_ASAP7_75t_L     g09512(.A(new_n9479), .B(new_n9768), .C(new_n9667), .Y(new_n9769));
  A2O1A1Ixp33_ASAP7_75t_L   g09513(.A1(new_n9473), .A2(new_n9477), .B(new_n9480), .C(new_n9667), .Y(new_n9770));
  NAND3xp33_ASAP7_75t_L     g09514(.A(new_n9770), .B(new_n9761), .C(new_n9767), .Y(new_n9771));
  NAND3xp33_ASAP7_75t_L     g09515(.A(new_n9771), .B(new_n9769), .C(new_n9665), .Y(new_n9772));
  AOI221xp5_ASAP7_75t_L     g09516(.A1(new_n9767), .A2(new_n9761), .B1(new_n9478), .B2(new_n9487), .C(new_n9666), .Y(new_n9773));
  O2A1O1Ixp33_ASAP7_75t_L   g09517(.A1(new_n9480), .A2(new_n9483), .B(new_n9667), .C(new_n9768), .Y(new_n9774));
  OAI21xp33_ASAP7_75t_L     g09518(.A1(new_n9773), .A2(new_n9774), .B(new_n9664), .Y(new_n9775));
  AOI21xp33_ASAP7_75t_L     g09519(.A1(new_n9775), .A2(new_n9772), .B(new_n9661), .Y(new_n9776));
  AOI21xp33_ASAP7_75t_L     g09520(.A1(new_n9385), .A2(new_n9489), .B(new_n9491), .Y(new_n9777));
  NAND2xp33_ASAP7_75t_L     g09521(.A(new_n9775), .B(new_n9772), .Y(new_n9778));
  NOR2xp33_ASAP7_75t_L      g09522(.A(new_n9777), .B(new_n9778), .Y(new_n9779));
  AOI22xp33_ASAP7_75t_L     g09523(.A1(new_n3633), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n3858), .Y(new_n9780));
  OAI221xp5_ASAP7_75t_L     g09524(.A1(new_n3853), .A2(new_n1929), .B1(new_n3856), .B2(new_n2075), .C(new_n9780), .Y(new_n9781));
  XNOR2x2_ASAP7_75t_L       g09525(.A(new_n3628), .B(new_n9781), .Y(new_n9782));
  NOR3xp33_ASAP7_75t_L      g09526(.A(new_n9779), .B(new_n9782), .C(new_n9776), .Y(new_n9783));
  NAND2xp33_ASAP7_75t_L     g09527(.A(new_n9777), .B(new_n9778), .Y(new_n9784));
  NAND3xp33_ASAP7_75t_L     g09528(.A(new_n9661), .B(new_n9772), .C(new_n9775), .Y(new_n9785));
  XNOR2x2_ASAP7_75t_L       g09529(.A(\a[35] ), .B(new_n9781), .Y(new_n9786));
  AOI21xp33_ASAP7_75t_L     g09530(.A1(new_n9784), .A2(new_n9785), .B(new_n9786), .Y(new_n9787));
  NAND2xp33_ASAP7_75t_L     g09531(.A(new_n9493), .B(new_n9490), .Y(new_n9788));
  MAJIxp5_ASAP7_75t_L       g09532(.A(new_n9499), .B(new_n9496), .C(new_n9788), .Y(new_n9789));
  NOR3xp33_ASAP7_75t_L      g09533(.A(new_n9789), .B(new_n9787), .C(new_n9783), .Y(new_n9790));
  OA21x2_ASAP7_75t_L        g09534(.A1(new_n9783), .A2(new_n9787), .B(new_n9789), .Y(new_n9791));
  AOI22xp33_ASAP7_75t_L     g09535(.A1(new_n3029), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n3258), .Y(new_n9792));
  OAI221xp5_ASAP7_75t_L     g09536(.A1(new_n3024), .A2(new_n2497), .B1(new_n3256), .B2(new_n2672), .C(new_n9792), .Y(new_n9793));
  XNOR2x2_ASAP7_75t_L       g09537(.A(\a[32] ), .B(new_n9793), .Y(new_n9794));
  INVx1_ASAP7_75t_L         g09538(.A(new_n9794), .Y(new_n9795));
  NOR3xp33_ASAP7_75t_L      g09539(.A(new_n9791), .B(new_n9795), .C(new_n9790), .Y(new_n9796));
  NAND3xp33_ASAP7_75t_L     g09540(.A(new_n9784), .B(new_n9785), .C(new_n9786), .Y(new_n9797));
  OAI21xp33_ASAP7_75t_L     g09541(.A1(new_n9776), .A2(new_n9779), .B(new_n9782), .Y(new_n9798));
  OR2x4_ASAP7_75t_L         g09542(.A(new_n9496), .B(new_n9788), .Y(new_n9799));
  NAND4xp25_ASAP7_75t_L     g09543(.A(new_n9507), .B(new_n9799), .C(new_n9798), .D(new_n9797), .Y(new_n9800));
  OAI21xp33_ASAP7_75t_L     g09544(.A1(new_n9787), .A2(new_n9783), .B(new_n9789), .Y(new_n9801));
  AOI21xp33_ASAP7_75t_L     g09545(.A1(new_n9800), .A2(new_n9801), .B(new_n9794), .Y(new_n9802));
  NOR2xp33_ASAP7_75t_L      g09546(.A(new_n9802), .B(new_n9796), .Y(new_n9803));
  NAND2xp33_ASAP7_75t_L     g09547(.A(new_n9660), .B(new_n9803), .Y(new_n9804));
  AOI31xp33_ASAP7_75t_L     g09548(.A1(new_n9510), .A2(new_n9506), .A3(new_n9199), .B(new_n9659), .Y(new_n9805));
  NAND3xp33_ASAP7_75t_L     g09549(.A(new_n9800), .B(new_n9801), .C(new_n9794), .Y(new_n9806));
  OAI21xp33_ASAP7_75t_L     g09550(.A1(new_n9790), .A2(new_n9791), .B(new_n9795), .Y(new_n9807));
  NAND2xp33_ASAP7_75t_L     g09551(.A(new_n9806), .B(new_n9807), .Y(new_n9808));
  NAND2xp33_ASAP7_75t_L     g09552(.A(new_n9805), .B(new_n9808), .Y(new_n9809));
  AOI22xp33_ASAP7_75t_L     g09553(.A1(new_n2552), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n2736), .Y(new_n9810));
  OAI221xp5_ASAP7_75t_L     g09554(.A1(new_n2547), .A2(new_n2982), .B1(new_n2734), .B2(new_n3187), .C(new_n9810), .Y(new_n9811));
  XNOR2x2_ASAP7_75t_L       g09555(.A(\a[29] ), .B(new_n9811), .Y(new_n9812));
  AOI21xp33_ASAP7_75t_L     g09556(.A1(new_n9804), .A2(new_n9809), .B(new_n9812), .Y(new_n9813));
  NOR2xp33_ASAP7_75t_L      g09557(.A(new_n9805), .B(new_n9808), .Y(new_n9814));
  NOR2xp33_ASAP7_75t_L      g09558(.A(new_n9660), .B(new_n9803), .Y(new_n9815));
  INVx1_ASAP7_75t_L         g09559(.A(new_n9812), .Y(new_n9816));
  NOR3xp33_ASAP7_75t_L      g09560(.A(new_n9815), .B(new_n9814), .C(new_n9816), .Y(new_n9817));
  OAI21xp33_ASAP7_75t_L     g09561(.A1(new_n9813), .A2(new_n9817), .B(new_n9658), .Y(new_n9818));
  OAI21xp33_ASAP7_75t_L     g09562(.A1(new_n9517), .A2(new_n9521), .B(new_n9522), .Y(new_n9819));
  OAI21xp33_ASAP7_75t_L     g09563(.A1(new_n9814), .A2(new_n9815), .B(new_n9816), .Y(new_n9820));
  NAND3xp33_ASAP7_75t_L     g09564(.A(new_n9804), .B(new_n9809), .C(new_n9812), .Y(new_n9821));
  NAND3xp33_ASAP7_75t_L     g09565(.A(new_n9819), .B(new_n9820), .C(new_n9821), .Y(new_n9822));
  AOI22xp33_ASAP7_75t_L     g09566(.A1(new_n2114), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n2259), .Y(new_n9823));
  OAI221xp5_ASAP7_75t_L     g09567(.A1(new_n2109), .A2(new_n3565), .B1(new_n2257), .B2(new_n3591), .C(new_n9823), .Y(new_n9824));
  XNOR2x2_ASAP7_75t_L       g09568(.A(\a[26] ), .B(new_n9824), .Y(new_n9825));
  NAND3xp33_ASAP7_75t_L     g09569(.A(new_n9822), .B(new_n9818), .C(new_n9825), .Y(new_n9826));
  AOI21xp33_ASAP7_75t_L     g09570(.A1(new_n9821), .A2(new_n9820), .B(new_n9819), .Y(new_n9827));
  NOR3xp33_ASAP7_75t_L      g09571(.A(new_n9658), .B(new_n9813), .C(new_n9817), .Y(new_n9828));
  INVx1_ASAP7_75t_L         g09572(.A(new_n9825), .Y(new_n9829));
  OAI21xp33_ASAP7_75t_L     g09573(.A1(new_n9828), .A2(new_n9827), .B(new_n9829), .Y(new_n9830));
  NAND2xp33_ASAP7_75t_L     g09574(.A(new_n9525), .B(new_n9519), .Y(new_n9831));
  NOR2xp33_ASAP7_75t_L      g09575(.A(new_n9528), .B(new_n9831), .Y(new_n9832));
  O2A1O1Ixp33_ASAP7_75t_L   g09576(.A1(new_n9225), .A2(new_n9235), .B(new_n9535), .C(new_n9832), .Y(new_n9833));
  NAND3xp33_ASAP7_75t_L     g09577(.A(new_n9833), .B(new_n9830), .C(new_n9826), .Y(new_n9834));
  NAND2xp33_ASAP7_75t_L     g09578(.A(new_n9826), .B(new_n9830), .Y(new_n9835));
  MAJIxp5_ASAP7_75t_L       g09579(.A(new_n9538), .B(new_n9831), .C(new_n9528), .Y(new_n9836));
  NAND2xp33_ASAP7_75t_L     g09580(.A(new_n9836), .B(new_n9835), .Y(new_n9837));
  AOI22xp33_ASAP7_75t_L     g09581(.A1(new_n1704), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1837), .Y(new_n9838));
  OAI221xp5_ASAP7_75t_L     g09582(.A1(new_n1699), .A2(new_n4216), .B1(new_n1827), .B2(new_n4431), .C(new_n9838), .Y(new_n9839));
  XNOR2x2_ASAP7_75t_L       g09583(.A(\a[23] ), .B(new_n9839), .Y(new_n9840));
  NAND3xp33_ASAP7_75t_L     g09584(.A(new_n9834), .B(new_n9837), .C(new_n9840), .Y(new_n9841));
  NOR2xp33_ASAP7_75t_L      g09585(.A(new_n9836), .B(new_n9835), .Y(new_n9842));
  AOI21xp33_ASAP7_75t_L     g09586(.A1(new_n9830), .A2(new_n9826), .B(new_n9833), .Y(new_n9843));
  INVx1_ASAP7_75t_L         g09587(.A(new_n9840), .Y(new_n9844));
  OAI21xp33_ASAP7_75t_L     g09588(.A1(new_n9842), .A2(new_n9843), .B(new_n9844), .Y(new_n9845));
  NOR3xp33_ASAP7_75t_L      g09589(.A(new_n9542), .B(new_n9541), .C(new_n9374), .Y(new_n9846));
  A2O1A1O1Ixp25_ASAP7_75t_L g09590(.A1(new_n9241), .A2(new_n9239), .B(new_n9370), .C(new_n9543), .D(new_n9846), .Y(new_n9847));
  AND3x1_ASAP7_75t_L        g09591(.A(new_n9847), .B(new_n9841), .C(new_n9845), .Y(new_n9848));
  AOI21xp33_ASAP7_75t_L     g09592(.A1(new_n9841), .A2(new_n9845), .B(new_n9847), .Y(new_n9849));
  NOR2xp33_ASAP7_75t_L      g09593(.A(new_n4848), .B(new_n1373), .Y(new_n9850));
  INVx1_ASAP7_75t_L         g09594(.A(new_n9850), .Y(new_n9851));
  NAND2xp33_ASAP7_75t_L     g09595(.A(new_n1365), .B(new_n4876), .Y(new_n9852));
  AOI22xp33_ASAP7_75t_L     g09596(.A1(new_n1360), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n1581), .Y(new_n9853));
  AND4x1_ASAP7_75t_L        g09597(.A(new_n9853), .B(new_n9852), .C(new_n9851), .D(\a[20] ), .Y(new_n9854));
  AOI31xp33_ASAP7_75t_L     g09598(.A1(new_n9852), .A2(new_n9851), .A3(new_n9853), .B(\a[20] ), .Y(new_n9855));
  NOR2xp33_ASAP7_75t_L      g09599(.A(new_n9855), .B(new_n9854), .Y(new_n9856));
  INVx1_ASAP7_75t_L         g09600(.A(new_n9856), .Y(new_n9857));
  NOR3xp33_ASAP7_75t_L      g09601(.A(new_n9848), .B(new_n9857), .C(new_n9849), .Y(new_n9858));
  NAND3xp33_ASAP7_75t_L     g09602(.A(new_n9847), .B(new_n9841), .C(new_n9845), .Y(new_n9859));
  AO21x2_ASAP7_75t_L        g09603(.A1(new_n9841), .A2(new_n9845), .B(new_n9847), .Y(new_n9860));
  AOI21xp33_ASAP7_75t_L     g09604(.A1(new_n9860), .A2(new_n9859), .B(new_n9856), .Y(new_n9861));
  NOR2xp33_ASAP7_75t_L      g09605(.A(new_n9861), .B(new_n9858), .Y(new_n9862));
  NAND2xp33_ASAP7_75t_L     g09606(.A(new_n9547), .B(new_n9545), .Y(new_n9863));
  MAJx2_ASAP7_75t_L         g09607(.A(new_n9557), .B(new_n9550), .C(new_n9863), .Y(new_n9864));
  NAND2xp33_ASAP7_75t_L     g09608(.A(new_n9862), .B(new_n9864), .Y(new_n9865));
  NAND3xp33_ASAP7_75t_L     g09609(.A(new_n9860), .B(new_n9859), .C(new_n9856), .Y(new_n9866));
  OAI21xp33_ASAP7_75t_L     g09610(.A1(new_n9849), .A2(new_n9848), .B(new_n9857), .Y(new_n9867));
  NAND2xp33_ASAP7_75t_L     g09611(.A(new_n9866), .B(new_n9867), .Y(new_n9868));
  NAND3xp33_ASAP7_75t_L     g09612(.A(new_n9545), .B(new_n9547), .C(new_n9554), .Y(new_n9869));
  A2O1A1Ixp33_ASAP7_75t_L   g09613(.A1(new_n9555), .A2(new_n9551), .B(new_n9557), .C(new_n9869), .Y(new_n9870));
  NAND2xp33_ASAP7_75t_L     g09614(.A(new_n9870), .B(new_n9868), .Y(new_n9871));
  OAI22xp33_ASAP7_75t_L     g09615(.A1(new_n1158), .A2(new_n5321), .B1(new_n5805), .B2(new_n1259), .Y(new_n9872));
  AOI221xp5_ASAP7_75t_L     g09616(.A1(\b[42] ), .A2(new_n1080), .B1(new_n1073), .B2(new_n5812), .C(new_n9872), .Y(new_n9873));
  XNOR2x2_ASAP7_75t_L       g09617(.A(new_n1071), .B(new_n9873), .Y(new_n9874));
  INVx1_ASAP7_75t_L         g09618(.A(new_n9874), .Y(new_n9875));
  AOI21xp33_ASAP7_75t_L     g09619(.A1(new_n9865), .A2(new_n9871), .B(new_n9875), .Y(new_n9876));
  NOR2xp33_ASAP7_75t_L      g09620(.A(new_n9870), .B(new_n9868), .Y(new_n9877));
  AOI21xp33_ASAP7_75t_L     g09621(.A1(new_n9559), .A2(new_n9869), .B(new_n9862), .Y(new_n9878));
  NOR3xp33_ASAP7_75t_L      g09622(.A(new_n9878), .B(new_n9874), .C(new_n9877), .Y(new_n9879));
  OA21x2_ASAP7_75t_L        g09623(.A1(new_n9876), .A2(new_n9879), .B(new_n9657), .Y(new_n9880));
  NOR3xp33_ASAP7_75t_L      g09624(.A(new_n9657), .B(new_n9876), .C(new_n9879), .Y(new_n9881));
  OA21x2_ASAP7_75t_L        g09625(.A1(new_n9881), .A2(new_n9880), .B(new_n9656), .Y(new_n9882));
  NOR3xp33_ASAP7_75t_L      g09626(.A(new_n9880), .B(new_n9656), .C(new_n9881), .Y(new_n9883));
  NOR3xp33_ASAP7_75t_L      g09627(.A(new_n9653), .B(new_n9882), .C(new_n9883), .Y(new_n9884));
  NOR2xp33_ASAP7_75t_L      g09628(.A(new_n9583), .B(new_n9581), .Y(new_n9885));
  MAJx2_ASAP7_75t_L         g09629(.A(new_n9585), .B(new_n9885), .C(new_n9576), .Y(new_n9886));
  OAI21xp33_ASAP7_75t_L     g09630(.A1(new_n9881), .A2(new_n9880), .B(new_n9656), .Y(new_n9887));
  INVx1_ASAP7_75t_L         g09631(.A(new_n9883), .Y(new_n9888));
  AOI21xp33_ASAP7_75t_L     g09632(.A1(new_n9888), .A2(new_n9887), .B(new_n9886), .Y(new_n9889));
  OAI21xp33_ASAP7_75t_L     g09633(.A1(new_n9884), .A2(new_n9889), .B(new_n9651), .Y(new_n9890));
  INVx1_ASAP7_75t_L         g09634(.A(new_n9651), .Y(new_n9891));
  NAND3xp33_ASAP7_75t_L     g09635(.A(new_n9888), .B(new_n9886), .C(new_n9887), .Y(new_n9892));
  OAI21xp33_ASAP7_75t_L     g09636(.A1(new_n9883), .A2(new_n9882), .B(new_n9653), .Y(new_n9893));
  NAND3xp33_ASAP7_75t_L     g09637(.A(new_n9892), .B(new_n9891), .C(new_n9893), .Y(new_n9894));
  NAND3xp33_ASAP7_75t_L     g09638(.A(new_n9648), .B(new_n9890), .C(new_n9894), .Y(new_n9895));
  AND2x2_ASAP7_75t_L        g09639(.A(new_n9588), .B(new_n9593), .Y(new_n9896));
  NOR2xp33_ASAP7_75t_L      g09640(.A(new_n9590), .B(new_n9647), .Y(new_n9897));
  INVx1_ASAP7_75t_L         g09641(.A(new_n9897), .Y(new_n9898));
  AOI21xp33_ASAP7_75t_L     g09642(.A1(new_n9892), .A2(new_n9893), .B(new_n9891), .Y(new_n9899));
  NOR3xp33_ASAP7_75t_L      g09643(.A(new_n9889), .B(new_n9884), .C(new_n9651), .Y(new_n9900));
  OAI221xp5_ASAP7_75t_L     g09644(.A1(new_n9900), .A2(new_n9899), .B1(new_n9896), .B2(new_n9596), .C(new_n9898), .Y(new_n9901));
  AOI21xp33_ASAP7_75t_L     g09645(.A1(new_n9901), .A2(new_n9895), .B(new_n9646), .Y(new_n9902));
  AND3x1_ASAP7_75t_L        g09646(.A(new_n9901), .B(new_n9895), .C(new_n9646), .Y(new_n9903));
  NOR3xp33_ASAP7_75t_L      g09647(.A(new_n9643), .B(new_n9902), .C(new_n9903), .Y(new_n9904));
  AO21x2_ASAP7_75t_L        g09648(.A1(new_n9895), .A2(new_n9901), .B(new_n9646), .Y(new_n9905));
  NAND3xp33_ASAP7_75t_L     g09649(.A(new_n9901), .B(new_n9895), .C(new_n9646), .Y(new_n9906));
  AOI221xp5_ASAP7_75t_L     g09650(.A1(new_n9607), .A2(new_n9348), .B1(new_n9905), .B2(new_n9906), .C(new_n9642), .Y(new_n9907));
  OAI21xp33_ASAP7_75t_L     g09651(.A1(new_n9907), .A2(new_n9904), .B(new_n9641), .Y(new_n9908));
  INVx1_ASAP7_75t_L         g09652(.A(new_n9641), .Y(new_n9909));
  NOR2xp33_ASAP7_75t_L      g09653(.A(new_n9902), .B(new_n9903), .Y(new_n9910));
  OAI21xp33_ASAP7_75t_L     g09654(.A1(new_n9604), .A2(new_n9642), .B(new_n9910), .Y(new_n9911));
  OAI21xp33_ASAP7_75t_L     g09655(.A1(new_n9902), .A2(new_n9903), .B(new_n9643), .Y(new_n9912));
  NAND3xp33_ASAP7_75t_L     g09656(.A(new_n9911), .B(new_n9909), .C(new_n9912), .Y(new_n9913));
  NAND3xp33_ASAP7_75t_L     g09657(.A(new_n9638), .B(new_n9908), .C(new_n9913), .Y(new_n9914));
  NOR2xp33_ASAP7_75t_L      g09658(.A(new_n9604), .B(new_n9608), .Y(new_n9915));
  MAJIxp5_ASAP7_75t_L       g09659(.A(new_n9340), .B(new_n9346), .C(new_n9915), .Y(new_n9916));
  NAND2xp33_ASAP7_75t_L     g09660(.A(new_n9908), .B(new_n9913), .Y(new_n9917));
  NAND2xp33_ASAP7_75t_L     g09661(.A(new_n9916), .B(new_n9917), .Y(new_n9918));
  NOR2xp33_ASAP7_75t_L      g09662(.A(\b[57] ), .B(\b[58] ), .Y(new_n9919));
  INVx1_ASAP7_75t_L         g09663(.A(\b[58] ), .Y(new_n9920));
  NOR2xp33_ASAP7_75t_L      g09664(.A(new_n9620), .B(new_n9920), .Y(new_n9921));
  NOR2xp33_ASAP7_75t_L      g09665(.A(new_n9919), .B(new_n9921), .Y(new_n9922));
  A2O1A1Ixp33_ASAP7_75t_L   g09666(.A1(\b[57] ), .A2(\b[56] ), .B(new_n9624), .C(new_n9922), .Y(new_n9923));
  OR3x1_ASAP7_75t_L         g09667(.A(new_n9624), .B(new_n9621), .C(new_n9922), .Y(new_n9924));
  NAND2xp33_ASAP7_75t_L     g09668(.A(new_n9923), .B(new_n9924), .Y(new_n9925));
  AOI22xp33_ASAP7_75t_L     g09669(.A1(\b[56] ), .A2(new_n282), .B1(\b[58] ), .B2(new_n303), .Y(new_n9926));
  OAI221xp5_ASAP7_75t_L     g09670(.A1(new_n291), .A2(new_n9620), .B1(new_n268), .B2(new_n9925), .C(new_n9926), .Y(new_n9927));
  INVx1_ASAP7_75t_L         g09671(.A(new_n9927), .Y(new_n9928));
  NAND2xp33_ASAP7_75t_L     g09672(.A(\a[2] ), .B(new_n9928), .Y(new_n9929));
  NAND2xp33_ASAP7_75t_L     g09673(.A(new_n262), .B(new_n9927), .Y(new_n9930));
  NAND2xp33_ASAP7_75t_L     g09674(.A(new_n9930), .B(new_n9929), .Y(new_n9931));
  INVx1_ASAP7_75t_L         g09675(.A(new_n9931), .Y(new_n9932));
  NAND3xp33_ASAP7_75t_L     g09676(.A(new_n9918), .B(new_n9914), .C(new_n9932), .Y(new_n9933));
  NOR2xp33_ASAP7_75t_L      g09677(.A(new_n9916), .B(new_n9917), .Y(new_n9934));
  AOI21xp33_ASAP7_75t_L     g09678(.A1(new_n9913), .A2(new_n9908), .B(new_n9638), .Y(new_n9935));
  OAI21xp33_ASAP7_75t_L     g09679(.A1(new_n9935), .A2(new_n9934), .B(new_n9931), .Y(new_n9936));
  NAND2xp33_ASAP7_75t_L     g09680(.A(new_n9933), .B(new_n9936), .Y(new_n9937));
  AO21x2_ASAP7_75t_L        g09681(.A1(new_n9633), .A2(new_n9339), .B(new_n9631), .Y(new_n9938));
  XOR2x2_ASAP7_75t_L        g09682(.A(new_n9938), .B(new_n9937), .Y(\f[58] ));
  NAND3xp33_ASAP7_75t_L     g09683(.A(new_n9918), .B(new_n9914), .C(new_n9931), .Y(new_n9940));
  INVx1_ASAP7_75t_L         g09684(.A(new_n9940), .Y(new_n9941));
  OAI21xp33_ASAP7_75t_L     g09685(.A1(new_n9916), .A2(new_n9917), .B(new_n9913), .Y(new_n9942));
  NAND2xp33_ASAP7_75t_L     g09686(.A(\b[58] ), .B(new_n272), .Y(new_n9943));
  INVx1_ASAP7_75t_L         g09687(.A(new_n9621), .Y(new_n9944));
  A2O1A1Ixp33_ASAP7_75t_L   g09688(.A1(new_n9328), .A2(new_n9618), .B(new_n9619), .C(new_n9944), .Y(new_n9945));
  NOR2xp33_ASAP7_75t_L      g09689(.A(\b[58] ), .B(\b[59] ), .Y(new_n9946));
  INVx1_ASAP7_75t_L         g09690(.A(\b[59] ), .Y(new_n9947));
  NOR2xp33_ASAP7_75t_L      g09691(.A(new_n9920), .B(new_n9947), .Y(new_n9948));
  NOR2xp33_ASAP7_75t_L      g09692(.A(new_n9946), .B(new_n9948), .Y(new_n9949));
  A2O1A1Ixp33_ASAP7_75t_L   g09693(.A1(new_n9945), .A2(new_n9922), .B(new_n9921), .C(new_n9949), .Y(new_n9950));
  O2A1O1Ixp33_ASAP7_75t_L   g09694(.A1(new_n9621), .A2(new_n9624), .B(new_n9922), .C(new_n9921), .Y(new_n9951));
  INVx1_ASAP7_75t_L         g09695(.A(new_n9949), .Y(new_n9952));
  NAND2xp33_ASAP7_75t_L     g09696(.A(new_n9952), .B(new_n9951), .Y(new_n9953));
  NAND3xp33_ASAP7_75t_L     g09697(.A(new_n9950), .B(new_n267), .C(new_n9953), .Y(new_n9954));
  AOI22xp33_ASAP7_75t_L     g09698(.A1(\b[57] ), .A2(new_n282), .B1(\b[59] ), .B2(new_n303), .Y(new_n9955));
  NAND4xp25_ASAP7_75t_L     g09699(.A(new_n9954), .B(\a[2] ), .C(new_n9943), .D(new_n9955), .Y(new_n9956));
  NAND2xp33_ASAP7_75t_L     g09700(.A(new_n9955), .B(new_n9954), .Y(new_n9957));
  A2O1A1Ixp33_ASAP7_75t_L   g09701(.A1(\b[58] ), .A2(new_n272), .B(new_n9957), .C(new_n262), .Y(new_n9958));
  NAND2xp33_ASAP7_75t_L     g09702(.A(new_n9956), .B(new_n9958), .Y(new_n9959));
  INVx1_ASAP7_75t_L         g09703(.A(new_n9959), .Y(new_n9960));
  A2O1A1O1Ixp25_ASAP7_75t_L g09704(.A1(new_n9348), .A2(new_n9607), .B(new_n9642), .C(new_n9905), .D(new_n9903), .Y(new_n9961));
  AOI22xp33_ASAP7_75t_L     g09705(.A1(new_n444), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n471), .Y(new_n9962));
  OAI21xp33_ASAP7_75t_L     g09706(.A1(new_n469), .A2(new_n8174), .B(new_n9962), .Y(new_n9963));
  AOI21xp33_ASAP7_75t_L     g09707(.A1(new_n447), .A2(\b[52] ), .B(new_n9963), .Y(new_n9964));
  NAND2xp33_ASAP7_75t_L     g09708(.A(\a[8] ), .B(new_n9964), .Y(new_n9965));
  A2O1A1Ixp33_ASAP7_75t_L   g09709(.A1(\b[52] ), .A2(new_n447), .B(new_n9963), .C(new_n435), .Y(new_n9966));
  AND2x2_ASAP7_75t_L        g09710(.A(new_n9966), .B(new_n9965), .Y(new_n9967));
  A2O1A1O1Ixp25_ASAP7_75t_L g09711(.A1(new_n9594), .A2(new_n9601), .B(new_n9897), .C(new_n9890), .D(new_n9900), .Y(new_n9968));
  AOI22xp33_ASAP7_75t_L     g09712(.A1(new_n811), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n900), .Y(new_n9969));
  OAI221xp5_ASAP7_75t_L     g09713(.A1(new_n904), .A2(new_n6568), .B1(new_n898), .B2(new_n6820), .C(new_n9969), .Y(new_n9970));
  XNOR2x2_ASAP7_75t_L       g09714(.A(new_n806), .B(new_n9970), .Y(new_n9971));
  INVx1_ASAP7_75t_L         g09715(.A(new_n9876), .Y(new_n9972));
  AOI22xp33_ASAP7_75t_L     g09716(.A1(new_n1076), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1253), .Y(new_n9973));
  OAI221xp5_ASAP7_75t_L     g09717(.A1(new_n1154), .A2(new_n5805), .B1(new_n1156), .B2(new_n5835), .C(new_n9973), .Y(new_n9974));
  XNOR2x2_ASAP7_75t_L       g09718(.A(\a[17] ), .B(new_n9974), .Y(new_n9975));
  INVx1_ASAP7_75t_L         g09719(.A(new_n9975), .Y(new_n9976));
  NAND3xp33_ASAP7_75t_L     g09720(.A(new_n9860), .B(new_n9857), .C(new_n9859), .Y(new_n9977));
  INVx1_ASAP7_75t_L         g09721(.A(new_n9977), .Y(new_n9978));
  OAI21xp33_ASAP7_75t_L     g09722(.A1(new_n9817), .A2(new_n9658), .B(new_n9820), .Y(new_n9979));
  NAND2xp33_ASAP7_75t_L     g09723(.A(\b[31] ), .B(new_n2553), .Y(new_n9980));
  NAND3xp33_ASAP7_75t_L     g09724(.A(new_n3210), .B(new_n2544), .C(new_n3213), .Y(new_n9981));
  AOI22xp33_ASAP7_75t_L     g09725(.A1(new_n2552), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n2736), .Y(new_n9982));
  AND4x1_ASAP7_75t_L        g09726(.A(new_n9982), .B(new_n9981), .C(new_n9980), .D(\a[29] ), .Y(new_n9983));
  AOI31xp33_ASAP7_75t_L     g09727(.A1(new_n9981), .A2(new_n9980), .A3(new_n9982), .B(\a[29] ), .Y(new_n9984));
  NOR2xp33_ASAP7_75t_L      g09728(.A(new_n9984), .B(new_n9983), .Y(new_n9985));
  NOR3xp33_ASAP7_75t_L      g09729(.A(new_n9791), .B(new_n9794), .C(new_n9790), .Y(new_n9986));
  INVx1_ASAP7_75t_L         g09730(.A(new_n9986), .Y(new_n9987));
  A2O1A1Ixp33_ASAP7_75t_L   g09731(.A1(new_n9806), .A2(new_n9807), .B(new_n9805), .C(new_n9987), .Y(new_n9988));
  NOR3xp33_ASAP7_75t_L      g09732(.A(new_n9774), .B(new_n9773), .C(new_n9664), .Y(new_n9989));
  A2O1A1O1Ixp25_ASAP7_75t_L g09733(.A1(new_n9489), .A2(new_n9385), .B(new_n9491), .C(new_n9775), .D(new_n9989), .Y(new_n9990));
  AOI22xp33_ASAP7_75t_L     g09734(.A1(new_n4283), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n4512), .Y(new_n9991));
  OAI221xp5_ASAP7_75t_L     g09735(.A1(new_n4277), .A2(new_n1774), .B1(new_n4499), .B2(new_n1915), .C(new_n9991), .Y(new_n9992));
  XNOR2x2_ASAP7_75t_L       g09736(.A(\a[38] ), .B(new_n9992), .Y(new_n9993));
  AOI22xp33_ASAP7_75t_L     g09737(.A1(new_n4920), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n5167), .Y(new_n9994));
  OAI221xp5_ASAP7_75t_L     g09738(.A1(new_n5154), .A2(new_n1432), .B1(new_n5158), .B2(new_n1547), .C(new_n9994), .Y(new_n9995));
  XNOR2x2_ASAP7_75t_L       g09739(.A(new_n4915), .B(new_n9995), .Y(new_n9996));
  NOR3xp33_ASAP7_75t_L      g09740(.A(new_n9753), .B(new_n9752), .C(new_n9671), .Y(new_n9997));
  NOR2xp33_ASAP7_75t_L      g09741(.A(new_n1030), .B(new_n5900), .Y(new_n9998));
  INVx1_ASAP7_75t_L         g09742(.A(new_n9998), .Y(new_n9999));
  NAND2xp33_ASAP7_75t_L     g09743(.A(new_n5621), .B(new_n3305), .Y(new_n10000));
  AOI22xp33_ASAP7_75t_L     g09744(.A1(new_n5624), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n5901), .Y(new_n10001));
  AND4x1_ASAP7_75t_L        g09745(.A(new_n10001), .B(new_n10000), .C(new_n9999), .D(\a[44] ), .Y(new_n10002));
  AOI31xp33_ASAP7_75t_L     g09746(.A1(new_n10000), .A2(new_n9999), .A3(new_n10001), .B(\a[44] ), .Y(new_n10003));
  INVx1_ASAP7_75t_L         g09747(.A(new_n9741), .Y(new_n10004));
  NAND2xp33_ASAP7_75t_L     g09748(.A(new_n9722), .B(new_n9728), .Y(new_n10005));
  MAJIxp5_ASAP7_75t_L       g09749(.A(new_n9735), .B(new_n9731), .C(new_n10005), .Y(new_n10006));
  AOI22xp33_ASAP7_75t_L     g09750(.A1(new_n7111), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n7391), .Y(new_n10007));
  OAI221xp5_ASAP7_75t_L     g09751(.A1(new_n8558), .A2(new_n617), .B1(new_n8237), .B2(new_n685), .C(new_n10007), .Y(new_n10008));
  XNOR2x2_ASAP7_75t_L       g09752(.A(\a[50] ), .B(new_n10008), .Y(new_n10009));
  A2O1A1O1Ixp25_ASAP7_75t_L g09753(.A1(new_n9450), .A2(new_n9441), .B(new_n9675), .C(new_n9717), .D(new_n9727), .Y(new_n10010));
  AOI22xp33_ASAP7_75t_L     g09754(.A1(new_n7960), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n8537), .Y(new_n10011));
  OAI221xp5_ASAP7_75t_L     g09755(.A1(new_n8817), .A2(new_n420), .B1(new_n7957), .B2(new_n494), .C(new_n10011), .Y(new_n10012));
  XNOR2x2_ASAP7_75t_L       g09756(.A(\a[53] ), .B(new_n10012), .Y(new_n10013));
  INVx1_ASAP7_75t_L         g09757(.A(new_n10013), .Y(new_n10014));
  A2O1A1O1Ixp25_ASAP7_75t_L g09758(.A1(new_n9680), .A2(new_n9413), .B(new_n9435), .C(new_n9714), .D(new_n9710), .Y(new_n10015));
  INVx1_ASAP7_75t_L         g09759(.A(new_n8828), .Y(new_n10016));
  NAND2xp33_ASAP7_75t_L     g09760(.A(\b[4] ), .B(new_n8835), .Y(new_n10017));
  AOI22xp33_ASAP7_75t_L     g09761(.A1(new_n8831), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n9115), .Y(new_n10018));
  OAI311xp33_ASAP7_75t_L    g09762(.A1(new_n357), .A2(new_n10016), .A3(new_n358), .B1(new_n10017), .C1(new_n10018), .Y(new_n10019));
  INVx1_ASAP7_75t_L         g09763(.A(new_n10019), .Y(new_n10020));
  NAND2xp33_ASAP7_75t_L     g09764(.A(\a[56] ), .B(new_n10020), .Y(new_n10021));
  NAND2xp33_ASAP7_75t_L     g09765(.A(new_n8826), .B(new_n10019), .Y(new_n10022));
  NAND2xp33_ASAP7_75t_L     g09766(.A(new_n10022), .B(new_n10021), .Y(new_n10023));
  INVx1_ASAP7_75t_L         g09767(.A(new_n9703), .Y(new_n10024));
  NOR2xp33_ASAP7_75t_L      g09768(.A(new_n280), .B(new_n9696), .Y(new_n10025));
  NAND3xp33_ASAP7_75t_L     g09769(.A(new_n9412), .B(new_n9695), .C(new_n9702), .Y(new_n10026));
  INVx1_ASAP7_75t_L         g09770(.A(new_n10026), .Y(new_n10027));
  AOI221xp5_ASAP7_75t_L     g09771(.A1(\b[2] ), .A2(new_n9700), .B1(\b[0] ), .B2(new_n10027), .C(new_n10025), .Y(new_n10028));
  OAI21xp33_ASAP7_75t_L     g09772(.A1(new_n261), .A2(new_n10024), .B(new_n10028), .Y(new_n10029));
  O2A1O1Ixp33_ASAP7_75t_L   g09773(.A1(new_n9413), .A2(new_n9705), .B(\a[59] ), .C(new_n10029), .Y(new_n10030));
  A2O1A1Ixp33_ASAP7_75t_L   g09774(.A1(\b[0] ), .A2(new_n9690), .B(new_n9705), .C(\a[59] ), .Y(new_n10031));
  O2A1O1Ixp33_ASAP7_75t_L   g09775(.A1(new_n10024), .A2(new_n261), .B(new_n10028), .C(new_n10031), .Y(new_n10032));
  NOR2xp33_ASAP7_75t_L      g09776(.A(new_n10030), .B(new_n10032), .Y(new_n10033));
  NOR2xp33_ASAP7_75t_L      g09777(.A(new_n10023), .B(new_n10033), .Y(new_n10034));
  OA21x2_ASAP7_75t_L        g09778(.A1(new_n261), .A2(new_n10024), .B(new_n10028), .Y(new_n10035));
  XNOR2x2_ASAP7_75t_L       g09779(.A(new_n10035), .B(new_n10031), .Y(new_n10036));
  AOI21xp33_ASAP7_75t_L     g09780(.A1(new_n10022), .A2(new_n10021), .B(new_n10036), .Y(new_n10037));
  OAI21xp33_ASAP7_75t_L     g09781(.A1(new_n10037), .A2(new_n10034), .B(new_n10015), .Y(new_n10038));
  A2O1A1Ixp33_ASAP7_75t_L   g09782(.A1(new_n9424), .A2(new_n9712), .B(new_n9707), .C(new_n9715), .Y(new_n10039));
  NAND3xp33_ASAP7_75t_L     g09783(.A(new_n10036), .B(new_n10022), .C(new_n10021), .Y(new_n10040));
  NAND2xp33_ASAP7_75t_L     g09784(.A(new_n10023), .B(new_n10033), .Y(new_n10041));
  NAND3xp33_ASAP7_75t_L     g09785(.A(new_n10039), .B(new_n10040), .C(new_n10041), .Y(new_n10042));
  AOI21xp33_ASAP7_75t_L     g09786(.A1(new_n10042), .A2(new_n10038), .B(new_n10014), .Y(new_n10043));
  AOI21xp33_ASAP7_75t_L     g09787(.A1(new_n10041), .A2(new_n10040), .B(new_n10039), .Y(new_n10044));
  NOR3xp33_ASAP7_75t_L      g09788(.A(new_n10015), .B(new_n10034), .C(new_n10037), .Y(new_n10045));
  NOR3xp33_ASAP7_75t_L      g09789(.A(new_n10045), .B(new_n10044), .C(new_n10013), .Y(new_n10046));
  NOR3xp33_ASAP7_75t_L      g09790(.A(new_n10010), .B(new_n10043), .C(new_n10046), .Y(new_n10047));
  INVx1_ASAP7_75t_L         g09791(.A(new_n9675), .Y(new_n10048));
  OAI211xp5_ASAP7_75t_L     g09792(.A1(new_n9723), .A2(new_n9724), .B(new_n9439), .C(new_n9128), .Y(new_n10049));
  A2O1A1Ixp33_ASAP7_75t_L   g09793(.A1(new_n10049), .A2(new_n10048), .B(new_n9726), .C(new_n9721), .Y(new_n10050));
  OAI21xp33_ASAP7_75t_L     g09794(.A1(new_n10044), .A2(new_n10045), .B(new_n10013), .Y(new_n10051));
  NAND3xp33_ASAP7_75t_L     g09795(.A(new_n10014), .B(new_n10038), .C(new_n10042), .Y(new_n10052));
  AOI21xp33_ASAP7_75t_L     g09796(.A1(new_n10052), .A2(new_n10051), .B(new_n10050), .Y(new_n10053));
  OAI21xp33_ASAP7_75t_L     g09797(.A1(new_n10047), .A2(new_n10053), .B(new_n10009), .Y(new_n10054));
  XNOR2x2_ASAP7_75t_L       g09798(.A(new_n7106), .B(new_n10008), .Y(new_n10055));
  NAND3xp33_ASAP7_75t_L     g09799(.A(new_n10050), .B(new_n10051), .C(new_n10052), .Y(new_n10056));
  OAI21xp33_ASAP7_75t_L     g09800(.A1(new_n10043), .A2(new_n10046), .B(new_n10010), .Y(new_n10057));
  NAND3xp33_ASAP7_75t_L     g09801(.A(new_n10056), .B(new_n10055), .C(new_n10057), .Y(new_n10058));
  NAND3xp33_ASAP7_75t_L     g09802(.A(new_n10006), .B(new_n10054), .C(new_n10058), .Y(new_n10059));
  NAND2xp33_ASAP7_75t_L     g09803(.A(new_n10058), .B(new_n10054), .Y(new_n10060));
  OAI211xp5_ASAP7_75t_L     g09804(.A1(new_n10005), .A2(new_n9731), .B(new_n10060), .C(new_n9743), .Y(new_n10061));
  AOI22xp33_ASAP7_75t_L     g09805(.A1(new_n6376), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n6648), .Y(new_n10062));
  OAI221xp5_ASAP7_75t_L     g09806(.A1(new_n6646), .A2(new_n784), .B1(new_n6636), .B2(new_n875), .C(new_n10062), .Y(new_n10063));
  XNOR2x2_ASAP7_75t_L       g09807(.A(\a[47] ), .B(new_n10063), .Y(new_n10064));
  NAND3xp33_ASAP7_75t_L     g09808(.A(new_n10061), .B(new_n10059), .C(new_n10064), .Y(new_n10065));
  O2A1O1Ixp33_ASAP7_75t_L   g09809(.A1(new_n10005), .A2(new_n9731), .B(new_n9743), .C(new_n10060), .Y(new_n10066));
  AOI21xp33_ASAP7_75t_L     g09810(.A1(new_n10058), .A2(new_n10054), .B(new_n10006), .Y(new_n10067));
  INVx1_ASAP7_75t_L         g09811(.A(new_n10064), .Y(new_n10068));
  OAI21xp33_ASAP7_75t_L     g09812(.A1(new_n10067), .A2(new_n10066), .B(new_n10068), .Y(new_n10069));
  AOI221xp5_ASAP7_75t_L     g09813(.A1(new_n9674), .A2(new_n9745), .B1(new_n10065), .B2(new_n10069), .C(new_n10004), .Y(new_n10070));
  NOR3xp33_ASAP7_75t_L      g09814(.A(new_n10066), .B(new_n10068), .C(new_n10067), .Y(new_n10071));
  AOI21xp33_ASAP7_75t_L     g09815(.A1(new_n10061), .A2(new_n10059), .B(new_n10064), .Y(new_n10072));
  OAI211xp5_ASAP7_75t_L     g09816(.A1(new_n9401), .A2(new_n9459), .B(new_n9745), .C(new_n9748), .Y(new_n10073));
  AOI211xp5_ASAP7_75t_L     g09817(.A1(new_n10073), .A2(new_n9741), .B(new_n10071), .C(new_n10072), .Y(new_n10074));
  OAI22xp33_ASAP7_75t_L     g09818(.A1(new_n10070), .A2(new_n10074), .B1(new_n10002), .B2(new_n10003), .Y(new_n10075));
  NOR2xp33_ASAP7_75t_L      g09819(.A(new_n10003), .B(new_n10002), .Y(new_n10076));
  OAI211xp5_ASAP7_75t_L     g09820(.A1(new_n10071), .A2(new_n10072), .B(new_n9741), .C(new_n10073), .Y(new_n10077));
  AO211x2_ASAP7_75t_L       g09821(.A1(new_n10073), .A2(new_n9741), .B(new_n10071), .C(new_n10072), .Y(new_n10078));
  NAND3xp33_ASAP7_75t_L     g09822(.A(new_n10078), .B(new_n10076), .C(new_n10077), .Y(new_n10079));
  NAND2xp33_ASAP7_75t_L     g09823(.A(new_n10075), .B(new_n10079), .Y(new_n10080));
  A2O1A1Ixp33_ASAP7_75t_L   g09824(.A1(new_n9764), .A2(new_n9763), .B(new_n9997), .C(new_n10080), .Y(new_n10081));
  A2O1A1O1Ixp25_ASAP7_75t_L g09825(.A1(new_n9468), .A2(new_n9471), .B(new_n9668), .C(new_n9754), .D(new_n9997), .Y(new_n10082));
  NAND3xp33_ASAP7_75t_L     g09826(.A(new_n10082), .B(new_n10075), .C(new_n10079), .Y(new_n10083));
  NAND3xp33_ASAP7_75t_L     g09827(.A(new_n10081), .B(new_n9996), .C(new_n10083), .Y(new_n10084));
  AO21x2_ASAP7_75t_L        g09828(.A1(new_n10083), .A2(new_n10081), .B(new_n9996), .Y(new_n10085));
  OAI211xp5_ASAP7_75t_L     g09829(.A1(new_n9480), .A2(new_n9483), .B(new_n9667), .C(new_n9767), .Y(new_n10086));
  AND4x1_ASAP7_75t_L        g09830(.A(new_n10086), .B(new_n10085), .C(new_n10084), .D(new_n9761), .Y(new_n10087));
  AOI22xp33_ASAP7_75t_L     g09831(.A1(new_n10085), .A2(new_n10084), .B1(new_n9761), .B2(new_n10086), .Y(new_n10088));
  NOR3xp33_ASAP7_75t_L      g09832(.A(new_n10087), .B(new_n10088), .C(new_n9993), .Y(new_n10089));
  INVx1_ASAP7_75t_L         g09833(.A(new_n9993), .Y(new_n10090));
  NAND4xp25_ASAP7_75t_L     g09834(.A(new_n10086), .B(new_n9761), .C(new_n10084), .D(new_n10085), .Y(new_n10091));
  A2O1A1O1Ixp25_ASAP7_75t_L g09835(.A1(new_n9164), .A2(new_n9166), .B(new_n9390), .C(new_n9478), .D(new_n9666), .Y(new_n10092));
  INVx1_ASAP7_75t_L         g09836(.A(new_n9761), .Y(new_n10093));
  NAND2xp33_ASAP7_75t_L     g09837(.A(new_n10084), .B(new_n10085), .Y(new_n10094));
  A2O1A1Ixp33_ASAP7_75t_L   g09838(.A1(new_n9767), .A2(new_n10092), .B(new_n10093), .C(new_n10094), .Y(new_n10095));
  AOI21xp33_ASAP7_75t_L     g09839(.A1(new_n10095), .A2(new_n10091), .B(new_n10090), .Y(new_n10096));
  OAI21xp33_ASAP7_75t_L     g09840(.A1(new_n10089), .A2(new_n10096), .B(new_n9990), .Y(new_n10097));
  NOR2xp33_ASAP7_75t_L      g09841(.A(new_n10089), .B(new_n10096), .Y(new_n10098));
  A2O1A1Ixp33_ASAP7_75t_L   g09842(.A1(new_n9775), .A2(new_n9661), .B(new_n9989), .C(new_n10098), .Y(new_n10099));
  AOI22xp33_ASAP7_75t_L     g09843(.A1(new_n3633), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n3858), .Y(new_n10100));
  OAI221xp5_ASAP7_75t_L     g09844(.A1(new_n3853), .A2(new_n2067), .B1(new_n3856), .B2(new_n2355), .C(new_n10100), .Y(new_n10101));
  XNOR2x2_ASAP7_75t_L       g09845(.A(\a[35] ), .B(new_n10101), .Y(new_n10102));
  NAND3xp33_ASAP7_75t_L     g09846(.A(new_n10099), .B(new_n10097), .C(new_n10102), .Y(new_n10103));
  NAND3xp33_ASAP7_75t_L     g09847(.A(new_n10095), .B(new_n10091), .C(new_n10090), .Y(new_n10104));
  OAI21xp33_ASAP7_75t_L     g09848(.A1(new_n10088), .A2(new_n10087), .B(new_n9993), .Y(new_n10105));
  AOI221xp5_ASAP7_75t_L     g09849(.A1(new_n9661), .A2(new_n9775), .B1(new_n10104), .B2(new_n10105), .C(new_n9989), .Y(new_n10106));
  NAND2xp33_ASAP7_75t_L     g09850(.A(new_n10105), .B(new_n10104), .Y(new_n10107));
  O2A1O1Ixp33_ASAP7_75t_L   g09851(.A1(new_n9777), .A2(new_n9778), .B(new_n9772), .C(new_n10107), .Y(new_n10108));
  INVx1_ASAP7_75t_L         g09852(.A(new_n10102), .Y(new_n10109));
  OAI21xp33_ASAP7_75t_L     g09853(.A1(new_n10106), .A2(new_n10108), .B(new_n10109), .Y(new_n10110));
  NOR3xp33_ASAP7_75t_L      g09854(.A(new_n9779), .B(new_n9786), .C(new_n9776), .Y(new_n10111));
  INVx1_ASAP7_75t_L         g09855(.A(new_n10111), .Y(new_n10112));
  AND4x1_ASAP7_75t_L        g09856(.A(new_n9801), .B(new_n10112), .C(new_n10103), .D(new_n10110), .Y(new_n10113));
  O2A1O1Ixp33_ASAP7_75t_L   g09857(.A1(new_n9787), .A2(new_n9783), .B(new_n9789), .C(new_n10111), .Y(new_n10114));
  AOI21xp33_ASAP7_75t_L     g09858(.A1(new_n10110), .A2(new_n10103), .B(new_n10114), .Y(new_n10115));
  AOI22xp33_ASAP7_75t_L     g09859(.A1(new_n3029), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n3258), .Y(new_n10116));
  OAI221xp5_ASAP7_75t_L     g09860(.A1(new_n3024), .A2(new_n2666), .B1(new_n3256), .B2(new_n2695), .C(new_n10116), .Y(new_n10117));
  XNOR2x2_ASAP7_75t_L       g09861(.A(\a[32] ), .B(new_n10117), .Y(new_n10118));
  OAI21xp33_ASAP7_75t_L     g09862(.A1(new_n10115), .A2(new_n10113), .B(new_n10118), .Y(new_n10119));
  NAND3xp33_ASAP7_75t_L     g09863(.A(new_n10114), .B(new_n10110), .C(new_n10103), .Y(new_n10120));
  AO22x1_ASAP7_75t_L        g09864(.A1(new_n10103), .A2(new_n10110), .B1(new_n10112), .B2(new_n9801), .Y(new_n10121));
  INVx1_ASAP7_75t_L         g09865(.A(new_n10118), .Y(new_n10122));
  NAND3xp33_ASAP7_75t_L     g09866(.A(new_n10121), .B(new_n10120), .C(new_n10122), .Y(new_n10123));
  AOI21xp33_ASAP7_75t_L     g09867(.A1(new_n10123), .A2(new_n10119), .B(new_n9988), .Y(new_n10124));
  O2A1O1Ixp33_ASAP7_75t_L   g09868(.A1(new_n9796), .A2(new_n9802), .B(new_n9660), .C(new_n9986), .Y(new_n10125));
  NAND2xp33_ASAP7_75t_L     g09869(.A(new_n10119), .B(new_n10123), .Y(new_n10126));
  NOR2xp33_ASAP7_75t_L      g09870(.A(new_n10126), .B(new_n10125), .Y(new_n10127));
  OAI21xp33_ASAP7_75t_L     g09871(.A1(new_n10124), .A2(new_n10127), .B(new_n9985), .Y(new_n10128));
  INVx1_ASAP7_75t_L         g09872(.A(new_n9985), .Y(new_n10129));
  NAND2xp33_ASAP7_75t_L     g09873(.A(new_n10126), .B(new_n10125), .Y(new_n10130));
  NAND3xp33_ASAP7_75t_L     g09874(.A(new_n9988), .B(new_n10119), .C(new_n10123), .Y(new_n10131));
  NAND3xp33_ASAP7_75t_L     g09875(.A(new_n10130), .B(new_n10131), .C(new_n10129), .Y(new_n10132));
  NAND3xp33_ASAP7_75t_L     g09876(.A(new_n9979), .B(new_n10128), .C(new_n10132), .Y(new_n10133));
  AOI21xp33_ASAP7_75t_L     g09877(.A1(new_n10130), .A2(new_n10131), .B(new_n10129), .Y(new_n10134));
  NOR3xp33_ASAP7_75t_L      g09878(.A(new_n10127), .B(new_n9985), .C(new_n10124), .Y(new_n10135));
  OAI221xp5_ASAP7_75t_L     g09879(.A1(new_n9817), .A2(new_n9658), .B1(new_n10134), .B2(new_n10135), .C(new_n9820), .Y(new_n10136));
  INVx1_ASAP7_75t_L         g09880(.A(new_n3811), .Y(new_n10137));
  AOI22xp33_ASAP7_75t_L     g09881(.A1(new_n2114), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n2259), .Y(new_n10138));
  OAI221xp5_ASAP7_75t_L     g09882(.A1(new_n2109), .A2(new_n3584), .B1(new_n2257), .B2(new_n10137), .C(new_n10138), .Y(new_n10139));
  XNOR2x2_ASAP7_75t_L       g09883(.A(\a[26] ), .B(new_n10139), .Y(new_n10140));
  NAND3xp33_ASAP7_75t_L     g09884(.A(new_n10133), .B(new_n10136), .C(new_n10140), .Y(new_n10141));
  AO21x2_ASAP7_75t_L        g09885(.A1(new_n10136), .A2(new_n10133), .B(new_n10140), .Y(new_n10142));
  NAND2xp33_ASAP7_75t_L     g09886(.A(new_n10141), .B(new_n10142), .Y(new_n10143));
  NOR3xp33_ASAP7_75t_L      g09887(.A(new_n9827), .B(new_n9828), .C(new_n9825), .Y(new_n10144));
  AO21x2_ASAP7_75t_L        g09888(.A1(new_n9836), .A2(new_n9835), .B(new_n10144), .Y(new_n10145));
  NOR2xp33_ASAP7_75t_L      g09889(.A(new_n10143), .B(new_n10145), .Y(new_n10146));
  AND2x2_ASAP7_75t_L        g09890(.A(new_n10141), .B(new_n10142), .Y(new_n10147));
  O2A1O1Ixp33_ASAP7_75t_L   g09891(.A1(new_n9832), .A2(new_n9541), .B(new_n9835), .C(new_n10144), .Y(new_n10148));
  NOR2xp33_ASAP7_75t_L      g09892(.A(new_n10148), .B(new_n10147), .Y(new_n10149));
  AOI22xp33_ASAP7_75t_L     g09893(.A1(new_n1704), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1837), .Y(new_n10150));
  OAI221xp5_ASAP7_75t_L     g09894(.A1(new_n1699), .A2(new_n4424), .B1(new_n1827), .B2(new_n4641), .C(new_n10150), .Y(new_n10151));
  XNOR2x2_ASAP7_75t_L       g09895(.A(new_n1689), .B(new_n10151), .Y(new_n10152));
  NOR3xp33_ASAP7_75t_L      g09896(.A(new_n10146), .B(new_n10149), .C(new_n10152), .Y(new_n10153));
  OA21x2_ASAP7_75t_L        g09897(.A1(new_n10149), .A2(new_n10146), .B(new_n10152), .Y(new_n10154));
  XNOR2x2_ASAP7_75t_L       g09898(.A(new_n9836), .B(new_n9835), .Y(new_n10155));
  MAJIxp5_ASAP7_75t_L       g09899(.A(new_n9847), .B(new_n9840), .C(new_n10155), .Y(new_n10156));
  NOR3xp33_ASAP7_75t_L      g09900(.A(new_n10156), .B(new_n10154), .C(new_n10153), .Y(new_n10157));
  OA21x2_ASAP7_75t_L        g09901(.A1(new_n10153), .A2(new_n10154), .B(new_n10156), .Y(new_n10158));
  AOI22xp33_ASAP7_75t_L     g09902(.A1(new_n1360), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1581), .Y(new_n10159));
  OAI221xp5_ASAP7_75t_L     g09903(.A1(new_n1373), .A2(new_n4869), .B1(new_n1359), .B2(new_n5327), .C(new_n10159), .Y(new_n10160));
  XNOR2x2_ASAP7_75t_L       g09904(.A(\a[20] ), .B(new_n10160), .Y(new_n10161));
  OAI21xp33_ASAP7_75t_L     g09905(.A1(new_n10157), .A2(new_n10158), .B(new_n10161), .Y(new_n10162));
  OR3x1_ASAP7_75t_L         g09906(.A(new_n10146), .B(new_n10149), .C(new_n10152), .Y(new_n10163));
  OAI21xp33_ASAP7_75t_L     g09907(.A1(new_n10149), .A2(new_n10146), .B(new_n10152), .Y(new_n10164));
  NAND3xp33_ASAP7_75t_L     g09908(.A(new_n9834), .B(new_n9837), .C(new_n9844), .Y(new_n10165));
  NAND4xp25_ASAP7_75t_L     g09909(.A(new_n9860), .B(new_n10163), .C(new_n10165), .D(new_n10164), .Y(new_n10166));
  OAI21xp33_ASAP7_75t_L     g09910(.A1(new_n10153), .A2(new_n10154), .B(new_n10156), .Y(new_n10167));
  INVx1_ASAP7_75t_L         g09911(.A(new_n10161), .Y(new_n10168));
  NAND3xp33_ASAP7_75t_L     g09912(.A(new_n10166), .B(new_n10167), .C(new_n10168), .Y(new_n10169));
  AOI221xp5_ASAP7_75t_L     g09913(.A1(new_n9868), .A2(new_n9870), .B1(new_n10169), .B2(new_n10162), .C(new_n9978), .Y(new_n10170));
  INVx1_ASAP7_75t_L         g09914(.A(new_n10170), .Y(new_n10171));
  AOI21xp33_ASAP7_75t_L     g09915(.A1(new_n10166), .A2(new_n10167), .B(new_n10168), .Y(new_n10172));
  NOR3xp33_ASAP7_75t_L      g09916(.A(new_n10158), .B(new_n10161), .C(new_n10157), .Y(new_n10173));
  NOR2xp33_ASAP7_75t_L      g09917(.A(new_n10172), .B(new_n10173), .Y(new_n10174));
  A2O1A1Ixp33_ASAP7_75t_L   g09918(.A1(new_n9870), .A2(new_n9868), .B(new_n9978), .C(new_n10174), .Y(new_n10175));
  NAND3xp33_ASAP7_75t_L     g09919(.A(new_n10171), .B(new_n10175), .C(new_n9976), .Y(new_n10176));
  NAND2xp33_ASAP7_75t_L     g09920(.A(new_n10169), .B(new_n10162), .Y(new_n10177));
  O2A1O1Ixp33_ASAP7_75t_L   g09921(.A1(new_n9862), .A2(new_n9864), .B(new_n9977), .C(new_n10177), .Y(new_n10178));
  OAI21xp33_ASAP7_75t_L     g09922(.A1(new_n10170), .A2(new_n10178), .B(new_n9975), .Y(new_n10179));
  NAND3xp33_ASAP7_75t_L     g09923(.A(new_n9865), .B(new_n9871), .C(new_n9875), .Y(new_n10180));
  OAI211xp5_ASAP7_75t_L     g09924(.A1(new_n9580), .A2(new_n9577), .B(new_n9579), .C(new_n10180), .Y(new_n10181));
  NAND4xp25_ASAP7_75t_L     g09925(.A(new_n10181), .B(new_n10176), .C(new_n10179), .D(new_n9972), .Y(new_n10182));
  NOR3xp33_ASAP7_75t_L      g09926(.A(new_n10178), .B(new_n10170), .C(new_n9975), .Y(new_n10183));
  AOI21xp33_ASAP7_75t_L     g09927(.A1(new_n10171), .A2(new_n10175), .B(new_n9976), .Y(new_n10184));
  AOI211xp5_ASAP7_75t_L     g09928(.A1(new_n9369), .A2(new_n9578), .B(new_n9571), .C(new_n9879), .Y(new_n10185));
  OAI22xp33_ASAP7_75t_L     g09929(.A1(new_n10185), .A2(new_n9876), .B1(new_n10183), .B2(new_n10184), .Y(new_n10186));
  AND3x1_ASAP7_75t_L        g09930(.A(new_n10186), .B(new_n10182), .C(new_n9971), .Y(new_n10187));
  AOI21xp33_ASAP7_75t_L     g09931(.A1(new_n10186), .A2(new_n10182), .B(new_n9971), .Y(new_n10188));
  NOR2xp33_ASAP7_75t_L      g09932(.A(new_n10188), .B(new_n10187), .Y(new_n10189));
  A2O1A1Ixp33_ASAP7_75t_L   g09933(.A1(new_n9887), .A2(new_n9886), .B(new_n9883), .C(new_n10189), .Y(new_n10190));
  OAI21xp33_ASAP7_75t_L     g09934(.A1(new_n9583), .A2(new_n9581), .B(new_n9576), .Y(new_n10191));
  NAND3xp33_ASAP7_75t_L     g09935(.A(new_n9573), .B(new_n9366), .C(new_n9574), .Y(new_n10192));
  NAND2xp33_ASAP7_75t_L     g09936(.A(new_n10192), .B(new_n10191), .Y(new_n10193));
  A2O1A1O1Ixp25_ASAP7_75t_L g09937(.A1(new_n9585), .A2(new_n10193), .B(new_n9652), .C(new_n9887), .D(new_n9883), .Y(new_n10194));
  OAI21xp33_ASAP7_75t_L     g09938(.A1(new_n10187), .A2(new_n10188), .B(new_n10194), .Y(new_n10195));
  NOR2xp33_ASAP7_75t_L      g09939(.A(new_n7317), .B(new_n821), .Y(new_n10196));
  INVx1_ASAP7_75t_L         g09940(.A(new_n10196), .Y(new_n10197));
  NAND2xp33_ASAP7_75t_L     g09941(.A(new_n578), .B(new_n7601), .Y(new_n10198));
  AOI22xp33_ASAP7_75t_L     g09942(.A1(\b[48] ), .A2(new_n651), .B1(\b[50] ), .B2(new_n581), .Y(new_n10199));
  NAND3xp33_ASAP7_75t_L     g09943(.A(new_n10198), .B(new_n10197), .C(new_n10199), .Y(new_n10200));
  XNOR2x2_ASAP7_75t_L       g09944(.A(\a[11] ), .B(new_n10200), .Y(new_n10201));
  NAND3xp33_ASAP7_75t_L     g09945(.A(new_n10190), .B(new_n10195), .C(new_n10201), .Y(new_n10202));
  AO21x2_ASAP7_75t_L        g09946(.A1(new_n10195), .A2(new_n10190), .B(new_n10201), .Y(new_n10203));
  AO21x2_ASAP7_75t_L        g09947(.A1(new_n10203), .A2(new_n10202), .B(new_n9968), .Y(new_n10204));
  NAND3xp33_ASAP7_75t_L     g09948(.A(new_n9968), .B(new_n10203), .C(new_n10202), .Y(new_n10205));
  AOI21xp33_ASAP7_75t_L     g09949(.A1(new_n10204), .A2(new_n10205), .B(new_n9967), .Y(new_n10206));
  NAND2xp33_ASAP7_75t_L     g09950(.A(new_n9966), .B(new_n9965), .Y(new_n10207));
  AOI21xp33_ASAP7_75t_L     g09951(.A1(new_n10203), .A2(new_n10202), .B(new_n9968), .Y(new_n10208));
  AND3x1_ASAP7_75t_L        g09952(.A(new_n9968), .B(new_n10203), .C(new_n10202), .Y(new_n10209));
  NOR3xp33_ASAP7_75t_L      g09953(.A(new_n10209), .B(new_n10208), .C(new_n10207), .Y(new_n10210));
  NOR3xp33_ASAP7_75t_L      g09954(.A(new_n9961), .B(new_n10206), .C(new_n10210), .Y(new_n10211));
  OAI21xp33_ASAP7_75t_L     g09955(.A1(new_n9902), .A2(new_n9643), .B(new_n9906), .Y(new_n10212));
  OAI21xp33_ASAP7_75t_L     g09956(.A1(new_n10208), .A2(new_n10209), .B(new_n10207), .Y(new_n10213));
  NAND3xp33_ASAP7_75t_L     g09957(.A(new_n10204), .B(new_n9967), .C(new_n10205), .Y(new_n10214));
  AOI21xp33_ASAP7_75t_L     g09958(.A1(new_n10214), .A2(new_n10213), .B(new_n10212), .Y(new_n10215));
  OAI22xp33_ASAP7_75t_L     g09959(.A1(new_n407), .A2(new_n8458), .B1(new_n9323), .B2(new_n343), .Y(new_n10216));
  AOI221xp5_ASAP7_75t_L     g09960(.A1(\b[55] ), .A2(new_n347), .B1(new_n341), .B2(new_n9332), .C(new_n10216), .Y(new_n10217));
  XNOR2x2_ASAP7_75t_L       g09961(.A(new_n338), .B(new_n10217), .Y(new_n10218));
  INVx1_ASAP7_75t_L         g09962(.A(new_n10218), .Y(new_n10219));
  OAI21xp33_ASAP7_75t_L     g09963(.A1(new_n10211), .A2(new_n10215), .B(new_n10219), .Y(new_n10220));
  NOR2xp33_ASAP7_75t_L      g09964(.A(new_n10206), .B(new_n10210), .Y(new_n10221));
  NAND2xp33_ASAP7_75t_L     g09965(.A(new_n10212), .B(new_n10221), .Y(new_n10222));
  OAI21xp33_ASAP7_75t_L     g09966(.A1(new_n10206), .A2(new_n10210), .B(new_n9961), .Y(new_n10223));
  NAND3xp33_ASAP7_75t_L     g09967(.A(new_n10222), .B(new_n10223), .C(new_n10218), .Y(new_n10224));
  NAND3xp33_ASAP7_75t_L     g09968(.A(new_n10224), .B(new_n10220), .C(new_n9960), .Y(new_n10225));
  AOI21xp33_ASAP7_75t_L     g09969(.A1(new_n10222), .A2(new_n10223), .B(new_n10218), .Y(new_n10226));
  NOR3xp33_ASAP7_75t_L      g09970(.A(new_n10215), .B(new_n10211), .C(new_n10219), .Y(new_n10227));
  OAI21xp33_ASAP7_75t_L     g09971(.A1(new_n10227), .A2(new_n10226), .B(new_n9959), .Y(new_n10228));
  NAND3xp33_ASAP7_75t_L     g09972(.A(new_n10228), .B(new_n10225), .C(new_n9942), .Y(new_n10229));
  NOR2xp33_ASAP7_75t_L      g09973(.A(new_n9907), .B(new_n9904), .Y(new_n10230));
  MAJIxp5_ASAP7_75t_L       g09974(.A(new_n9638), .B(new_n9909), .C(new_n10230), .Y(new_n10231));
  NOR3xp33_ASAP7_75t_L      g09975(.A(new_n10226), .B(new_n10227), .C(new_n9959), .Y(new_n10232));
  AOI21xp33_ASAP7_75t_L     g09976(.A1(new_n10224), .A2(new_n10220), .B(new_n9960), .Y(new_n10233));
  OAI21xp33_ASAP7_75t_L     g09977(.A1(new_n10233), .A2(new_n10232), .B(new_n10231), .Y(new_n10234));
  NAND2xp33_ASAP7_75t_L     g09978(.A(new_n10229), .B(new_n10234), .Y(new_n10235));
  A2O1A1Ixp33_ASAP7_75t_L   g09979(.A1(new_n9937), .A2(new_n9938), .B(new_n9941), .C(new_n10235), .Y(new_n10236));
  NOR3xp33_ASAP7_75t_L      g09980(.A(new_n9934), .B(new_n9935), .C(new_n9931), .Y(new_n10237));
  AOI21xp33_ASAP7_75t_L     g09981(.A1(new_n9918), .A2(new_n9914), .B(new_n9932), .Y(new_n10238));
  O2A1O1Ixp33_ASAP7_75t_L   g09982(.A1(new_n10237), .A2(new_n10238), .B(new_n9938), .C(new_n9941), .Y(new_n10239));
  NOR3xp33_ASAP7_75t_L      g09983(.A(new_n10232), .B(new_n10233), .C(new_n10231), .Y(new_n10240));
  AOI21xp33_ASAP7_75t_L     g09984(.A1(new_n10228), .A2(new_n10225), .B(new_n9942), .Y(new_n10241));
  NOR2xp33_ASAP7_75t_L      g09985(.A(new_n10241), .B(new_n10240), .Y(new_n10242));
  NAND2xp33_ASAP7_75t_L     g09986(.A(new_n10242), .B(new_n10239), .Y(new_n10243));
  AND2x2_ASAP7_75t_L        g09987(.A(new_n10236), .B(new_n10243), .Y(\f[59] ));
  NAND2xp33_ASAP7_75t_L     g09988(.A(new_n10225), .B(new_n10228), .Y(new_n10245));
  A2O1A1Ixp33_ASAP7_75t_L   g09989(.A1(new_n10230), .A2(new_n9909), .B(new_n9934), .C(new_n10245), .Y(new_n10246));
  NAND2xp33_ASAP7_75t_L     g09990(.A(\b[59] ), .B(new_n272), .Y(new_n10247));
  INVx1_ASAP7_75t_L         g09991(.A(new_n9948), .Y(new_n10248));
  NOR2xp33_ASAP7_75t_L      g09992(.A(\b[59] ), .B(\b[60] ), .Y(new_n10249));
  INVx1_ASAP7_75t_L         g09993(.A(\b[60] ), .Y(new_n10250));
  NOR2xp33_ASAP7_75t_L      g09994(.A(new_n9947), .B(new_n10250), .Y(new_n10251));
  NOR2xp33_ASAP7_75t_L      g09995(.A(new_n10249), .B(new_n10251), .Y(new_n10252));
  INVx1_ASAP7_75t_L         g09996(.A(new_n10252), .Y(new_n10253));
  O2A1O1Ixp33_ASAP7_75t_L   g09997(.A1(new_n9952), .A2(new_n9951), .B(new_n10248), .C(new_n10253), .Y(new_n10254));
  INVx1_ASAP7_75t_L         g09998(.A(new_n9921), .Y(new_n10255));
  A2O1A1Ixp33_ASAP7_75t_L   g09999(.A1(new_n9923), .A2(new_n10255), .B(new_n9946), .C(new_n10248), .Y(new_n10256));
  NOR2xp33_ASAP7_75t_L      g10000(.A(new_n10252), .B(new_n10256), .Y(new_n10257));
  NOR2xp33_ASAP7_75t_L      g10001(.A(new_n10254), .B(new_n10257), .Y(new_n10258));
  NAND2xp33_ASAP7_75t_L     g10002(.A(new_n267), .B(new_n10258), .Y(new_n10259));
  AOI22xp33_ASAP7_75t_L     g10003(.A1(\b[58] ), .A2(new_n282), .B1(\b[60] ), .B2(new_n303), .Y(new_n10260));
  NAND4xp25_ASAP7_75t_L     g10004(.A(new_n10259), .B(\a[2] ), .C(new_n10247), .D(new_n10260), .Y(new_n10261));
  NAND2xp33_ASAP7_75t_L     g10005(.A(new_n10260), .B(new_n10259), .Y(new_n10262));
  A2O1A1Ixp33_ASAP7_75t_L   g10006(.A1(\b[59] ), .A2(new_n272), .B(new_n10262), .C(new_n262), .Y(new_n10263));
  NAND2xp33_ASAP7_75t_L     g10007(.A(new_n10261), .B(new_n10263), .Y(new_n10264));
  AOI22xp33_ASAP7_75t_L     g10008(.A1(new_n344), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n370), .Y(new_n10265));
  OAI221xp5_ASAP7_75t_L     g10009(.A1(new_n429), .A2(new_n9323), .B1(new_n366), .B2(new_n9627), .C(new_n10265), .Y(new_n10266));
  XNOR2x2_ASAP7_75t_L       g10010(.A(new_n338), .B(new_n10266), .Y(new_n10267));
  NAND3xp33_ASAP7_75t_L     g10011(.A(new_n10204), .B(new_n10207), .C(new_n10205), .Y(new_n10268));
  A2O1A1Ixp33_ASAP7_75t_L   g10012(.A1(new_n10213), .A2(new_n10214), .B(new_n9961), .C(new_n10268), .Y(new_n10269));
  AOI22xp33_ASAP7_75t_L     g10013(.A1(new_n444), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n471), .Y(new_n10270));
  OAI221xp5_ASAP7_75t_L     g10014(.A1(new_n468), .A2(new_n8165), .B1(new_n469), .B2(new_n8465), .C(new_n10270), .Y(new_n10271));
  XNOR2x2_ASAP7_75t_L       g10015(.A(\a[8] ), .B(new_n10271), .Y(new_n10272));
  NAND2xp33_ASAP7_75t_L     g10016(.A(new_n10195), .B(new_n10190), .Y(new_n10273));
  NOR2xp33_ASAP7_75t_L      g10017(.A(new_n7593), .B(new_n821), .Y(new_n10274));
  NOR2xp33_ASAP7_75t_L      g10018(.A(new_n577), .B(new_n7623), .Y(new_n10275));
  AOI22xp33_ASAP7_75t_L     g10019(.A1(\b[49] ), .A2(new_n651), .B1(\b[51] ), .B2(new_n581), .Y(new_n10276));
  INVx1_ASAP7_75t_L         g10020(.A(new_n10276), .Y(new_n10277));
  NOR4xp25_ASAP7_75t_L      g10021(.A(new_n10275), .B(new_n574), .C(new_n10277), .D(new_n10274), .Y(new_n10278));
  NOR2xp33_ASAP7_75t_L      g10022(.A(new_n10277), .B(new_n10275), .Y(new_n10279));
  O2A1O1Ixp33_ASAP7_75t_L   g10023(.A1(new_n7593), .A2(new_n821), .B(new_n10279), .C(\a[11] ), .Y(new_n10280));
  NOR2xp33_ASAP7_75t_L      g10024(.A(new_n10278), .B(new_n10280), .Y(new_n10281));
  INVx1_ASAP7_75t_L         g10025(.A(new_n10187), .Y(new_n10282));
  OAI21xp33_ASAP7_75t_L     g10026(.A1(new_n10188), .A2(new_n10194), .B(new_n10282), .Y(new_n10283));
  AOI22xp33_ASAP7_75t_L     g10027(.A1(new_n811), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n900), .Y(new_n10284));
  OAI221xp5_ASAP7_75t_L     g10028(.A1(new_n904), .A2(new_n6812), .B1(new_n898), .B2(new_n6837), .C(new_n10284), .Y(new_n10285));
  XNOR2x2_ASAP7_75t_L       g10029(.A(\a[14] ), .B(new_n10285), .Y(new_n10286));
  INVx1_ASAP7_75t_L         g10030(.A(new_n10286), .Y(new_n10287));
  AOI31xp33_ASAP7_75t_L     g10031(.A1(new_n10181), .A2(new_n9972), .A3(new_n10179), .B(new_n10183), .Y(new_n10288));
  NAND2xp33_ASAP7_75t_L     g10032(.A(\b[44] ), .B(new_n1080), .Y(new_n10289));
  NAND2xp33_ASAP7_75t_L     g10033(.A(new_n1073), .B(new_n7066), .Y(new_n10290));
  AOI22xp33_ASAP7_75t_L     g10034(.A1(new_n1076), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n1253), .Y(new_n10291));
  AND4x1_ASAP7_75t_L        g10035(.A(new_n10291), .B(new_n10290), .C(new_n10289), .D(\a[17] ), .Y(new_n10292));
  AOI31xp33_ASAP7_75t_L     g10036(.A1(new_n10290), .A2(new_n10289), .A3(new_n10291), .B(\a[17] ), .Y(new_n10293));
  NOR2xp33_ASAP7_75t_L      g10037(.A(new_n10293), .B(new_n10292), .Y(new_n10294));
  INVx1_ASAP7_75t_L         g10038(.A(new_n10294), .Y(new_n10295));
  INVx1_ASAP7_75t_L         g10039(.A(new_n10140), .Y(new_n10296));
  AND3x1_ASAP7_75t_L        g10040(.A(new_n10133), .B(new_n10136), .C(new_n10296), .Y(new_n10297));
  A2O1A1O1Ixp25_ASAP7_75t_L g10041(.A1(new_n9836), .A2(new_n9835), .B(new_n10144), .C(new_n10143), .D(new_n10297), .Y(new_n10298));
  AOI22xp33_ASAP7_75t_L     g10042(.A1(new_n2114), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n2259), .Y(new_n10299));
  OAI221xp5_ASAP7_75t_L     g10043(.A1(new_n2109), .A2(new_n3804), .B1(new_n2257), .B2(new_n4223), .C(new_n10299), .Y(new_n10300));
  XNOR2x2_ASAP7_75t_L       g10044(.A(\a[26] ), .B(new_n10300), .Y(new_n10301));
  INVx1_ASAP7_75t_L         g10045(.A(new_n10301), .Y(new_n10302));
  INVx1_ASAP7_75t_L         g10046(.A(new_n10084), .Y(new_n10303));
  AO31x2_ASAP7_75t_L        g10047(.A1(new_n10086), .A2(new_n9761), .A3(new_n10085), .B(new_n10303), .Y(new_n10304));
  AOI22xp33_ASAP7_75t_L     g10048(.A1(new_n4920), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n5167), .Y(new_n10305));
  OAI221xp5_ASAP7_75t_L     g10049(.A1(new_n5154), .A2(new_n1539), .B1(new_n5158), .B2(new_n1662), .C(new_n10305), .Y(new_n10306));
  XNOR2x2_ASAP7_75t_L       g10050(.A(\a[41] ), .B(new_n10306), .Y(new_n10307));
  INVx1_ASAP7_75t_L         g10051(.A(new_n10307), .Y(new_n10308));
  A2O1A1Ixp33_ASAP7_75t_L   g10052(.A1(new_n9475), .A2(new_n9465), .B(new_n9756), .C(new_n9751), .Y(new_n10309));
  NOR3xp33_ASAP7_75t_L      g10053(.A(new_n10070), .B(new_n10074), .C(new_n10076), .Y(new_n10310));
  OAI22xp33_ASAP7_75t_L     g10054(.A1(new_n5895), .A2(new_n1030), .B1(new_n1313), .B2(new_n5894), .Y(new_n10311));
  AOI221xp5_ASAP7_75t_L     g10055(.A1(new_n5628), .A2(\b[17] ), .B1(new_n5621), .B2(new_n1319), .C(new_n10311), .Y(new_n10312));
  XNOR2x2_ASAP7_75t_L       g10056(.A(new_n5619), .B(new_n10312), .Y(new_n10313));
  INVx1_ASAP7_75t_L         g10057(.A(new_n10313), .Y(new_n10314));
  NOR3xp33_ASAP7_75t_L      g10058(.A(new_n10066), .B(new_n10067), .C(new_n10064), .Y(new_n10315));
  INVx1_ASAP7_75t_L         g10059(.A(new_n10315), .Y(new_n10316));
  AOI22xp33_ASAP7_75t_L     g10060(.A1(new_n6376), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n6648), .Y(new_n10317));
  OAI221xp5_ASAP7_75t_L     g10061(.A1(new_n6646), .A2(new_n869), .B1(new_n6636), .B2(new_n950), .C(new_n10317), .Y(new_n10318));
  XNOR2x2_ASAP7_75t_L       g10062(.A(\a[47] ), .B(new_n10318), .Y(new_n10319));
  NOR2xp33_ASAP7_75t_L      g10063(.A(new_n9731), .B(new_n10005), .Y(new_n10320));
  NOR3xp33_ASAP7_75t_L      g10064(.A(new_n10053), .B(new_n10047), .C(new_n10009), .Y(new_n10321));
  O2A1O1Ixp33_ASAP7_75t_L   g10065(.A1(new_n10320), .A2(new_n9737), .B(new_n10054), .C(new_n10321), .Y(new_n10322));
  AOI22xp33_ASAP7_75t_L     g10066(.A1(new_n7111), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n7391), .Y(new_n10323));
  OAI221xp5_ASAP7_75t_L     g10067(.A1(new_n8558), .A2(new_n679), .B1(new_n8237), .B2(new_n768), .C(new_n10323), .Y(new_n10324));
  XNOR2x2_ASAP7_75t_L       g10068(.A(\a[50] ), .B(new_n10324), .Y(new_n10325));
  INVx1_ASAP7_75t_L         g10069(.A(new_n10325), .Y(new_n10326));
  A2O1A1Ixp33_ASAP7_75t_L   g10070(.A1(new_n9722), .A2(new_n9721), .B(new_n10043), .C(new_n10052), .Y(new_n10327));
  NAND5xp2_ASAP7_75t_L      g10071(.A(\a[59] ), .B(new_n9701), .C(new_n9698), .D(new_n9704), .E(new_n9416), .Y(new_n10328));
  INVx1_ASAP7_75t_L         g10072(.A(\a[60] ), .Y(new_n10329));
  NAND2xp33_ASAP7_75t_L     g10073(.A(\a[59] ), .B(new_n10329), .Y(new_n10330));
  NAND2xp33_ASAP7_75t_L     g10074(.A(\a[60] ), .B(new_n9693), .Y(new_n10331));
  AND2x2_ASAP7_75t_L        g10075(.A(new_n10330), .B(new_n10331), .Y(new_n10332));
  NOR2xp33_ASAP7_75t_L      g10076(.A(new_n258), .B(new_n10332), .Y(new_n10333));
  OAI21xp33_ASAP7_75t_L     g10077(.A1(new_n10328), .A2(new_n10029), .B(new_n10333), .Y(new_n10334));
  INVx1_ASAP7_75t_L         g10078(.A(new_n10328), .Y(new_n10335));
  INVx1_ASAP7_75t_L         g10079(.A(new_n10333), .Y(new_n10336));
  NAND3xp33_ASAP7_75t_L     g10080(.A(new_n10035), .B(new_n10335), .C(new_n10336), .Y(new_n10337));
  OAI22xp33_ASAP7_75t_L     g10081(.A1(new_n10026), .A2(new_n261), .B1(new_n298), .B2(new_n9699), .Y(new_n10338));
  AOI221xp5_ASAP7_75t_L     g10082(.A1(\b[2] ), .A2(new_n9703), .B1(new_n406), .B2(new_n9697), .C(new_n10338), .Y(new_n10339));
  XNOR2x2_ASAP7_75t_L       g10083(.A(new_n9693), .B(new_n10339), .Y(new_n10340));
  AO21x2_ASAP7_75t_L        g10084(.A1(new_n10334), .A2(new_n10337), .B(new_n10340), .Y(new_n10341));
  NAND3xp33_ASAP7_75t_L     g10085(.A(new_n10337), .B(new_n10340), .C(new_n10334), .Y(new_n10342));
  INVx1_ASAP7_75t_L         g10086(.A(new_n8835), .Y(new_n10343));
  AOI22xp33_ASAP7_75t_L     g10087(.A1(new_n8831), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n9115), .Y(new_n10344));
  OAI221xp5_ASAP7_75t_L     g10088(.A1(new_n10343), .A2(new_n354), .B1(new_n10016), .B2(new_n390), .C(new_n10344), .Y(new_n10345));
  NOR2xp33_ASAP7_75t_L      g10089(.A(new_n8826), .B(new_n10345), .Y(new_n10346));
  INVx1_ASAP7_75t_L         g10090(.A(new_n10346), .Y(new_n10347));
  NAND2xp33_ASAP7_75t_L     g10091(.A(new_n8826), .B(new_n10345), .Y(new_n10348));
  NAND4xp25_ASAP7_75t_L     g10092(.A(new_n10347), .B(new_n10341), .C(new_n10342), .D(new_n10348), .Y(new_n10349));
  AOI21xp33_ASAP7_75t_L     g10093(.A1(new_n10337), .A2(new_n10334), .B(new_n10340), .Y(new_n10350));
  AND3x1_ASAP7_75t_L        g10094(.A(new_n10337), .B(new_n10340), .C(new_n10334), .Y(new_n10351));
  INVx1_ASAP7_75t_L         g10095(.A(new_n10348), .Y(new_n10352));
  OAI22xp33_ASAP7_75t_L     g10096(.A1(new_n10346), .A2(new_n10352), .B1(new_n10350), .B2(new_n10351), .Y(new_n10353));
  NAND2xp33_ASAP7_75t_L     g10097(.A(new_n10349), .B(new_n10353), .Y(new_n10354));
  OAI21xp33_ASAP7_75t_L     g10098(.A1(new_n10037), .A2(new_n10039), .B(new_n10040), .Y(new_n10355));
  NOR2xp33_ASAP7_75t_L      g10099(.A(new_n10355), .B(new_n10354), .Y(new_n10356));
  AOI21xp33_ASAP7_75t_L     g10100(.A1(new_n10015), .A2(new_n10041), .B(new_n10034), .Y(new_n10357));
  AOI21xp33_ASAP7_75t_L     g10101(.A1(new_n10353), .A2(new_n10349), .B(new_n10357), .Y(new_n10358));
  AOI22xp33_ASAP7_75t_L     g10102(.A1(new_n7960), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n8537), .Y(new_n10359));
  OAI221xp5_ASAP7_75t_L     g10103(.A1(new_n8817), .A2(new_n488), .B1(new_n7957), .B2(new_n548), .C(new_n10359), .Y(new_n10360));
  NOR2xp33_ASAP7_75t_L      g10104(.A(new_n7954), .B(new_n10360), .Y(new_n10361));
  AND2x2_ASAP7_75t_L        g10105(.A(new_n7954), .B(new_n10360), .Y(new_n10362));
  OAI22xp33_ASAP7_75t_L     g10106(.A1(new_n10356), .A2(new_n10358), .B1(new_n10362), .B2(new_n10361), .Y(new_n10363));
  NAND3xp33_ASAP7_75t_L     g10107(.A(new_n10357), .B(new_n10353), .C(new_n10349), .Y(new_n10364));
  A2O1A1Ixp33_ASAP7_75t_L   g10108(.A1(new_n10041), .A2(new_n10015), .B(new_n10034), .C(new_n10354), .Y(new_n10365));
  XNOR2x2_ASAP7_75t_L       g10109(.A(\a[53] ), .B(new_n10360), .Y(new_n10366));
  NAND3xp33_ASAP7_75t_L     g10110(.A(new_n10365), .B(new_n10364), .C(new_n10366), .Y(new_n10367));
  NAND3xp33_ASAP7_75t_L     g10111(.A(new_n10327), .B(new_n10363), .C(new_n10367), .Y(new_n10368));
  AOI21xp33_ASAP7_75t_L     g10112(.A1(new_n10367), .A2(new_n10363), .B(new_n10327), .Y(new_n10369));
  INVx1_ASAP7_75t_L         g10113(.A(new_n10369), .Y(new_n10370));
  AOI21xp33_ASAP7_75t_L     g10114(.A1(new_n10370), .A2(new_n10368), .B(new_n10326), .Y(new_n10371));
  NAND2xp33_ASAP7_75t_L     g10115(.A(new_n10367), .B(new_n10363), .Y(new_n10372));
  O2A1O1Ixp33_ASAP7_75t_L   g10116(.A1(new_n10010), .A2(new_n10043), .B(new_n10052), .C(new_n10372), .Y(new_n10373));
  NOR3xp33_ASAP7_75t_L      g10117(.A(new_n10373), .B(new_n10369), .C(new_n10325), .Y(new_n10374));
  NOR3xp33_ASAP7_75t_L      g10118(.A(new_n10371), .B(new_n10322), .C(new_n10374), .Y(new_n10375));
  AO21x2_ASAP7_75t_L        g10119(.A1(new_n10054), .A2(new_n10006), .B(new_n10321), .Y(new_n10376));
  OAI21xp33_ASAP7_75t_L     g10120(.A1(new_n10369), .A2(new_n10373), .B(new_n10325), .Y(new_n10377));
  NAND3xp33_ASAP7_75t_L     g10121(.A(new_n10370), .B(new_n10368), .C(new_n10326), .Y(new_n10378));
  AOI21xp33_ASAP7_75t_L     g10122(.A1(new_n10378), .A2(new_n10377), .B(new_n10376), .Y(new_n10379));
  NOR3xp33_ASAP7_75t_L      g10123(.A(new_n10375), .B(new_n10379), .C(new_n10319), .Y(new_n10380));
  INVx1_ASAP7_75t_L         g10124(.A(new_n10319), .Y(new_n10381));
  NAND3xp33_ASAP7_75t_L     g10125(.A(new_n10376), .B(new_n10378), .C(new_n10377), .Y(new_n10382));
  OAI21xp33_ASAP7_75t_L     g10126(.A1(new_n10374), .A2(new_n10371), .B(new_n10322), .Y(new_n10383));
  AOI21xp33_ASAP7_75t_L     g10127(.A1(new_n10383), .A2(new_n10382), .B(new_n10381), .Y(new_n10384));
  AOI211xp5_ASAP7_75t_L     g10128(.A1(new_n10077), .A2(new_n10316), .B(new_n10380), .C(new_n10384), .Y(new_n10385));
  NAND3xp33_ASAP7_75t_L     g10129(.A(new_n10381), .B(new_n10383), .C(new_n10382), .Y(new_n10386));
  OAI21xp33_ASAP7_75t_L     g10130(.A1(new_n10379), .A2(new_n10375), .B(new_n10319), .Y(new_n10387));
  AOI211xp5_ASAP7_75t_L     g10131(.A1(new_n10386), .A2(new_n10387), .B(new_n10315), .C(new_n10070), .Y(new_n10388));
  OAI21xp33_ASAP7_75t_L     g10132(.A1(new_n10388), .A2(new_n10385), .B(new_n10314), .Y(new_n10389));
  OAI211xp5_ASAP7_75t_L     g10133(.A1(new_n10315), .A2(new_n10070), .B(new_n10386), .C(new_n10387), .Y(new_n10390));
  OAI211xp5_ASAP7_75t_L     g10134(.A1(new_n10380), .A2(new_n10384), .B(new_n10077), .C(new_n10316), .Y(new_n10391));
  NAND3xp33_ASAP7_75t_L     g10135(.A(new_n10390), .B(new_n10313), .C(new_n10391), .Y(new_n10392));
  NAND2xp33_ASAP7_75t_L     g10136(.A(new_n10392), .B(new_n10389), .Y(new_n10393));
  A2O1A1Ixp33_ASAP7_75t_L   g10137(.A1(new_n10080), .A2(new_n10309), .B(new_n10310), .C(new_n10393), .Y(new_n10394));
  INVx1_ASAP7_75t_L         g10138(.A(new_n10310), .Y(new_n10395));
  A2O1A1Ixp33_ASAP7_75t_L   g10139(.A1(new_n10075), .A2(new_n10079), .B(new_n10082), .C(new_n10395), .Y(new_n10396));
  NOR2xp33_ASAP7_75t_L      g10140(.A(new_n10396), .B(new_n10393), .Y(new_n10397));
  INVx1_ASAP7_75t_L         g10141(.A(new_n10397), .Y(new_n10398));
  NAND3xp33_ASAP7_75t_L     g10142(.A(new_n10398), .B(new_n10394), .C(new_n10308), .Y(new_n10399));
  AOI21xp33_ASAP7_75t_L     g10143(.A1(new_n10390), .A2(new_n10391), .B(new_n10313), .Y(new_n10400));
  NOR3xp33_ASAP7_75t_L      g10144(.A(new_n10385), .B(new_n10314), .C(new_n10388), .Y(new_n10401));
  NOR2xp33_ASAP7_75t_L      g10145(.A(new_n10400), .B(new_n10401), .Y(new_n10402));
  A2O1A1O1Ixp25_ASAP7_75t_L g10146(.A1(new_n10075), .A2(new_n10079), .B(new_n10082), .C(new_n10395), .D(new_n10402), .Y(new_n10403));
  OAI21xp33_ASAP7_75t_L     g10147(.A1(new_n10397), .A2(new_n10403), .B(new_n10307), .Y(new_n10404));
  NAND3xp33_ASAP7_75t_L     g10148(.A(new_n10304), .B(new_n10399), .C(new_n10404), .Y(new_n10405));
  AOI31xp33_ASAP7_75t_L     g10149(.A1(new_n10086), .A2(new_n9761), .A3(new_n10085), .B(new_n10303), .Y(new_n10406));
  NAND2xp33_ASAP7_75t_L     g10150(.A(new_n10404), .B(new_n10399), .Y(new_n10407));
  NAND2xp33_ASAP7_75t_L     g10151(.A(new_n10406), .B(new_n10407), .Y(new_n10408));
  OAI22xp33_ASAP7_75t_L     g10152(.A1(new_n4501), .A2(new_n1774), .B1(new_n1929), .B2(new_n4275), .Y(new_n10409));
  AOI221xp5_ASAP7_75t_L     g10153(.A1(new_n4285), .A2(\b[23] ), .B1(new_n4274), .B2(new_n1935), .C(new_n10409), .Y(new_n10410));
  XNOR2x2_ASAP7_75t_L       g10154(.A(new_n4268), .B(new_n10410), .Y(new_n10411));
  NAND3xp33_ASAP7_75t_L     g10155(.A(new_n10408), .B(new_n10405), .C(new_n10411), .Y(new_n10412));
  NOR2xp33_ASAP7_75t_L      g10156(.A(new_n10406), .B(new_n10407), .Y(new_n10413));
  AOI21xp33_ASAP7_75t_L     g10157(.A1(new_n10404), .A2(new_n10399), .B(new_n10304), .Y(new_n10414));
  INVx1_ASAP7_75t_L         g10158(.A(new_n10411), .Y(new_n10415));
  OAI21xp33_ASAP7_75t_L     g10159(.A1(new_n10414), .A2(new_n10413), .B(new_n10415), .Y(new_n10416));
  A2O1A1O1Ixp25_ASAP7_75t_L g10160(.A1(new_n9775), .A2(new_n9661), .B(new_n9989), .C(new_n10105), .D(new_n10089), .Y(new_n10417));
  NAND3xp33_ASAP7_75t_L     g10161(.A(new_n10417), .B(new_n10416), .C(new_n10412), .Y(new_n10418));
  NOR3xp33_ASAP7_75t_L      g10162(.A(new_n10413), .B(new_n10414), .C(new_n10415), .Y(new_n10419));
  AOI21xp33_ASAP7_75t_L     g10163(.A1(new_n10408), .A2(new_n10405), .B(new_n10411), .Y(new_n10420));
  OAI21xp33_ASAP7_75t_L     g10164(.A1(new_n10096), .A2(new_n9990), .B(new_n10104), .Y(new_n10421));
  OAI21xp33_ASAP7_75t_L     g10165(.A1(new_n10419), .A2(new_n10420), .B(new_n10421), .Y(new_n10422));
  NAND2xp33_ASAP7_75t_L     g10166(.A(\b[26] ), .B(new_n3639), .Y(new_n10423));
  NAND2xp33_ASAP7_75t_L     g10167(.A(new_n3630), .B(new_n2504), .Y(new_n10424));
  AOI22xp33_ASAP7_75t_L     g10168(.A1(new_n3633), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n3858), .Y(new_n10425));
  NAND4xp25_ASAP7_75t_L     g10169(.A(new_n10424), .B(\a[35] ), .C(new_n10423), .D(new_n10425), .Y(new_n10426));
  NAND2xp33_ASAP7_75t_L     g10170(.A(new_n10425), .B(new_n10424), .Y(new_n10427));
  A2O1A1Ixp33_ASAP7_75t_L   g10171(.A1(\b[26] ), .A2(new_n3639), .B(new_n10427), .C(new_n3628), .Y(new_n10428));
  NAND2xp33_ASAP7_75t_L     g10172(.A(new_n10426), .B(new_n10428), .Y(new_n10429));
  INVx1_ASAP7_75t_L         g10173(.A(new_n10429), .Y(new_n10430));
  NAND3xp33_ASAP7_75t_L     g10174(.A(new_n10422), .B(new_n10418), .C(new_n10430), .Y(new_n10431));
  NOR3xp33_ASAP7_75t_L      g10175(.A(new_n10421), .B(new_n10420), .C(new_n10419), .Y(new_n10432));
  AOI21xp33_ASAP7_75t_L     g10176(.A1(new_n10416), .A2(new_n10412), .B(new_n10417), .Y(new_n10433));
  OAI21xp33_ASAP7_75t_L     g10177(.A1(new_n10433), .A2(new_n10432), .B(new_n10429), .Y(new_n10434));
  NAND2xp33_ASAP7_75t_L     g10178(.A(new_n10431), .B(new_n10434), .Y(new_n10435));
  NAND3xp33_ASAP7_75t_L     g10179(.A(new_n10099), .B(new_n10097), .C(new_n10109), .Y(new_n10436));
  A2O1A1Ixp33_ASAP7_75t_L   g10180(.A1(new_n10110), .A2(new_n10103), .B(new_n10114), .C(new_n10436), .Y(new_n10437));
  NOR2xp33_ASAP7_75t_L      g10181(.A(new_n10435), .B(new_n10437), .Y(new_n10438));
  NAND2xp33_ASAP7_75t_L     g10182(.A(new_n10097), .B(new_n10099), .Y(new_n10439));
  NOR3xp33_ASAP7_75t_L      g10183(.A(new_n10432), .B(new_n10433), .C(new_n10429), .Y(new_n10440));
  AOI21xp33_ASAP7_75t_L     g10184(.A1(new_n10422), .A2(new_n10418), .B(new_n10430), .Y(new_n10441));
  NOR2xp33_ASAP7_75t_L      g10185(.A(new_n10441), .B(new_n10440), .Y(new_n10442));
  O2A1O1Ixp33_ASAP7_75t_L   g10186(.A1(new_n10439), .A2(new_n10102), .B(new_n10121), .C(new_n10442), .Y(new_n10443));
  AOI22xp33_ASAP7_75t_L     g10187(.A1(new_n3029), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n3258), .Y(new_n10444));
  OAI221xp5_ASAP7_75t_L     g10188(.A1(new_n3024), .A2(new_n2688), .B1(new_n3256), .B2(new_n2990), .C(new_n10444), .Y(new_n10445));
  XNOR2x2_ASAP7_75t_L       g10189(.A(\a[32] ), .B(new_n10445), .Y(new_n10446));
  OAI21xp33_ASAP7_75t_L     g10190(.A1(new_n10438), .A2(new_n10443), .B(new_n10446), .Y(new_n10447));
  NAND3xp33_ASAP7_75t_L     g10191(.A(new_n10442), .B(new_n10121), .C(new_n10436), .Y(new_n10448));
  NAND2xp33_ASAP7_75t_L     g10192(.A(new_n10435), .B(new_n10437), .Y(new_n10449));
  INVx1_ASAP7_75t_L         g10193(.A(new_n10446), .Y(new_n10450));
  NAND3xp33_ASAP7_75t_L     g10194(.A(new_n10448), .B(new_n10449), .C(new_n10450), .Y(new_n10451));
  OAI211xp5_ASAP7_75t_L     g10195(.A1(new_n9805), .A2(new_n9803), .B(new_n9987), .C(new_n10123), .Y(new_n10452));
  NAND4xp25_ASAP7_75t_L     g10196(.A(new_n10452), .B(new_n10447), .C(new_n10119), .D(new_n10451), .Y(new_n10453));
  INVx1_ASAP7_75t_L         g10197(.A(new_n10119), .Y(new_n10454));
  AOI21xp33_ASAP7_75t_L     g10198(.A1(new_n10448), .A2(new_n10449), .B(new_n10450), .Y(new_n10455));
  NOR3xp33_ASAP7_75t_L      g10199(.A(new_n10443), .B(new_n10446), .C(new_n10438), .Y(new_n10456));
  NOR3xp33_ASAP7_75t_L      g10200(.A(new_n10113), .B(new_n10115), .C(new_n10118), .Y(new_n10457));
  AOI211xp5_ASAP7_75t_L     g10201(.A1(new_n9808), .A2(new_n9660), .B(new_n9986), .C(new_n10457), .Y(new_n10458));
  OAI22xp33_ASAP7_75t_L     g10202(.A1(new_n10458), .A2(new_n10454), .B1(new_n10455), .B2(new_n10456), .Y(new_n10459));
  NOR2xp33_ASAP7_75t_L      g10203(.A(new_n3207), .B(new_n2547), .Y(new_n10460));
  NOR2xp33_ASAP7_75t_L      g10204(.A(new_n2734), .B(new_n3572), .Y(new_n10461));
  AOI22xp33_ASAP7_75t_L     g10205(.A1(new_n2552), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n2736), .Y(new_n10462));
  INVx1_ASAP7_75t_L         g10206(.A(new_n10462), .Y(new_n10463));
  NOR4xp25_ASAP7_75t_L      g10207(.A(new_n10461), .B(new_n2538), .C(new_n10463), .D(new_n10460), .Y(new_n10464));
  NOR2xp33_ASAP7_75t_L      g10208(.A(new_n10463), .B(new_n10461), .Y(new_n10465));
  O2A1O1Ixp33_ASAP7_75t_L   g10209(.A1(new_n3207), .A2(new_n2547), .B(new_n10465), .C(\a[29] ), .Y(new_n10466));
  NOR2xp33_ASAP7_75t_L      g10210(.A(new_n10464), .B(new_n10466), .Y(new_n10467));
  NAND3xp33_ASAP7_75t_L     g10211(.A(new_n10459), .B(new_n10453), .C(new_n10467), .Y(new_n10468));
  NOR4xp25_ASAP7_75t_L      g10212(.A(new_n10458), .B(new_n10456), .C(new_n10455), .D(new_n10454), .Y(new_n10469));
  AOI22xp33_ASAP7_75t_L     g10213(.A1(new_n10447), .A2(new_n10451), .B1(new_n10452), .B2(new_n10119), .Y(new_n10470));
  OR2x4_ASAP7_75t_L         g10214(.A(new_n10464), .B(new_n10466), .Y(new_n10471));
  OAI21xp33_ASAP7_75t_L     g10215(.A1(new_n10470), .A2(new_n10469), .B(new_n10471), .Y(new_n10472));
  NAND2xp33_ASAP7_75t_L     g10216(.A(new_n10468), .B(new_n10472), .Y(new_n10473));
  A2O1A1Ixp33_ASAP7_75t_L   g10217(.A1(new_n10128), .A2(new_n9979), .B(new_n10135), .C(new_n10473), .Y(new_n10474));
  A2O1A1O1Ixp25_ASAP7_75t_L g10218(.A1(new_n9821), .A2(new_n9819), .B(new_n9813), .C(new_n10128), .D(new_n10135), .Y(new_n10475));
  NAND3xp33_ASAP7_75t_L     g10219(.A(new_n10475), .B(new_n10468), .C(new_n10472), .Y(new_n10476));
  NAND3xp33_ASAP7_75t_L     g10220(.A(new_n10474), .B(new_n10302), .C(new_n10476), .Y(new_n10477));
  AOI21xp33_ASAP7_75t_L     g10221(.A1(new_n10472), .A2(new_n10468), .B(new_n10475), .Y(new_n10478));
  AND3x1_ASAP7_75t_L        g10222(.A(new_n10475), .B(new_n10472), .C(new_n10468), .Y(new_n10479));
  OAI21xp33_ASAP7_75t_L     g10223(.A1(new_n10478), .A2(new_n10479), .B(new_n10301), .Y(new_n10480));
  NAND2xp33_ASAP7_75t_L     g10224(.A(new_n10477), .B(new_n10480), .Y(new_n10481));
  NAND2xp33_ASAP7_75t_L     g10225(.A(new_n10481), .B(new_n10298), .Y(new_n10482));
  AND2x2_ASAP7_75t_L        g10226(.A(new_n10477), .B(new_n10480), .Y(new_n10483));
  A2O1A1Ixp33_ASAP7_75t_L   g10227(.A1(new_n10145), .A2(new_n10143), .B(new_n10297), .C(new_n10483), .Y(new_n10484));
  AOI22xp33_ASAP7_75t_L     g10228(.A1(new_n1704), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1837), .Y(new_n10485));
  OAI221xp5_ASAP7_75t_L     g10229(.A1(new_n1699), .A2(new_n4632), .B1(new_n1827), .B2(new_n4858), .C(new_n10485), .Y(new_n10486));
  NOR2xp33_ASAP7_75t_L      g10230(.A(new_n1689), .B(new_n10486), .Y(new_n10487));
  AND2x2_ASAP7_75t_L        g10231(.A(new_n1689), .B(new_n10486), .Y(new_n10488));
  NOR2xp33_ASAP7_75t_L      g10232(.A(new_n10487), .B(new_n10488), .Y(new_n10489));
  NAND3xp33_ASAP7_75t_L     g10233(.A(new_n10484), .B(new_n10482), .C(new_n10489), .Y(new_n10490));
  INVx1_ASAP7_75t_L         g10234(.A(new_n10297), .Y(new_n10491));
  A2O1A1Ixp33_ASAP7_75t_L   g10235(.A1(new_n10142), .A2(new_n10141), .B(new_n10148), .C(new_n10491), .Y(new_n10492));
  NOR2xp33_ASAP7_75t_L      g10236(.A(new_n10483), .B(new_n10492), .Y(new_n10493));
  O2A1O1Ixp33_ASAP7_75t_L   g10237(.A1(new_n10147), .A2(new_n10148), .B(new_n10491), .C(new_n10481), .Y(new_n10494));
  OAI22xp33_ASAP7_75t_L     g10238(.A1(new_n10493), .A2(new_n10494), .B1(new_n10488), .B2(new_n10487), .Y(new_n10495));
  NOR2xp33_ASAP7_75t_L      g10239(.A(new_n10149), .B(new_n10146), .Y(new_n10496));
  MAJIxp5_ASAP7_75t_L       g10240(.A(new_n10156), .B(new_n10152), .C(new_n10496), .Y(new_n10497));
  NAND3xp33_ASAP7_75t_L     g10241(.A(new_n10497), .B(new_n10495), .C(new_n10490), .Y(new_n10498));
  AO21x2_ASAP7_75t_L        g10242(.A1(new_n10490), .A2(new_n10495), .B(new_n10497), .Y(new_n10499));
  NOR2xp33_ASAP7_75t_L      g10243(.A(new_n5321), .B(new_n1373), .Y(new_n10500));
  INVx1_ASAP7_75t_L         g10244(.A(new_n10500), .Y(new_n10501));
  NAND3xp33_ASAP7_75t_L     g10245(.A(new_n5343), .B(new_n1365), .C(new_n5345), .Y(new_n10502));
  AOI22xp33_ASAP7_75t_L     g10246(.A1(new_n1360), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n1581), .Y(new_n10503));
  NAND4xp25_ASAP7_75t_L     g10247(.A(new_n10502), .B(\a[20] ), .C(new_n10501), .D(new_n10503), .Y(new_n10504));
  AOI31xp33_ASAP7_75t_L     g10248(.A1(new_n10502), .A2(new_n10501), .A3(new_n10503), .B(\a[20] ), .Y(new_n10505));
  INVx1_ASAP7_75t_L         g10249(.A(new_n10505), .Y(new_n10506));
  NAND2xp33_ASAP7_75t_L     g10250(.A(new_n10504), .B(new_n10506), .Y(new_n10507));
  AOI21xp33_ASAP7_75t_L     g10251(.A1(new_n10499), .A2(new_n10498), .B(new_n10507), .Y(new_n10508));
  NAND2xp33_ASAP7_75t_L     g10252(.A(new_n10152), .B(new_n10496), .Y(new_n10509));
  AND4x1_ASAP7_75t_L        g10253(.A(new_n10167), .B(new_n10509), .C(new_n10490), .D(new_n10495), .Y(new_n10510));
  AOI21xp33_ASAP7_75t_L     g10254(.A1(new_n10495), .A2(new_n10490), .B(new_n10497), .Y(new_n10511));
  INVx1_ASAP7_75t_L         g10255(.A(new_n10507), .Y(new_n10512));
  NOR3xp33_ASAP7_75t_L      g10256(.A(new_n10510), .B(new_n10511), .C(new_n10512), .Y(new_n10513));
  AOI211xp5_ASAP7_75t_L     g10257(.A1(new_n9868), .A2(new_n9870), .B(new_n9978), .C(new_n10173), .Y(new_n10514));
  NOR4xp25_ASAP7_75t_L      g10258(.A(new_n10514), .B(new_n10508), .C(new_n10513), .D(new_n10172), .Y(new_n10515));
  OAI21xp33_ASAP7_75t_L     g10259(.A1(new_n10511), .A2(new_n10510), .B(new_n10512), .Y(new_n10516));
  NAND3xp33_ASAP7_75t_L     g10260(.A(new_n10499), .B(new_n10498), .C(new_n10507), .Y(new_n10517));
  OAI211xp5_ASAP7_75t_L     g10261(.A1(new_n9862), .A2(new_n9864), .B(new_n9977), .C(new_n10169), .Y(new_n10518));
  AOI22xp33_ASAP7_75t_L     g10262(.A1(new_n10517), .A2(new_n10516), .B1(new_n10162), .B2(new_n10518), .Y(new_n10519));
  OAI21xp33_ASAP7_75t_L     g10263(.A1(new_n10515), .A2(new_n10519), .B(new_n10295), .Y(new_n10520));
  NAND4xp25_ASAP7_75t_L     g10264(.A(new_n10518), .B(new_n10162), .C(new_n10516), .D(new_n10517), .Y(new_n10521));
  OAI22xp33_ASAP7_75t_L     g10265(.A1(new_n10514), .A2(new_n10172), .B1(new_n10508), .B2(new_n10513), .Y(new_n10522));
  NAND3xp33_ASAP7_75t_L     g10266(.A(new_n10521), .B(new_n10522), .C(new_n10294), .Y(new_n10523));
  AOI21xp33_ASAP7_75t_L     g10267(.A1(new_n10523), .A2(new_n10520), .B(new_n10288), .Y(new_n10524));
  OAI31xp33_ASAP7_75t_L     g10268(.A1(new_n10185), .A2(new_n10184), .A3(new_n9876), .B(new_n10176), .Y(new_n10525));
  NAND2xp33_ASAP7_75t_L     g10269(.A(new_n10523), .B(new_n10520), .Y(new_n10526));
  NOR2xp33_ASAP7_75t_L      g10270(.A(new_n10526), .B(new_n10525), .Y(new_n10527));
  OAI21xp33_ASAP7_75t_L     g10271(.A1(new_n10524), .A2(new_n10527), .B(new_n10287), .Y(new_n10528));
  NAND2xp33_ASAP7_75t_L     g10272(.A(new_n10526), .B(new_n10525), .Y(new_n10529));
  NAND4xp25_ASAP7_75t_L     g10273(.A(new_n10182), .B(new_n10520), .C(new_n10523), .D(new_n10176), .Y(new_n10530));
  NAND3xp33_ASAP7_75t_L     g10274(.A(new_n10529), .B(new_n10286), .C(new_n10530), .Y(new_n10531));
  NAND2xp33_ASAP7_75t_L     g10275(.A(new_n10531), .B(new_n10528), .Y(new_n10532));
  NAND2xp33_ASAP7_75t_L     g10276(.A(new_n10283), .B(new_n10532), .Y(new_n10533));
  AO21x2_ASAP7_75t_L        g10277(.A1(new_n10182), .A2(new_n10186), .B(new_n9971), .Y(new_n10534));
  A2O1A1O1Ixp25_ASAP7_75t_L g10278(.A1(new_n9887), .A2(new_n9886), .B(new_n9883), .C(new_n10534), .D(new_n10187), .Y(new_n10535));
  NAND3xp33_ASAP7_75t_L     g10279(.A(new_n10535), .B(new_n10528), .C(new_n10531), .Y(new_n10536));
  AOI21xp33_ASAP7_75t_L     g10280(.A1(new_n10533), .A2(new_n10536), .B(new_n10281), .Y(new_n10537));
  INVx1_ASAP7_75t_L         g10281(.A(new_n10281), .Y(new_n10538));
  AOI21xp33_ASAP7_75t_L     g10282(.A1(new_n10531), .A2(new_n10528), .B(new_n10535), .Y(new_n10539));
  NOR2xp33_ASAP7_75t_L      g10283(.A(new_n10283), .B(new_n10532), .Y(new_n10540));
  NOR3xp33_ASAP7_75t_L      g10284(.A(new_n10540), .B(new_n10538), .C(new_n10539), .Y(new_n10541));
  NOR2xp33_ASAP7_75t_L      g10285(.A(new_n10537), .B(new_n10541), .Y(new_n10542));
  O2A1O1Ixp33_ASAP7_75t_L   g10286(.A1(new_n10273), .A2(new_n10201), .B(new_n10204), .C(new_n10542), .Y(new_n10543));
  MAJIxp5_ASAP7_75t_L       g10287(.A(new_n9968), .B(new_n10201), .C(new_n10273), .Y(new_n10544));
  OAI21xp33_ASAP7_75t_L     g10288(.A1(new_n10539), .A2(new_n10540), .B(new_n10538), .Y(new_n10545));
  NAND3xp33_ASAP7_75t_L     g10289(.A(new_n10533), .B(new_n10281), .C(new_n10536), .Y(new_n10546));
  NAND2xp33_ASAP7_75t_L     g10290(.A(new_n10546), .B(new_n10545), .Y(new_n10547));
  NOR2xp33_ASAP7_75t_L      g10291(.A(new_n10544), .B(new_n10547), .Y(new_n10548));
  OR3x1_ASAP7_75t_L         g10292(.A(new_n10543), .B(new_n10272), .C(new_n10548), .Y(new_n10549));
  OAI21xp33_ASAP7_75t_L     g10293(.A1(new_n10548), .A2(new_n10543), .B(new_n10272), .Y(new_n10550));
  NAND3xp33_ASAP7_75t_L     g10294(.A(new_n10269), .B(new_n10549), .C(new_n10550), .Y(new_n10551));
  NOR3xp33_ASAP7_75t_L      g10295(.A(new_n10543), .B(new_n10548), .C(new_n10272), .Y(new_n10552));
  OA21x2_ASAP7_75t_L        g10296(.A1(new_n10548), .A2(new_n10543), .B(new_n10272), .Y(new_n10553));
  OAI221xp5_ASAP7_75t_L     g10297(.A1(new_n10221), .A2(new_n9961), .B1(new_n10552), .B2(new_n10553), .C(new_n10268), .Y(new_n10554));
  NAND3xp33_ASAP7_75t_L     g10298(.A(new_n10554), .B(new_n10551), .C(new_n10267), .Y(new_n10555));
  AO21x2_ASAP7_75t_L        g10299(.A1(new_n10551), .A2(new_n10554), .B(new_n10267), .Y(new_n10556));
  NAND3xp33_ASAP7_75t_L     g10300(.A(new_n10556), .B(new_n10555), .C(new_n10264), .Y(new_n10557));
  INVx1_ASAP7_75t_L         g10301(.A(new_n10264), .Y(new_n10558));
  AND3x1_ASAP7_75t_L        g10302(.A(new_n10554), .B(new_n10551), .C(new_n10267), .Y(new_n10559));
  AOI21xp33_ASAP7_75t_L     g10303(.A1(new_n10554), .A2(new_n10551), .B(new_n10267), .Y(new_n10560));
  OAI21xp33_ASAP7_75t_L     g10304(.A1(new_n10560), .A2(new_n10559), .B(new_n10558), .Y(new_n10561));
  NAND4xp25_ASAP7_75t_L     g10305(.A(new_n10561), .B(new_n10557), .C(new_n10224), .D(new_n10225), .Y(new_n10562));
  NOR3xp33_ASAP7_75t_L      g10306(.A(new_n10559), .B(new_n10560), .C(new_n10558), .Y(new_n10563));
  AOI21xp33_ASAP7_75t_L     g10307(.A1(new_n10556), .A2(new_n10555), .B(new_n10264), .Y(new_n10564));
  OAI22xp33_ASAP7_75t_L     g10308(.A1(new_n10563), .A2(new_n10564), .B1(new_n10227), .B2(new_n10232), .Y(new_n10565));
  NAND2xp33_ASAP7_75t_L     g10309(.A(new_n10562), .B(new_n10565), .Y(new_n10566));
  O2A1O1Ixp33_ASAP7_75t_L   g10310(.A1(new_n10239), .A2(new_n10242), .B(new_n10246), .C(new_n10566), .Y(new_n10567));
  OAI21xp33_ASAP7_75t_L     g10311(.A1(new_n10237), .A2(new_n10238), .B(new_n9938), .Y(new_n10568));
  A2O1A1Ixp33_ASAP7_75t_L   g10312(.A1(new_n10568), .A2(new_n9940), .B(new_n10242), .C(new_n10246), .Y(new_n10569));
  AOI21xp33_ASAP7_75t_L     g10313(.A1(new_n10565), .A2(new_n10562), .B(new_n10569), .Y(new_n10570));
  NOR2xp33_ASAP7_75t_L      g10314(.A(new_n10567), .B(new_n10570), .Y(\f[60] ));
  INVx1_ASAP7_75t_L         g10315(.A(new_n10562), .Y(new_n10572));
  NOR3xp33_ASAP7_75t_L      g10316(.A(new_n10540), .B(new_n10539), .C(new_n10281), .Y(new_n10573));
  AOI22xp33_ASAP7_75t_L     g10317(.A1(\b[50] ), .A2(new_n651), .B1(\b[52] ), .B2(new_n581), .Y(new_n10574));
  OAI221xp5_ASAP7_75t_L     g10318(.A1(new_n821), .A2(new_n7616), .B1(new_n577), .B2(new_n7906), .C(new_n10574), .Y(new_n10575));
  XNOR2x2_ASAP7_75t_L       g10319(.A(\a[11] ), .B(new_n10575), .Y(new_n10576));
  INVx1_ASAP7_75t_L         g10320(.A(new_n10576), .Y(new_n10577));
  NOR3xp33_ASAP7_75t_L      g10321(.A(new_n10527), .B(new_n10524), .C(new_n10286), .Y(new_n10578));
  INVx1_ASAP7_75t_L         g10322(.A(new_n10578), .Y(new_n10579));
  A2O1A1Ixp33_ASAP7_75t_L   g10323(.A1(new_n10528), .A2(new_n10531), .B(new_n10535), .C(new_n10579), .Y(new_n10580));
  AOI22xp33_ASAP7_75t_L     g10324(.A1(new_n811), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n900), .Y(new_n10581));
  OAI221xp5_ASAP7_75t_L     g10325(.A1(new_n904), .A2(new_n6830), .B1(new_n898), .B2(new_n7323), .C(new_n10581), .Y(new_n10582));
  NOR2xp33_ASAP7_75t_L      g10326(.A(new_n806), .B(new_n10582), .Y(new_n10583));
  AND2x2_ASAP7_75t_L        g10327(.A(new_n806), .B(new_n10582), .Y(new_n10584));
  NOR2xp33_ASAP7_75t_L      g10328(.A(new_n10583), .B(new_n10584), .Y(new_n10585));
  NOR3xp33_ASAP7_75t_L      g10329(.A(new_n10519), .B(new_n10515), .C(new_n10294), .Y(new_n10586));
  AOI21xp33_ASAP7_75t_L     g10330(.A1(new_n10525), .A2(new_n10526), .B(new_n10586), .Y(new_n10587));
  AOI22xp33_ASAP7_75t_L     g10331(.A1(new_n1076), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n1253), .Y(new_n10588));
  OAI221xp5_ASAP7_75t_L     g10332(.A1(new_n1154), .A2(new_n6321), .B1(new_n1156), .B2(new_n6573), .C(new_n10588), .Y(new_n10589));
  XNOR2x2_ASAP7_75t_L       g10333(.A(\a[17] ), .B(new_n10589), .Y(new_n10590));
  OAI31xp33_ASAP7_75t_L     g10334(.A1(new_n10514), .A2(new_n10508), .A3(new_n10172), .B(new_n10517), .Y(new_n10591));
  NAND3xp33_ASAP7_75t_L     g10335(.A(new_n10471), .B(new_n10459), .C(new_n10453), .Y(new_n10592));
  A2O1A1Ixp33_ASAP7_75t_L   g10336(.A1(new_n10468), .A2(new_n10472), .B(new_n10475), .C(new_n10592), .Y(new_n10593));
  AOI31xp33_ASAP7_75t_L     g10337(.A1(new_n10452), .A2(new_n10447), .A3(new_n10119), .B(new_n10456), .Y(new_n10594));
  NOR3xp33_ASAP7_75t_L      g10338(.A(new_n10403), .B(new_n10397), .C(new_n10307), .Y(new_n10595));
  O2A1O1Ixp33_ASAP7_75t_L   g10339(.A1(new_n10303), .A2(new_n10087), .B(new_n10404), .C(new_n10595), .Y(new_n10596));
  AOI22xp33_ASAP7_75t_L     g10340(.A1(new_n4920), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n5167), .Y(new_n10597));
  OAI221xp5_ASAP7_75t_L     g10341(.A1(new_n5154), .A2(new_n1655), .B1(new_n5158), .B2(new_n1780), .C(new_n10597), .Y(new_n10598));
  XNOR2x2_ASAP7_75t_L       g10342(.A(\a[41] ), .B(new_n10598), .Y(new_n10599));
  INVx1_ASAP7_75t_L         g10343(.A(new_n10599), .Y(new_n10600));
  NOR3xp33_ASAP7_75t_L      g10344(.A(new_n10385), .B(new_n10388), .C(new_n10313), .Y(new_n10601));
  O2A1O1Ixp33_ASAP7_75t_L   g10345(.A1(new_n10400), .A2(new_n10401), .B(new_n10396), .C(new_n10601), .Y(new_n10602));
  A2O1A1Ixp33_ASAP7_75t_L   g10346(.A1(new_n10077), .A2(new_n10316), .B(new_n10384), .C(new_n10386), .Y(new_n10603));
  AOI22xp33_ASAP7_75t_L     g10347(.A1(new_n6376), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n6648), .Y(new_n10604));
  OAI221xp5_ASAP7_75t_L     g10348(.A1(new_n6646), .A2(new_n942), .B1(new_n6636), .B2(new_n1035), .C(new_n10604), .Y(new_n10605));
  XNOR2x2_ASAP7_75t_L       g10349(.A(\a[47] ), .B(new_n10605), .Y(new_n10606));
  INVx1_ASAP7_75t_L         g10350(.A(new_n10606), .Y(new_n10607));
  A2O1A1O1Ixp25_ASAP7_75t_L g10351(.A1(new_n10054), .A2(new_n10006), .B(new_n10321), .C(new_n10377), .D(new_n10374), .Y(new_n10608));
  OAI211xp5_ASAP7_75t_L     g10352(.A1(new_n10346), .A2(new_n10352), .B(new_n10342), .C(new_n10341), .Y(new_n10609));
  A2O1A1Ixp33_ASAP7_75t_L   g10353(.A1(new_n10353), .A2(new_n10349), .B(new_n10355), .C(new_n10609), .Y(new_n10610));
  AOI22xp33_ASAP7_75t_L     g10354(.A1(new_n8831), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n9115), .Y(new_n10611));
  OAI221xp5_ASAP7_75t_L     g10355(.A1(new_n10343), .A2(new_n418), .B1(new_n10016), .B2(new_n425), .C(new_n10611), .Y(new_n10612));
  XNOR2x2_ASAP7_75t_L       g10356(.A(new_n8826), .B(new_n10612), .Y(new_n10613));
  NOR3xp33_ASAP7_75t_L      g10357(.A(new_n10029), .B(new_n10336), .C(new_n10328), .Y(new_n10614));
  INVx1_ASAP7_75t_L         g10358(.A(new_n10614), .Y(new_n10615));
  A2O1A1Ixp33_ASAP7_75t_L   g10359(.A1(new_n10337), .A2(new_n10334), .B(new_n10340), .C(new_n10615), .Y(new_n10616));
  OAI22xp33_ASAP7_75t_L     g10360(.A1(new_n10026), .A2(new_n276), .B1(new_n324), .B2(new_n9699), .Y(new_n10617));
  AOI221xp5_ASAP7_75t_L     g10361(.A1(new_n9703), .A2(\b[3] ), .B1(new_n9697), .B2(new_n329), .C(new_n10617), .Y(new_n10618));
  NAND2xp33_ASAP7_75t_L     g10362(.A(\a[59] ), .B(new_n10618), .Y(new_n10619));
  AO21x2_ASAP7_75t_L        g10363(.A1(new_n329), .A2(new_n9697), .B(new_n10617), .Y(new_n10620));
  A2O1A1Ixp33_ASAP7_75t_L   g10364(.A1(\b[3] ), .A2(new_n9703), .B(new_n10620), .C(new_n9693), .Y(new_n10621));
  INVx1_ASAP7_75t_L         g10365(.A(\a[62] ), .Y(new_n10622));
  NOR2xp33_ASAP7_75t_L      g10366(.A(new_n10622), .B(new_n10336), .Y(new_n10623));
  NAND2xp33_ASAP7_75t_L     g10367(.A(new_n10331), .B(new_n10330), .Y(new_n10624));
  INVx1_ASAP7_75t_L         g10368(.A(\a[61] ), .Y(new_n10625));
  NAND2xp33_ASAP7_75t_L     g10369(.A(\a[62] ), .B(new_n10625), .Y(new_n10626));
  NAND2xp33_ASAP7_75t_L     g10370(.A(\a[61] ), .B(new_n10622), .Y(new_n10627));
  NAND2xp33_ASAP7_75t_L     g10371(.A(new_n10627), .B(new_n10626), .Y(new_n10628));
  NAND2xp33_ASAP7_75t_L     g10372(.A(new_n10628), .B(new_n10624), .Y(new_n10629));
  NAND3xp33_ASAP7_75t_L     g10373(.A(new_n10624), .B(new_n10626), .C(new_n10627), .Y(new_n10630));
  XNOR2x2_ASAP7_75t_L       g10374(.A(\a[61] ), .B(\a[60] ), .Y(new_n10631));
  NOR2xp33_ASAP7_75t_L      g10375(.A(new_n10631), .B(new_n10624), .Y(new_n10632));
  NAND2xp33_ASAP7_75t_L     g10376(.A(\b[0] ), .B(new_n10632), .Y(new_n10633));
  OAI221xp5_ASAP7_75t_L     g10377(.A1(new_n10629), .A2(new_n270), .B1(new_n261), .B2(new_n10630), .C(new_n10633), .Y(new_n10634));
  XNOR2x2_ASAP7_75t_L       g10378(.A(new_n10623), .B(new_n10634), .Y(new_n10635));
  NAND3xp33_ASAP7_75t_L     g10379(.A(new_n10621), .B(new_n10635), .C(new_n10619), .Y(new_n10636));
  AOI21xp33_ASAP7_75t_L     g10380(.A1(new_n10621), .A2(new_n10619), .B(new_n10635), .Y(new_n10637));
  INVx1_ASAP7_75t_L         g10381(.A(new_n10637), .Y(new_n10638));
  NAND3xp33_ASAP7_75t_L     g10382(.A(new_n10616), .B(new_n10636), .C(new_n10638), .Y(new_n10639));
  INVx1_ASAP7_75t_L         g10383(.A(new_n10636), .Y(new_n10640));
  OAI211xp5_ASAP7_75t_L     g10384(.A1(new_n10640), .A2(new_n10637), .B(new_n10341), .C(new_n10615), .Y(new_n10641));
  AOI21xp33_ASAP7_75t_L     g10385(.A1(new_n10639), .A2(new_n10641), .B(new_n10613), .Y(new_n10642));
  INVx1_ASAP7_75t_L         g10386(.A(new_n10642), .Y(new_n10643));
  NAND3xp33_ASAP7_75t_L     g10387(.A(new_n10639), .B(new_n10641), .C(new_n10613), .Y(new_n10644));
  NAND3xp33_ASAP7_75t_L     g10388(.A(new_n10610), .B(new_n10643), .C(new_n10644), .Y(new_n10645));
  NAND2xp33_ASAP7_75t_L     g10389(.A(new_n10354), .B(new_n10357), .Y(new_n10646));
  INVx1_ASAP7_75t_L         g10390(.A(new_n10644), .Y(new_n10647));
  OAI211xp5_ASAP7_75t_L     g10391(.A1(new_n10642), .A2(new_n10647), .B(new_n10646), .C(new_n10609), .Y(new_n10648));
  AOI22xp33_ASAP7_75t_L     g10392(.A1(new_n7960), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n8537), .Y(new_n10649));
  OAI221xp5_ASAP7_75t_L     g10393(.A1(new_n8817), .A2(new_n540), .B1(new_n7957), .B2(new_n624), .C(new_n10649), .Y(new_n10650));
  XNOR2x2_ASAP7_75t_L       g10394(.A(\a[53] ), .B(new_n10650), .Y(new_n10651));
  NAND3xp33_ASAP7_75t_L     g10395(.A(new_n10648), .B(new_n10645), .C(new_n10651), .Y(new_n10652));
  AO21x2_ASAP7_75t_L        g10396(.A1(new_n10645), .A2(new_n10648), .B(new_n10651), .Y(new_n10653));
  AOI21xp33_ASAP7_75t_L     g10397(.A1(new_n10365), .A2(new_n10364), .B(new_n10366), .Y(new_n10654));
  A2O1A1O1Ixp25_ASAP7_75t_L g10398(.A1(new_n10051), .A2(new_n10050), .B(new_n10046), .C(new_n10367), .D(new_n10654), .Y(new_n10655));
  NAND3xp33_ASAP7_75t_L     g10399(.A(new_n10653), .B(new_n10655), .C(new_n10652), .Y(new_n10656));
  AO21x2_ASAP7_75t_L        g10400(.A1(new_n10652), .A2(new_n10653), .B(new_n10655), .Y(new_n10657));
  AOI22xp33_ASAP7_75t_L     g10401(.A1(new_n7111), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n7391), .Y(new_n10658));
  OAI221xp5_ASAP7_75t_L     g10402(.A1(new_n8558), .A2(new_n760), .B1(new_n8237), .B2(new_n790), .C(new_n10658), .Y(new_n10659));
  XNOR2x2_ASAP7_75t_L       g10403(.A(\a[50] ), .B(new_n10659), .Y(new_n10660));
  INVx1_ASAP7_75t_L         g10404(.A(new_n10660), .Y(new_n10661));
  AOI21xp33_ASAP7_75t_L     g10405(.A1(new_n10657), .A2(new_n10656), .B(new_n10661), .Y(new_n10662));
  NAND3xp33_ASAP7_75t_L     g10406(.A(new_n10657), .B(new_n10656), .C(new_n10661), .Y(new_n10663));
  INVx1_ASAP7_75t_L         g10407(.A(new_n10663), .Y(new_n10664));
  OAI21xp33_ASAP7_75t_L     g10408(.A1(new_n10662), .A2(new_n10664), .B(new_n10608), .Y(new_n10665));
  A2O1A1Ixp33_ASAP7_75t_L   g10409(.A1(new_n10059), .A2(new_n10058), .B(new_n10371), .C(new_n10378), .Y(new_n10666));
  INVx1_ASAP7_75t_L         g10410(.A(new_n10662), .Y(new_n10667));
  NAND3xp33_ASAP7_75t_L     g10411(.A(new_n10666), .B(new_n10667), .C(new_n10663), .Y(new_n10668));
  NAND3xp33_ASAP7_75t_L     g10412(.A(new_n10668), .B(new_n10665), .C(new_n10607), .Y(new_n10669));
  AOI21xp33_ASAP7_75t_L     g10413(.A1(new_n10663), .A2(new_n10667), .B(new_n10666), .Y(new_n10670));
  NOR3xp33_ASAP7_75t_L      g10414(.A(new_n10608), .B(new_n10664), .C(new_n10662), .Y(new_n10671));
  OAI21xp33_ASAP7_75t_L     g10415(.A1(new_n10671), .A2(new_n10670), .B(new_n10606), .Y(new_n10672));
  AOI21xp33_ASAP7_75t_L     g10416(.A1(new_n10672), .A2(new_n10669), .B(new_n10603), .Y(new_n10673));
  O2A1O1Ixp33_ASAP7_75t_L   g10417(.A1(new_n10315), .A2(new_n10070), .B(new_n10387), .C(new_n10380), .Y(new_n10674));
  NAND2xp33_ASAP7_75t_L     g10418(.A(new_n10669), .B(new_n10672), .Y(new_n10675));
  NOR2xp33_ASAP7_75t_L      g10419(.A(new_n10674), .B(new_n10675), .Y(new_n10676));
  AOI22xp33_ASAP7_75t_L     g10420(.A1(new_n5624), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n5901), .Y(new_n10677));
  OAI221xp5_ASAP7_75t_L     g10421(.A1(new_n5900), .A2(new_n1313), .B1(new_n5892), .B2(new_n1438), .C(new_n10677), .Y(new_n10678));
  XNOR2x2_ASAP7_75t_L       g10422(.A(\a[44] ), .B(new_n10678), .Y(new_n10679));
  OAI21xp33_ASAP7_75t_L     g10423(.A1(new_n10673), .A2(new_n10676), .B(new_n10679), .Y(new_n10680));
  NAND2xp33_ASAP7_75t_L     g10424(.A(new_n10674), .B(new_n10675), .Y(new_n10681));
  NAND3xp33_ASAP7_75t_L     g10425(.A(new_n10603), .B(new_n10669), .C(new_n10672), .Y(new_n10682));
  INVx1_ASAP7_75t_L         g10426(.A(new_n10679), .Y(new_n10683));
  NAND3xp33_ASAP7_75t_L     g10427(.A(new_n10681), .B(new_n10682), .C(new_n10683), .Y(new_n10684));
  NAND2xp33_ASAP7_75t_L     g10428(.A(new_n10684), .B(new_n10680), .Y(new_n10685));
  NAND2xp33_ASAP7_75t_L     g10429(.A(new_n10602), .B(new_n10685), .Y(new_n10686));
  A2O1A1O1Ixp25_ASAP7_75t_L g10430(.A1(new_n9763), .A2(new_n9764), .B(new_n9997), .C(new_n10080), .D(new_n10310), .Y(new_n10687));
  INVx1_ASAP7_75t_L         g10431(.A(new_n10601), .Y(new_n10688));
  A2O1A1Ixp33_ASAP7_75t_L   g10432(.A1(new_n10389), .A2(new_n10392), .B(new_n10687), .C(new_n10688), .Y(new_n10689));
  NAND3xp33_ASAP7_75t_L     g10433(.A(new_n10689), .B(new_n10680), .C(new_n10684), .Y(new_n10690));
  NAND3xp33_ASAP7_75t_L     g10434(.A(new_n10690), .B(new_n10686), .C(new_n10600), .Y(new_n10691));
  AOI21xp33_ASAP7_75t_L     g10435(.A1(new_n10684), .A2(new_n10680), .B(new_n10689), .Y(new_n10692));
  O2A1O1Ixp33_ASAP7_75t_L   g10436(.A1(new_n10687), .A2(new_n10402), .B(new_n10688), .C(new_n10685), .Y(new_n10693));
  OAI21xp33_ASAP7_75t_L     g10437(.A1(new_n10692), .A2(new_n10693), .B(new_n10599), .Y(new_n10694));
  NAND2xp33_ASAP7_75t_L     g10438(.A(new_n10691), .B(new_n10694), .Y(new_n10695));
  NAND2xp33_ASAP7_75t_L     g10439(.A(new_n10695), .B(new_n10596), .Y(new_n10696));
  AOI21xp33_ASAP7_75t_L     g10440(.A1(new_n10398), .A2(new_n10394), .B(new_n10308), .Y(new_n10697));
  A2O1A1Ixp33_ASAP7_75t_L   g10441(.A1(new_n10091), .A2(new_n10084), .B(new_n10697), .C(new_n10399), .Y(new_n10698));
  NAND3xp33_ASAP7_75t_L     g10442(.A(new_n10698), .B(new_n10691), .C(new_n10694), .Y(new_n10699));
  AOI22xp33_ASAP7_75t_L     g10443(.A1(new_n4283), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n4512), .Y(new_n10700));
  OAI221xp5_ASAP7_75t_L     g10444(.A1(new_n4277), .A2(new_n1929), .B1(new_n4499), .B2(new_n2075), .C(new_n10700), .Y(new_n10701));
  XNOR2x2_ASAP7_75t_L       g10445(.A(\a[38] ), .B(new_n10701), .Y(new_n10702));
  NAND3xp33_ASAP7_75t_L     g10446(.A(new_n10696), .B(new_n10699), .C(new_n10702), .Y(new_n10703));
  AO21x2_ASAP7_75t_L        g10447(.A1(new_n10699), .A2(new_n10696), .B(new_n10702), .Y(new_n10704));
  NAND3xp33_ASAP7_75t_L     g10448(.A(new_n10408), .B(new_n10405), .C(new_n10415), .Y(new_n10705));
  NAND4xp25_ASAP7_75t_L     g10449(.A(new_n10422), .B(new_n10705), .C(new_n10704), .D(new_n10703), .Y(new_n10706));
  AND3x1_ASAP7_75t_L        g10450(.A(new_n10696), .B(new_n10702), .C(new_n10699), .Y(new_n10707));
  AOI21xp33_ASAP7_75t_L     g10451(.A1(new_n10696), .A2(new_n10699), .B(new_n10702), .Y(new_n10708));
  A2O1A1Ixp33_ASAP7_75t_L   g10452(.A1(new_n10416), .A2(new_n10412), .B(new_n10417), .C(new_n10705), .Y(new_n10709));
  OAI21xp33_ASAP7_75t_L     g10453(.A1(new_n10708), .A2(new_n10707), .B(new_n10709), .Y(new_n10710));
  AOI22xp33_ASAP7_75t_L     g10454(.A1(new_n3633), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n3858), .Y(new_n10711));
  OAI221xp5_ASAP7_75t_L     g10455(.A1(new_n3853), .A2(new_n2497), .B1(new_n3856), .B2(new_n2672), .C(new_n10711), .Y(new_n10712));
  XNOR2x2_ASAP7_75t_L       g10456(.A(\a[35] ), .B(new_n10712), .Y(new_n10713));
  NAND3xp33_ASAP7_75t_L     g10457(.A(new_n10706), .B(new_n10710), .C(new_n10713), .Y(new_n10714));
  NOR3xp33_ASAP7_75t_L      g10458(.A(new_n10709), .B(new_n10707), .C(new_n10708), .Y(new_n10715));
  AOI22xp33_ASAP7_75t_L     g10459(.A1(new_n10703), .A2(new_n10704), .B1(new_n10705), .B2(new_n10422), .Y(new_n10716));
  INVx1_ASAP7_75t_L         g10460(.A(new_n10713), .Y(new_n10717));
  OAI21xp33_ASAP7_75t_L     g10461(.A1(new_n10716), .A2(new_n10715), .B(new_n10717), .Y(new_n10718));
  NAND2xp33_ASAP7_75t_L     g10462(.A(new_n10714), .B(new_n10718), .Y(new_n10719));
  NOR3xp33_ASAP7_75t_L      g10463(.A(new_n10432), .B(new_n10430), .C(new_n10433), .Y(new_n10720));
  INVx1_ASAP7_75t_L         g10464(.A(new_n10720), .Y(new_n10721));
  A2O1A1Ixp33_ASAP7_75t_L   g10465(.A1(new_n10121), .A2(new_n10436), .B(new_n10442), .C(new_n10721), .Y(new_n10722));
  NOR2xp33_ASAP7_75t_L      g10466(.A(new_n10719), .B(new_n10722), .Y(new_n10723));
  O2A1O1Ixp33_ASAP7_75t_L   g10467(.A1(new_n10440), .A2(new_n10441), .B(new_n10437), .C(new_n10720), .Y(new_n10724));
  AOI21xp33_ASAP7_75t_L     g10468(.A1(new_n10718), .A2(new_n10714), .B(new_n10724), .Y(new_n10725));
  AOI22xp33_ASAP7_75t_L     g10469(.A1(new_n3029), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n3258), .Y(new_n10726));
  OAI221xp5_ASAP7_75t_L     g10470(.A1(new_n3024), .A2(new_n2982), .B1(new_n3256), .B2(new_n3187), .C(new_n10726), .Y(new_n10727));
  XNOR2x2_ASAP7_75t_L       g10471(.A(\a[32] ), .B(new_n10727), .Y(new_n10728));
  INVx1_ASAP7_75t_L         g10472(.A(new_n10728), .Y(new_n10729));
  NOR3xp33_ASAP7_75t_L      g10473(.A(new_n10723), .B(new_n10725), .C(new_n10729), .Y(new_n10730));
  NAND3xp33_ASAP7_75t_L     g10474(.A(new_n10724), .B(new_n10718), .C(new_n10714), .Y(new_n10731));
  A2O1A1Ixp33_ASAP7_75t_L   g10475(.A1(new_n10435), .A2(new_n10437), .B(new_n10720), .C(new_n10719), .Y(new_n10732));
  AOI21xp33_ASAP7_75t_L     g10476(.A1(new_n10731), .A2(new_n10732), .B(new_n10728), .Y(new_n10733));
  NOR3xp33_ASAP7_75t_L      g10477(.A(new_n10594), .B(new_n10730), .C(new_n10733), .Y(new_n10734));
  OAI31xp33_ASAP7_75t_L     g10478(.A1(new_n10458), .A2(new_n10455), .A3(new_n10454), .B(new_n10451), .Y(new_n10735));
  NAND3xp33_ASAP7_75t_L     g10479(.A(new_n10731), .B(new_n10732), .C(new_n10728), .Y(new_n10736));
  OAI21xp33_ASAP7_75t_L     g10480(.A1(new_n10725), .A2(new_n10723), .B(new_n10729), .Y(new_n10737));
  AOI21xp33_ASAP7_75t_L     g10481(.A1(new_n10737), .A2(new_n10736), .B(new_n10735), .Y(new_n10738));
  AOI22xp33_ASAP7_75t_L     g10482(.A1(new_n2552), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n2736), .Y(new_n10739));
  OAI221xp5_ASAP7_75t_L     g10483(.A1(new_n2547), .A2(new_n3565), .B1(new_n2734), .B2(new_n3591), .C(new_n10739), .Y(new_n10740));
  XNOR2x2_ASAP7_75t_L       g10484(.A(\a[29] ), .B(new_n10740), .Y(new_n10741));
  INVx1_ASAP7_75t_L         g10485(.A(new_n10741), .Y(new_n10742));
  OAI21xp33_ASAP7_75t_L     g10486(.A1(new_n10738), .A2(new_n10734), .B(new_n10742), .Y(new_n10743));
  NAND3xp33_ASAP7_75t_L     g10487(.A(new_n10735), .B(new_n10736), .C(new_n10737), .Y(new_n10744));
  OAI21xp33_ASAP7_75t_L     g10488(.A1(new_n10733), .A2(new_n10730), .B(new_n10594), .Y(new_n10745));
  NAND3xp33_ASAP7_75t_L     g10489(.A(new_n10744), .B(new_n10741), .C(new_n10745), .Y(new_n10746));
  AOI21xp33_ASAP7_75t_L     g10490(.A1(new_n10746), .A2(new_n10743), .B(new_n10593), .Y(new_n10747));
  AND2x2_ASAP7_75t_L        g10491(.A(new_n10468), .B(new_n10472), .Y(new_n10748));
  NAND2xp33_ASAP7_75t_L     g10492(.A(new_n10746), .B(new_n10743), .Y(new_n10749));
  O2A1O1Ixp33_ASAP7_75t_L   g10493(.A1(new_n10475), .A2(new_n10748), .B(new_n10592), .C(new_n10749), .Y(new_n10750));
  AOI22xp33_ASAP7_75t_L     g10494(.A1(new_n2114), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n2259), .Y(new_n10751));
  OAI221xp5_ASAP7_75t_L     g10495(.A1(new_n2109), .A2(new_n4216), .B1(new_n2257), .B2(new_n4431), .C(new_n10751), .Y(new_n10752));
  XNOR2x2_ASAP7_75t_L       g10496(.A(\a[26] ), .B(new_n10752), .Y(new_n10753));
  INVx1_ASAP7_75t_L         g10497(.A(new_n10753), .Y(new_n10754));
  NOR3xp33_ASAP7_75t_L      g10498(.A(new_n10750), .B(new_n10754), .C(new_n10747), .Y(new_n10755));
  AOI21xp33_ASAP7_75t_L     g10499(.A1(new_n10744), .A2(new_n10745), .B(new_n10741), .Y(new_n10756));
  NOR3xp33_ASAP7_75t_L      g10500(.A(new_n10734), .B(new_n10738), .C(new_n10742), .Y(new_n10757));
  OAI221xp5_ASAP7_75t_L     g10501(.A1(new_n10757), .A2(new_n10756), .B1(new_n10475), .B2(new_n10748), .C(new_n10592), .Y(new_n10758));
  NAND3xp33_ASAP7_75t_L     g10502(.A(new_n10593), .B(new_n10743), .C(new_n10746), .Y(new_n10759));
  AOI21xp33_ASAP7_75t_L     g10503(.A1(new_n10759), .A2(new_n10758), .B(new_n10753), .Y(new_n10760));
  NOR2xp33_ASAP7_75t_L      g10504(.A(new_n10760), .B(new_n10755), .Y(new_n10761));
  INVx1_ASAP7_75t_L         g10505(.A(new_n10477), .Y(new_n10762));
  A2O1A1O1Ixp25_ASAP7_75t_L g10506(.A1(new_n10143), .A2(new_n10145), .B(new_n10297), .C(new_n10480), .D(new_n10762), .Y(new_n10763));
  NAND2xp33_ASAP7_75t_L     g10507(.A(new_n10763), .B(new_n10761), .Y(new_n10764));
  NAND3xp33_ASAP7_75t_L     g10508(.A(new_n10759), .B(new_n10758), .C(new_n10753), .Y(new_n10765));
  OAI21xp33_ASAP7_75t_L     g10509(.A1(new_n10747), .A2(new_n10750), .B(new_n10754), .Y(new_n10766));
  NAND2xp33_ASAP7_75t_L     g10510(.A(new_n10765), .B(new_n10766), .Y(new_n10767));
  A2O1A1Ixp33_ASAP7_75t_L   g10511(.A1(new_n10483), .A2(new_n10492), .B(new_n10762), .C(new_n10767), .Y(new_n10768));
  NOR2xp33_ASAP7_75t_L      g10512(.A(new_n4848), .B(new_n1699), .Y(new_n10769));
  INVx1_ASAP7_75t_L         g10513(.A(new_n10769), .Y(new_n10770));
  NAND2xp33_ASAP7_75t_L     g10514(.A(new_n1695), .B(new_n4876), .Y(new_n10771));
  AOI22xp33_ASAP7_75t_L     g10515(.A1(new_n1704), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n1837), .Y(new_n10772));
  AND4x1_ASAP7_75t_L        g10516(.A(new_n10772), .B(new_n10771), .C(new_n10770), .D(\a[23] ), .Y(new_n10773));
  AOI31xp33_ASAP7_75t_L     g10517(.A1(new_n10771), .A2(new_n10770), .A3(new_n10772), .B(\a[23] ), .Y(new_n10774));
  NOR2xp33_ASAP7_75t_L      g10518(.A(new_n10774), .B(new_n10773), .Y(new_n10775));
  NAND3xp33_ASAP7_75t_L     g10519(.A(new_n10768), .B(new_n10764), .C(new_n10775), .Y(new_n10776));
  NOR3xp33_ASAP7_75t_L      g10520(.A(new_n10494), .B(new_n10767), .C(new_n10762), .Y(new_n10777));
  NOR2xp33_ASAP7_75t_L      g10521(.A(new_n10763), .B(new_n10761), .Y(new_n10778));
  INVx1_ASAP7_75t_L         g10522(.A(new_n10775), .Y(new_n10779));
  OAI21xp33_ASAP7_75t_L     g10523(.A1(new_n10778), .A2(new_n10777), .B(new_n10779), .Y(new_n10780));
  NAND2xp33_ASAP7_75t_L     g10524(.A(new_n10776), .B(new_n10780), .Y(new_n10781));
  OAI211xp5_ASAP7_75t_L     g10525(.A1(new_n10487), .A2(new_n10488), .B(new_n10484), .C(new_n10482), .Y(new_n10782));
  A2O1A1Ixp33_ASAP7_75t_L   g10526(.A1(new_n10495), .A2(new_n10490), .B(new_n10497), .C(new_n10782), .Y(new_n10783));
  NOR2xp33_ASAP7_75t_L      g10527(.A(new_n10783), .B(new_n10781), .Y(new_n10784));
  NOR3xp33_ASAP7_75t_L      g10528(.A(new_n10777), .B(new_n10779), .C(new_n10778), .Y(new_n10785));
  AOI21xp33_ASAP7_75t_L     g10529(.A1(new_n10768), .A2(new_n10764), .B(new_n10775), .Y(new_n10786));
  NOR2xp33_ASAP7_75t_L      g10530(.A(new_n10786), .B(new_n10785), .Y(new_n10787));
  A2O1A1O1Ixp25_ASAP7_75t_L g10531(.A1(new_n10495), .A2(new_n10490), .B(new_n10497), .C(new_n10782), .D(new_n10787), .Y(new_n10788));
  AOI22xp33_ASAP7_75t_L     g10532(.A1(new_n1360), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n1581), .Y(new_n10789));
  INVx1_ASAP7_75t_L         g10533(.A(new_n10789), .Y(new_n10790));
  AOI221xp5_ASAP7_75t_L     g10534(.A1(\b[42] ), .A2(new_n1362), .B1(new_n1365), .B2(new_n5812), .C(new_n10790), .Y(new_n10791));
  XNOR2x2_ASAP7_75t_L       g10535(.A(new_n1356), .B(new_n10791), .Y(new_n10792));
  OAI21xp33_ASAP7_75t_L     g10536(.A1(new_n10784), .A2(new_n10788), .B(new_n10792), .Y(new_n10793));
  NAND3xp33_ASAP7_75t_L     g10537(.A(new_n10787), .B(new_n10499), .C(new_n10782), .Y(new_n10794));
  NAND2xp33_ASAP7_75t_L     g10538(.A(new_n10783), .B(new_n10781), .Y(new_n10795));
  INVx1_ASAP7_75t_L         g10539(.A(new_n10792), .Y(new_n10796));
  NAND3xp33_ASAP7_75t_L     g10540(.A(new_n10794), .B(new_n10796), .C(new_n10795), .Y(new_n10797));
  AOI21xp33_ASAP7_75t_L     g10541(.A1(new_n10793), .A2(new_n10797), .B(new_n10591), .Y(new_n10798));
  AOI31xp33_ASAP7_75t_L     g10542(.A1(new_n10518), .A2(new_n10516), .A3(new_n10162), .B(new_n10513), .Y(new_n10799));
  AOI21xp33_ASAP7_75t_L     g10543(.A1(new_n10794), .A2(new_n10795), .B(new_n10796), .Y(new_n10800));
  NOR3xp33_ASAP7_75t_L      g10544(.A(new_n10788), .B(new_n10792), .C(new_n10784), .Y(new_n10801));
  NOR3xp33_ASAP7_75t_L      g10545(.A(new_n10799), .B(new_n10800), .C(new_n10801), .Y(new_n10802));
  OAI21xp33_ASAP7_75t_L     g10546(.A1(new_n10798), .A2(new_n10802), .B(new_n10590), .Y(new_n10803));
  INVx1_ASAP7_75t_L         g10547(.A(new_n10590), .Y(new_n10804));
  OAI21xp33_ASAP7_75t_L     g10548(.A1(new_n10800), .A2(new_n10801), .B(new_n10799), .Y(new_n10805));
  NAND3xp33_ASAP7_75t_L     g10549(.A(new_n10591), .B(new_n10793), .C(new_n10797), .Y(new_n10806));
  NAND3xp33_ASAP7_75t_L     g10550(.A(new_n10806), .B(new_n10805), .C(new_n10804), .Y(new_n10807));
  NAND2xp33_ASAP7_75t_L     g10551(.A(new_n10807), .B(new_n10803), .Y(new_n10808));
  NOR2xp33_ASAP7_75t_L      g10552(.A(new_n10587), .B(new_n10808), .Y(new_n10809));
  INVx1_ASAP7_75t_L         g10553(.A(new_n10586), .Y(new_n10810));
  A2O1A1Ixp33_ASAP7_75t_L   g10554(.A1(new_n10520), .A2(new_n10523), .B(new_n10288), .C(new_n10810), .Y(new_n10811));
  AOI21xp33_ASAP7_75t_L     g10555(.A1(new_n10807), .A2(new_n10803), .B(new_n10811), .Y(new_n10812));
  OAI21xp33_ASAP7_75t_L     g10556(.A1(new_n10812), .A2(new_n10809), .B(new_n10585), .Y(new_n10813));
  NAND3xp33_ASAP7_75t_L     g10557(.A(new_n10811), .B(new_n10803), .C(new_n10807), .Y(new_n10814));
  NAND2xp33_ASAP7_75t_L     g10558(.A(new_n10587), .B(new_n10808), .Y(new_n10815));
  OAI211xp5_ASAP7_75t_L     g10559(.A1(new_n10583), .A2(new_n10584), .B(new_n10815), .C(new_n10814), .Y(new_n10816));
  NAND3xp33_ASAP7_75t_L     g10560(.A(new_n10580), .B(new_n10813), .C(new_n10816), .Y(new_n10817));
  AOI21xp33_ASAP7_75t_L     g10561(.A1(new_n10532), .A2(new_n10283), .B(new_n10578), .Y(new_n10818));
  NAND2xp33_ASAP7_75t_L     g10562(.A(new_n10813), .B(new_n10816), .Y(new_n10819));
  NAND2xp33_ASAP7_75t_L     g10563(.A(new_n10818), .B(new_n10819), .Y(new_n10820));
  AOI21xp33_ASAP7_75t_L     g10564(.A1(new_n10820), .A2(new_n10817), .B(new_n10577), .Y(new_n10821));
  NOR2xp33_ASAP7_75t_L      g10565(.A(new_n10818), .B(new_n10819), .Y(new_n10822));
  AOI21xp33_ASAP7_75t_L     g10566(.A1(new_n10816), .A2(new_n10813), .B(new_n10580), .Y(new_n10823));
  NOR3xp33_ASAP7_75t_L      g10567(.A(new_n10822), .B(new_n10823), .C(new_n10576), .Y(new_n10824));
  NOR2xp33_ASAP7_75t_L      g10568(.A(new_n10821), .B(new_n10824), .Y(new_n10825));
  A2O1A1Ixp33_ASAP7_75t_L   g10569(.A1(new_n10547), .A2(new_n10544), .B(new_n10573), .C(new_n10825), .Y(new_n10826));
  O2A1O1Ixp33_ASAP7_75t_L   g10570(.A1(new_n10537), .A2(new_n10541), .B(new_n10544), .C(new_n10573), .Y(new_n10827));
  OAI21xp33_ASAP7_75t_L     g10571(.A1(new_n10821), .A2(new_n10824), .B(new_n10827), .Y(new_n10828));
  AOI22xp33_ASAP7_75t_L     g10572(.A1(new_n444), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n471), .Y(new_n10829));
  OAI221xp5_ASAP7_75t_L     g10573(.A1(new_n468), .A2(new_n8458), .B1(new_n469), .B2(new_n8768), .C(new_n10829), .Y(new_n10830));
  XNOR2x2_ASAP7_75t_L       g10574(.A(\a[8] ), .B(new_n10830), .Y(new_n10831));
  NAND3xp33_ASAP7_75t_L     g10575(.A(new_n10826), .B(new_n10828), .C(new_n10831), .Y(new_n10832));
  AO21x2_ASAP7_75t_L        g10576(.A1(new_n10828), .A2(new_n10826), .B(new_n10831), .Y(new_n10833));
  AOI21xp33_ASAP7_75t_L     g10577(.A1(new_n10269), .A2(new_n10550), .B(new_n10552), .Y(new_n10834));
  AND3x1_ASAP7_75t_L        g10578(.A(new_n10834), .B(new_n10832), .C(new_n10833), .Y(new_n10835));
  AOI21xp33_ASAP7_75t_L     g10579(.A1(new_n10832), .A2(new_n10833), .B(new_n10834), .Y(new_n10836));
  AOI22xp33_ASAP7_75t_L     g10580(.A1(new_n344), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n370), .Y(new_n10837));
  OAI221xp5_ASAP7_75t_L     g10581(.A1(new_n429), .A2(new_n9620), .B1(new_n366), .B2(new_n9925), .C(new_n10837), .Y(new_n10838));
  XNOR2x2_ASAP7_75t_L       g10582(.A(\a[5] ), .B(new_n10838), .Y(new_n10839));
  OAI21xp33_ASAP7_75t_L     g10583(.A1(new_n10836), .A2(new_n10835), .B(new_n10839), .Y(new_n10840));
  NAND3xp33_ASAP7_75t_L     g10584(.A(new_n10834), .B(new_n10832), .C(new_n10833), .Y(new_n10841));
  NAND2xp33_ASAP7_75t_L     g10585(.A(new_n10832), .B(new_n10833), .Y(new_n10842));
  A2O1A1Ixp33_ASAP7_75t_L   g10586(.A1(new_n10550), .A2(new_n10269), .B(new_n10552), .C(new_n10842), .Y(new_n10843));
  INVx1_ASAP7_75t_L         g10587(.A(new_n10839), .Y(new_n10844));
  NAND3xp33_ASAP7_75t_L     g10588(.A(new_n10843), .B(new_n10841), .C(new_n10844), .Y(new_n10845));
  NOR2xp33_ASAP7_75t_L      g10589(.A(\b[60] ), .B(\b[61] ), .Y(new_n10846));
  INVx1_ASAP7_75t_L         g10590(.A(\b[61] ), .Y(new_n10847));
  NOR2xp33_ASAP7_75t_L      g10591(.A(new_n10250), .B(new_n10847), .Y(new_n10848));
  NOR2xp33_ASAP7_75t_L      g10592(.A(new_n10846), .B(new_n10848), .Y(new_n10849));
  A2O1A1Ixp33_ASAP7_75t_L   g10593(.A1(new_n10256), .A2(new_n10252), .B(new_n10251), .C(new_n10849), .Y(new_n10850));
  A2O1A1O1Ixp25_ASAP7_75t_L g10594(.A1(new_n9944), .A2(new_n9625), .B(new_n9919), .C(new_n10255), .D(new_n9952), .Y(new_n10851));
  O2A1O1Ixp33_ASAP7_75t_L   g10595(.A1(new_n9948), .A2(new_n10851), .B(new_n10252), .C(new_n10251), .Y(new_n10852));
  INVx1_ASAP7_75t_L         g10596(.A(new_n10849), .Y(new_n10853));
  NAND2xp33_ASAP7_75t_L     g10597(.A(new_n10853), .B(new_n10852), .Y(new_n10854));
  NAND2xp33_ASAP7_75t_L     g10598(.A(new_n10850), .B(new_n10854), .Y(new_n10855));
  AOI22xp33_ASAP7_75t_L     g10599(.A1(\b[59] ), .A2(new_n282), .B1(\b[61] ), .B2(new_n303), .Y(new_n10856));
  OAI221xp5_ASAP7_75t_L     g10600(.A1(new_n291), .A2(new_n10250), .B1(new_n268), .B2(new_n10855), .C(new_n10856), .Y(new_n10857));
  XNOR2x2_ASAP7_75t_L       g10601(.A(\a[2] ), .B(new_n10857), .Y(new_n10858));
  NAND3xp33_ASAP7_75t_L     g10602(.A(new_n10845), .B(new_n10840), .C(new_n10858), .Y(new_n10859));
  AOI21xp33_ASAP7_75t_L     g10603(.A1(new_n10843), .A2(new_n10841), .B(new_n10844), .Y(new_n10860));
  NOR3xp33_ASAP7_75t_L      g10604(.A(new_n10835), .B(new_n10836), .C(new_n10839), .Y(new_n10861));
  INVx1_ASAP7_75t_L         g10605(.A(new_n10858), .Y(new_n10862));
  OAI21xp33_ASAP7_75t_L     g10606(.A1(new_n10861), .A2(new_n10860), .B(new_n10862), .Y(new_n10863));
  A2O1A1Ixp33_ASAP7_75t_L   g10607(.A1(new_n10261), .A2(new_n10263), .B(new_n10560), .C(new_n10555), .Y(new_n10864));
  INVx1_ASAP7_75t_L         g10608(.A(new_n10864), .Y(new_n10865));
  NAND3xp33_ASAP7_75t_L     g10609(.A(new_n10863), .B(new_n10859), .C(new_n10865), .Y(new_n10866));
  INVx1_ASAP7_75t_L         g10610(.A(new_n10866), .Y(new_n10867));
  AOI21xp33_ASAP7_75t_L     g10611(.A1(new_n10863), .A2(new_n10859), .B(new_n10865), .Y(new_n10868));
  NOR2xp33_ASAP7_75t_L      g10612(.A(new_n10868), .B(new_n10867), .Y(new_n10869));
  A2O1A1Ixp33_ASAP7_75t_L   g10613(.A1(new_n10565), .A2(new_n10569), .B(new_n10572), .C(new_n10869), .Y(new_n10870));
  INVx1_ASAP7_75t_L         g10614(.A(new_n10870), .Y(new_n10871));
  A2O1A1Ixp33_ASAP7_75t_L   g10615(.A1(new_n10236), .A2(new_n10246), .B(new_n10566), .C(new_n10562), .Y(new_n10872));
  NOR2xp33_ASAP7_75t_L      g10616(.A(new_n10872), .B(new_n10869), .Y(new_n10873));
  NOR2xp33_ASAP7_75t_L      g10617(.A(new_n10873), .B(new_n10871), .Y(\f[61] ));
  OAI21xp33_ASAP7_75t_L     g10618(.A1(new_n10823), .A2(new_n10822), .B(new_n10576), .Y(new_n10875));
  A2O1A1O1Ixp25_ASAP7_75t_L g10619(.A1(new_n10544), .A2(new_n10547), .B(new_n10573), .C(new_n10875), .D(new_n10824), .Y(new_n10876));
  OAI22xp33_ASAP7_75t_L     g10620(.A1(new_n706), .A2(new_n7616), .B1(new_n8165), .B2(new_n580), .Y(new_n10877));
  AOI221xp5_ASAP7_75t_L     g10621(.A1(\b[52] ), .A2(new_n584), .B1(new_n578), .B2(new_n8173), .C(new_n10877), .Y(new_n10878));
  XNOR2x2_ASAP7_75t_L       g10622(.A(new_n574), .B(new_n10878), .Y(new_n10879));
  NOR3xp33_ASAP7_75t_L      g10623(.A(new_n10809), .B(new_n10812), .C(new_n10585), .Y(new_n10880));
  A2O1A1O1Ixp25_ASAP7_75t_L g10624(.A1(new_n10283), .A2(new_n10532), .B(new_n10578), .C(new_n10813), .D(new_n10880), .Y(new_n10881));
  NOR3xp33_ASAP7_75t_L      g10625(.A(new_n10802), .B(new_n10798), .C(new_n10590), .Y(new_n10882));
  A2O1A1O1Ixp25_ASAP7_75t_L g10626(.A1(new_n10526), .A2(new_n10525), .B(new_n10586), .C(new_n10803), .D(new_n10882), .Y(new_n10883));
  NOR2xp33_ASAP7_75t_L      g10627(.A(new_n6568), .B(new_n1154), .Y(new_n10884));
  INVx1_ASAP7_75t_L         g10628(.A(new_n10884), .Y(new_n10885));
  NAND2xp33_ASAP7_75t_L     g10629(.A(new_n1073), .B(new_n8186), .Y(new_n10886));
  AOI22xp33_ASAP7_75t_L     g10630(.A1(new_n1076), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1253), .Y(new_n10887));
  NAND4xp25_ASAP7_75t_L     g10631(.A(new_n10886), .B(\a[17] ), .C(new_n10885), .D(new_n10887), .Y(new_n10888));
  NAND2xp33_ASAP7_75t_L     g10632(.A(new_n10887), .B(new_n10886), .Y(new_n10889));
  A2O1A1Ixp33_ASAP7_75t_L   g10633(.A1(\b[46] ), .A2(new_n1080), .B(new_n10889), .C(new_n1071), .Y(new_n10890));
  AND2x2_ASAP7_75t_L        g10634(.A(new_n10888), .B(new_n10890), .Y(new_n10891));
  AOI22xp33_ASAP7_75t_L     g10635(.A1(new_n1360), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1581), .Y(new_n10892));
  OAI221xp5_ASAP7_75t_L     g10636(.A1(new_n1373), .A2(new_n5805), .B1(new_n1359), .B2(new_n5835), .C(new_n10892), .Y(new_n10893));
  XNOR2x2_ASAP7_75t_L       g10637(.A(\a[20] ), .B(new_n10893), .Y(new_n10894));
  NAND3xp33_ASAP7_75t_L     g10638(.A(new_n10768), .B(new_n10764), .C(new_n10779), .Y(new_n10895));
  INVx1_ASAP7_75t_L         g10639(.A(new_n10895), .Y(new_n10896));
  AOI21xp33_ASAP7_75t_L     g10640(.A1(new_n10593), .A2(new_n10746), .B(new_n10756), .Y(new_n10897));
  AOI22xp33_ASAP7_75t_L     g10641(.A1(new_n2552), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n2736), .Y(new_n10898));
  OAI221xp5_ASAP7_75t_L     g10642(.A1(new_n2547), .A2(new_n3584), .B1(new_n2734), .B2(new_n10137), .C(new_n10898), .Y(new_n10899));
  XNOR2x2_ASAP7_75t_L       g10643(.A(\a[29] ), .B(new_n10899), .Y(new_n10900));
  NAND2xp33_ASAP7_75t_L     g10644(.A(new_n10732), .B(new_n10731), .Y(new_n10901));
  MAJIxp5_ASAP7_75t_L       g10645(.A(new_n10594), .B(new_n10728), .C(new_n10901), .Y(new_n10902));
  NOR3xp33_ASAP7_75t_L      g10646(.A(new_n10693), .B(new_n10692), .C(new_n10599), .Y(new_n10903));
  A2O1A1O1Ixp25_ASAP7_75t_L g10647(.A1(new_n10404), .A2(new_n10304), .B(new_n10595), .C(new_n10694), .D(new_n10903), .Y(new_n10904));
  NOR2xp33_ASAP7_75t_L      g10648(.A(new_n1774), .B(new_n5154), .Y(new_n10905));
  INVx1_ASAP7_75t_L         g10649(.A(new_n10905), .Y(new_n10906));
  NAND3xp33_ASAP7_75t_L     g10650(.A(new_n1912), .B(new_n1914), .C(new_n4917), .Y(new_n10907));
  AOI22xp33_ASAP7_75t_L     g10651(.A1(new_n4920), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n5167), .Y(new_n10908));
  AND4x1_ASAP7_75t_L        g10652(.A(new_n10908), .B(new_n10907), .C(new_n10906), .D(\a[41] ), .Y(new_n10909));
  AOI31xp33_ASAP7_75t_L     g10653(.A1(new_n10907), .A2(new_n10906), .A3(new_n10908), .B(\a[41] ), .Y(new_n10910));
  NOR2xp33_ASAP7_75t_L      g10654(.A(new_n10910), .B(new_n10909), .Y(new_n10911));
  INVx1_ASAP7_75t_L         g10655(.A(new_n10911), .Y(new_n10912));
  AOI22xp33_ASAP7_75t_L     g10656(.A1(new_n5624), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n5901), .Y(new_n10913));
  OAI221xp5_ASAP7_75t_L     g10657(.A1(new_n5900), .A2(new_n1432), .B1(new_n5892), .B2(new_n1547), .C(new_n10913), .Y(new_n10914));
  XNOR2x2_ASAP7_75t_L       g10658(.A(\a[44] ), .B(new_n10914), .Y(new_n10915));
  INVx1_ASAP7_75t_L         g10659(.A(new_n10915), .Y(new_n10916));
  NOR3xp33_ASAP7_75t_L      g10660(.A(new_n10670), .B(new_n10671), .C(new_n10606), .Y(new_n10917));
  AOI22xp33_ASAP7_75t_L     g10661(.A1(new_n6376), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n6648), .Y(new_n10918));
  OAI221xp5_ASAP7_75t_L     g10662(.A1(new_n6646), .A2(new_n1030), .B1(new_n6636), .B2(new_n1209), .C(new_n10918), .Y(new_n10919));
  XNOR2x2_ASAP7_75t_L       g10663(.A(\a[47] ), .B(new_n10919), .Y(new_n10920));
  INVx1_ASAP7_75t_L         g10664(.A(new_n10920), .Y(new_n10921));
  NAND2xp33_ASAP7_75t_L     g10665(.A(new_n10645), .B(new_n10648), .Y(new_n10922));
  MAJIxp5_ASAP7_75t_L       g10666(.A(new_n10655), .B(new_n10651), .C(new_n10922), .Y(new_n10923));
  AOI22xp33_ASAP7_75t_L     g10667(.A1(new_n7960), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n8537), .Y(new_n10924));
  OAI221xp5_ASAP7_75t_L     g10668(.A1(new_n8817), .A2(new_n617), .B1(new_n7957), .B2(new_n685), .C(new_n10924), .Y(new_n10925));
  XNOR2x2_ASAP7_75t_L       g10669(.A(new_n7954), .B(new_n10925), .Y(new_n10926));
  A2O1A1Ixp33_ASAP7_75t_L   g10670(.A1(new_n10646), .A2(new_n10609), .B(new_n10642), .C(new_n10644), .Y(new_n10927));
  AOI22xp33_ASAP7_75t_L     g10671(.A1(new_n8831), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n9115), .Y(new_n10928));
  OAI221xp5_ASAP7_75t_L     g10672(.A1(new_n10343), .A2(new_n420), .B1(new_n10016), .B2(new_n494), .C(new_n10928), .Y(new_n10929));
  XNOR2x2_ASAP7_75t_L       g10673(.A(\a[56] ), .B(new_n10929), .Y(new_n10930));
  O2A1O1Ixp33_ASAP7_75t_L   g10674(.A1(new_n10614), .A2(new_n10350), .B(new_n10636), .C(new_n10637), .Y(new_n10931));
  OAI22xp33_ASAP7_75t_L     g10675(.A1(new_n10026), .A2(new_n298), .B1(new_n354), .B2(new_n9699), .Y(new_n10932));
  AOI221xp5_ASAP7_75t_L     g10676(.A1(new_n9703), .A2(\b[4] ), .B1(new_n9697), .B2(new_n359), .C(new_n10932), .Y(new_n10933));
  NAND2xp33_ASAP7_75t_L     g10677(.A(\a[59] ), .B(new_n10933), .Y(new_n10934));
  AO21x2_ASAP7_75t_L        g10678(.A1(new_n9697), .A2(new_n359), .B(new_n10932), .Y(new_n10935));
  A2O1A1Ixp33_ASAP7_75t_L   g10679(.A1(\b[4] ), .A2(new_n9703), .B(new_n10935), .C(new_n9693), .Y(new_n10936));
  INVx1_ASAP7_75t_L         g10680(.A(new_n10632), .Y(new_n10937));
  INVx1_ASAP7_75t_L         g10681(.A(new_n10630), .Y(new_n10938));
  AND3x1_ASAP7_75t_L        g10682(.A(new_n10332), .B(new_n10631), .C(new_n10628), .Y(new_n10939));
  AOI22xp33_ASAP7_75t_L     g10683(.A1(new_n10938), .A2(\b[2] ), .B1(\b[0] ), .B2(new_n10939), .Y(new_n10940));
  OAI221xp5_ASAP7_75t_L     g10684(.A1(new_n10629), .A2(new_n280), .B1(new_n261), .B2(new_n10937), .C(new_n10940), .Y(new_n10941));
  O2A1O1Ixp33_ASAP7_75t_L   g10685(.A1(new_n10333), .A2(new_n10634), .B(\a[62] ), .C(new_n10941), .Y(new_n10942));
  A2O1A1Ixp33_ASAP7_75t_L   g10686(.A1(\b[0] ), .A2(new_n10624), .B(new_n10634), .C(\a[62] ), .Y(new_n10943));
  OA21x2_ASAP7_75t_L        g10687(.A1(new_n280), .A2(new_n10629), .B(new_n10940), .Y(new_n10944));
  O2A1O1Ixp33_ASAP7_75t_L   g10688(.A1(new_n10937), .A2(new_n261), .B(new_n10944), .C(new_n10943), .Y(new_n10945));
  OAI211xp5_ASAP7_75t_L     g10689(.A1(new_n10942), .A2(new_n10945), .B(new_n10936), .C(new_n10934), .Y(new_n10946));
  NAND2xp33_ASAP7_75t_L     g10690(.A(new_n10934), .B(new_n10936), .Y(new_n10947));
  NOR2xp33_ASAP7_75t_L      g10691(.A(new_n10942), .B(new_n10945), .Y(new_n10948));
  NAND2xp33_ASAP7_75t_L     g10692(.A(new_n10948), .B(new_n10947), .Y(new_n10949));
  NAND2xp33_ASAP7_75t_L     g10693(.A(new_n10946), .B(new_n10949), .Y(new_n10950));
  NAND2xp33_ASAP7_75t_L     g10694(.A(new_n10950), .B(new_n10931), .Y(new_n10951));
  A2O1A1Ixp33_ASAP7_75t_L   g10695(.A1(new_n10341), .A2(new_n10615), .B(new_n10640), .C(new_n10638), .Y(new_n10952));
  NAND3xp33_ASAP7_75t_L     g10696(.A(new_n10952), .B(new_n10946), .C(new_n10949), .Y(new_n10953));
  NAND2xp33_ASAP7_75t_L     g10697(.A(new_n10951), .B(new_n10953), .Y(new_n10954));
  NAND2xp33_ASAP7_75t_L     g10698(.A(new_n10930), .B(new_n10954), .Y(new_n10955));
  INVx1_ASAP7_75t_L         g10699(.A(new_n10930), .Y(new_n10956));
  AOI21xp33_ASAP7_75t_L     g10700(.A1(new_n10949), .A2(new_n10946), .B(new_n10952), .Y(new_n10957));
  A2O1A1O1Ixp25_ASAP7_75t_L g10701(.A1(new_n10615), .A2(new_n10341), .B(new_n10640), .C(new_n10638), .D(new_n10950), .Y(new_n10958));
  NOR2xp33_ASAP7_75t_L      g10702(.A(new_n10957), .B(new_n10958), .Y(new_n10959));
  NAND2xp33_ASAP7_75t_L     g10703(.A(new_n10956), .B(new_n10959), .Y(new_n10960));
  NAND3xp33_ASAP7_75t_L     g10704(.A(new_n10927), .B(new_n10955), .C(new_n10960), .Y(new_n10961));
  NOR2xp33_ASAP7_75t_L      g10705(.A(new_n10956), .B(new_n10959), .Y(new_n10962));
  NOR2xp33_ASAP7_75t_L      g10706(.A(new_n10930), .B(new_n10954), .Y(new_n10963));
  OAI211xp5_ASAP7_75t_L     g10707(.A1(new_n10963), .A2(new_n10962), .B(new_n10645), .C(new_n10644), .Y(new_n10964));
  AO21x2_ASAP7_75t_L        g10708(.A1(new_n10961), .A2(new_n10964), .B(new_n10926), .Y(new_n10965));
  NAND3xp33_ASAP7_75t_L     g10709(.A(new_n10964), .B(new_n10961), .C(new_n10926), .Y(new_n10966));
  NAND3xp33_ASAP7_75t_L     g10710(.A(new_n10965), .B(new_n10923), .C(new_n10966), .Y(new_n10967));
  AO21x2_ASAP7_75t_L        g10711(.A1(new_n10966), .A2(new_n10965), .B(new_n10923), .Y(new_n10968));
  AOI22xp33_ASAP7_75t_L     g10712(.A1(new_n7111), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n7391), .Y(new_n10969));
  OAI221xp5_ASAP7_75t_L     g10713(.A1(new_n8558), .A2(new_n784), .B1(new_n8237), .B2(new_n875), .C(new_n10969), .Y(new_n10970));
  XNOR2x2_ASAP7_75t_L       g10714(.A(\a[50] ), .B(new_n10970), .Y(new_n10971));
  NAND3xp33_ASAP7_75t_L     g10715(.A(new_n10968), .B(new_n10967), .C(new_n10971), .Y(new_n10972));
  AO21x2_ASAP7_75t_L        g10716(.A1(new_n10967), .A2(new_n10968), .B(new_n10971), .Y(new_n10973));
  OAI21xp33_ASAP7_75t_L     g10717(.A1(new_n10664), .A2(new_n10666), .B(new_n10667), .Y(new_n10974));
  AOI21xp33_ASAP7_75t_L     g10718(.A1(new_n10973), .A2(new_n10972), .B(new_n10974), .Y(new_n10975));
  AND3x1_ASAP7_75t_L        g10719(.A(new_n10968), .B(new_n10971), .C(new_n10967), .Y(new_n10976));
  AOI21xp33_ASAP7_75t_L     g10720(.A1(new_n10968), .A2(new_n10967), .B(new_n10971), .Y(new_n10977));
  AOI21xp33_ASAP7_75t_L     g10721(.A1(new_n10608), .A2(new_n10663), .B(new_n10662), .Y(new_n10978));
  NOR3xp33_ASAP7_75t_L      g10722(.A(new_n10978), .B(new_n10977), .C(new_n10976), .Y(new_n10979));
  OAI21xp33_ASAP7_75t_L     g10723(.A1(new_n10975), .A2(new_n10979), .B(new_n10921), .Y(new_n10980));
  OAI21xp33_ASAP7_75t_L     g10724(.A1(new_n10976), .A2(new_n10977), .B(new_n10978), .Y(new_n10981));
  NAND3xp33_ASAP7_75t_L     g10725(.A(new_n10974), .B(new_n10973), .C(new_n10972), .Y(new_n10982));
  NAND3xp33_ASAP7_75t_L     g10726(.A(new_n10982), .B(new_n10981), .C(new_n10920), .Y(new_n10983));
  NAND2xp33_ASAP7_75t_L     g10727(.A(new_n10983), .B(new_n10980), .Y(new_n10984));
  A2O1A1Ixp33_ASAP7_75t_L   g10728(.A1(new_n10672), .A2(new_n10603), .B(new_n10917), .C(new_n10984), .Y(new_n10985));
  A2O1A1Ixp33_ASAP7_75t_L   g10729(.A1(new_n9743), .A2(new_n9742), .B(new_n9744), .C(new_n10073), .Y(new_n10986));
  A2O1A1Ixp33_ASAP7_75t_L   g10730(.A1(new_n10069), .A2(new_n10065), .B(new_n10986), .C(new_n10316), .Y(new_n10987));
  A2O1A1O1Ixp25_ASAP7_75t_L g10731(.A1(new_n10387), .A2(new_n10987), .B(new_n10380), .C(new_n10672), .D(new_n10917), .Y(new_n10988));
  NAND3xp33_ASAP7_75t_L     g10732(.A(new_n10988), .B(new_n10980), .C(new_n10983), .Y(new_n10989));
  NAND3xp33_ASAP7_75t_L     g10733(.A(new_n10985), .B(new_n10916), .C(new_n10989), .Y(new_n10990));
  AOI21xp33_ASAP7_75t_L     g10734(.A1(new_n10983), .A2(new_n10980), .B(new_n10988), .Y(new_n10991));
  A2O1A1Ixp33_ASAP7_75t_L   g10735(.A1(new_n10386), .A2(new_n10390), .B(new_n10675), .C(new_n10669), .Y(new_n10992));
  NOR2xp33_ASAP7_75t_L      g10736(.A(new_n10984), .B(new_n10992), .Y(new_n10993));
  OAI21xp33_ASAP7_75t_L     g10737(.A1(new_n10991), .A2(new_n10993), .B(new_n10915), .Y(new_n10994));
  OAI211xp5_ASAP7_75t_L     g10738(.A1(new_n10687), .A2(new_n10402), .B(new_n10688), .C(new_n10684), .Y(new_n10995));
  NAND4xp25_ASAP7_75t_L     g10739(.A(new_n10995), .B(new_n10994), .C(new_n10990), .D(new_n10680), .Y(new_n10996));
  INVx1_ASAP7_75t_L         g10740(.A(new_n10680), .Y(new_n10997));
  NOR3xp33_ASAP7_75t_L      g10741(.A(new_n10993), .B(new_n10991), .C(new_n10915), .Y(new_n10998));
  AOI21xp33_ASAP7_75t_L     g10742(.A1(new_n10985), .A2(new_n10989), .B(new_n10916), .Y(new_n10999));
  NOR2xp33_ASAP7_75t_L      g10743(.A(new_n10673), .B(new_n10676), .Y(new_n11000));
  AOI221xp5_ASAP7_75t_L     g10744(.A1(new_n10393), .A2(new_n10396), .B1(new_n11000), .B2(new_n10683), .C(new_n10601), .Y(new_n11001));
  OAI22xp33_ASAP7_75t_L     g10745(.A1(new_n11001), .A2(new_n10997), .B1(new_n10998), .B2(new_n10999), .Y(new_n11002));
  NAND3xp33_ASAP7_75t_L     g10746(.A(new_n11002), .B(new_n10996), .C(new_n10912), .Y(new_n11003));
  NOR4xp25_ASAP7_75t_L      g10747(.A(new_n11001), .B(new_n10999), .C(new_n10998), .D(new_n10997), .Y(new_n11004));
  AOI22xp33_ASAP7_75t_L     g10748(.A1(new_n10994), .A2(new_n10990), .B1(new_n10680), .B2(new_n10995), .Y(new_n11005));
  OAI21xp33_ASAP7_75t_L     g10749(.A1(new_n11005), .A2(new_n11004), .B(new_n10911), .Y(new_n11006));
  NAND2xp33_ASAP7_75t_L     g10750(.A(new_n11003), .B(new_n11006), .Y(new_n11007));
  NAND2xp33_ASAP7_75t_L     g10751(.A(new_n10904), .B(new_n11007), .Y(new_n11008));
  NOR3xp33_ASAP7_75t_L      g10752(.A(new_n11004), .B(new_n11005), .C(new_n10911), .Y(new_n11009));
  AOI21xp33_ASAP7_75t_L     g10753(.A1(new_n11002), .A2(new_n10996), .B(new_n10912), .Y(new_n11010));
  NOR2xp33_ASAP7_75t_L      g10754(.A(new_n11010), .B(new_n11009), .Y(new_n11011));
  A2O1A1Ixp33_ASAP7_75t_L   g10755(.A1(new_n10694), .A2(new_n10698), .B(new_n10903), .C(new_n11011), .Y(new_n11012));
  AOI22xp33_ASAP7_75t_L     g10756(.A1(new_n4283), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n4512), .Y(new_n11013));
  OAI221xp5_ASAP7_75t_L     g10757(.A1(new_n4277), .A2(new_n2067), .B1(new_n4499), .B2(new_n2355), .C(new_n11013), .Y(new_n11014));
  XNOR2x2_ASAP7_75t_L       g10758(.A(\a[38] ), .B(new_n11014), .Y(new_n11015));
  NAND3xp33_ASAP7_75t_L     g10759(.A(new_n11012), .B(new_n11008), .C(new_n11015), .Y(new_n11016));
  AOI221xp5_ASAP7_75t_L     g10760(.A1(new_n11006), .A2(new_n11003), .B1(new_n10694), .B2(new_n10698), .C(new_n10903), .Y(new_n11017));
  O2A1O1Ixp33_ASAP7_75t_L   g10761(.A1(new_n10596), .A2(new_n10695), .B(new_n10691), .C(new_n11007), .Y(new_n11018));
  INVx1_ASAP7_75t_L         g10762(.A(new_n11015), .Y(new_n11019));
  OAI21xp33_ASAP7_75t_L     g10763(.A1(new_n11017), .A2(new_n11018), .B(new_n11019), .Y(new_n11020));
  AND2x2_ASAP7_75t_L        g10764(.A(new_n11020), .B(new_n11016), .Y(new_n11021));
  INVx1_ASAP7_75t_L         g10765(.A(new_n10702), .Y(new_n11022));
  AND3x1_ASAP7_75t_L        g10766(.A(new_n11022), .B(new_n10699), .C(new_n10696), .Y(new_n11023));
  O2A1O1Ixp33_ASAP7_75t_L   g10767(.A1(new_n10708), .A2(new_n10707), .B(new_n10709), .C(new_n11023), .Y(new_n11024));
  NAND2xp33_ASAP7_75t_L     g10768(.A(new_n11024), .B(new_n11021), .Y(new_n11025));
  NAND2xp33_ASAP7_75t_L     g10769(.A(new_n10703), .B(new_n10704), .Y(new_n11026));
  NAND2xp33_ASAP7_75t_L     g10770(.A(new_n11020), .B(new_n11016), .Y(new_n11027));
  A2O1A1Ixp33_ASAP7_75t_L   g10771(.A1(new_n11026), .A2(new_n10709), .B(new_n11023), .C(new_n11027), .Y(new_n11028));
  AOI22xp33_ASAP7_75t_L     g10772(.A1(new_n3633), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n3858), .Y(new_n11029));
  OAI221xp5_ASAP7_75t_L     g10773(.A1(new_n3853), .A2(new_n2666), .B1(new_n3856), .B2(new_n2695), .C(new_n11029), .Y(new_n11030));
  XNOR2x2_ASAP7_75t_L       g10774(.A(\a[35] ), .B(new_n11030), .Y(new_n11031));
  NAND3xp33_ASAP7_75t_L     g10775(.A(new_n11025), .B(new_n11028), .C(new_n11031), .Y(new_n11032));
  NOR3xp33_ASAP7_75t_L      g10776(.A(new_n10716), .B(new_n11027), .C(new_n11023), .Y(new_n11033));
  NOR2xp33_ASAP7_75t_L      g10777(.A(new_n11024), .B(new_n11021), .Y(new_n11034));
  INVx1_ASAP7_75t_L         g10778(.A(new_n11031), .Y(new_n11035));
  OAI21xp33_ASAP7_75t_L     g10779(.A1(new_n11033), .A2(new_n11034), .B(new_n11035), .Y(new_n11036));
  NAND2xp33_ASAP7_75t_L     g10780(.A(new_n11032), .B(new_n11036), .Y(new_n11037));
  NOR3xp33_ASAP7_75t_L      g10781(.A(new_n10715), .B(new_n10716), .C(new_n10713), .Y(new_n11038));
  INVx1_ASAP7_75t_L         g10782(.A(new_n11038), .Y(new_n11039));
  A2O1A1Ixp33_ASAP7_75t_L   g10783(.A1(new_n10718), .A2(new_n10714), .B(new_n10724), .C(new_n11039), .Y(new_n11040));
  NOR2xp33_ASAP7_75t_L      g10784(.A(new_n11037), .B(new_n11040), .Y(new_n11041));
  NOR3xp33_ASAP7_75t_L      g10785(.A(new_n11034), .B(new_n11033), .C(new_n11035), .Y(new_n11042));
  AOI21xp33_ASAP7_75t_L     g10786(.A1(new_n11025), .A2(new_n11028), .B(new_n11031), .Y(new_n11043));
  NOR2xp33_ASAP7_75t_L      g10787(.A(new_n11043), .B(new_n11042), .Y(new_n11044));
  A2O1A1O1Ixp25_ASAP7_75t_L g10788(.A1(new_n10437), .A2(new_n10435), .B(new_n10720), .C(new_n10719), .D(new_n11038), .Y(new_n11045));
  NOR2xp33_ASAP7_75t_L      g10789(.A(new_n11045), .B(new_n11044), .Y(new_n11046));
  NAND2xp33_ASAP7_75t_L     g10790(.A(new_n3213), .B(new_n3210), .Y(new_n11047));
  AOI22xp33_ASAP7_75t_L     g10791(.A1(new_n3029), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n3258), .Y(new_n11048));
  OAI221xp5_ASAP7_75t_L     g10792(.A1(new_n3024), .A2(new_n3180), .B1(new_n3256), .B2(new_n11047), .C(new_n11048), .Y(new_n11049));
  XNOR2x2_ASAP7_75t_L       g10793(.A(\a[32] ), .B(new_n11049), .Y(new_n11050));
  OAI21xp33_ASAP7_75t_L     g10794(.A1(new_n11046), .A2(new_n11041), .B(new_n11050), .Y(new_n11051));
  NAND2xp33_ASAP7_75t_L     g10795(.A(new_n11045), .B(new_n11044), .Y(new_n11052));
  A2O1A1Ixp33_ASAP7_75t_L   g10796(.A1(new_n10719), .A2(new_n10722), .B(new_n11038), .C(new_n11037), .Y(new_n11053));
  INVx1_ASAP7_75t_L         g10797(.A(new_n11050), .Y(new_n11054));
  NAND3xp33_ASAP7_75t_L     g10798(.A(new_n11053), .B(new_n11052), .C(new_n11054), .Y(new_n11055));
  AOI21xp33_ASAP7_75t_L     g10799(.A1(new_n11055), .A2(new_n11051), .B(new_n10902), .Y(new_n11056));
  XNOR2x2_ASAP7_75t_L       g10800(.A(new_n10719), .B(new_n10724), .Y(new_n11057));
  MAJIxp5_ASAP7_75t_L       g10801(.A(new_n10735), .B(new_n10729), .C(new_n11057), .Y(new_n11058));
  AOI21xp33_ASAP7_75t_L     g10802(.A1(new_n11053), .A2(new_n11052), .B(new_n11054), .Y(new_n11059));
  NOR3xp33_ASAP7_75t_L      g10803(.A(new_n11041), .B(new_n11046), .C(new_n11050), .Y(new_n11060));
  NOR3xp33_ASAP7_75t_L      g10804(.A(new_n11058), .B(new_n11059), .C(new_n11060), .Y(new_n11061));
  NOR3xp33_ASAP7_75t_L      g10805(.A(new_n11061), .B(new_n10900), .C(new_n11056), .Y(new_n11062));
  INVx1_ASAP7_75t_L         g10806(.A(new_n10900), .Y(new_n11063));
  OAI21xp33_ASAP7_75t_L     g10807(.A1(new_n11060), .A2(new_n11059), .B(new_n11058), .Y(new_n11064));
  NAND3xp33_ASAP7_75t_L     g10808(.A(new_n10902), .B(new_n11051), .C(new_n11055), .Y(new_n11065));
  AOI21xp33_ASAP7_75t_L     g10809(.A1(new_n11065), .A2(new_n11064), .B(new_n11063), .Y(new_n11066));
  OAI21xp33_ASAP7_75t_L     g10810(.A1(new_n11062), .A2(new_n11066), .B(new_n10897), .Y(new_n11067));
  AO21x2_ASAP7_75t_L        g10811(.A1(new_n10746), .A2(new_n10593), .B(new_n10756), .Y(new_n11068));
  NAND3xp33_ASAP7_75t_L     g10812(.A(new_n11065), .B(new_n11064), .C(new_n11063), .Y(new_n11069));
  OAI21xp33_ASAP7_75t_L     g10813(.A1(new_n11056), .A2(new_n11061), .B(new_n10900), .Y(new_n11070));
  NAND3xp33_ASAP7_75t_L     g10814(.A(new_n11068), .B(new_n11069), .C(new_n11070), .Y(new_n11071));
  OAI22xp33_ASAP7_75t_L     g10815(.A1(new_n2269), .A2(new_n4216), .B1(new_n4632), .B2(new_n2107), .Y(new_n11072));
  AOI221xp5_ASAP7_75t_L     g10816(.A1(\b[37] ), .A2(new_n2115), .B1(new_n2106), .B2(new_n4640), .C(new_n11072), .Y(new_n11073));
  XNOR2x2_ASAP7_75t_L       g10817(.A(new_n2100), .B(new_n11073), .Y(new_n11074));
  NAND3xp33_ASAP7_75t_L     g10818(.A(new_n11071), .B(new_n11067), .C(new_n11074), .Y(new_n11075));
  AOI221xp5_ASAP7_75t_L     g10819(.A1(new_n10593), .A2(new_n10746), .B1(new_n11069), .B2(new_n11070), .C(new_n10756), .Y(new_n11076));
  NOR3xp33_ASAP7_75t_L      g10820(.A(new_n10897), .B(new_n11062), .C(new_n11066), .Y(new_n11077));
  INVx1_ASAP7_75t_L         g10821(.A(new_n11074), .Y(new_n11078));
  OAI21xp33_ASAP7_75t_L     g10822(.A1(new_n11076), .A2(new_n11077), .B(new_n11078), .Y(new_n11079));
  NAND2xp33_ASAP7_75t_L     g10823(.A(new_n11079), .B(new_n11075), .Y(new_n11080));
  NAND3xp33_ASAP7_75t_L     g10824(.A(new_n10759), .B(new_n10758), .C(new_n10754), .Y(new_n11081));
  A2O1A1Ixp33_ASAP7_75t_L   g10825(.A1(new_n10766), .A2(new_n10765), .B(new_n10763), .C(new_n11081), .Y(new_n11082));
  NOR2xp33_ASAP7_75t_L      g10826(.A(new_n11080), .B(new_n11082), .Y(new_n11083));
  NOR3xp33_ASAP7_75t_L      g10827(.A(new_n11077), .B(new_n11078), .C(new_n11076), .Y(new_n11084));
  AOI21xp33_ASAP7_75t_L     g10828(.A1(new_n11071), .A2(new_n11067), .B(new_n11074), .Y(new_n11085));
  NOR2xp33_ASAP7_75t_L      g10829(.A(new_n11084), .B(new_n11085), .Y(new_n11086));
  AOI21xp33_ASAP7_75t_L     g10830(.A1(new_n10768), .A2(new_n11081), .B(new_n11086), .Y(new_n11087));
  AOI22xp33_ASAP7_75t_L     g10831(.A1(new_n1704), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1837), .Y(new_n11088));
  OAI221xp5_ASAP7_75t_L     g10832(.A1(new_n1699), .A2(new_n4869), .B1(new_n1827), .B2(new_n5327), .C(new_n11088), .Y(new_n11089));
  XNOR2x2_ASAP7_75t_L       g10833(.A(\a[23] ), .B(new_n11089), .Y(new_n11090));
  OAI21xp33_ASAP7_75t_L     g10834(.A1(new_n11083), .A2(new_n11087), .B(new_n11090), .Y(new_n11091));
  NAND3xp33_ASAP7_75t_L     g10835(.A(new_n11086), .B(new_n10768), .C(new_n11081), .Y(new_n11092));
  NAND2xp33_ASAP7_75t_L     g10836(.A(new_n11080), .B(new_n11082), .Y(new_n11093));
  INVx1_ASAP7_75t_L         g10837(.A(new_n11090), .Y(new_n11094));
  NAND3xp33_ASAP7_75t_L     g10838(.A(new_n11092), .B(new_n11093), .C(new_n11094), .Y(new_n11095));
  AOI221xp5_ASAP7_75t_L     g10839(.A1(new_n10781), .A2(new_n10783), .B1(new_n11091), .B2(new_n11095), .C(new_n10896), .Y(new_n11096));
  O2A1O1Ixp33_ASAP7_75t_L   g10840(.A1(new_n10785), .A2(new_n10786), .B(new_n10783), .C(new_n10896), .Y(new_n11097));
  NAND2xp33_ASAP7_75t_L     g10841(.A(new_n11095), .B(new_n11091), .Y(new_n11098));
  NOR2xp33_ASAP7_75t_L      g10842(.A(new_n11098), .B(new_n11097), .Y(new_n11099));
  NOR3xp33_ASAP7_75t_L      g10843(.A(new_n11099), .B(new_n11096), .C(new_n10894), .Y(new_n11100));
  INVx1_ASAP7_75t_L         g10844(.A(new_n10894), .Y(new_n11101));
  INVx1_ASAP7_75t_L         g10845(.A(new_n11096), .Y(new_n11102));
  AOI21xp33_ASAP7_75t_L     g10846(.A1(new_n11092), .A2(new_n11093), .B(new_n11094), .Y(new_n11103));
  NOR3xp33_ASAP7_75t_L      g10847(.A(new_n11087), .B(new_n11083), .C(new_n11090), .Y(new_n11104));
  NOR2xp33_ASAP7_75t_L      g10848(.A(new_n11103), .B(new_n11104), .Y(new_n11105));
  A2O1A1Ixp33_ASAP7_75t_L   g10849(.A1(new_n10783), .A2(new_n10781), .B(new_n10896), .C(new_n11105), .Y(new_n11106));
  AOI21xp33_ASAP7_75t_L     g10850(.A1(new_n11102), .A2(new_n11106), .B(new_n11101), .Y(new_n11107));
  OAI21xp33_ASAP7_75t_L     g10851(.A1(new_n10801), .A2(new_n10591), .B(new_n10793), .Y(new_n11108));
  NOR3xp33_ASAP7_75t_L      g10852(.A(new_n11108), .B(new_n11107), .C(new_n11100), .Y(new_n11109));
  NAND3xp33_ASAP7_75t_L     g10853(.A(new_n11102), .B(new_n11106), .C(new_n11101), .Y(new_n11110));
  OAI21xp33_ASAP7_75t_L     g10854(.A1(new_n11096), .A2(new_n11099), .B(new_n10894), .Y(new_n11111));
  OAI311xp33_ASAP7_75t_L    g10855(.A1(new_n10172), .A2(new_n10508), .A3(new_n10514), .B1(new_n10517), .C1(new_n10797), .Y(new_n11112));
  AOI22xp33_ASAP7_75t_L     g10856(.A1(new_n11112), .A2(new_n10793), .B1(new_n11111), .B2(new_n11110), .Y(new_n11113));
  NOR3xp33_ASAP7_75t_L      g10857(.A(new_n10891), .B(new_n11109), .C(new_n11113), .Y(new_n11114));
  NAND2xp33_ASAP7_75t_L     g10858(.A(new_n10888), .B(new_n10890), .Y(new_n11115));
  NAND4xp25_ASAP7_75t_L     g10859(.A(new_n11110), .B(new_n11112), .C(new_n10793), .D(new_n11111), .Y(new_n11116));
  OAI21xp33_ASAP7_75t_L     g10860(.A1(new_n11100), .A2(new_n11107), .B(new_n11108), .Y(new_n11117));
  AOI21xp33_ASAP7_75t_L     g10861(.A1(new_n11117), .A2(new_n11116), .B(new_n11115), .Y(new_n11118));
  OR3x1_ASAP7_75t_L         g10862(.A(new_n10883), .B(new_n11114), .C(new_n11118), .Y(new_n11119));
  NAND3xp33_ASAP7_75t_L     g10863(.A(new_n11117), .B(new_n11116), .C(new_n11115), .Y(new_n11120));
  OAI21xp33_ASAP7_75t_L     g10864(.A1(new_n11113), .A2(new_n11109), .B(new_n10891), .Y(new_n11121));
  NAND2xp33_ASAP7_75t_L     g10865(.A(new_n11120), .B(new_n11121), .Y(new_n11122));
  NAND2xp33_ASAP7_75t_L     g10866(.A(new_n10883), .B(new_n11122), .Y(new_n11123));
  NAND2xp33_ASAP7_75t_L     g10867(.A(\b[48] ), .B(new_n900), .Y(new_n11124));
  OAI221xp5_ASAP7_75t_L     g10868(.A1(new_n977), .A2(new_n7593), .B1(new_n898), .B2(new_n7602), .C(new_n11124), .Y(new_n11125));
  AOI21xp33_ASAP7_75t_L     g10869(.A1(new_n815), .A2(\b[49] ), .B(new_n11125), .Y(new_n11126));
  NAND2xp33_ASAP7_75t_L     g10870(.A(\a[14] ), .B(new_n11126), .Y(new_n11127));
  A2O1A1Ixp33_ASAP7_75t_L   g10871(.A1(\b[49] ), .A2(new_n815), .B(new_n11125), .C(new_n806), .Y(new_n11128));
  AND2x2_ASAP7_75t_L        g10872(.A(new_n11128), .B(new_n11127), .Y(new_n11129));
  NAND3xp33_ASAP7_75t_L     g10873(.A(new_n11129), .B(new_n11119), .C(new_n11123), .Y(new_n11130));
  NOR2xp33_ASAP7_75t_L      g10874(.A(new_n10883), .B(new_n11122), .Y(new_n11131));
  AOI221xp5_ASAP7_75t_L     g10875(.A1(new_n10811), .A2(new_n10803), .B1(new_n11120), .B2(new_n11121), .C(new_n10882), .Y(new_n11132));
  NAND2xp33_ASAP7_75t_L     g10876(.A(new_n11128), .B(new_n11127), .Y(new_n11133));
  OAI21xp33_ASAP7_75t_L     g10877(.A1(new_n11132), .A2(new_n11131), .B(new_n11133), .Y(new_n11134));
  AOI21xp33_ASAP7_75t_L     g10878(.A1(new_n11134), .A2(new_n11130), .B(new_n10881), .Y(new_n11135));
  INVx1_ASAP7_75t_L         g10879(.A(new_n10881), .Y(new_n11136));
  NAND2xp33_ASAP7_75t_L     g10880(.A(new_n11134), .B(new_n11130), .Y(new_n11137));
  NOR2xp33_ASAP7_75t_L      g10881(.A(new_n11137), .B(new_n11136), .Y(new_n11138));
  NOR3xp33_ASAP7_75t_L      g10882(.A(new_n11138), .B(new_n11135), .C(new_n10879), .Y(new_n11139));
  INVx1_ASAP7_75t_L         g10883(.A(new_n10879), .Y(new_n11140));
  NAND2xp33_ASAP7_75t_L     g10884(.A(new_n11137), .B(new_n11136), .Y(new_n11141));
  NAND3xp33_ASAP7_75t_L     g10885(.A(new_n10881), .B(new_n11130), .C(new_n11134), .Y(new_n11142));
  AOI21xp33_ASAP7_75t_L     g10886(.A1(new_n11141), .A2(new_n11142), .B(new_n11140), .Y(new_n11143));
  NOR3xp33_ASAP7_75t_L      g10887(.A(new_n10876), .B(new_n11139), .C(new_n11143), .Y(new_n11144));
  OA21x2_ASAP7_75t_L        g10888(.A1(new_n11139), .A2(new_n11143), .B(new_n10876), .Y(new_n11145));
  AOI22xp33_ASAP7_75t_L     g10889(.A1(new_n444), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n471), .Y(new_n11146));
  OAI221xp5_ASAP7_75t_L     g10890(.A1(new_n468), .A2(new_n8762), .B1(new_n469), .B2(new_n9331), .C(new_n11146), .Y(new_n11147));
  XNOR2x2_ASAP7_75t_L       g10891(.A(\a[8] ), .B(new_n11147), .Y(new_n11148));
  OAI21xp33_ASAP7_75t_L     g10892(.A1(new_n11144), .A2(new_n11145), .B(new_n11148), .Y(new_n11149));
  OR3x1_ASAP7_75t_L         g10893(.A(new_n11145), .B(new_n11144), .C(new_n11148), .Y(new_n11150));
  NOR2xp33_ASAP7_75t_L      g10894(.A(new_n9920), .B(new_n429), .Y(new_n11151));
  NAND2xp33_ASAP7_75t_L     g10895(.A(new_n9953), .B(new_n9950), .Y(new_n11152));
  NAND2xp33_ASAP7_75t_L     g10896(.A(\b[57] ), .B(new_n370), .Y(new_n11153));
  OAI221xp5_ASAP7_75t_L     g10897(.A1(new_n343), .A2(new_n9947), .B1(new_n366), .B2(new_n11152), .C(new_n11153), .Y(new_n11154));
  NOR3xp33_ASAP7_75t_L      g10898(.A(new_n11154), .B(new_n11151), .C(new_n338), .Y(new_n11155));
  OA21x2_ASAP7_75t_L        g10899(.A1(new_n11151), .A2(new_n11154), .B(new_n338), .Y(new_n11156));
  NOR2xp33_ASAP7_75t_L      g10900(.A(new_n11155), .B(new_n11156), .Y(new_n11157));
  NAND3xp33_ASAP7_75t_L     g10901(.A(new_n11150), .B(new_n11149), .C(new_n11157), .Y(new_n11158));
  OA21x2_ASAP7_75t_L        g10902(.A1(new_n11144), .A2(new_n11145), .B(new_n11148), .Y(new_n11159));
  NOR3xp33_ASAP7_75t_L      g10903(.A(new_n11145), .B(new_n11148), .C(new_n11144), .Y(new_n11160));
  OR2x4_ASAP7_75t_L         g10904(.A(new_n11155), .B(new_n11156), .Y(new_n11161));
  OAI21xp33_ASAP7_75t_L     g10905(.A1(new_n11160), .A2(new_n11159), .B(new_n11161), .Y(new_n11162));
  NAND2xp33_ASAP7_75t_L     g10906(.A(new_n10828), .B(new_n10826), .Y(new_n11163));
  MAJx2_ASAP7_75t_L         g10907(.A(new_n10834), .B(new_n10831), .C(new_n11163), .Y(new_n11164));
  NAND3xp33_ASAP7_75t_L     g10908(.A(new_n11164), .B(new_n11162), .C(new_n11158), .Y(new_n11165));
  NOR3xp33_ASAP7_75t_L      g10909(.A(new_n11161), .B(new_n11159), .C(new_n11160), .Y(new_n11166));
  AOI21xp33_ASAP7_75t_L     g10910(.A1(new_n11150), .A2(new_n11149), .B(new_n11157), .Y(new_n11167));
  MAJIxp5_ASAP7_75t_L       g10911(.A(new_n10834), .B(new_n10831), .C(new_n11163), .Y(new_n11168));
  OAI21xp33_ASAP7_75t_L     g10912(.A1(new_n11166), .A2(new_n11167), .B(new_n11168), .Y(new_n11169));
  NAND2xp33_ASAP7_75t_L     g10913(.A(\b[61] ), .B(new_n272), .Y(new_n11170));
  NOR2xp33_ASAP7_75t_L      g10914(.A(\b[61] ), .B(\b[62] ), .Y(new_n11171));
  INVx1_ASAP7_75t_L         g10915(.A(\b[62] ), .Y(new_n11172));
  NOR2xp33_ASAP7_75t_L      g10916(.A(new_n10847), .B(new_n11172), .Y(new_n11173));
  NOR2xp33_ASAP7_75t_L      g10917(.A(new_n11171), .B(new_n11173), .Y(new_n11174));
  INVx1_ASAP7_75t_L         g10918(.A(new_n11174), .Y(new_n11175));
  O2A1O1Ixp33_ASAP7_75t_L   g10919(.A1(new_n10250), .A2(new_n10847), .B(new_n10850), .C(new_n11175), .Y(new_n11176));
  A2O1A1O1Ixp25_ASAP7_75t_L g10920(.A1(new_n10252), .A2(new_n10256), .B(new_n10251), .C(new_n10849), .D(new_n10848), .Y(new_n11177));
  NAND2xp33_ASAP7_75t_L     g10921(.A(new_n11175), .B(new_n11177), .Y(new_n11178));
  INVx1_ASAP7_75t_L         g10922(.A(new_n11178), .Y(new_n11179));
  NOR2xp33_ASAP7_75t_L      g10923(.A(new_n11176), .B(new_n11179), .Y(new_n11180));
  NAND2xp33_ASAP7_75t_L     g10924(.A(new_n267), .B(new_n11180), .Y(new_n11181));
  AOI22xp33_ASAP7_75t_L     g10925(.A1(\b[60] ), .A2(new_n282), .B1(\b[62] ), .B2(new_n303), .Y(new_n11182));
  AND4x1_ASAP7_75t_L        g10926(.A(new_n11182), .B(new_n11181), .C(new_n11170), .D(\a[2] ), .Y(new_n11183));
  AOI31xp33_ASAP7_75t_L     g10927(.A1(new_n11181), .A2(new_n11170), .A3(new_n11182), .B(\a[2] ), .Y(new_n11184));
  OR2x4_ASAP7_75t_L         g10928(.A(new_n11184), .B(new_n11183), .Y(new_n11185));
  AOI21xp33_ASAP7_75t_L     g10929(.A1(new_n11165), .A2(new_n11169), .B(new_n11185), .Y(new_n11186));
  NOR3xp33_ASAP7_75t_L      g10930(.A(new_n11167), .B(new_n11166), .C(new_n11168), .Y(new_n11187));
  AOI21xp33_ASAP7_75t_L     g10931(.A1(new_n11162), .A2(new_n11158), .B(new_n11164), .Y(new_n11188));
  NOR2xp33_ASAP7_75t_L      g10932(.A(new_n11184), .B(new_n11183), .Y(new_n11189));
  NOR3xp33_ASAP7_75t_L      g10933(.A(new_n11187), .B(new_n11188), .C(new_n11189), .Y(new_n11190));
  OAI21xp33_ASAP7_75t_L     g10934(.A1(new_n10862), .A2(new_n10861), .B(new_n10840), .Y(new_n11191));
  NOR3xp33_ASAP7_75t_L      g10935(.A(new_n11190), .B(new_n11186), .C(new_n11191), .Y(new_n11192));
  OAI21xp33_ASAP7_75t_L     g10936(.A1(new_n11188), .A2(new_n11187), .B(new_n11189), .Y(new_n11193));
  NAND3xp33_ASAP7_75t_L     g10937(.A(new_n11185), .B(new_n11165), .C(new_n11169), .Y(new_n11194));
  AOI21xp33_ASAP7_75t_L     g10938(.A1(new_n10845), .A2(new_n10858), .B(new_n10860), .Y(new_n11195));
  AOI21xp33_ASAP7_75t_L     g10939(.A1(new_n11194), .A2(new_n11193), .B(new_n11195), .Y(new_n11196));
  NOR2xp33_ASAP7_75t_L      g10940(.A(new_n11196), .B(new_n11192), .Y(new_n11197));
  A2O1A1Ixp33_ASAP7_75t_L   g10941(.A1(new_n10872), .A2(new_n10866), .B(new_n10868), .C(new_n11197), .Y(new_n11198));
  A2O1A1O1Ixp25_ASAP7_75t_L g10942(.A1(new_n10565), .A2(new_n10569), .B(new_n10572), .C(new_n10866), .D(new_n10868), .Y(new_n11199));
  NAND3xp33_ASAP7_75t_L     g10943(.A(new_n11195), .B(new_n11194), .C(new_n11193), .Y(new_n11200));
  OAI21xp33_ASAP7_75t_L     g10944(.A1(new_n11186), .A2(new_n11190), .B(new_n11191), .Y(new_n11201));
  NAND2xp33_ASAP7_75t_L     g10945(.A(new_n11200), .B(new_n11201), .Y(new_n11202));
  NAND2xp33_ASAP7_75t_L     g10946(.A(new_n11202), .B(new_n11199), .Y(new_n11203));
  AND2x2_ASAP7_75t_L        g10947(.A(new_n11198), .B(new_n11203), .Y(\f[62] ));
  NAND3xp33_ASAP7_75t_L     g10948(.A(new_n11119), .B(new_n11123), .C(new_n11133), .Y(new_n11205));
  A2O1A1Ixp33_ASAP7_75t_L   g10949(.A1(new_n11130), .A2(new_n11134), .B(new_n10881), .C(new_n11205), .Y(new_n11206));
  OAI22xp33_ASAP7_75t_L     g10950(.A1(new_n978), .A2(new_n7317), .B1(new_n7616), .B2(new_n977), .Y(new_n11207));
  AOI221xp5_ASAP7_75t_L     g10951(.A1(\b[50] ), .A2(new_n815), .B1(new_n808), .B2(new_n7622), .C(new_n11207), .Y(new_n11208));
  XNOR2x2_ASAP7_75t_L       g10952(.A(new_n806), .B(new_n11208), .Y(new_n11209));
  INVx1_ASAP7_75t_L         g10953(.A(new_n11209), .Y(new_n11210));
  OAI21xp33_ASAP7_75t_L     g10954(.A1(new_n11118), .A2(new_n10883), .B(new_n11120), .Y(new_n11211));
  AOI22xp33_ASAP7_75t_L     g10955(.A1(new_n1076), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1253), .Y(new_n11212));
  OAI221xp5_ASAP7_75t_L     g10956(.A1(new_n1154), .A2(new_n6812), .B1(new_n1156), .B2(new_n6837), .C(new_n11212), .Y(new_n11213));
  XNOR2x2_ASAP7_75t_L       g10957(.A(\a[17] ), .B(new_n11213), .Y(new_n11214));
  AOI31xp33_ASAP7_75t_L     g10958(.A1(new_n11112), .A2(new_n11111), .A3(new_n10793), .B(new_n11100), .Y(new_n11215));
  AOI22xp33_ASAP7_75t_L     g10959(.A1(new_n1360), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n1581), .Y(new_n11216));
  OAI221xp5_ASAP7_75t_L     g10960(.A1(new_n1373), .A2(new_n5829), .B1(new_n1359), .B2(new_n6329), .C(new_n11216), .Y(new_n11217));
  XNOR2x2_ASAP7_75t_L       g10961(.A(\a[20] ), .B(new_n11217), .Y(new_n11218));
  INVx1_ASAP7_75t_L         g10962(.A(new_n11218), .Y(new_n11219));
  AOI22xp33_ASAP7_75t_L     g10963(.A1(new_n1704), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n1837), .Y(new_n11220));
  OAI221xp5_ASAP7_75t_L     g10964(.A1(new_n1699), .A2(new_n5321), .B1(new_n1827), .B2(new_n5346), .C(new_n11220), .Y(new_n11221));
  XNOR2x2_ASAP7_75t_L       g10965(.A(\a[23] ), .B(new_n11221), .Y(new_n11222));
  INVx1_ASAP7_75t_L         g10966(.A(new_n11222), .Y(new_n11223));
  NOR3xp33_ASAP7_75t_L      g10967(.A(new_n11077), .B(new_n11074), .C(new_n11076), .Y(new_n11224));
  INVx1_ASAP7_75t_L         g10968(.A(new_n11224), .Y(new_n11225));
  A2O1A1Ixp33_ASAP7_75t_L   g10969(.A1(new_n10759), .A2(new_n10743), .B(new_n11066), .C(new_n11069), .Y(new_n11226));
  AOI22xp33_ASAP7_75t_L     g10970(.A1(new_n2552), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n2736), .Y(new_n11227));
  OAI221xp5_ASAP7_75t_L     g10971(.A1(new_n2547), .A2(new_n3804), .B1(new_n2734), .B2(new_n4223), .C(new_n11227), .Y(new_n11228));
  XNOR2x2_ASAP7_75t_L       g10972(.A(\a[29] ), .B(new_n11228), .Y(new_n11229));
  INVx1_ASAP7_75t_L         g10973(.A(new_n11229), .Y(new_n11230));
  NOR2xp33_ASAP7_75t_L      g10974(.A(new_n11033), .B(new_n11034), .Y(new_n11231));
  AOI22xp33_ASAP7_75t_L     g10975(.A1(new_n5624), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n5901), .Y(new_n11232));
  OAI221xp5_ASAP7_75t_L     g10976(.A1(new_n5900), .A2(new_n1539), .B1(new_n5892), .B2(new_n1662), .C(new_n11232), .Y(new_n11233));
  XNOR2x2_ASAP7_75t_L       g10977(.A(\a[44] ), .B(new_n11233), .Y(new_n11234));
  NOR2xp33_ASAP7_75t_L      g10978(.A(new_n10975), .B(new_n10979), .Y(new_n11235));
  NAND2xp33_ASAP7_75t_L     g10979(.A(new_n10921), .B(new_n11235), .Y(new_n11236));
  AND3x1_ASAP7_75t_L        g10980(.A(new_n10961), .B(new_n10964), .C(new_n10926), .Y(new_n11237));
  AOI21xp33_ASAP7_75t_L     g10981(.A1(new_n10965), .A2(new_n10923), .B(new_n11237), .Y(new_n11238));
  INVx1_ASAP7_75t_L         g10982(.A(new_n11238), .Y(new_n11239));
  AOI22xp33_ASAP7_75t_L     g10983(.A1(new_n7960), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n8537), .Y(new_n11240));
  OAI221xp5_ASAP7_75t_L     g10984(.A1(new_n8817), .A2(new_n679), .B1(new_n7957), .B2(new_n768), .C(new_n11240), .Y(new_n11241));
  XNOR2x2_ASAP7_75t_L       g10985(.A(new_n7954), .B(new_n11241), .Y(new_n11242));
  A2O1A1O1Ixp25_ASAP7_75t_L g10986(.A1(new_n10643), .A2(new_n10610), .B(new_n10647), .C(new_n10955), .D(new_n10963), .Y(new_n11243));
  AOI22xp33_ASAP7_75t_L     g10987(.A1(new_n9700), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n10027), .Y(new_n11244));
  OAI221xp5_ASAP7_75t_L     g10988(.A1(new_n10024), .A2(new_n354), .B1(new_n9696), .B2(new_n390), .C(new_n11244), .Y(new_n11245));
  XNOR2x2_ASAP7_75t_L       g10989(.A(\a[59] ), .B(new_n11245), .Y(new_n11246));
  NOR2xp33_ASAP7_75t_L      g10990(.A(\a[63] ), .B(new_n10622), .Y(new_n11247));
  INVx1_ASAP7_75t_L         g10991(.A(\a[63] ), .Y(new_n11248));
  NOR2xp33_ASAP7_75t_L      g10992(.A(\a[62] ), .B(new_n11248), .Y(new_n11249));
  A2O1A1Ixp33_ASAP7_75t_L   g10993(.A1(new_n10330), .A2(new_n10331), .B(new_n258), .C(\a[62] ), .Y(new_n11250));
  OR3x1_ASAP7_75t_L         g10994(.A(new_n10941), .B(new_n10634), .C(new_n11250), .Y(new_n11251));
  O2A1O1Ixp33_ASAP7_75t_L   g10995(.A1(new_n11247), .A2(new_n11249), .B(\b[0] ), .C(new_n11251), .Y(new_n11252));
  NOR2xp33_ASAP7_75t_L      g10996(.A(new_n11247), .B(new_n11249), .Y(new_n11253));
  NOR3xp33_ASAP7_75t_L      g10997(.A(new_n10941), .B(new_n11250), .C(new_n10634), .Y(new_n11254));
  NOR3xp33_ASAP7_75t_L      g10998(.A(new_n11254), .B(new_n11253), .C(new_n258), .Y(new_n11255));
  INVx1_ASAP7_75t_L         g10999(.A(new_n10629), .Y(new_n11256));
  NAND3xp33_ASAP7_75t_L     g11000(.A(new_n10332), .B(new_n10628), .C(new_n10631), .Y(new_n11257));
  OAI22xp33_ASAP7_75t_L     g11001(.A1(new_n11257), .A2(new_n261), .B1(new_n298), .B2(new_n10630), .Y(new_n11258));
  AOI221xp5_ASAP7_75t_L     g11002(.A1(\b[2] ), .A2(new_n10632), .B1(new_n406), .B2(new_n11256), .C(new_n11258), .Y(new_n11259));
  XNOR2x2_ASAP7_75t_L       g11003(.A(\a[62] ), .B(new_n11259), .Y(new_n11260));
  OA21x2_ASAP7_75t_L        g11004(.A1(new_n11255), .A2(new_n11252), .B(new_n11260), .Y(new_n11261));
  NOR3xp33_ASAP7_75t_L      g11005(.A(new_n11252), .B(new_n11255), .C(new_n11260), .Y(new_n11262));
  OAI21xp33_ASAP7_75t_L     g11006(.A1(new_n11262), .A2(new_n11261), .B(new_n11246), .Y(new_n11263));
  INVx1_ASAP7_75t_L         g11007(.A(new_n11246), .Y(new_n11264));
  NOR2xp33_ASAP7_75t_L      g11008(.A(new_n11262), .B(new_n11261), .Y(new_n11265));
  NAND2xp33_ASAP7_75t_L     g11009(.A(new_n11264), .B(new_n11265), .Y(new_n11266));
  NOR2xp33_ASAP7_75t_L      g11010(.A(new_n10948), .B(new_n10947), .Y(new_n11267));
  AOI21xp33_ASAP7_75t_L     g11011(.A1(new_n10931), .A2(new_n10949), .B(new_n11267), .Y(new_n11268));
  NAND3xp33_ASAP7_75t_L     g11012(.A(new_n11266), .B(new_n11263), .C(new_n11268), .Y(new_n11269));
  AO21x2_ASAP7_75t_L        g11013(.A1(new_n11263), .A2(new_n11266), .B(new_n11268), .Y(new_n11270));
  AOI22xp33_ASAP7_75t_L     g11014(.A1(new_n8831), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n9115), .Y(new_n11271));
  OAI221xp5_ASAP7_75t_L     g11015(.A1(new_n10343), .A2(new_n488), .B1(new_n10016), .B2(new_n548), .C(new_n11271), .Y(new_n11272));
  NOR2xp33_ASAP7_75t_L      g11016(.A(new_n8826), .B(new_n11272), .Y(new_n11273));
  AND2x2_ASAP7_75t_L        g11017(.A(new_n8826), .B(new_n11272), .Y(new_n11274));
  NOR2xp33_ASAP7_75t_L      g11018(.A(new_n11273), .B(new_n11274), .Y(new_n11275));
  NAND3xp33_ASAP7_75t_L     g11019(.A(new_n11270), .B(new_n11269), .C(new_n11275), .Y(new_n11276));
  AOI21xp33_ASAP7_75t_L     g11020(.A1(new_n11270), .A2(new_n11269), .B(new_n11275), .Y(new_n11277));
  INVx1_ASAP7_75t_L         g11021(.A(new_n11277), .Y(new_n11278));
  AO21x2_ASAP7_75t_L        g11022(.A1(new_n11276), .A2(new_n11278), .B(new_n11243), .Y(new_n11279));
  NAND3xp33_ASAP7_75t_L     g11023(.A(new_n11278), .B(new_n11276), .C(new_n11243), .Y(new_n11280));
  AO21x2_ASAP7_75t_L        g11024(.A1(new_n11280), .A2(new_n11279), .B(new_n11242), .Y(new_n11281));
  NAND3xp33_ASAP7_75t_L     g11025(.A(new_n11279), .B(new_n11280), .C(new_n11242), .Y(new_n11282));
  NAND3xp33_ASAP7_75t_L     g11026(.A(new_n11239), .B(new_n11281), .C(new_n11282), .Y(new_n11283));
  AOI21xp33_ASAP7_75t_L     g11027(.A1(new_n11279), .A2(new_n11280), .B(new_n11242), .Y(new_n11284));
  AND3x1_ASAP7_75t_L        g11028(.A(new_n11279), .B(new_n11280), .C(new_n11242), .Y(new_n11285));
  OAI21xp33_ASAP7_75t_L     g11029(.A1(new_n11284), .A2(new_n11285), .B(new_n11238), .Y(new_n11286));
  AOI22xp33_ASAP7_75t_L     g11030(.A1(new_n7111), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n7391), .Y(new_n11287));
  OAI221xp5_ASAP7_75t_L     g11031(.A1(new_n8558), .A2(new_n869), .B1(new_n8237), .B2(new_n950), .C(new_n11287), .Y(new_n11288));
  XNOR2x2_ASAP7_75t_L       g11032(.A(\a[50] ), .B(new_n11288), .Y(new_n11289));
  NAND3xp33_ASAP7_75t_L     g11033(.A(new_n11283), .B(new_n11286), .C(new_n11289), .Y(new_n11290));
  NOR3xp33_ASAP7_75t_L      g11034(.A(new_n11285), .B(new_n11284), .C(new_n11238), .Y(new_n11291));
  AOI21xp33_ASAP7_75t_L     g11035(.A1(new_n11281), .A2(new_n11282), .B(new_n11239), .Y(new_n11292));
  INVx1_ASAP7_75t_L         g11036(.A(new_n11289), .Y(new_n11293));
  OAI21xp33_ASAP7_75t_L     g11037(.A1(new_n11292), .A2(new_n11291), .B(new_n11293), .Y(new_n11294));
  INVx1_ASAP7_75t_L         g11038(.A(new_n10971), .Y(new_n11295));
  AND3x1_ASAP7_75t_L        g11039(.A(new_n10968), .B(new_n11295), .C(new_n10967), .Y(new_n11296));
  O2A1O1Ixp33_ASAP7_75t_L   g11040(.A1(new_n10976), .A2(new_n10977), .B(new_n10978), .C(new_n11296), .Y(new_n11297));
  NAND3xp33_ASAP7_75t_L     g11041(.A(new_n11297), .B(new_n11294), .C(new_n11290), .Y(new_n11298));
  AO21x2_ASAP7_75t_L        g11042(.A1(new_n11290), .A2(new_n11294), .B(new_n11297), .Y(new_n11299));
  AOI22xp33_ASAP7_75t_L     g11043(.A1(new_n6376), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n6648), .Y(new_n11300));
  OAI221xp5_ASAP7_75t_L     g11044(.A1(new_n6646), .A2(new_n1201), .B1(new_n6636), .B2(new_n1320), .C(new_n11300), .Y(new_n11301));
  XNOR2x2_ASAP7_75t_L       g11045(.A(new_n6371), .B(new_n11301), .Y(new_n11302));
  AO21x2_ASAP7_75t_L        g11046(.A1(new_n11298), .A2(new_n11299), .B(new_n11302), .Y(new_n11303));
  NAND3xp33_ASAP7_75t_L     g11047(.A(new_n11299), .B(new_n11298), .C(new_n11302), .Y(new_n11304));
  NAND2xp33_ASAP7_75t_L     g11048(.A(new_n11304), .B(new_n11303), .Y(new_n11305));
  A2O1A1O1Ixp25_ASAP7_75t_L g11049(.A1(new_n10980), .A2(new_n10983), .B(new_n10988), .C(new_n11236), .D(new_n11305), .Y(new_n11306));
  A2O1A1Ixp33_ASAP7_75t_L   g11050(.A1(new_n10980), .A2(new_n10983), .B(new_n10988), .C(new_n11236), .Y(new_n11307));
  AOI21xp33_ASAP7_75t_L     g11051(.A1(new_n11303), .A2(new_n11304), .B(new_n11307), .Y(new_n11308));
  OR3x1_ASAP7_75t_L         g11052(.A(new_n11306), .B(new_n11234), .C(new_n11308), .Y(new_n11309));
  OAI21xp33_ASAP7_75t_L     g11053(.A1(new_n11308), .A2(new_n11306), .B(new_n11234), .Y(new_n11310));
  OAI211xp5_ASAP7_75t_L     g11054(.A1(new_n11004), .A2(new_n10998), .B(new_n11309), .C(new_n11310), .Y(new_n11311));
  NOR3xp33_ASAP7_75t_L      g11055(.A(new_n11306), .B(new_n11308), .C(new_n11234), .Y(new_n11312));
  OA21x2_ASAP7_75t_L        g11056(.A1(new_n11308), .A2(new_n11306), .B(new_n11234), .Y(new_n11313));
  OAI211xp5_ASAP7_75t_L     g11057(.A1(new_n11312), .A2(new_n11313), .B(new_n10996), .C(new_n10990), .Y(new_n11314));
  AOI22xp33_ASAP7_75t_L     g11058(.A1(new_n4920), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n5167), .Y(new_n11315));
  OAI221xp5_ASAP7_75t_L     g11059(.A1(new_n5154), .A2(new_n1909), .B1(new_n5158), .B2(new_n2477), .C(new_n11315), .Y(new_n11316));
  XNOR2x2_ASAP7_75t_L       g11060(.A(\a[41] ), .B(new_n11316), .Y(new_n11317));
  NAND3xp33_ASAP7_75t_L     g11061(.A(new_n11314), .B(new_n11311), .C(new_n11317), .Y(new_n11318));
  AO21x2_ASAP7_75t_L        g11062(.A1(new_n11311), .A2(new_n11314), .B(new_n11317), .Y(new_n11319));
  A2O1A1O1Ixp25_ASAP7_75t_L g11063(.A1(new_n10694), .A2(new_n10698), .B(new_n10903), .C(new_n11006), .D(new_n11009), .Y(new_n11320));
  NAND3xp33_ASAP7_75t_L     g11064(.A(new_n11319), .B(new_n11318), .C(new_n11320), .Y(new_n11321));
  INVx1_ASAP7_75t_L         g11065(.A(new_n11321), .Y(new_n11322));
  AOI21xp33_ASAP7_75t_L     g11066(.A1(new_n11319), .A2(new_n11318), .B(new_n11320), .Y(new_n11323));
  AOI22xp33_ASAP7_75t_L     g11067(.A1(new_n4283), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n4512), .Y(new_n11324));
  OAI221xp5_ASAP7_75t_L     g11068(.A1(new_n4277), .A2(new_n2348), .B1(new_n4499), .B2(new_n2505), .C(new_n11324), .Y(new_n11325));
  XNOR2x2_ASAP7_75t_L       g11069(.A(\a[38] ), .B(new_n11325), .Y(new_n11326));
  INVx1_ASAP7_75t_L         g11070(.A(new_n11326), .Y(new_n11327));
  NOR3xp33_ASAP7_75t_L      g11071(.A(new_n11322), .B(new_n11323), .C(new_n11327), .Y(new_n11328));
  INVx1_ASAP7_75t_L         g11072(.A(new_n11323), .Y(new_n11329));
  AOI21xp33_ASAP7_75t_L     g11073(.A1(new_n11329), .A2(new_n11321), .B(new_n11326), .Y(new_n11330));
  NOR2xp33_ASAP7_75t_L      g11074(.A(new_n11328), .B(new_n11330), .Y(new_n11331));
  NOR2xp33_ASAP7_75t_L      g11075(.A(new_n11017), .B(new_n11018), .Y(new_n11332));
  NAND2xp33_ASAP7_75t_L     g11076(.A(new_n11019), .B(new_n11332), .Y(new_n11333));
  NAND3xp33_ASAP7_75t_L     g11077(.A(new_n11331), .B(new_n11028), .C(new_n11333), .Y(new_n11334));
  NAND3xp33_ASAP7_75t_L     g11078(.A(new_n11329), .B(new_n11321), .C(new_n11326), .Y(new_n11335));
  OAI21xp33_ASAP7_75t_L     g11079(.A1(new_n11323), .A2(new_n11322), .B(new_n11327), .Y(new_n11336));
  NAND2xp33_ASAP7_75t_L     g11080(.A(new_n11336), .B(new_n11335), .Y(new_n11337));
  A2O1A1Ixp33_ASAP7_75t_L   g11081(.A1(new_n11019), .A2(new_n11332), .B(new_n11034), .C(new_n11337), .Y(new_n11338));
  AOI22xp33_ASAP7_75t_L     g11082(.A1(new_n3633), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n3858), .Y(new_n11339));
  OAI221xp5_ASAP7_75t_L     g11083(.A1(new_n3853), .A2(new_n2688), .B1(new_n3856), .B2(new_n2990), .C(new_n11339), .Y(new_n11340));
  XNOR2x2_ASAP7_75t_L       g11084(.A(\a[35] ), .B(new_n11340), .Y(new_n11341));
  INVx1_ASAP7_75t_L         g11085(.A(new_n11341), .Y(new_n11342));
  AOI21xp33_ASAP7_75t_L     g11086(.A1(new_n11334), .A2(new_n11338), .B(new_n11342), .Y(new_n11343));
  A2O1A1Ixp33_ASAP7_75t_L   g11087(.A1(new_n11020), .A2(new_n11016), .B(new_n11024), .C(new_n11333), .Y(new_n11344));
  NOR2xp33_ASAP7_75t_L      g11088(.A(new_n11344), .B(new_n11337), .Y(new_n11345));
  O2A1O1Ixp33_ASAP7_75t_L   g11089(.A1(new_n11024), .A2(new_n11021), .B(new_n11333), .C(new_n11331), .Y(new_n11346));
  NOR3xp33_ASAP7_75t_L      g11090(.A(new_n11346), .B(new_n11341), .C(new_n11345), .Y(new_n11347));
  NOR2xp33_ASAP7_75t_L      g11091(.A(new_n11343), .B(new_n11347), .Y(new_n11348));
  A2O1A1Ixp33_ASAP7_75t_L   g11092(.A1(new_n11035), .A2(new_n11231), .B(new_n11046), .C(new_n11348), .Y(new_n11349));
  OAI21xp33_ASAP7_75t_L     g11093(.A1(new_n11345), .A2(new_n11346), .B(new_n11341), .Y(new_n11350));
  NAND3xp33_ASAP7_75t_L     g11094(.A(new_n11334), .B(new_n11338), .C(new_n11342), .Y(new_n11351));
  NAND2xp33_ASAP7_75t_L     g11095(.A(new_n11351), .B(new_n11350), .Y(new_n11352));
  NAND2xp33_ASAP7_75t_L     g11096(.A(new_n11035), .B(new_n11231), .Y(new_n11353));
  NAND3xp33_ASAP7_75t_L     g11097(.A(new_n11352), .B(new_n11053), .C(new_n11353), .Y(new_n11354));
  AOI22xp33_ASAP7_75t_L     g11098(.A1(new_n3029), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n3258), .Y(new_n11355));
  OAI221xp5_ASAP7_75t_L     g11099(.A1(new_n3024), .A2(new_n3207), .B1(new_n3256), .B2(new_n3572), .C(new_n11355), .Y(new_n11356));
  XNOR2x2_ASAP7_75t_L       g11100(.A(\a[32] ), .B(new_n11356), .Y(new_n11357));
  NAND3xp33_ASAP7_75t_L     g11101(.A(new_n11349), .B(new_n11354), .C(new_n11357), .Y(new_n11358));
  O2A1O1Ixp33_ASAP7_75t_L   g11102(.A1(new_n11045), .A2(new_n11044), .B(new_n11353), .C(new_n11352), .Y(new_n11359));
  A2O1A1Ixp33_ASAP7_75t_L   g11103(.A1(new_n11036), .A2(new_n11032), .B(new_n11045), .C(new_n11353), .Y(new_n11360));
  NOR2xp33_ASAP7_75t_L      g11104(.A(new_n11360), .B(new_n11348), .Y(new_n11361));
  INVx1_ASAP7_75t_L         g11105(.A(new_n11357), .Y(new_n11362));
  OAI21xp33_ASAP7_75t_L     g11106(.A1(new_n11361), .A2(new_n11359), .B(new_n11362), .Y(new_n11363));
  OAI21xp33_ASAP7_75t_L     g11107(.A1(new_n11060), .A2(new_n10902), .B(new_n11051), .Y(new_n11364));
  AO21x2_ASAP7_75t_L        g11108(.A1(new_n11363), .A2(new_n11358), .B(new_n11364), .Y(new_n11365));
  NAND3xp33_ASAP7_75t_L     g11109(.A(new_n11358), .B(new_n11363), .C(new_n11364), .Y(new_n11366));
  NAND3xp33_ASAP7_75t_L     g11110(.A(new_n11365), .B(new_n11366), .C(new_n11230), .Y(new_n11367));
  AOI21xp33_ASAP7_75t_L     g11111(.A1(new_n11358), .A2(new_n11363), .B(new_n11364), .Y(new_n11368));
  AND3x1_ASAP7_75t_L        g11112(.A(new_n11358), .B(new_n11363), .C(new_n11364), .Y(new_n11369));
  OAI21xp33_ASAP7_75t_L     g11113(.A1(new_n11368), .A2(new_n11369), .B(new_n11229), .Y(new_n11370));
  AOI21xp33_ASAP7_75t_L     g11114(.A1(new_n11370), .A2(new_n11367), .B(new_n11226), .Y(new_n11371));
  A2O1A1O1Ixp25_ASAP7_75t_L g11115(.A1(new_n10593), .A2(new_n10746), .B(new_n10756), .C(new_n11070), .D(new_n11062), .Y(new_n11372));
  NOR3xp33_ASAP7_75t_L      g11116(.A(new_n11369), .B(new_n11368), .C(new_n11229), .Y(new_n11373));
  AOI21xp33_ASAP7_75t_L     g11117(.A1(new_n11365), .A2(new_n11366), .B(new_n11230), .Y(new_n11374));
  NOR3xp33_ASAP7_75t_L      g11118(.A(new_n11373), .B(new_n11374), .C(new_n11372), .Y(new_n11375));
  AOI22xp33_ASAP7_75t_L     g11119(.A1(new_n2114), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n2259), .Y(new_n11376));
  OAI221xp5_ASAP7_75t_L     g11120(.A1(new_n2109), .A2(new_n4632), .B1(new_n2257), .B2(new_n4858), .C(new_n11376), .Y(new_n11377));
  XNOR2x2_ASAP7_75t_L       g11121(.A(\a[26] ), .B(new_n11377), .Y(new_n11378));
  OAI21xp33_ASAP7_75t_L     g11122(.A1(new_n11371), .A2(new_n11375), .B(new_n11378), .Y(new_n11379));
  OAI21xp33_ASAP7_75t_L     g11123(.A1(new_n11374), .A2(new_n11373), .B(new_n11372), .Y(new_n11380));
  NAND3xp33_ASAP7_75t_L     g11124(.A(new_n11226), .B(new_n11367), .C(new_n11370), .Y(new_n11381));
  INVx1_ASAP7_75t_L         g11125(.A(new_n11378), .Y(new_n11382));
  NAND3xp33_ASAP7_75t_L     g11126(.A(new_n11381), .B(new_n11380), .C(new_n11382), .Y(new_n11383));
  NAND2xp33_ASAP7_75t_L     g11127(.A(new_n11383), .B(new_n11379), .Y(new_n11384));
  A2O1A1O1Ixp25_ASAP7_75t_L g11128(.A1(new_n10768), .A2(new_n11081), .B(new_n11086), .C(new_n11225), .D(new_n11384), .Y(new_n11385));
  A2O1A1Ixp33_ASAP7_75t_L   g11129(.A1(new_n10768), .A2(new_n11081), .B(new_n11086), .C(new_n11225), .Y(new_n11386));
  AOI21xp33_ASAP7_75t_L     g11130(.A1(new_n11383), .A2(new_n11379), .B(new_n11386), .Y(new_n11387));
  OAI21xp33_ASAP7_75t_L     g11131(.A1(new_n11387), .A2(new_n11385), .B(new_n11223), .Y(new_n11388));
  NAND3xp33_ASAP7_75t_L     g11132(.A(new_n11386), .B(new_n11379), .C(new_n11383), .Y(new_n11389));
  O2A1O1Ixp33_ASAP7_75t_L   g11133(.A1(new_n11084), .A2(new_n11085), .B(new_n11082), .C(new_n11224), .Y(new_n11390));
  NAND2xp33_ASAP7_75t_L     g11134(.A(new_n11384), .B(new_n11390), .Y(new_n11391));
  NAND3xp33_ASAP7_75t_L     g11135(.A(new_n11389), .B(new_n11222), .C(new_n11391), .Y(new_n11392));
  AOI221xp5_ASAP7_75t_L     g11136(.A1(new_n11095), .A2(new_n11097), .B1(new_n11392), .B2(new_n11388), .C(new_n11103), .Y(new_n11393));
  A2O1A1Ixp33_ASAP7_75t_L   g11137(.A1(new_n10499), .A2(new_n10782), .B(new_n10787), .C(new_n10895), .Y(new_n11394));
  NAND2xp33_ASAP7_75t_L     g11138(.A(new_n11392), .B(new_n11388), .Y(new_n11395));
  O2A1O1Ixp33_ASAP7_75t_L   g11139(.A1(new_n11394), .A2(new_n11104), .B(new_n11091), .C(new_n11395), .Y(new_n11396));
  OAI21xp33_ASAP7_75t_L     g11140(.A1(new_n11393), .A2(new_n11396), .B(new_n11219), .Y(new_n11397));
  AOI21xp33_ASAP7_75t_L     g11141(.A1(new_n11097), .A2(new_n11095), .B(new_n11103), .Y(new_n11398));
  NAND2xp33_ASAP7_75t_L     g11142(.A(new_n11398), .B(new_n11395), .Y(new_n11399));
  AOI21xp33_ASAP7_75t_L     g11143(.A1(new_n11389), .A2(new_n11391), .B(new_n11222), .Y(new_n11400));
  NOR3xp33_ASAP7_75t_L      g11144(.A(new_n11385), .B(new_n11387), .C(new_n11223), .Y(new_n11401));
  NOR2xp33_ASAP7_75t_L      g11145(.A(new_n11400), .B(new_n11401), .Y(new_n11402));
  A2O1A1Ixp33_ASAP7_75t_L   g11146(.A1(new_n11095), .A2(new_n11097), .B(new_n11103), .C(new_n11402), .Y(new_n11403));
  NAND3xp33_ASAP7_75t_L     g11147(.A(new_n11403), .B(new_n11399), .C(new_n11218), .Y(new_n11404));
  AO21x2_ASAP7_75t_L        g11148(.A1(new_n11404), .A2(new_n11397), .B(new_n11215), .Y(new_n11405));
  NAND3xp33_ASAP7_75t_L     g11149(.A(new_n11215), .B(new_n11404), .C(new_n11397), .Y(new_n11406));
  AOI21xp33_ASAP7_75t_L     g11150(.A1(new_n11405), .A2(new_n11406), .B(new_n11214), .Y(new_n11407));
  AND3x1_ASAP7_75t_L        g11151(.A(new_n11405), .B(new_n11406), .C(new_n11214), .Y(new_n11408));
  OAI21xp33_ASAP7_75t_L     g11152(.A1(new_n11407), .A2(new_n11408), .B(new_n11211), .Y(new_n11409));
  A2O1A1O1Ixp25_ASAP7_75t_L g11153(.A1(new_n10803), .A2(new_n10811), .B(new_n10882), .C(new_n11121), .D(new_n11114), .Y(new_n11410));
  AO21x2_ASAP7_75t_L        g11154(.A1(new_n11406), .A2(new_n11405), .B(new_n11214), .Y(new_n11411));
  NAND3xp33_ASAP7_75t_L     g11155(.A(new_n11405), .B(new_n11214), .C(new_n11406), .Y(new_n11412));
  NAND3xp33_ASAP7_75t_L     g11156(.A(new_n11410), .B(new_n11411), .C(new_n11412), .Y(new_n11413));
  NAND3xp33_ASAP7_75t_L     g11157(.A(new_n11413), .B(new_n11409), .C(new_n11210), .Y(new_n11414));
  AOI21xp33_ASAP7_75t_L     g11158(.A1(new_n11411), .A2(new_n11412), .B(new_n11410), .Y(new_n11415));
  NOR3xp33_ASAP7_75t_L      g11159(.A(new_n11211), .B(new_n11408), .C(new_n11407), .Y(new_n11416));
  OAI21xp33_ASAP7_75t_L     g11160(.A1(new_n11415), .A2(new_n11416), .B(new_n11209), .Y(new_n11417));
  AND2x2_ASAP7_75t_L        g11161(.A(new_n11414), .B(new_n11417), .Y(new_n11418));
  NAND2xp33_ASAP7_75t_L     g11162(.A(new_n11206), .B(new_n11418), .Y(new_n11419));
  NAND2xp33_ASAP7_75t_L     g11163(.A(new_n11414), .B(new_n11417), .Y(new_n11420));
  NAND3xp33_ASAP7_75t_L     g11164(.A(new_n11141), .B(new_n11205), .C(new_n11420), .Y(new_n11421));
  OAI22xp33_ASAP7_75t_L     g11165(.A1(new_n706), .A2(new_n7900), .B1(new_n8458), .B2(new_n580), .Y(new_n11422));
  AOI221xp5_ASAP7_75t_L     g11166(.A1(\b[53] ), .A2(new_n584), .B1(new_n578), .B2(new_n8464), .C(new_n11422), .Y(new_n11423));
  XNOR2x2_ASAP7_75t_L       g11167(.A(new_n574), .B(new_n11423), .Y(new_n11424));
  NAND3xp33_ASAP7_75t_L     g11168(.A(new_n11421), .B(new_n11419), .C(new_n11424), .Y(new_n11425));
  A2O1A1O1Ixp25_ASAP7_75t_L g11169(.A1(new_n11130), .A2(new_n11134), .B(new_n10881), .C(new_n11205), .D(new_n11420), .Y(new_n11426));
  NOR2xp33_ASAP7_75t_L      g11170(.A(new_n11206), .B(new_n11418), .Y(new_n11427));
  INVx1_ASAP7_75t_L         g11171(.A(new_n11424), .Y(new_n11428));
  OAI21xp33_ASAP7_75t_L     g11172(.A1(new_n11426), .A2(new_n11427), .B(new_n11428), .Y(new_n11429));
  NAND2xp33_ASAP7_75t_L     g11173(.A(new_n11429), .B(new_n11425), .Y(new_n11430));
  NAND3xp33_ASAP7_75t_L     g11174(.A(new_n11141), .B(new_n11140), .C(new_n11142), .Y(new_n11431));
  OAI21xp33_ASAP7_75t_L     g11175(.A1(new_n11143), .A2(new_n10876), .B(new_n11431), .Y(new_n11432));
  NOR2xp33_ASAP7_75t_L      g11176(.A(new_n11432), .B(new_n11430), .Y(new_n11433));
  AO21x2_ASAP7_75t_L        g11177(.A1(new_n10544), .A2(new_n10547), .B(new_n10573), .Y(new_n11434));
  OAI21xp33_ASAP7_75t_L     g11178(.A1(new_n11135), .A2(new_n11138), .B(new_n10879), .Y(new_n11435));
  A2O1A1O1Ixp25_ASAP7_75t_L g11179(.A1(new_n10875), .A2(new_n11434), .B(new_n10824), .C(new_n11435), .D(new_n11139), .Y(new_n11436));
  AOI21xp33_ASAP7_75t_L     g11180(.A1(new_n11429), .A2(new_n11425), .B(new_n11436), .Y(new_n11437));
  AOI22xp33_ASAP7_75t_L     g11181(.A1(new_n444), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n471), .Y(new_n11438));
  OAI221xp5_ASAP7_75t_L     g11182(.A1(new_n468), .A2(new_n9323), .B1(new_n469), .B2(new_n9627), .C(new_n11438), .Y(new_n11439));
  XNOR2x2_ASAP7_75t_L       g11183(.A(\a[8] ), .B(new_n11439), .Y(new_n11440));
  INVx1_ASAP7_75t_L         g11184(.A(new_n11440), .Y(new_n11441));
  NOR3xp33_ASAP7_75t_L      g11185(.A(new_n11433), .B(new_n11437), .C(new_n11441), .Y(new_n11442));
  NAND3xp33_ASAP7_75t_L     g11186(.A(new_n11436), .B(new_n11429), .C(new_n11425), .Y(new_n11443));
  NAND2xp33_ASAP7_75t_L     g11187(.A(new_n11432), .B(new_n11430), .Y(new_n11444));
  AOI21xp33_ASAP7_75t_L     g11188(.A1(new_n11444), .A2(new_n11443), .B(new_n11440), .Y(new_n11445));
  INVx1_ASAP7_75t_L         g11189(.A(new_n10258), .Y(new_n11446));
  AOI22xp33_ASAP7_75t_L     g11190(.A1(new_n344), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n370), .Y(new_n11447));
  OAI21xp33_ASAP7_75t_L     g11191(.A1(new_n366), .A2(new_n11446), .B(new_n11447), .Y(new_n11448));
  AOI21xp33_ASAP7_75t_L     g11192(.A1(new_n347), .A2(\b[59] ), .B(new_n11448), .Y(new_n11449));
  NAND2xp33_ASAP7_75t_L     g11193(.A(\a[5] ), .B(new_n11449), .Y(new_n11450));
  A2O1A1Ixp33_ASAP7_75t_L   g11194(.A1(\b[59] ), .A2(new_n347), .B(new_n11448), .C(new_n338), .Y(new_n11451));
  AND2x2_ASAP7_75t_L        g11195(.A(new_n11451), .B(new_n11450), .Y(new_n11452));
  OAI21xp33_ASAP7_75t_L     g11196(.A1(new_n11445), .A2(new_n11442), .B(new_n11452), .Y(new_n11453));
  NAND3xp33_ASAP7_75t_L     g11197(.A(new_n11444), .B(new_n11443), .C(new_n11440), .Y(new_n11454));
  OAI21xp33_ASAP7_75t_L     g11198(.A1(new_n11437), .A2(new_n11433), .B(new_n11441), .Y(new_n11455));
  NAND2xp33_ASAP7_75t_L     g11199(.A(new_n11451), .B(new_n11450), .Y(new_n11456));
  NAND3xp33_ASAP7_75t_L     g11200(.A(new_n11455), .B(new_n11456), .C(new_n11454), .Y(new_n11457));
  NAND2xp33_ASAP7_75t_L     g11201(.A(new_n11149), .B(new_n11158), .Y(new_n11458));
  NAND3xp33_ASAP7_75t_L     g11202(.A(new_n11453), .B(new_n11457), .C(new_n11458), .Y(new_n11459));
  AOI21xp33_ASAP7_75t_L     g11203(.A1(new_n11455), .A2(new_n11454), .B(new_n11456), .Y(new_n11460));
  NOR3xp33_ASAP7_75t_L      g11204(.A(new_n11452), .B(new_n11445), .C(new_n11442), .Y(new_n11461));
  O2A1O1Ixp33_ASAP7_75t_L   g11205(.A1(new_n11144), .A2(new_n11145), .B(new_n11148), .C(new_n11166), .Y(new_n11462));
  OAI21xp33_ASAP7_75t_L     g11206(.A1(new_n11460), .A2(new_n11461), .B(new_n11462), .Y(new_n11463));
  INVx1_ASAP7_75t_L         g11207(.A(new_n10251), .Y(new_n11464));
  A2O1A1Ixp33_ASAP7_75t_L   g11208(.A1(new_n9950), .A2(new_n10248), .B(new_n10249), .C(new_n11464), .Y(new_n11465));
  A2O1A1O1Ixp25_ASAP7_75t_L g11209(.A1(new_n10849), .A2(new_n11465), .B(new_n10848), .C(new_n11174), .D(new_n11173), .Y(new_n11466));
  NOR2xp33_ASAP7_75t_L      g11210(.A(\b[63] ), .B(new_n11172), .Y(new_n11467));
  INVx1_ASAP7_75t_L         g11211(.A(\b[63] ), .Y(new_n11468));
  NOR2xp33_ASAP7_75t_L      g11212(.A(\b[62] ), .B(new_n11468), .Y(new_n11469));
  OAI21xp33_ASAP7_75t_L     g11213(.A1(new_n11467), .A2(new_n11469), .B(new_n11466), .Y(new_n11470));
  INVx1_ASAP7_75t_L         g11214(.A(new_n11177), .Y(new_n11471));
  NOR2xp33_ASAP7_75t_L      g11215(.A(new_n11467), .B(new_n11469), .Y(new_n11472));
  A2O1A1Ixp33_ASAP7_75t_L   g11216(.A1(new_n11471), .A2(new_n11174), .B(new_n11173), .C(new_n11472), .Y(new_n11473));
  NOR2xp33_ASAP7_75t_L      g11217(.A(new_n11172), .B(new_n291), .Y(new_n11474));
  AOI221xp5_ASAP7_75t_L     g11218(.A1(\b[61] ), .A2(new_n282), .B1(\b[63] ), .B2(new_n303), .C(new_n11474), .Y(new_n11475));
  A2O1A1Ixp33_ASAP7_75t_L   g11219(.A1(new_n11470), .A2(new_n11473), .B(new_n268), .C(new_n11475), .Y(new_n11476));
  NOR2xp33_ASAP7_75t_L      g11220(.A(new_n262), .B(new_n11476), .Y(new_n11477));
  A2O1A1O1Ixp25_ASAP7_75t_L g11221(.A1(new_n11473), .A2(new_n11470), .B(new_n268), .C(new_n11475), .D(\a[2] ), .Y(new_n11478));
  NOR2xp33_ASAP7_75t_L      g11222(.A(new_n11478), .B(new_n11477), .Y(new_n11479));
  NAND3xp33_ASAP7_75t_L     g11223(.A(new_n11463), .B(new_n11459), .C(new_n11479), .Y(new_n11480));
  NOR3xp33_ASAP7_75t_L      g11224(.A(new_n11461), .B(new_n11460), .C(new_n11462), .Y(new_n11481));
  AOI21xp33_ASAP7_75t_L     g11225(.A1(new_n11453), .A2(new_n11457), .B(new_n11458), .Y(new_n11482));
  INVx1_ASAP7_75t_L         g11226(.A(new_n11479), .Y(new_n11483));
  OAI21xp33_ASAP7_75t_L     g11227(.A1(new_n11482), .A2(new_n11481), .B(new_n11483), .Y(new_n11484));
  O2A1O1Ixp33_ASAP7_75t_L   g11228(.A1(new_n11183), .A2(new_n11184), .B(new_n11165), .C(new_n11188), .Y(new_n11485));
  AO21x2_ASAP7_75t_L        g11229(.A1(new_n11480), .A2(new_n11484), .B(new_n11485), .Y(new_n11486));
  NAND3xp33_ASAP7_75t_L     g11230(.A(new_n11484), .B(new_n11480), .C(new_n11485), .Y(new_n11487));
  NAND2xp33_ASAP7_75t_L     g11231(.A(new_n11487), .B(new_n11486), .Y(new_n11488));
  O2A1O1Ixp33_ASAP7_75t_L   g11232(.A1(new_n11199), .A2(new_n11196), .B(new_n11200), .C(new_n11488), .Y(new_n11489));
  OAI21xp33_ASAP7_75t_L     g11233(.A1(new_n11202), .A2(new_n11199), .B(new_n11200), .Y(new_n11490));
  AOI21xp33_ASAP7_75t_L     g11234(.A1(new_n11484), .A2(new_n11480), .B(new_n11485), .Y(new_n11491));
  AND3x1_ASAP7_75t_L        g11235(.A(new_n11484), .B(new_n11485), .C(new_n11480), .Y(new_n11492));
  NOR2xp33_ASAP7_75t_L      g11236(.A(new_n11491), .B(new_n11492), .Y(new_n11493));
  NOR2xp33_ASAP7_75t_L      g11237(.A(new_n11493), .B(new_n11490), .Y(new_n11494));
  NOR2xp33_ASAP7_75t_L      g11238(.A(new_n11489), .B(new_n11494), .Y(\f[63] ));
  A2O1A1Ixp33_ASAP7_75t_L   g11239(.A1(new_n11198), .A2(new_n11200), .B(new_n11488), .C(new_n11486), .Y(new_n11496));
  INVx1_ASAP7_75t_L         g11240(.A(new_n11173), .Y(new_n11497));
  INVx1_ASAP7_75t_L         g11241(.A(new_n11176), .Y(new_n11498));
  OAI21xp33_ASAP7_75t_L     g11242(.A1(\b[62] ), .A2(new_n11468), .B(new_n11466), .Y(new_n11499));
  A2O1A1Ixp33_ASAP7_75t_L   g11243(.A1(new_n11498), .A2(new_n11497), .B(new_n11467), .C(new_n11499), .Y(new_n11500));
  NAND2xp33_ASAP7_75t_L     g11244(.A(\b[63] ), .B(new_n272), .Y(new_n11501));
  OAI221xp5_ASAP7_75t_L     g11245(.A1(new_n283), .A2(new_n11172), .B1(new_n268), .B2(new_n11500), .C(new_n11501), .Y(new_n11502));
  XNOR2x2_ASAP7_75t_L       g11246(.A(\a[2] ), .B(new_n11502), .Y(new_n11503));
  NOR3xp33_ASAP7_75t_L      g11247(.A(new_n11433), .B(new_n11437), .C(new_n11440), .Y(new_n11504));
  O2A1O1Ixp33_ASAP7_75t_L   g11248(.A1(new_n11445), .A2(new_n11442), .B(new_n11456), .C(new_n11504), .Y(new_n11505));
  XNOR2x2_ASAP7_75t_L       g11249(.A(new_n11206), .B(new_n11420), .Y(new_n11506));
  NAND2xp33_ASAP7_75t_L     g11250(.A(new_n11428), .B(new_n11506), .Y(new_n11507));
  A2O1A1Ixp33_ASAP7_75t_L   g11251(.A1(new_n11429), .A2(new_n11425), .B(new_n11436), .C(new_n11507), .Y(new_n11508));
  AOI22xp33_ASAP7_75t_L     g11252(.A1(\b[53] ), .A2(new_n651), .B1(\b[55] ), .B2(new_n581), .Y(new_n11509));
  OAI221xp5_ASAP7_75t_L     g11253(.A1(new_n821), .A2(new_n8458), .B1(new_n577), .B2(new_n8768), .C(new_n11509), .Y(new_n11510));
  XNOR2x2_ASAP7_75t_L       g11254(.A(\a[11] ), .B(new_n11510), .Y(new_n11511));
  INVx1_ASAP7_75t_L         g11255(.A(new_n11205), .Y(new_n11512));
  INVx1_ASAP7_75t_L         g11256(.A(new_n11414), .Y(new_n11513));
  A2O1A1O1Ixp25_ASAP7_75t_L g11257(.A1(new_n11137), .A2(new_n11136), .B(new_n11512), .C(new_n11417), .D(new_n11513), .Y(new_n11514));
  AOI22xp33_ASAP7_75t_L     g11258(.A1(new_n811), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n900), .Y(new_n11515));
  OAI221xp5_ASAP7_75t_L     g11259(.A1(new_n904), .A2(new_n7616), .B1(new_n898), .B2(new_n7906), .C(new_n11515), .Y(new_n11516));
  INVx1_ASAP7_75t_L         g11260(.A(new_n11516), .Y(new_n11517));
  NAND2xp33_ASAP7_75t_L     g11261(.A(\a[14] ), .B(new_n11517), .Y(new_n11518));
  NAND2xp33_ASAP7_75t_L     g11262(.A(new_n806), .B(new_n11516), .Y(new_n11519));
  NAND2xp33_ASAP7_75t_L     g11263(.A(new_n11519), .B(new_n11518), .Y(new_n11520));
  NAND2xp33_ASAP7_75t_L     g11264(.A(new_n11406), .B(new_n11405), .Y(new_n11521));
  MAJIxp5_ASAP7_75t_L       g11265(.A(new_n11410), .B(new_n11214), .C(new_n11521), .Y(new_n11522));
  AOI22xp33_ASAP7_75t_L     g11266(.A1(new_n1076), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1253), .Y(new_n11523));
  OAI221xp5_ASAP7_75t_L     g11267(.A1(new_n1154), .A2(new_n6830), .B1(new_n1156), .B2(new_n7323), .C(new_n11523), .Y(new_n11524));
  XNOR2x2_ASAP7_75t_L       g11268(.A(\a[17] ), .B(new_n11524), .Y(new_n11525));
  NAND3xp33_ASAP7_75t_L     g11269(.A(new_n11403), .B(new_n11399), .C(new_n11219), .Y(new_n11526));
  A2O1A1Ixp33_ASAP7_75t_L   g11270(.A1(new_n11404), .A2(new_n11397), .B(new_n11215), .C(new_n11526), .Y(new_n11527));
  AOI22xp33_ASAP7_75t_L     g11271(.A1(new_n1360), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n1581), .Y(new_n11528));
  OAI221xp5_ASAP7_75t_L     g11272(.A1(new_n1373), .A2(new_n6321), .B1(new_n1359), .B2(new_n6573), .C(new_n11528), .Y(new_n11529));
  XNOR2x2_ASAP7_75t_L       g11273(.A(\a[20] ), .B(new_n11529), .Y(new_n11530));
  NOR3xp33_ASAP7_75t_L      g11274(.A(new_n11385), .B(new_n11387), .C(new_n11222), .Y(new_n11531));
  MAJIxp5_ASAP7_75t_L       g11275(.A(new_n11268), .B(new_n11264), .C(new_n11265), .Y(new_n11532));
  INVx1_ASAP7_75t_L         g11276(.A(new_n11253), .Y(new_n11533));
  NOR2xp33_ASAP7_75t_L      g11277(.A(new_n10622), .B(new_n11248), .Y(new_n11534));
  INVx1_ASAP7_75t_L         g11278(.A(new_n11534), .Y(new_n11535));
  NOR2xp33_ASAP7_75t_L      g11279(.A(new_n258), .B(new_n11535), .Y(new_n11536));
  OAI22xp33_ASAP7_75t_L     g11280(.A1(new_n11257), .A2(new_n276), .B1(new_n324), .B2(new_n10630), .Y(new_n11537));
  AOI21xp33_ASAP7_75t_L     g11281(.A1(new_n329), .A2(new_n11256), .B(new_n11537), .Y(new_n11538));
  OA211x2_ASAP7_75t_L       g11282(.A1(new_n10937), .A2(new_n298), .B(new_n11538), .C(\a[62] ), .Y(new_n11539));
  O2A1O1Ixp33_ASAP7_75t_L   g11283(.A1(new_n298), .A2(new_n10937), .B(new_n11538), .C(\a[62] ), .Y(new_n11540));
  NOR2xp33_ASAP7_75t_L      g11284(.A(new_n11540), .B(new_n11539), .Y(new_n11541));
  A2O1A1Ixp33_ASAP7_75t_L   g11285(.A1(new_n11533), .A2(\b[1] ), .B(new_n11536), .C(new_n11541), .Y(new_n11542));
  O2A1O1Ixp33_ASAP7_75t_L   g11286(.A1(new_n11247), .A2(new_n11249), .B(\b[1] ), .C(new_n11536), .Y(new_n11543));
  OAI21xp33_ASAP7_75t_L     g11287(.A1(new_n11540), .A2(new_n11539), .B(new_n11543), .Y(new_n11544));
  NOR3xp33_ASAP7_75t_L      g11288(.A(new_n11251), .B(new_n11253), .C(new_n258), .Y(new_n11545));
  O2A1O1Ixp33_ASAP7_75t_L   g11289(.A1(new_n11255), .A2(new_n11252), .B(new_n11260), .C(new_n11545), .Y(new_n11546));
  NAND3xp33_ASAP7_75t_L     g11290(.A(new_n11546), .B(new_n11544), .C(new_n11542), .Y(new_n11547));
  AO21x2_ASAP7_75t_L        g11291(.A1(new_n11542), .A2(new_n11544), .B(new_n11546), .Y(new_n11548));
  AOI22xp33_ASAP7_75t_L     g11292(.A1(new_n9700), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n10027), .Y(new_n11549));
  OAI221xp5_ASAP7_75t_L     g11293(.A1(new_n10024), .A2(new_n418), .B1(new_n9696), .B2(new_n425), .C(new_n11549), .Y(new_n11550));
  XNOR2x2_ASAP7_75t_L       g11294(.A(new_n9693), .B(new_n11550), .Y(new_n11551));
  AOI21xp33_ASAP7_75t_L     g11295(.A1(new_n11548), .A2(new_n11547), .B(new_n11551), .Y(new_n11552));
  NAND3xp33_ASAP7_75t_L     g11296(.A(new_n11548), .B(new_n11547), .C(new_n11551), .Y(new_n11553));
  INVx1_ASAP7_75t_L         g11297(.A(new_n11553), .Y(new_n11554));
  NOR3xp33_ASAP7_75t_L      g11298(.A(new_n11554), .B(new_n11532), .C(new_n11552), .Y(new_n11555));
  INVx1_ASAP7_75t_L         g11299(.A(new_n11555), .Y(new_n11556));
  OAI21xp33_ASAP7_75t_L     g11300(.A1(new_n11552), .A2(new_n11554), .B(new_n11532), .Y(new_n11557));
  AOI22xp33_ASAP7_75t_L     g11301(.A1(new_n8831), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n9115), .Y(new_n11558));
  OAI221xp5_ASAP7_75t_L     g11302(.A1(new_n10343), .A2(new_n540), .B1(new_n10016), .B2(new_n624), .C(new_n11558), .Y(new_n11559));
  XNOR2x2_ASAP7_75t_L       g11303(.A(\a[56] ), .B(new_n11559), .Y(new_n11560));
  NAND3xp33_ASAP7_75t_L     g11304(.A(new_n11556), .B(new_n11557), .C(new_n11560), .Y(new_n11561));
  OA21x2_ASAP7_75t_L        g11305(.A1(new_n11552), .A2(new_n11554), .B(new_n11532), .Y(new_n11562));
  INVx1_ASAP7_75t_L         g11306(.A(new_n11560), .Y(new_n11563));
  OAI21xp33_ASAP7_75t_L     g11307(.A1(new_n11555), .A2(new_n11562), .B(new_n11563), .Y(new_n11564));
  NAND2xp33_ASAP7_75t_L     g11308(.A(new_n11269), .B(new_n11270), .Y(new_n11565));
  MAJx2_ASAP7_75t_L         g11309(.A(new_n11243), .B(new_n11565), .C(new_n11275), .Y(new_n11566));
  NAND3xp33_ASAP7_75t_L     g11310(.A(new_n11566), .B(new_n11561), .C(new_n11564), .Y(new_n11567));
  INVx1_ASAP7_75t_L         g11311(.A(new_n11567), .Y(new_n11568));
  AOI21xp33_ASAP7_75t_L     g11312(.A1(new_n11561), .A2(new_n11564), .B(new_n11566), .Y(new_n11569));
  AOI22xp33_ASAP7_75t_L     g11313(.A1(new_n7960), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n8537), .Y(new_n11570));
  OAI221xp5_ASAP7_75t_L     g11314(.A1(new_n8817), .A2(new_n760), .B1(new_n7957), .B2(new_n790), .C(new_n11570), .Y(new_n11571));
  XNOR2x2_ASAP7_75t_L       g11315(.A(new_n7954), .B(new_n11571), .Y(new_n11572));
  INVx1_ASAP7_75t_L         g11316(.A(new_n11572), .Y(new_n11573));
  OAI21xp33_ASAP7_75t_L     g11317(.A1(new_n11569), .A2(new_n11568), .B(new_n11573), .Y(new_n11574));
  INVx1_ASAP7_75t_L         g11318(.A(new_n11569), .Y(new_n11575));
  NAND3xp33_ASAP7_75t_L     g11319(.A(new_n11575), .B(new_n11567), .C(new_n11572), .Y(new_n11576));
  A2O1A1Ixp33_ASAP7_75t_L   g11320(.A1(new_n10967), .A2(new_n10966), .B(new_n11284), .C(new_n11282), .Y(new_n11577));
  NAND3xp33_ASAP7_75t_L     g11321(.A(new_n11574), .B(new_n11576), .C(new_n11577), .Y(new_n11578));
  AOI21xp33_ASAP7_75t_L     g11322(.A1(new_n11575), .A2(new_n11567), .B(new_n11572), .Y(new_n11579));
  NOR3xp33_ASAP7_75t_L      g11323(.A(new_n11568), .B(new_n11569), .C(new_n11573), .Y(new_n11580));
  A2O1A1O1Ixp25_ASAP7_75t_L g11324(.A1(new_n10965), .A2(new_n10923), .B(new_n11237), .C(new_n11281), .D(new_n11285), .Y(new_n11581));
  OAI21xp33_ASAP7_75t_L     g11325(.A1(new_n11579), .A2(new_n11580), .B(new_n11581), .Y(new_n11582));
  AOI22xp33_ASAP7_75t_L     g11326(.A1(new_n7111), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n7391), .Y(new_n11583));
  OAI221xp5_ASAP7_75t_L     g11327(.A1(new_n8558), .A2(new_n942), .B1(new_n8237), .B2(new_n1035), .C(new_n11583), .Y(new_n11584));
  XNOR2x2_ASAP7_75t_L       g11328(.A(\a[50] ), .B(new_n11584), .Y(new_n11585));
  NAND3xp33_ASAP7_75t_L     g11329(.A(new_n11582), .B(new_n11578), .C(new_n11585), .Y(new_n11586));
  NOR3xp33_ASAP7_75t_L      g11330(.A(new_n11581), .B(new_n11580), .C(new_n11579), .Y(new_n11587));
  AOI21xp33_ASAP7_75t_L     g11331(.A1(new_n11574), .A2(new_n11576), .B(new_n11577), .Y(new_n11588));
  INVx1_ASAP7_75t_L         g11332(.A(new_n11585), .Y(new_n11589));
  OAI21xp33_ASAP7_75t_L     g11333(.A1(new_n11588), .A2(new_n11587), .B(new_n11589), .Y(new_n11590));
  AND2x2_ASAP7_75t_L        g11334(.A(new_n11586), .B(new_n11590), .Y(new_n11591));
  NOR2xp33_ASAP7_75t_L      g11335(.A(new_n11292), .B(new_n11291), .Y(new_n11592));
  NAND2xp33_ASAP7_75t_L     g11336(.A(new_n11293), .B(new_n11592), .Y(new_n11593));
  A2O1A1Ixp33_ASAP7_75t_L   g11337(.A1(new_n11294), .A2(new_n11290), .B(new_n11297), .C(new_n11593), .Y(new_n11594));
  INVx1_ASAP7_75t_L         g11338(.A(new_n11594), .Y(new_n11595));
  NAND2xp33_ASAP7_75t_L     g11339(.A(new_n11591), .B(new_n11595), .Y(new_n11596));
  AOI21xp33_ASAP7_75t_L     g11340(.A1(new_n11294), .A2(new_n11290), .B(new_n11297), .Y(new_n11597));
  NAND2xp33_ASAP7_75t_L     g11341(.A(new_n11586), .B(new_n11590), .Y(new_n11598));
  A2O1A1Ixp33_ASAP7_75t_L   g11342(.A1(new_n11293), .A2(new_n11592), .B(new_n11597), .C(new_n11598), .Y(new_n11599));
  AOI22xp33_ASAP7_75t_L     g11343(.A1(new_n6376), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n6648), .Y(new_n11600));
  OAI221xp5_ASAP7_75t_L     g11344(.A1(new_n6646), .A2(new_n1313), .B1(new_n6636), .B2(new_n1438), .C(new_n11600), .Y(new_n11601));
  XNOR2x2_ASAP7_75t_L       g11345(.A(\a[47] ), .B(new_n11601), .Y(new_n11602));
  INVx1_ASAP7_75t_L         g11346(.A(new_n11602), .Y(new_n11603));
  AOI21xp33_ASAP7_75t_L     g11347(.A1(new_n11596), .A2(new_n11599), .B(new_n11603), .Y(new_n11604));
  NOR2xp33_ASAP7_75t_L      g11348(.A(new_n11594), .B(new_n11598), .Y(new_n11605));
  NOR2xp33_ASAP7_75t_L      g11349(.A(new_n11591), .B(new_n11595), .Y(new_n11606));
  NOR3xp33_ASAP7_75t_L      g11350(.A(new_n11606), .B(new_n11605), .C(new_n11602), .Y(new_n11607));
  AND3x1_ASAP7_75t_L        g11351(.A(new_n11299), .B(new_n11302), .C(new_n11298), .Y(new_n11608));
  A2O1A1O1Ixp25_ASAP7_75t_L g11352(.A1(new_n11235), .A2(new_n10921), .B(new_n10991), .C(new_n11303), .D(new_n11608), .Y(new_n11609));
  NOR3xp33_ASAP7_75t_L      g11353(.A(new_n11607), .B(new_n11604), .C(new_n11609), .Y(new_n11610));
  OA21x2_ASAP7_75t_L        g11354(.A1(new_n11604), .A2(new_n11607), .B(new_n11609), .Y(new_n11611));
  AOI22xp33_ASAP7_75t_L     g11355(.A1(new_n5624), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n5901), .Y(new_n11612));
  OAI221xp5_ASAP7_75t_L     g11356(.A1(new_n5900), .A2(new_n1655), .B1(new_n5892), .B2(new_n1780), .C(new_n11612), .Y(new_n11613));
  XNOR2x2_ASAP7_75t_L       g11357(.A(new_n5619), .B(new_n11613), .Y(new_n11614));
  NOR3xp33_ASAP7_75t_L      g11358(.A(new_n11611), .B(new_n11614), .C(new_n11610), .Y(new_n11615));
  OA21x2_ASAP7_75t_L        g11359(.A1(new_n11610), .A2(new_n11611), .B(new_n11614), .Y(new_n11616));
  A2O1A1Ixp33_ASAP7_75t_L   g11360(.A1(new_n10990), .A2(new_n10996), .B(new_n11313), .C(new_n11309), .Y(new_n11617));
  OR3x1_ASAP7_75t_L         g11361(.A(new_n11617), .B(new_n11615), .C(new_n11616), .Y(new_n11618));
  OAI21xp33_ASAP7_75t_L     g11362(.A1(new_n11615), .A2(new_n11616), .B(new_n11617), .Y(new_n11619));
  AOI22xp33_ASAP7_75t_L     g11363(.A1(new_n4920), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n5167), .Y(new_n11620));
  OAI221xp5_ASAP7_75t_L     g11364(.A1(new_n5154), .A2(new_n1929), .B1(new_n5158), .B2(new_n2075), .C(new_n11620), .Y(new_n11621));
  XNOR2x2_ASAP7_75t_L       g11365(.A(\a[41] ), .B(new_n11621), .Y(new_n11622));
  NAND3xp33_ASAP7_75t_L     g11366(.A(new_n11618), .B(new_n11619), .C(new_n11622), .Y(new_n11623));
  NOR3xp33_ASAP7_75t_L      g11367(.A(new_n11617), .B(new_n11616), .C(new_n11615), .Y(new_n11624));
  OA21x2_ASAP7_75t_L        g11368(.A1(new_n11615), .A2(new_n11616), .B(new_n11617), .Y(new_n11625));
  INVx1_ASAP7_75t_L         g11369(.A(new_n11622), .Y(new_n11626));
  OAI21xp33_ASAP7_75t_L     g11370(.A1(new_n11624), .A2(new_n11625), .B(new_n11626), .Y(new_n11627));
  NAND2xp33_ASAP7_75t_L     g11371(.A(new_n11627), .B(new_n11623), .Y(new_n11628));
  NAND2xp33_ASAP7_75t_L     g11372(.A(new_n11311), .B(new_n11314), .Y(new_n11629));
  OR2x4_ASAP7_75t_L         g11373(.A(new_n11317), .B(new_n11629), .Y(new_n11630));
  A2O1A1Ixp33_ASAP7_75t_L   g11374(.A1(new_n11319), .A2(new_n11318), .B(new_n11320), .C(new_n11630), .Y(new_n11631));
  NOR2xp33_ASAP7_75t_L      g11375(.A(new_n11628), .B(new_n11631), .Y(new_n11632));
  AOI22xp33_ASAP7_75t_L     g11376(.A1(new_n11623), .A2(new_n11627), .B1(new_n11630), .B2(new_n11329), .Y(new_n11633));
  AOI22xp33_ASAP7_75t_L     g11377(.A1(new_n4283), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n4512), .Y(new_n11634));
  OAI221xp5_ASAP7_75t_L     g11378(.A1(new_n4277), .A2(new_n2497), .B1(new_n4499), .B2(new_n2672), .C(new_n11634), .Y(new_n11635));
  XNOR2x2_ASAP7_75t_L       g11379(.A(\a[38] ), .B(new_n11635), .Y(new_n11636));
  INVx1_ASAP7_75t_L         g11380(.A(new_n11636), .Y(new_n11637));
  NOR3xp33_ASAP7_75t_L      g11381(.A(new_n11632), .B(new_n11633), .C(new_n11637), .Y(new_n11638));
  NAND4xp25_ASAP7_75t_L     g11382(.A(new_n11329), .B(new_n11630), .C(new_n11627), .D(new_n11623), .Y(new_n11639));
  NAND2xp33_ASAP7_75t_L     g11383(.A(new_n11628), .B(new_n11631), .Y(new_n11640));
  AOI21xp33_ASAP7_75t_L     g11384(.A1(new_n11640), .A2(new_n11639), .B(new_n11636), .Y(new_n11641));
  NOR2xp33_ASAP7_75t_L      g11385(.A(new_n11641), .B(new_n11638), .Y(new_n11642));
  NOR3xp33_ASAP7_75t_L      g11386(.A(new_n11322), .B(new_n11323), .C(new_n11326), .Y(new_n11643));
  O2A1O1Ixp33_ASAP7_75t_L   g11387(.A1(new_n11328), .A2(new_n11330), .B(new_n11344), .C(new_n11643), .Y(new_n11644));
  NAND2xp33_ASAP7_75t_L     g11388(.A(new_n11644), .B(new_n11642), .Y(new_n11645));
  NAND3xp33_ASAP7_75t_L     g11389(.A(new_n11640), .B(new_n11639), .C(new_n11636), .Y(new_n11646));
  OAI21xp33_ASAP7_75t_L     g11390(.A1(new_n11633), .A2(new_n11632), .B(new_n11637), .Y(new_n11647));
  NAND2xp33_ASAP7_75t_L     g11391(.A(new_n11646), .B(new_n11647), .Y(new_n11648));
  A2O1A1Ixp33_ASAP7_75t_L   g11392(.A1(new_n11337), .A2(new_n11344), .B(new_n11643), .C(new_n11648), .Y(new_n11649));
  AOI22xp33_ASAP7_75t_L     g11393(.A1(new_n3633), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n3858), .Y(new_n11650));
  OAI221xp5_ASAP7_75t_L     g11394(.A1(new_n3853), .A2(new_n2982), .B1(new_n3856), .B2(new_n3187), .C(new_n11650), .Y(new_n11651));
  XNOR2x2_ASAP7_75t_L       g11395(.A(\a[35] ), .B(new_n11651), .Y(new_n11652));
  INVx1_ASAP7_75t_L         g11396(.A(new_n11652), .Y(new_n11653));
  AO21x2_ASAP7_75t_L        g11397(.A1(new_n11645), .A2(new_n11649), .B(new_n11653), .Y(new_n11654));
  NAND3xp33_ASAP7_75t_L     g11398(.A(new_n11649), .B(new_n11645), .C(new_n11653), .Y(new_n11655));
  A2O1A1O1Ixp25_ASAP7_75t_L g11399(.A1(new_n11035), .A2(new_n11231), .B(new_n11046), .C(new_n11350), .D(new_n11347), .Y(new_n11656));
  INVx1_ASAP7_75t_L         g11400(.A(new_n11656), .Y(new_n11657));
  NAND3xp33_ASAP7_75t_L     g11401(.A(new_n11657), .B(new_n11655), .C(new_n11654), .Y(new_n11658));
  NAND2xp33_ASAP7_75t_L     g11402(.A(new_n11655), .B(new_n11654), .Y(new_n11659));
  NAND2xp33_ASAP7_75t_L     g11403(.A(new_n11656), .B(new_n11659), .Y(new_n11660));
  AOI22xp33_ASAP7_75t_L     g11404(.A1(new_n3029), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n3258), .Y(new_n11661));
  OAI221xp5_ASAP7_75t_L     g11405(.A1(new_n3024), .A2(new_n3565), .B1(new_n3256), .B2(new_n3591), .C(new_n11661), .Y(new_n11662));
  XNOR2x2_ASAP7_75t_L       g11406(.A(\a[32] ), .B(new_n11662), .Y(new_n11663));
  NAND3xp33_ASAP7_75t_L     g11407(.A(new_n11658), .B(new_n11660), .C(new_n11663), .Y(new_n11664));
  INVx1_ASAP7_75t_L         g11408(.A(new_n11360), .Y(new_n11665));
  O2A1O1Ixp33_ASAP7_75t_L   g11409(.A1(new_n11343), .A2(new_n11665), .B(new_n11351), .C(new_n11659), .Y(new_n11666));
  AOI21xp33_ASAP7_75t_L     g11410(.A1(new_n11654), .A2(new_n11655), .B(new_n11657), .Y(new_n11667));
  INVx1_ASAP7_75t_L         g11411(.A(new_n11663), .Y(new_n11668));
  OAI21xp33_ASAP7_75t_L     g11412(.A1(new_n11667), .A2(new_n11666), .B(new_n11668), .Y(new_n11669));
  NOR2xp33_ASAP7_75t_L      g11413(.A(new_n11361), .B(new_n11359), .Y(new_n11670));
  AOI21xp33_ASAP7_75t_L     g11414(.A1(new_n11058), .A2(new_n11055), .B(new_n11059), .Y(new_n11671));
  MAJIxp5_ASAP7_75t_L       g11415(.A(new_n11670), .B(new_n11362), .C(new_n11671), .Y(new_n11672));
  NAND3xp33_ASAP7_75t_L     g11416(.A(new_n11669), .B(new_n11664), .C(new_n11672), .Y(new_n11673));
  AO21x2_ASAP7_75t_L        g11417(.A1(new_n11664), .A2(new_n11669), .B(new_n11672), .Y(new_n11674));
  AOI22xp33_ASAP7_75t_L     g11418(.A1(new_n2552), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n2736), .Y(new_n11675));
  OAI221xp5_ASAP7_75t_L     g11419(.A1(new_n2547), .A2(new_n4216), .B1(new_n2734), .B2(new_n4431), .C(new_n11675), .Y(new_n11676));
  XNOR2x2_ASAP7_75t_L       g11420(.A(\a[29] ), .B(new_n11676), .Y(new_n11677));
  NAND3xp33_ASAP7_75t_L     g11421(.A(new_n11674), .B(new_n11673), .C(new_n11677), .Y(new_n11678));
  AO21x2_ASAP7_75t_L        g11422(.A1(new_n11673), .A2(new_n11674), .B(new_n11677), .Y(new_n11679));
  A2O1A1O1Ixp25_ASAP7_75t_L g11423(.A1(new_n11068), .A2(new_n11070), .B(new_n11062), .C(new_n11370), .D(new_n11373), .Y(new_n11680));
  NAND3xp33_ASAP7_75t_L     g11424(.A(new_n11679), .B(new_n11678), .C(new_n11680), .Y(new_n11681));
  AND3x1_ASAP7_75t_L        g11425(.A(new_n11674), .B(new_n11673), .C(new_n11677), .Y(new_n11682));
  AOI21xp33_ASAP7_75t_L     g11426(.A1(new_n11674), .A2(new_n11673), .B(new_n11677), .Y(new_n11683));
  A2O1A1Ixp33_ASAP7_75t_L   g11427(.A1(new_n11071), .A2(new_n11069), .B(new_n11374), .C(new_n11367), .Y(new_n11684));
  OAI21xp33_ASAP7_75t_L     g11428(.A1(new_n11683), .A2(new_n11682), .B(new_n11684), .Y(new_n11685));
  INVx1_ASAP7_75t_L         g11429(.A(new_n4876), .Y(new_n11686));
  AOI22xp33_ASAP7_75t_L     g11430(.A1(new_n2114), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n2259), .Y(new_n11687));
  OAI221xp5_ASAP7_75t_L     g11431(.A1(new_n2109), .A2(new_n4848), .B1(new_n2257), .B2(new_n11686), .C(new_n11687), .Y(new_n11688));
  XNOR2x2_ASAP7_75t_L       g11432(.A(\a[26] ), .B(new_n11688), .Y(new_n11689));
  NAND3xp33_ASAP7_75t_L     g11433(.A(new_n11685), .B(new_n11681), .C(new_n11689), .Y(new_n11690));
  AO21x2_ASAP7_75t_L        g11434(.A1(new_n11681), .A2(new_n11685), .B(new_n11689), .Y(new_n11691));
  NAND2xp33_ASAP7_75t_L     g11435(.A(new_n11690), .B(new_n11691), .Y(new_n11692));
  INVx1_ASAP7_75t_L         g11436(.A(new_n11383), .Y(new_n11693));
  A2O1A1O1Ixp25_ASAP7_75t_L g11437(.A1(new_n11080), .A2(new_n11082), .B(new_n11224), .C(new_n11379), .D(new_n11693), .Y(new_n11694));
  NAND2xp33_ASAP7_75t_L     g11438(.A(new_n11694), .B(new_n11692), .Y(new_n11695));
  OAI211xp5_ASAP7_75t_L     g11439(.A1(new_n11693), .A2(new_n11385), .B(new_n11690), .C(new_n11691), .Y(new_n11696));
  AOI22xp33_ASAP7_75t_L     g11440(.A1(new_n1704), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n1837), .Y(new_n11697));
  OAI221xp5_ASAP7_75t_L     g11441(.A1(new_n1699), .A2(new_n5338), .B1(new_n1827), .B2(new_n6338), .C(new_n11697), .Y(new_n11698));
  XNOR2x2_ASAP7_75t_L       g11442(.A(\a[23] ), .B(new_n11698), .Y(new_n11699));
  AO21x2_ASAP7_75t_L        g11443(.A1(new_n11696), .A2(new_n11695), .B(new_n11699), .Y(new_n11700));
  NAND3xp33_ASAP7_75t_L     g11444(.A(new_n11695), .B(new_n11696), .C(new_n11699), .Y(new_n11701));
  OAI211xp5_ASAP7_75t_L     g11445(.A1(new_n11531), .A2(new_n11393), .B(new_n11700), .C(new_n11701), .Y(new_n11702));
  O2A1O1Ixp33_ASAP7_75t_L   g11446(.A1(new_n11400), .A2(new_n11401), .B(new_n11398), .C(new_n11531), .Y(new_n11703));
  NAND2xp33_ASAP7_75t_L     g11447(.A(new_n11701), .B(new_n11700), .Y(new_n11704));
  NAND2xp33_ASAP7_75t_L     g11448(.A(new_n11703), .B(new_n11704), .Y(new_n11705));
  AOI21xp33_ASAP7_75t_L     g11449(.A1(new_n11705), .A2(new_n11702), .B(new_n11530), .Y(new_n11706));
  INVx1_ASAP7_75t_L         g11450(.A(new_n11530), .Y(new_n11707));
  NOR2xp33_ASAP7_75t_L      g11451(.A(new_n11703), .B(new_n11704), .Y(new_n11708));
  AOI211xp5_ASAP7_75t_L     g11452(.A1(new_n11700), .A2(new_n11701), .B(new_n11531), .C(new_n11393), .Y(new_n11709));
  NOR3xp33_ASAP7_75t_L      g11453(.A(new_n11708), .B(new_n11709), .C(new_n11707), .Y(new_n11710));
  OAI21xp33_ASAP7_75t_L     g11454(.A1(new_n11706), .A2(new_n11710), .B(new_n11527), .Y(new_n11711));
  OAI21xp33_ASAP7_75t_L     g11455(.A1(new_n11709), .A2(new_n11708), .B(new_n11707), .Y(new_n11712));
  NAND3xp33_ASAP7_75t_L     g11456(.A(new_n11705), .B(new_n11702), .C(new_n11530), .Y(new_n11713));
  NAND4xp25_ASAP7_75t_L     g11457(.A(new_n11405), .B(new_n11712), .C(new_n11713), .D(new_n11526), .Y(new_n11714));
  AOI21xp33_ASAP7_75t_L     g11458(.A1(new_n11714), .A2(new_n11711), .B(new_n11525), .Y(new_n11715));
  INVx1_ASAP7_75t_L         g11459(.A(new_n11525), .Y(new_n11716));
  AOI22xp33_ASAP7_75t_L     g11460(.A1(new_n11712), .A2(new_n11713), .B1(new_n11526), .B2(new_n11405), .Y(new_n11717));
  NOR3xp33_ASAP7_75t_L      g11461(.A(new_n11710), .B(new_n11706), .C(new_n11527), .Y(new_n11718));
  NOR3xp33_ASAP7_75t_L      g11462(.A(new_n11717), .B(new_n11718), .C(new_n11716), .Y(new_n11719));
  OAI21xp33_ASAP7_75t_L     g11463(.A1(new_n11715), .A2(new_n11719), .B(new_n11522), .Y(new_n11720));
  OR2x4_ASAP7_75t_L         g11464(.A(new_n11214), .B(new_n11521), .Y(new_n11721));
  OAI21xp33_ASAP7_75t_L     g11465(.A1(new_n11718), .A2(new_n11717), .B(new_n11716), .Y(new_n11722));
  NAND3xp33_ASAP7_75t_L     g11466(.A(new_n11714), .B(new_n11711), .C(new_n11525), .Y(new_n11723));
  NAND4xp25_ASAP7_75t_L     g11467(.A(new_n11409), .B(new_n11721), .C(new_n11722), .D(new_n11723), .Y(new_n11724));
  NAND3xp33_ASAP7_75t_L     g11468(.A(new_n11724), .B(new_n11720), .C(new_n11520), .Y(new_n11725));
  INVx1_ASAP7_75t_L         g11469(.A(new_n11520), .Y(new_n11726));
  AOI22xp33_ASAP7_75t_L     g11470(.A1(new_n11722), .A2(new_n11723), .B1(new_n11721), .B2(new_n11409), .Y(new_n11727));
  NOR3xp33_ASAP7_75t_L      g11471(.A(new_n11522), .B(new_n11719), .C(new_n11715), .Y(new_n11728));
  OAI21xp33_ASAP7_75t_L     g11472(.A1(new_n11727), .A2(new_n11728), .B(new_n11726), .Y(new_n11729));
  NAND2xp33_ASAP7_75t_L     g11473(.A(new_n11725), .B(new_n11729), .Y(new_n11730));
  NOR2xp33_ASAP7_75t_L      g11474(.A(new_n11514), .B(new_n11730), .Y(new_n11731));
  AOI221xp5_ASAP7_75t_L     g11475(.A1(new_n11206), .A2(new_n11417), .B1(new_n11725), .B2(new_n11729), .C(new_n11513), .Y(new_n11732));
  NOR3xp33_ASAP7_75t_L      g11476(.A(new_n11731), .B(new_n11732), .C(new_n11511), .Y(new_n11733));
  INVx1_ASAP7_75t_L         g11477(.A(new_n11511), .Y(new_n11734));
  AO21x2_ASAP7_75t_L        g11478(.A1(new_n11417), .A2(new_n11206), .B(new_n11513), .Y(new_n11735));
  NOR3xp33_ASAP7_75t_L      g11479(.A(new_n11728), .B(new_n11727), .C(new_n11726), .Y(new_n11736));
  AOI21xp33_ASAP7_75t_L     g11480(.A1(new_n11724), .A2(new_n11720), .B(new_n11520), .Y(new_n11737));
  NOR2xp33_ASAP7_75t_L      g11481(.A(new_n11737), .B(new_n11736), .Y(new_n11738));
  NAND2xp33_ASAP7_75t_L     g11482(.A(new_n11738), .B(new_n11735), .Y(new_n11739));
  NAND2xp33_ASAP7_75t_L     g11483(.A(new_n11514), .B(new_n11730), .Y(new_n11740));
  AOI21xp33_ASAP7_75t_L     g11484(.A1(new_n11739), .A2(new_n11740), .B(new_n11734), .Y(new_n11741));
  NOR2xp33_ASAP7_75t_L      g11485(.A(new_n11733), .B(new_n11741), .Y(new_n11742));
  NAND2xp33_ASAP7_75t_L     g11486(.A(new_n11508), .B(new_n11742), .Y(new_n11743));
  MAJIxp5_ASAP7_75t_L       g11487(.A(new_n11432), .B(new_n11506), .C(new_n11428), .Y(new_n11744));
  OAI21xp33_ASAP7_75t_L     g11488(.A1(new_n11733), .A2(new_n11741), .B(new_n11744), .Y(new_n11745));
  AOI22xp33_ASAP7_75t_L     g11489(.A1(new_n444), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n471), .Y(new_n11746));
  OAI221xp5_ASAP7_75t_L     g11490(.A1(new_n468), .A2(new_n9620), .B1(new_n469), .B2(new_n9925), .C(new_n11746), .Y(new_n11747));
  XNOR2x2_ASAP7_75t_L       g11491(.A(\a[8] ), .B(new_n11747), .Y(new_n11748));
  NAND3xp33_ASAP7_75t_L     g11492(.A(new_n11743), .B(new_n11745), .C(new_n11748), .Y(new_n11749));
  NOR3xp33_ASAP7_75t_L      g11493(.A(new_n11744), .B(new_n11733), .C(new_n11741), .Y(new_n11750));
  INVx1_ASAP7_75t_L         g11494(.A(new_n11507), .Y(new_n11751));
  NAND3xp33_ASAP7_75t_L     g11495(.A(new_n11739), .B(new_n11734), .C(new_n11740), .Y(new_n11752));
  OAI21xp33_ASAP7_75t_L     g11496(.A1(new_n11732), .A2(new_n11731), .B(new_n11511), .Y(new_n11753));
  AOI221xp5_ASAP7_75t_L     g11497(.A1(new_n11752), .A2(new_n11753), .B1(new_n11432), .B2(new_n11430), .C(new_n11751), .Y(new_n11754));
  INVx1_ASAP7_75t_L         g11498(.A(new_n11748), .Y(new_n11755));
  OAI21xp33_ASAP7_75t_L     g11499(.A1(new_n11754), .A2(new_n11750), .B(new_n11755), .Y(new_n11756));
  NOR2xp33_ASAP7_75t_L      g11500(.A(new_n10250), .B(new_n429), .Y(new_n11757));
  INVx1_ASAP7_75t_L         g11501(.A(new_n11757), .Y(new_n11758));
  AND2x2_ASAP7_75t_L        g11502(.A(new_n10850), .B(new_n10854), .Y(new_n11759));
  NAND2xp33_ASAP7_75t_L     g11503(.A(new_n341), .B(new_n11759), .Y(new_n11760));
  AOI22xp33_ASAP7_75t_L     g11504(.A1(new_n344), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n370), .Y(new_n11761));
  AND4x1_ASAP7_75t_L        g11505(.A(new_n11761), .B(new_n11760), .C(new_n11758), .D(\a[5] ), .Y(new_n11762));
  AOI31xp33_ASAP7_75t_L     g11506(.A1(new_n11760), .A2(new_n11758), .A3(new_n11761), .B(\a[5] ), .Y(new_n11763));
  NOR2xp33_ASAP7_75t_L      g11507(.A(new_n11763), .B(new_n11762), .Y(new_n11764));
  AOI21xp33_ASAP7_75t_L     g11508(.A1(new_n11749), .A2(new_n11756), .B(new_n11764), .Y(new_n11765));
  NOR3xp33_ASAP7_75t_L      g11509(.A(new_n11750), .B(new_n11754), .C(new_n11755), .Y(new_n11766));
  AOI21xp33_ASAP7_75t_L     g11510(.A1(new_n11743), .A2(new_n11745), .B(new_n11748), .Y(new_n11767));
  OR2x4_ASAP7_75t_L         g11511(.A(new_n11763), .B(new_n11762), .Y(new_n11768));
  NOR3xp33_ASAP7_75t_L      g11512(.A(new_n11767), .B(new_n11766), .C(new_n11768), .Y(new_n11769));
  NOR3xp33_ASAP7_75t_L      g11513(.A(new_n11769), .B(new_n11765), .C(new_n11505), .Y(new_n11770));
  NOR2xp33_ASAP7_75t_L      g11514(.A(new_n11437), .B(new_n11433), .Y(new_n11771));
  NAND2xp33_ASAP7_75t_L     g11515(.A(new_n11441), .B(new_n11771), .Y(new_n11772));
  A2O1A1Ixp33_ASAP7_75t_L   g11516(.A1(new_n11455), .A2(new_n11454), .B(new_n11452), .C(new_n11772), .Y(new_n11773));
  OAI21xp33_ASAP7_75t_L     g11517(.A1(new_n11766), .A2(new_n11767), .B(new_n11768), .Y(new_n11774));
  NAND3xp33_ASAP7_75t_L     g11518(.A(new_n11749), .B(new_n11756), .C(new_n11764), .Y(new_n11775));
  AOI21xp33_ASAP7_75t_L     g11519(.A1(new_n11774), .A2(new_n11775), .B(new_n11773), .Y(new_n11776));
  NOR3xp33_ASAP7_75t_L      g11520(.A(new_n11770), .B(new_n11776), .C(new_n11503), .Y(new_n11777));
  INVx1_ASAP7_75t_L         g11521(.A(new_n11503), .Y(new_n11778));
  NAND3xp33_ASAP7_75t_L     g11522(.A(new_n11774), .B(new_n11773), .C(new_n11775), .Y(new_n11779));
  OAI21xp33_ASAP7_75t_L     g11523(.A1(new_n11765), .A2(new_n11769), .B(new_n11505), .Y(new_n11780));
  AOI21xp33_ASAP7_75t_L     g11524(.A1(new_n11780), .A2(new_n11779), .B(new_n11778), .Y(new_n11781));
  OAI21xp33_ASAP7_75t_L     g11525(.A1(new_n11483), .A2(new_n11482), .B(new_n11459), .Y(new_n11782));
  NOR3xp33_ASAP7_75t_L      g11526(.A(new_n11777), .B(new_n11781), .C(new_n11782), .Y(new_n11783));
  NAND3xp33_ASAP7_75t_L     g11527(.A(new_n11780), .B(new_n11779), .C(new_n11778), .Y(new_n11784));
  OAI21xp33_ASAP7_75t_L     g11528(.A1(new_n11776), .A2(new_n11770), .B(new_n11503), .Y(new_n11785));
  INVx1_ASAP7_75t_L         g11529(.A(new_n11782), .Y(new_n11786));
  AOI21xp33_ASAP7_75t_L     g11530(.A1(new_n11785), .A2(new_n11784), .B(new_n11786), .Y(new_n11787));
  NOR2xp33_ASAP7_75t_L      g11531(.A(new_n11787), .B(new_n11783), .Y(new_n11788));
  XOR2x2_ASAP7_75t_L        g11532(.A(new_n11788), .B(new_n11496), .Y(\f[64] ));
  NOR3xp33_ASAP7_75t_L      g11533(.A(new_n11717), .B(new_n11718), .C(new_n11525), .Y(new_n11790));
  O2A1O1Ixp33_ASAP7_75t_L   g11534(.A1(new_n11715), .A2(new_n11719), .B(new_n11522), .C(new_n11790), .Y(new_n11791));
  INVx1_ASAP7_75t_L         g11535(.A(new_n11791), .Y(new_n11792));
  AOI22xp33_ASAP7_75t_L     g11536(.A1(new_n1076), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1253), .Y(new_n11793));
  OAI221xp5_ASAP7_75t_L     g11537(.A1(new_n1154), .A2(new_n7317), .B1(new_n1156), .B2(new_n7602), .C(new_n11793), .Y(new_n11794));
  XNOR2x2_ASAP7_75t_L       g11538(.A(new_n1071), .B(new_n11794), .Y(new_n11795));
  INVx1_ASAP7_75t_L         g11539(.A(new_n11795), .Y(new_n11796));
  NAND3xp33_ASAP7_75t_L     g11540(.A(new_n11705), .B(new_n11702), .C(new_n11707), .Y(new_n11797));
  AOI22xp33_ASAP7_75t_L     g11541(.A1(new_n1360), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1581), .Y(new_n11798));
  OAI221xp5_ASAP7_75t_L     g11542(.A1(new_n1373), .A2(new_n6568), .B1(new_n1359), .B2(new_n6820), .C(new_n11798), .Y(new_n11799));
  XNOR2x2_ASAP7_75t_L       g11543(.A(\a[20] ), .B(new_n11799), .Y(new_n11800));
  INVx1_ASAP7_75t_L         g11544(.A(new_n11800), .Y(new_n11801));
  AOI22xp33_ASAP7_75t_L     g11545(.A1(new_n1704), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1837), .Y(new_n11802));
  OAI221xp5_ASAP7_75t_L     g11546(.A1(new_n1699), .A2(new_n5805), .B1(new_n1827), .B2(new_n5835), .C(new_n11802), .Y(new_n11803));
  XNOR2x2_ASAP7_75t_L       g11547(.A(\a[23] ), .B(new_n11803), .Y(new_n11804));
  INVx1_ASAP7_75t_L         g11548(.A(new_n11804), .Y(new_n11805));
  NAND2xp33_ASAP7_75t_L     g11549(.A(new_n11681), .B(new_n11685), .Y(new_n11806));
  MAJIxp5_ASAP7_75t_L       g11550(.A(new_n11694), .B(new_n11689), .C(new_n11806), .Y(new_n11807));
  NAND3xp33_ASAP7_75t_L     g11551(.A(new_n11660), .B(new_n11658), .C(new_n11668), .Y(new_n11808));
  A2O1A1Ixp33_ASAP7_75t_L   g11552(.A1(new_n11669), .A2(new_n11664), .B(new_n11672), .C(new_n11808), .Y(new_n11809));
  AOI22xp33_ASAP7_75t_L     g11553(.A1(new_n3029), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n3258), .Y(new_n11810));
  OAI221xp5_ASAP7_75t_L     g11554(.A1(new_n3024), .A2(new_n3584), .B1(new_n3256), .B2(new_n10137), .C(new_n11810), .Y(new_n11811));
  XNOR2x2_ASAP7_75t_L       g11555(.A(\a[32] ), .B(new_n11811), .Y(new_n11812));
  INVx1_ASAP7_75t_L         g11556(.A(new_n11812), .Y(new_n11813));
  INVx1_ASAP7_75t_L         g11557(.A(new_n11655), .Y(new_n11814));
  A2O1A1O1Ixp25_ASAP7_75t_L g11558(.A1(new_n11350), .A2(new_n11360), .B(new_n11347), .C(new_n11654), .D(new_n11814), .Y(new_n11815));
  OR2x4_ASAP7_75t_L         g11559(.A(new_n11610), .B(new_n11611), .Y(new_n11816));
  INVx1_ASAP7_75t_L         g11560(.A(new_n11614), .Y(new_n11817));
  NOR2xp33_ASAP7_75t_L      g11561(.A(new_n11817), .B(new_n11816), .Y(new_n11818));
  AOI22xp33_ASAP7_75t_L     g11562(.A1(new_n5624), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n5901), .Y(new_n11819));
  OAI221xp5_ASAP7_75t_L     g11563(.A1(new_n5900), .A2(new_n1774), .B1(new_n5892), .B2(new_n1915), .C(new_n11819), .Y(new_n11820));
  XNOR2x2_ASAP7_75t_L       g11564(.A(\a[44] ), .B(new_n11820), .Y(new_n11821));
  INVx1_ASAP7_75t_L         g11565(.A(new_n11821), .Y(new_n11822));
  NAND2xp33_ASAP7_75t_L     g11566(.A(new_n11599), .B(new_n11596), .Y(new_n11823));
  MAJIxp5_ASAP7_75t_L       g11567(.A(new_n11823), .B(new_n11602), .C(new_n11609), .Y(new_n11824));
  NOR3xp33_ASAP7_75t_L      g11568(.A(new_n11587), .B(new_n11588), .C(new_n11585), .Y(new_n11825));
  AOI22xp33_ASAP7_75t_L     g11569(.A1(new_n7111), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n7391), .Y(new_n11826));
  OAI221xp5_ASAP7_75t_L     g11570(.A1(new_n8558), .A2(new_n1030), .B1(new_n8237), .B2(new_n1209), .C(new_n11826), .Y(new_n11827));
  XNOR2x2_ASAP7_75t_L       g11571(.A(\a[50] ), .B(new_n11827), .Y(new_n11828));
  INVx1_ASAP7_75t_L         g11572(.A(new_n11828), .Y(new_n11829));
  A2O1A1Ixp33_ASAP7_75t_L   g11573(.A1(new_n11283), .A2(new_n11282), .B(new_n11579), .C(new_n11576), .Y(new_n11830));
  NOR2xp33_ASAP7_75t_L      g11574(.A(new_n11555), .B(new_n11562), .Y(new_n11831));
  NAND2xp33_ASAP7_75t_L     g11575(.A(new_n11563), .B(new_n11831), .Y(new_n11832));
  AOI22xp33_ASAP7_75t_L     g11576(.A1(new_n8831), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n9115), .Y(new_n11833));
  OAI221xp5_ASAP7_75t_L     g11577(.A1(new_n10343), .A2(new_n617), .B1(new_n10016), .B2(new_n685), .C(new_n11833), .Y(new_n11834));
  XNOR2x2_ASAP7_75t_L       g11578(.A(\a[56] ), .B(new_n11834), .Y(new_n11835));
  A2O1A1Ixp33_ASAP7_75t_L   g11579(.A1(new_n11269), .A2(new_n11266), .B(new_n11552), .C(new_n11553), .Y(new_n11836));
  NOR2xp33_ASAP7_75t_L      g11580(.A(new_n261), .B(new_n11535), .Y(new_n11837));
  O2A1O1Ixp33_ASAP7_75t_L   g11581(.A1(new_n11247), .A2(new_n11249), .B(\b[2] ), .C(new_n11837), .Y(new_n11838));
  NAND2xp33_ASAP7_75t_L     g11582(.A(new_n11256), .B(new_n359), .Y(new_n11839));
  AOI22xp33_ASAP7_75t_L     g11583(.A1(\b[3] ), .A2(new_n10939), .B1(\b[5] ), .B2(new_n10938), .Y(new_n11840));
  OAI211xp5_ASAP7_75t_L     g11584(.A1(new_n10937), .A2(new_n324), .B(new_n11839), .C(new_n11840), .Y(new_n11841));
  XNOR2x2_ASAP7_75t_L       g11585(.A(new_n10622), .B(new_n11841), .Y(new_n11842));
  XNOR2x2_ASAP7_75t_L       g11586(.A(new_n11838), .B(new_n11842), .Y(new_n11843));
  OAI21xp33_ASAP7_75t_L     g11587(.A1(new_n11543), .A2(new_n11541), .B(new_n11548), .Y(new_n11844));
  NOR2xp33_ASAP7_75t_L      g11588(.A(new_n11843), .B(new_n11844), .Y(new_n11845));
  AND2x2_ASAP7_75t_L        g11589(.A(new_n11843), .B(new_n11844), .Y(new_n11846));
  AOI22xp33_ASAP7_75t_L     g11590(.A1(new_n9700), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n10027), .Y(new_n11847));
  OAI221xp5_ASAP7_75t_L     g11591(.A1(new_n10024), .A2(new_n420), .B1(new_n9696), .B2(new_n494), .C(new_n11847), .Y(new_n11848));
  XNOR2x2_ASAP7_75t_L       g11592(.A(\a[59] ), .B(new_n11848), .Y(new_n11849));
  OAI21xp33_ASAP7_75t_L     g11593(.A1(new_n11845), .A2(new_n11846), .B(new_n11849), .Y(new_n11850));
  OR3x1_ASAP7_75t_L         g11594(.A(new_n11846), .B(new_n11845), .C(new_n11849), .Y(new_n11851));
  AOI21xp33_ASAP7_75t_L     g11595(.A1(new_n11851), .A2(new_n11850), .B(new_n11836), .Y(new_n11852));
  INVx1_ASAP7_75t_L         g11596(.A(new_n11836), .Y(new_n11853));
  OA21x2_ASAP7_75t_L        g11597(.A1(new_n11845), .A2(new_n11846), .B(new_n11849), .Y(new_n11854));
  NOR3xp33_ASAP7_75t_L      g11598(.A(new_n11846), .B(new_n11849), .C(new_n11845), .Y(new_n11855));
  NOR3xp33_ASAP7_75t_L      g11599(.A(new_n11853), .B(new_n11854), .C(new_n11855), .Y(new_n11856));
  OAI21xp33_ASAP7_75t_L     g11600(.A1(new_n11856), .A2(new_n11852), .B(new_n11835), .Y(new_n11857));
  INVx1_ASAP7_75t_L         g11601(.A(new_n11835), .Y(new_n11858));
  OAI21xp33_ASAP7_75t_L     g11602(.A1(new_n11855), .A2(new_n11854), .B(new_n11853), .Y(new_n11859));
  NAND3xp33_ASAP7_75t_L     g11603(.A(new_n11851), .B(new_n11850), .C(new_n11836), .Y(new_n11860));
  NAND3xp33_ASAP7_75t_L     g11604(.A(new_n11860), .B(new_n11859), .C(new_n11858), .Y(new_n11861));
  NAND2xp33_ASAP7_75t_L     g11605(.A(new_n11861), .B(new_n11857), .Y(new_n11862));
  A2O1A1O1Ixp25_ASAP7_75t_L g11606(.A1(new_n11564), .A2(new_n11561), .B(new_n11566), .C(new_n11832), .D(new_n11862), .Y(new_n11863));
  A2O1A1Ixp33_ASAP7_75t_L   g11607(.A1(new_n11564), .A2(new_n11561), .B(new_n11566), .C(new_n11832), .Y(new_n11864));
  AOI21xp33_ASAP7_75t_L     g11608(.A1(new_n11860), .A2(new_n11859), .B(new_n11858), .Y(new_n11865));
  NOR3xp33_ASAP7_75t_L      g11609(.A(new_n11852), .B(new_n11856), .C(new_n11835), .Y(new_n11866));
  NOR2xp33_ASAP7_75t_L      g11610(.A(new_n11865), .B(new_n11866), .Y(new_n11867));
  NOR2xp33_ASAP7_75t_L      g11611(.A(new_n11864), .B(new_n11867), .Y(new_n11868));
  AOI22xp33_ASAP7_75t_L     g11612(.A1(new_n7960), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n8537), .Y(new_n11869));
  OAI221xp5_ASAP7_75t_L     g11613(.A1(new_n8817), .A2(new_n784), .B1(new_n7957), .B2(new_n875), .C(new_n11869), .Y(new_n11870));
  XNOR2x2_ASAP7_75t_L       g11614(.A(\a[53] ), .B(new_n11870), .Y(new_n11871));
  INVx1_ASAP7_75t_L         g11615(.A(new_n11871), .Y(new_n11872));
  NOR3xp33_ASAP7_75t_L      g11616(.A(new_n11863), .B(new_n11868), .C(new_n11872), .Y(new_n11873));
  A2O1A1Ixp33_ASAP7_75t_L   g11617(.A1(new_n11563), .A2(new_n11831), .B(new_n11569), .C(new_n11867), .Y(new_n11874));
  NAND3xp33_ASAP7_75t_L     g11618(.A(new_n11862), .B(new_n11832), .C(new_n11575), .Y(new_n11875));
  AOI21xp33_ASAP7_75t_L     g11619(.A1(new_n11874), .A2(new_n11875), .B(new_n11871), .Y(new_n11876));
  OAI21xp33_ASAP7_75t_L     g11620(.A1(new_n11876), .A2(new_n11873), .B(new_n11830), .Y(new_n11877));
  O2A1O1Ixp33_ASAP7_75t_L   g11621(.A1(new_n11285), .A2(new_n11291), .B(new_n11574), .C(new_n11580), .Y(new_n11878));
  NAND3xp33_ASAP7_75t_L     g11622(.A(new_n11874), .B(new_n11875), .C(new_n11871), .Y(new_n11879));
  OAI21xp33_ASAP7_75t_L     g11623(.A1(new_n11868), .A2(new_n11863), .B(new_n11872), .Y(new_n11880));
  NAND3xp33_ASAP7_75t_L     g11624(.A(new_n11880), .B(new_n11879), .C(new_n11878), .Y(new_n11881));
  NAND3xp33_ASAP7_75t_L     g11625(.A(new_n11877), .B(new_n11881), .C(new_n11829), .Y(new_n11882));
  AOI21xp33_ASAP7_75t_L     g11626(.A1(new_n11880), .A2(new_n11879), .B(new_n11878), .Y(new_n11883));
  NOR3xp33_ASAP7_75t_L      g11627(.A(new_n11873), .B(new_n11876), .C(new_n11830), .Y(new_n11884));
  OAI21xp33_ASAP7_75t_L     g11628(.A1(new_n11883), .A2(new_n11884), .B(new_n11828), .Y(new_n11885));
  AOI221xp5_ASAP7_75t_L     g11629(.A1(new_n11598), .A2(new_n11594), .B1(new_n11882), .B2(new_n11885), .C(new_n11825), .Y(new_n11886));
  A2O1A1O1Ixp25_ASAP7_75t_L g11630(.A1(new_n11293), .A2(new_n11592), .B(new_n11597), .C(new_n11598), .D(new_n11825), .Y(new_n11887));
  NAND2xp33_ASAP7_75t_L     g11631(.A(new_n11882), .B(new_n11885), .Y(new_n11888));
  NOR2xp33_ASAP7_75t_L      g11632(.A(new_n11887), .B(new_n11888), .Y(new_n11889));
  AOI22xp33_ASAP7_75t_L     g11633(.A1(new_n6376), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n6648), .Y(new_n11890));
  OAI221xp5_ASAP7_75t_L     g11634(.A1(new_n6646), .A2(new_n1432), .B1(new_n6636), .B2(new_n1547), .C(new_n11890), .Y(new_n11891));
  XNOR2x2_ASAP7_75t_L       g11635(.A(\a[47] ), .B(new_n11891), .Y(new_n11892));
  INVx1_ASAP7_75t_L         g11636(.A(new_n11892), .Y(new_n11893));
  NOR3xp33_ASAP7_75t_L      g11637(.A(new_n11889), .B(new_n11893), .C(new_n11886), .Y(new_n11894));
  NAND2xp33_ASAP7_75t_L     g11638(.A(new_n11887), .B(new_n11888), .Y(new_n11895));
  OAI211xp5_ASAP7_75t_L     g11639(.A1(new_n11825), .A2(new_n11606), .B(new_n11882), .C(new_n11885), .Y(new_n11896));
  AOI21xp33_ASAP7_75t_L     g11640(.A1(new_n11896), .A2(new_n11895), .B(new_n11892), .Y(new_n11897));
  OAI21xp33_ASAP7_75t_L     g11641(.A1(new_n11894), .A2(new_n11897), .B(new_n11824), .Y(new_n11898));
  MAJx2_ASAP7_75t_L         g11642(.A(new_n11823), .B(new_n11602), .C(new_n11609), .Y(new_n11899));
  NAND3xp33_ASAP7_75t_L     g11643(.A(new_n11896), .B(new_n11895), .C(new_n11892), .Y(new_n11900));
  OAI21xp33_ASAP7_75t_L     g11644(.A1(new_n11886), .A2(new_n11889), .B(new_n11893), .Y(new_n11901));
  NAND3xp33_ASAP7_75t_L     g11645(.A(new_n11899), .B(new_n11900), .C(new_n11901), .Y(new_n11902));
  NAND3xp33_ASAP7_75t_L     g11646(.A(new_n11898), .B(new_n11902), .C(new_n11822), .Y(new_n11903));
  AOI21xp33_ASAP7_75t_L     g11647(.A1(new_n11900), .A2(new_n11901), .B(new_n11899), .Y(new_n11904));
  NOR3xp33_ASAP7_75t_L      g11648(.A(new_n11897), .B(new_n11894), .C(new_n11824), .Y(new_n11905));
  OAI21xp33_ASAP7_75t_L     g11649(.A1(new_n11904), .A2(new_n11905), .B(new_n11821), .Y(new_n11906));
  AOI211xp5_ASAP7_75t_L     g11650(.A1(new_n11903), .A2(new_n11906), .B(new_n11818), .C(new_n11625), .Y(new_n11907));
  NAND2xp33_ASAP7_75t_L     g11651(.A(new_n11903), .B(new_n11906), .Y(new_n11908));
  O2A1O1Ixp33_ASAP7_75t_L   g11652(.A1(new_n11816), .A2(new_n11817), .B(new_n11619), .C(new_n11908), .Y(new_n11909));
  AOI22xp33_ASAP7_75t_L     g11653(.A1(new_n4920), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n5167), .Y(new_n11910));
  OAI221xp5_ASAP7_75t_L     g11654(.A1(new_n5154), .A2(new_n2067), .B1(new_n5158), .B2(new_n2355), .C(new_n11910), .Y(new_n11911));
  XNOR2x2_ASAP7_75t_L       g11655(.A(\a[41] ), .B(new_n11911), .Y(new_n11912));
  INVx1_ASAP7_75t_L         g11656(.A(new_n11912), .Y(new_n11913));
  NOR3xp33_ASAP7_75t_L      g11657(.A(new_n11909), .B(new_n11907), .C(new_n11913), .Y(new_n11914));
  OAI211xp5_ASAP7_75t_L     g11658(.A1(new_n11816), .A2(new_n11817), .B(new_n11908), .C(new_n11619), .Y(new_n11915));
  OAI211xp5_ASAP7_75t_L     g11659(.A1(new_n11818), .A2(new_n11625), .B(new_n11903), .C(new_n11906), .Y(new_n11916));
  AOI21xp33_ASAP7_75t_L     g11660(.A1(new_n11915), .A2(new_n11916), .B(new_n11912), .Y(new_n11917));
  NOR2xp33_ASAP7_75t_L      g11661(.A(new_n11914), .B(new_n11917), .Y(new_n11918));
  NOR3xp33_ASAP7_75t_L      g11662(.A(new_n11625), .B(new_n11622), .C(new_n11624), .Y(new_n11919));
  INVx1_ASAP7_75t_L         g11663(.A(new_n11919), .Y(new_n11920));
  NAND3xp33_ASAP7_75t_L     g11664(.A(new_n11918), .B(new_n11640), .C(new_n11920), .Y(new_n11921));
  NAND3xp33_ASAP7_75t_L     g11665(.A(new_n11915), .B(new_n11916), .C(new_n11912), .Y(new_n11922));
  OAI21xp33_ASAP7_75t_L     g11666(.A1(new_n11907), .A2(new_n11909), .B(new_n11913), .Y(new_n11923));
  NAND2xp33_ASAP7_75t_L     g11667(.A(new_n11922), .B(new_n11923), .Y(new_n11924));
  A2O1A1Ixp33_ASAP7_75t_L   g11668(.A1(new_n11628), .A2(new_n11631), .B(new_n11919), .C(new_n11924), .Y(new_n11925));
  AOI22xp33_ASAP7_75t_L     g11669(.A1(new_n4283), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n4512), .Y(new_n11926));
  OAI221xp5_ASAP7_75t_L     g11670(.A1(new_n4277), .A2(new_n2666), .B1(new_n4499), .B2(new_n2695), .C(new_n11926), .Y(new_n11927));
  XNOR2x2_ASAP7_75t_L       g11671(.A(\a[38] ), .B(new_n11927), .Y(new_n11928));
  NAND3xp33_ASAP7_75t_L     g11672(.A(new_n11921), .B(new_n11925), .C(new_n11928), .Y(new_n11929));
  NOR3xp33_ASAP7_75t_L      g11673(.A(new_n11924), .B(new_n11919), .C(new_n11633), .Y(new_n11930));
  AOI21xp33_ASAP7_75t_L     g11674(.A1(new_n11640), .A2(new_n11920), .B(new_n11918), .Y(new_n11931));
  INVx1_ASAP7_75t_L         g11675(.A(new_n11928), .Y(new_n11932));
  OAI21xp33_ASAP7_75t_L     g11676(.A1(new_n11931), .A2(new_n11930), .B(new_n11932), .Y(new_n11933));
  NAND2xp33_ASAP7_75t_L     g11677(.A(new_n11929), .B(new_n11933), .Y(new_n11934));
  NAND3xp33_ASAP7_75t_L     g11678(.A(new_n11640), .B(new_n11639), .C(new_n11637), .Y(new_n11935));
  A2O1A1Ixp33_ASAP7_75t_L   g11679(.A1(new_n11647), .A2(new_n11646), .B(new_n11644), .C(new_n11935), .Y(new_n11936));
  NOR2xp33_ASAP7_75t_L      g11680(.A(new_n11936), .B(new_n11934), .Y(new_n11937));
  NOR3xp33_ASAP7_75t_L      g11681(.A(new_n11930), .B(new_n11931), .C(new_n11932), .Y(new_n11938));
  AOI21xp33_ASAP7_75t_L     g11682(.A1(new_n11921), .A2(new_n11925), .B(new_n11928), .Y(new_n11939));
  NOR2xp33_ASAP7_75t_L      g11683(.A(new_n11939), .B(new_n11938), .Y(new_n11940));
  O2A1O1Ixp33_ASAP7_75t_L   g11684(.A1(new_n11644), .A2(new_n11642), .B(new_n11935), .C(new_n11940), .Y(new_n11941));
  AOI22xp33_ASAP7_75t_L     g11685(.A1(new_n3633), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n3858), .Y(new_n11942));
  OAI221xp5_ASAP7_75t_L     g11686(.A1(new_n3853), .A2(new_n3180), .B1(new_n3856), .B2(new_n11047), .C(new_n11942), .Y(new_n11943));
  XNOR2x2_ASAP7_75t_L       g11687(.A(\a[35] ), .B(new_n11943), .Y(new_n11944));
  OAI21xp33_ASAP7_75t_L     g11688(.A1(new_n11937), .A2(new_n11941), .B(new_n11944), .Y(new_n11945));
  INVx1_ASAP7_75t_L         g11689(.A(new_n11936), .Y(new_n11946));
  NAND2xp33_ASAP7_75t_L     g11690(.A(new_n11946), .B(new_n11940), .Y(new_n11947));
  NAND2xp33_ASAP7_75t_L     g11691(.A(new_n11936), .B(new_n11934), .Y(new_n11948));
  INVx1_ASAP7_75t_L         g11692(.A(new_n11944), .Y(new_n11949));
  NAND3xp33_ASAP7_75t_L     g11693(.A(new_n11947), .B(new_n11948), .C(new_n11949), .Y(new_n11950));
  NAND2xp33_ASAP7_75t_L     g11694(.A(new_n11950), .B(new_n11945), .Y(new_n11951));
  NAND2xp33_ASAP7_75t_L     g11695(.A(new_n11815), .B(new_n11951), .Y(new_n11952));
  INVx1_ASAP7_75t_L         g11696(.A(new_n11654), .Y(new_n11953));
  A2O1A1Ixp33_ASAP7_75t_L   g11697(.A1(new_n11349), .A2(new_n11351), .B(new_n11953), .C(new_n11655), .Y(new_n11954));
  NAND3xp33_ASAP7_75t_L     g11698(.A(new_n11954), .B(new_n11945), .C(new_n11950), .Y(new_n11955));
  NAND3xp33_ASAP7_75t_L     g11699(.A(new_n11952), .B(new_n11955), .C(new_n11813), .Y(new_n11956));
  AOI21xp33_ASAP7_75t_L     g11700(.A1(new_n11945), .A2(new_n11950), .B(new_n11954), .Y(new_n11957));
  NOR2xp33_ASAP7_75t_L      g11701(.A(new_n11815), .B(new_n11951), .Y(new_n11958));
  OAI21xp33_ASAP7_75t_L     g11702(.A1(new_n11957), .A2(new_n11958), .B(new_n11812), .Y(new_n11959));
  AOI21xp33_ASAP7_75t_L     g11703(.A1(new_n11959), .A2(new_n11956), .B(new_n11809), .Y(new_n11960));
  INVx1_ASAP7_75t_L         g11704(.A(new_n11809), .Y(new_n11961));
  NAND2xp33_ASAP7_75t_L     g11705(.A(new_n11956), .B(new_n11959), .Y(new_n11962));
  NOR2xp33_ASAP7_75t_L      g11706(.A(new_n11961), .B(new_n11962), .Y(new_n11963));
  AOI22xp33_ASAP7_75t_L     g11707(.A1(new_n2552), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n2736), .Y(new_n11964));
  OAI221xp5_ASAP7_75t_L     g11708(.A1(new_n2547), .A2(new_n4424), .B1(new_n2734), .B2(new_n4641), .C(new_n11964), .Y(new_n11965));
  XNOR2x2_ASAP7_75t_L       g11709(.A(\a[29] ), .B(new_n11965), .Y(new_n11966));
  INVx1_ASAP7_75t_L         g11710(.A(new_n11966), .Y(new_n11967));
  NOR3xp33_ASAP7_75t_L      g11711(.A(new_n11963), .B(new_n11967), .C(new_n11960), .Y(new_n11968));
  NAND2xp33_ASAP7_75t_L     g11712(.A(new_n11961), .B(new_n11962), .Y(new_n11969));
  NAND3xp33_ASAP7_75t_L     g11713(.A(new_n11809), .B(new_n11956), .C(new_n11959), .Y(new_n11970));
  AOI21xp33_ASAP7_75t_L     g11714(.A1(new_n11969), .A2(new_n11970), .B(new_n11966), .Y(new_n11971));
  INVx1_ASAP7_75t_L         g11715(.A(new_n11677), .Y(new_n11972));
  NAND3xp33_ASAP7_75t_L     g11716(.A(new_n11674), .B(new_n11673), .C(new_n11972), .Y(new_n11973));
  A2O1A1Ixp33_ASAP7_75t_L   g11717(.A1(new_n11679), .A2(new_n11678), .B(new_n11680), .C(new_n11973), .Y(new_n11974));
  NOR3xp33_ASAP7_75t_L      g11718(.A(new_n11968), .B(new_n11971), .C(new_n11974), .Y(new_n11975));
  NAND3xp33_ASAP7_75t_L     g11719(.A(new_n11969), .B(new_n11970), .C(new_n11966), .Y(new_n11976));
  OAI21xp33_ASAP7_75t_L     g11720(.A1(new_n11960), .A2(new_n11963), .B(new_n11967), .Y(new_n11977));
  AOI22xp33_ASAP7_75t_L     g11721(.A1(new_n11685), .A2(new_n11973), .B1(new_n11976), .B2(new_n11977), .Y(new_n11978));
  AOI22xp33_ASAP7_75t_L     g11722(.A1(new_n2114), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n2259), .Y(new_n11979));
  OAI221xp5_ASAP7_75t_L     g11723(.A1(new_n2109), .A2(new_n4869), .B1(new_n2257), .B2(new_n5327), .C(new_n11979), .Y(new_n11980));
  XNOR2x2_ASAP7_75t_L       g11724(.A(\a[26] ), .B(new_n11980), .Y(new_n11981));
  OAI21xp33_ASAP7_75t_L     g11725(.A1(new_n11978), .A2(new_n11975), .B(new_n11981), .Y(new_n11982));
  NAND4xp25_ASAP7_75t_L     g11726(.A(new_n11977), .B(new_n11976), .C(new_n11685), .D(new_n11973), .Y(new_n11983));
  OAI21xp33_ASAP7_75t_L     g11727(.A1(new_n11971), .A2(new_n11968), .B(new_n11974), .Y(new_n11984));
  INVx1_ASAP7_75t_L         g11728(.A(new_n11981), .Y(new_n11985));
  NAND3xp33_ASAP7_75t_L     g11729(.A(new_n11984), .B(new_n11983), .C(new_n11985), .Y(new_n11986));
  AOI21xp33_ASAP7_75t_L     g11730(.A1(new_n11982), .A2(new_n11986), .B(new_n11807), .Y(new_n11987));
  INVx1_ASAP7_75t_L         g11731(.A(new_n11987), .Y(new_n11988));
  NAND3xp33_ASAP7_75t_L     g11732(.A(new_n11982), .B(new_n11986), .C(new_n11807), .Y(new_n11989));
  NAND3xp33_ASAP7_75t_L     g11733(.A(new_n11988), .B(new_n11805), .C(new_n11989), .Y(new_n11990));
  INVx1_ASAP7_75t_L         g11734(.A(new_n11989), .Y(new_n11991));
  OAI21xp33_ASAP7_75t_L     g11735(.A1(new_n11987), .A2(new_n11991), .B(new_n11804), .Y(new_n11992));
  NAND2xp33_ASAP7_75t_L     g11736(.A(new_n11990), .B(new_n11992), .Y(new_n11993));
  O2A1O1Ixp33_ASAP7_75t_L   g11737(.A1(new_n11703), .A2(new_n11704), .B(new_n11700), .C(new_n11993), .Y(new_n11994));
  A2O1A1Ixp33_ASAP7_75t_L   g11738(.A1(new_n11696), .A2(new_n11695), .B(new_n11699), .C(new_n11702), .Y(new_n11995));
  NOR3xp33_ASAP7_75t_L      g11739(.A(new_n11991), .B(new_n11987), .C(new_n11804), .Y(new_n11996));
  AOI21xp33_ASAP7_75t_L     g11740(.A1(new_n11988), .A2(new_n11989), .B(new_n11805), .Y(new_n11997));
  NOR2xp33_ASAP7_75t_L      g11741(.A(new_n11997), .B(new_n11996), .Y(new_n11998));
  NOR2xp33_ASAP7_75t_L      g11742(.A(new_n11998), .B(new_n11995), .Y(new_n11999));
  OAI21xp33_ASAP7_75t_L     g11743(.A1(new_n11994), .A2(new_n11999), .B(new_n11801), .Y(new_n12000));
  NAND2xp33_ASAP7_75t_L     g11744(.A(new_n11696), .B(new_n11695), .Y(new_n12001));
  INVx1_ASAP7_75t_L         g11745(.A(new_n11699), .Y(new_n12002));
  A2O1A1Ixp33_ASAP7_75t_L   g11746(.A1(new_n12002), .A2(new_n12001), .B(new_n11708), .C(new_n11998), .Y(new_n12003));
  NAND3xp33_ASAP7_75t_L     g11747(.A(new_n11993), .B(new_n11702), .C(new_n11700), .Y(new_n12004));
  NAND3xp33_ASAP7_75t_L     g11748(.A(new_n12003), .B(new_n11800), .C(new_n12004), .Y(new_n12005));
  AOI22xp33_ASAP7_75t_L     g11749(.A1(new_n11797), .A2(new_n11711), .B1(new_n12005), .B2(new_n12000), .Y(new_n12006));
  NAND4xp25_ASAP7_75t_L     g11750(.A(new_n12000), .B(new_n12005), .C(new_n11711), .D(new_n11797), .Y(new_n12007));
  INVx1_ASAP7_75t_L         g11751(.A(new_n12007), .Y(new_n12008));
  OAI21xp33_ASAP7_75t_L     g11752(.A1(new_n12006), .A2(new_n12008), .B(new_n11796), .Y(new_n12009));
  INVx1_ASAP7_75t_L         g11753(.A(new_n12006), .Y(new_n12010));
  NAND3xp33_ASAP7_75t_L     g11754(.A(new_n12010), .B(new_n11795), .C(new_n12007), .Y(new_n12011));
  NAND3xp33_ASAP7_75t_L     g11755(.A(new_n11792), .B(new_n12009), .C(new_n12011), .Y(new_n12012));
  AOI21xp33_ASAP7_75t_L     g11756(.A1(new_n12011), .A2(new_n12009), .B(new_n11792), .Y(new_n12013));
  INVx1_ASAP7_75t_L         g11757(.A(new_n12013), .Y(new_n12014));
  AOI22xp33_ASAP7_75t_L     g11758(.A1(new_n811), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n900), .Y(new_n12015));
  OAI221xp5_ASAP7_75t_L     g11759(.A1(new_n904), .A2(new_n7900), .B1(new_n898), .B2(new_n8174), .C(new_n12015), .Y(new_n12016));
  XNOR2x2_ASAP7_75t_L       g11760(.A(\a[14] ), .B(new_n12016), .Y(new_n12017));
  NAND3xp33_ASAP7_75t_L     g11761(.A(new_n12014), .B(new_n12012), .C(new_n12017), .Y(new_n12018));
  INVx1_ASAP7_75t_L         g11762(.A(new_n12012), .Y(new_n12019));
  INVx1_ASAP7_75t_L         g11763(.A(new_n12017), .Y(new_n12020));
  OAI21xp33_ASAP7_75t_L     g11764(.A1(new_n12013), .A2(new_n12019), .B(new_n12020), .Y(new_n12021));
  A2O1A1O1Ixp25_ASAP7_75t_L g11765(.A1(new_n11417), .A2(new_n11206), .B(new_n11513), .C(new_n11729), .D(new_n11736), .Y(new_n12022));
  AND3x1_ASAP7_75t_L        g11766(.A(new_n12021), .B(new_n12018), .C(new_n12022), .Y(new_n12023));
  AOI21xp33_ASAP7_75t_L     g11767(.A1(new_n12021), .A2(new_n12018), .B(new_n12022), .Y(new_n12024));
  AOI22xp33_ASAP7_75t_L     g11768(.A1(\b[54] ), .A2(new_n651), .B1(\b[56] ), .B2(new_n581), .Y(new_n12025));
  OAI221xp5_ASAP7_75t_L     g11769(.A1(new_n821), .A2(new_n8762), .B1(new_n577), .B2(new_n9331), .C(new_n12025), .Y(new_n12026));
  XNOR2x2_ASAP7_75t_L       g11770(.A(\a[11] ), .B(new_n12026), .Y(new_n12027));
  OAI21xp33_ASAP7_75t_L     g11771(.A1(new_n12024), .A2(new_n12023), .B(new_n12027), .Y(new_n12028));
  NAND3xp33_ASAP7_75t_L     g11772(.A(new_n12021), .B(new_n12018), .C(new_n12022), .Y(new_n12029));
  AO21x2_ASAP7_75t_L        g11773(.A1(new_n12018), .A2(new_n12021), .B(new_n12022), .Y(new_n12030));
  INVx1_ASAP7_75t_L         g11774(.A(new_n12027), .Y(new_n12031));
  NAND3xp33_ASAP7_75t_L     g11775(.A(new_n12030), .B(new_n12029), .C(new_n12031), .Y(new_n12032));
  AOI22xp33_ASAP7_75t_L     g11776(.A1(new_n444), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n471), .Y(new_n12033));
  OAI221xp5_ASAP7_75t_L     g11777(.A1(new_n468), .A2(new_n9920), .B1(new_n469), .B2(new_n11152), .C(new_n12033), .Y(new_n12034));
  XNOR2x2_ASAP7_75t_L       g11778(.A(\a[8] ), .B(new_n12034), .Y(new_n12035));
  NAND3xp33_ASAP7_75t_L     g11779(.A(new_n12028), .B(new_n12032), .C(new_n12035), .Y(new_n12036));
  AOI21xp33_ASAP7_75t_L     g11780(.A1(new_n12030), .A2(new_n12029), .B(new_n12031), .Y(new_n12037));
  NOR3xp33_ASAP7_75t_L      g11781(.A(new_n12023), .B(new_n12024), .C(new_n12027), .Y(new_n12038));
  INVx1_ASAP7_75t_L         g11782(.A(new_n12035), .Y(new_n12039));
  OAI21xp33_ASAP7_75t_L     g11783(.A1(new_n12037), .A2(new_n12038), .B(new_n12039), .Y(new_n12040));
  A2O1A1O1Ixp25_ASAP7_75t_L g11784(.A1(new_n11432), .A2(new_n11430), .B(new_n11751), .C(new_n11753), .D(new_n11733), .Y(new_n12041));
  NAND3xp33_ASAP7_75t_L     g11785(.A(new_n12040), .B(new_n12036), .C(new_n12041), .Y(new_n12042));
  NOR3xp33_ASAP7_75t_L      g11786(.A(new_n12038), .B(new_n12037), .C(new_n12039), .Y(new_n12043));
  AOI21xp33_ASAP7_75t_L     g11787(.A1(new_n12028), .A2(new_n12032), .B(new_n12035), .Y(new_n12044));
  INVx1_ASAP7_75t_L         g11788(.A(new_n12041), .Y(new_n12045));
  OAI21xp33_ASAP7_75t_L     g11789(.A1(new_n12044), .A2(new_n12043), .B(new_n12045), .Y(new_n12046));
  NAND2xp33_ASAP7_75t_L     g11790(.A(new_n11178), .B(new_n11498), .Y(new_n12047));
  AOI22xp33_ASAP7_75t_L     g11791(.A1(new_n344), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n370), .Y(new_n12048));
  OAI221xp5_ASAP7_75t_L     g11792(.A1(new_n429), .A2(new_n10847), .B1(new_n366), .B2(new_n12047), .C(new_n12048), .Y(new_n12049));
  XNOR2x2_ASAP7_75t_L       g11793(.A(\a[5] ), .B(new_n12049), .Y(new_n12050));
  NAND3xp33_ASAP7_75t_L     g11794(.A(new_n12046), .B(new_n12042), .C(new_n12050), .Y(new_n12051));
  NOR3xp33_ASAP7_75t_L      g11795(.A(new_n12043), .B(new_n12044), .C(new_n12045), .Y(new_n12052));
  AOI21xp33_ASAP7_75t_L     g11796(.A1(new_n12040), .A2(new_n12036), .B(new_n12041), .Y(new_n12053));
  INVx1_ASAP7_75t_L         g11797(.A(new_n12050), .Y(new_n12054));
  OAI21xp33_ASAP7_75t_L     g11798(.A1(new_n12053), .A2(new_n12052), .B(new_n12054), .Y(new_n12055));
  NAND3xp33_ASAP7_75t_L     g11799(.A(new_n11743), .B(new_n11745), .C(new_n11755), .Y(new_n12056));
  A2O1A1Ixp33_ASAP7_75t_L   g11800(.A1(new_n11749), .A2(new_n11756), .B(new_n11764), .C(new_n12056), .Y(new_n12057));
  NAND2xp33_ASAP7_75t_L     g11801(.A(\b[63] ), .B(new_n267), .Y(new_n12058));
  A2O1A1O1Ixp25_ASAP7_75t_L g11802(.A1(new_n10250), .A2(new_n10852), .B(new_n10847), .C(new_n11172), .D(new_n12058), .Y(new_n12059));
  A2O1A1O1Ixp25_ASAP7_75t_L g11803(.A1(\b[59] ), .A2(new_n10256), .B(\b[60] ), .C(\b[61] ), .D(\b[62] ), .Y(new_n12060));
  INVx1_ASAP7_75t_L         g11804(.A(new_n12060), .Y(new_n12061));
  A2O1A1O1Ixp25_ASAP7_75t_L g11805(.A1(new_n267), .A2(new_n12061), .B(new_n282), .C(\b[63] ), .D(new_n262), .Y(new_n12062));
  A2O1A1Ixp33_ASAP7_75t_L   g11806(.A1(new_n262), .A2(new_n12059), .B(new_n12062), .C(new_n12057), .Y(new_n12063));
  AOI21xp33_ASAP7_75t_L     g11807(.A1(new_n12059), .A2(new_n262), .B(new_n12062), .Y(new_n12064));
  NAND3xp33_ASAP7_75t_L     g11808(.A(new_n11774), .B(new_n12056), .C(new_n12064), .Y(new_n12065));
  AOI22xp33_ASAP7_75t_L     g11809(.A1(new_n12063), .A2(new_n12065), .B1(new_n12051), .B2(new_n12055), .Y(new_n12066));
  NAND4xp25_ASAP7_75t_L     g11810(.A(new_n12055), .B(new_n12063), .C(new_n12051), .D(new_n12065), .Y(new_n12067));
  INVx1_ASAP7_75t_L         g11811(.A(new_n12067), .Y(new_n12068));
  NAND2xp33_ASAP7_75t_L     g11812(.A(new_n11779), .B(new_n11784), .Y(new_n12069));
  NOR3xp33_ASAP7_75t_L      g11813(.A(new_n12068), .B(new_n12069), .C(new_n12066), .Y(new_n12070));
  INVx1_ASAP7_75t_L         g11814(.A(new_n12066), .Y(new_n12071));
  NOR2xp33_ASAP7_75t_L      g11815(.A(new_n11770), .B(new_n11777), .Y(new_n12072));
  AOI21xp33_ASAP7_75t_L     g11816(.A1(new_n12071), .A2(new_n12067), .B(new_n12072), .Y(new_n12073));
  NOR2xp33_ASAP7_75t_L      g11817(.A(new_n12073), .B(new_n12070), .Y(new_n12074));
  A2O1A1Ixp33_ASAP7_75t_L   g11818(.A1(new_n11496), .A2(new_n11788), .B(new_n11783), .C(new_n12074), .Y(new_n12075));
  NAND3xp33_ASAP7_75t_L     g11819(.A(new_n12072), .B(new_n12071), .C(new_n12067), .Y(new_n12076));
  OAI21xp33_ASAP7_75t_L     g11820(.A1(new_n12066), .A2(new_n12068), .B(new_n12069), .Y(new_n12077));
  NAND2xp33_ASAP7_75t_L     g11821(.A(new_n12077), .B(new_n12076), .Y(new_n12078));
  A2O1A1O1Ixp25_ASAP7_75t_L g11822(.A1(new_n11493), .A2(new_n11490), .B(new_n11491), .C(new_n11788), .D(new_n11783), .Y(new_n12079));
  NAND2xp33_ASAP7_75t_L     g11823(.A(new_n12078), .B(new_n12079), .Y(new_n12080));
  AND2x2_ASAP7_75t_L        g11824(.A(new_n12075), .B(new_n12080), .Y(\f[65] ));
  NAND2xp33_ASAP7_75t_L     g11825(.A(new_n12065), .B(new_n12067), .Y(new_n12082));
  AOI22xp33_ASAP7_75t_L     g11826(.A1(\b[55] ), .A2(new_n651), .B1(\b[57] ), .B2(new_n581), .Y(new_n12083));
  OAI221xp5_ASAP7_75t_L     g11827(.A1(new_n821), .A2(new_n9323), .B1(new_n577), .B2(new_n9627), .C(new_n12083), .Y(new_n12084));
  XNOR2x2_ASAP7_75t_L       g11828(.A(new_n574), .B(new_n12084), .Y(new_n12085));
  NAND3xp33_ASAP7_75t_L     g11829(.A(new_n12014), .B(new_n12012), .C(new_n12020), .Y(new_n12086));
  A2O1A1Ixp33_ASAP7_75t_L   g11830(.A1(new_n12021), .A2(new_n12018), .B(new_n12022), .C(new_n12086), .Y(new_n12087));
  NOR2xp33_ASAP7_75t_L      g11831(.A(new_n12085), .B(new_n12087), .Y(new_n12088));
  INVx1_ASAP7_75t_L         g11832(.A(new_n12088), .Y(new_n12089));
  NAND2xp33_ASAP7_75t_L     g11833(.A(new_n12085), .B(new_n12087), .Y(new_n12090));
  INVx1_ASAP7_75t_L         g11834(.A(new_n12011), .Y(new_n12091));
  NAND2xp33_ASAP7_75t_L     g11835(.A(\b[53] ), .B(new_n815), .Y(new_n12092));
  OAI221xp5_ASAP7_75t_L     g11836(.A1(new_n977), .A2(new_n8458), .B1(new_n7900), .B2(new_n978), .C(new_n12092), .Y(new_n12093));
  AOI21xp33_ASAP7_75t_L     g11837(.A1(new_n8464), .A2(new_n808), .B(new_n12093), .Y(new_n12094));
  NAND2xp33_ASAP7_75t_L     g11838(.A(\a[14] ), .B(new_n12094), .Y(new_n12095));
  A2O1A1Ixp33_ASAP7_75t_L   g11839(.A1(new_n8464), .A2(new_n808), .B(new_n12093), .C(new_n806), .Y(new_n12096));
  AND2x2_ASAP7_75t_L        g11840(.A(new_n12096), .B(new_n12095), .Y(new_n12097));
  A2O1A1Ixp33_ASAP7_75t_L   g11841(.A1(new_n11792), .A2(new_n12009), .B(new_n12091), .C(new_n12097), .Y(new_n12098));
  O2A1O1Ixp33_ASAP7_75t_L   g11842(.A1(new_n11727), .A2(new_n11790), .B(new_n12009), .C(new_n12091), .Y(new_n12099));
  INVx1_ASAP7_75t_L         g11843(.A(new_n12097), .Y(new_n12100));
  NAND2xp33_ASAP7_75t_L     g11844(.A(new_n12100), .B(new_n12099), .Y(new_n12101));
  NAND2xp33_ASAP7_75t_L     g11845(.A(new_n12098), .B(new_n12101), .Y(new_n12102));
  NOR2xp33_ASAP7_75t_L      g11846(.A(new_n11994), .B(new_n11999), .Y(new_n12103));
  AOI22xp33_ASAP7_75t_L     g11847(.A1(new_n1076), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1253), .Y(new_n12104));
  OAI221xp5_ASAP7_75t_L     g11848(.A1(new_n1154), .A2(new_n7593), .B1(new_n1156), .B2(new_n7623), .C(new_n12104), .Y(new_n12105));
  XNOR2x2_ASAP7_75t_L       g11849(.A(\a[17] ), .B(new_n12105), .Y(new_n12106));
  INVx1_ASAP7_75t_L         g11850(.A(new_n12106), .Y(new_n12107));
  AOI211xp5_ASAP7_75t_L     g11851(.A1(new_n12103), .A2(new_n11801), .B(new_n12107), .C(new_n12006), .Y(new_n12108));
  A2O1A1Ixp33_ASAP7_75t_L   g11852(.A1(new_n12103), .A2(new_n11801), .B(new_n12006), .C(new_n12107), .Y(new_n12109));
  INVx1_ASAP7_75t_L         g11853(.A(new_n12109), .Y(new_n12110));
  NOR2xp33_ASAP7_75t_L      g11854(.A(new_n12108), .B(new_n12110), .Y(new_n12111));
  AOI22xp33_ASAP7_75t_L     g11855(.A1(new_n1360), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1581), .Y(new_n12112));
  OAI221xp5_ASAP7_75t_L     g11856(.A1(new_n1373), .A2(new_n6812), .B1(new_n1359), .B2(new_n6837), .C(new_n12112), .Y(new_n12113));
  XNOR2x2_ASAP7_75t_L       g11857(.A(\a[20] ), .B(new_n12113), .Y(new_n12114));
  A2O1A1O1Ixp25_ASAP7_75t_L g11858(.A1(new_n12002), .A2(new_n12001), .B(new_n11708), .C(new_n11992), .D(new_n11996), .Y(new_n12115));
  NAND2xp33_ASAP7_75t_L     g11859(.A(new_n12114), .B(new_n12115), .Y(new_n12116));
  A2O1A1O1Ixp25_ASAP7_75t_L g11860(.A1(new_n11700), .A2(new_n11702), .B(new_n11997), .C(new_n11990), .D(new_n12114), .Y(new_n12117));
  INVx1_ASAP7_75t_L         g11861(.A(new_n12117), .Y(new_n12118));
  NAND2xp33_ASAP7_75t_L     g11862(.A(new_n12118), .B(new_n12116), .Y(new_n12119));
  AOI22xp33_ASAP7_75t_L     g11863(.A1(new_n1704), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n1837), .Y(new_n12120));
  OAI221xp5_ASAP7_75t_L     g11864(.A1(new_n1699), .A2(new_n5829), .B1(new_n1827), .B2(new_n6329), .C(new_n12120), .Y(new_n12121));
  XNOR2x2_ASAP7_75t_L       g11865(.A(\a[23] ), .B(new_n12121), .Y(new_n12122));
  INVx1_ASAP7_75t_L         g11866(.A(new_n12122), .Y(new_n12123));
  NOR3xp33_ASAP7_75t_L      g11867(.A(new_n11975), .B(new_n11978), .C(new_n11981), .Y(new_n12124));
  NOR2xp33_ASAP7_75t_L      g11868(.A(new_n11807), .B(new_n12124), .Y(new_n12125));
  O2A1O1Ixp33_ASAP7_75t_L   g11869(.A1(new_n11975), .A2(new_n11978), .B(new_n11981), .C(new_n12125), .Y(new_n12126));
  INVx1_ASAP7_75t_L         g11870(.A(new_n12126), .Y(new_n12127));
  NOR2xp33_ASAP7_75t_L      g11871(.A(new_n12123), .B(new_n12127), .Y(new_n12128));
  O2A1O1Ixp33_ASAP7_75t_L   g11872(.A1(new_n11807), .A2(new_n12124), .B(new_n11982), .C(new_n12122), .Y(new_n12129));
  NOR2xp33_ASAP7_75t_L      g11873(.A(new_n12129), .B(new_n12128), .Y(new_n12130));
  NAND2xp33_ASAP7_75t_L     g11874(.A(new_n11970), .B(new_n11969), .Y(new_n12131));
  AOI22xp33_ASAP7_75t_L     g11875(.A1(new_n2114), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n2259), .Y(new_n12132));
  OAI221xp5_ASAP7_75t_L     g11876(.A1(new_n2109), .A2(new_n5321), .B1(new_n2257), .B2(new_n5346), .C(new_n12132), .Y(new_n12133));
  XNOR2x2_ASAP7_75t_L       g11877(.A(\a[26] ), .B(new_n12133), .Y(new_n12134));
  OAI211xp5_ASAP7_75t_L     g11878(.A1(new_n11966), .A2(new_n12131), .B(new_n11984), .C(new_n12134), .Y(new_n12135));
  O2A1O1Ixp33_ASAP7_75t_L   g11879(.A1(new_n12131), .A2(new_n11966), .B(new_n11984), .C(new_n12134), .Y(new_n12136));
  INVx1_ASAP7_75t_L         g11880(.A(new_n12136), .Y(new_n12137));
  AOI21xp33_ASAP7_75t_L     g11881(.A1(new_n11952), .A2(new_n11955), .B(new_n11813), .Y(new_n12138));
  NAND2xp33_ASAP7_75t_L     g11882(.A(\b[38] ), .B(new_n2553), .Y(new_n12139));
  OAI221xp5_ASAP7_75t_L     g11883(.A1(new_n2545), .A2(new_n4848), .B1(new_n4424), .B2(new_n2747), .C(new_n12139), .Y(new_n12140));
  AOI21xp33_ASAP7_75t_L     g11884(.A1(new_n5352), .A2(new_n2544), .B(new_n12140), .Y(new_n12141));
  NAND2xp33_ASAP7_75t_L     g11885(.A(\a[29] ), .B(new_n12141), .Y(new_n12142));
  A2O1A1Ixp33_ASAP7_75t_L   g11886(.A1(new_n5352), .A2(new_n2544), .B(new_n12140), .C(new_n2538), .Y(new_n12143));
  AND2x2_ASAP7_75t_L        g11887(.A(new_n12143), .B(new_n12142), .Y(new_n12144));
  A2O1A1O1Ixp25_ASAP7_75t_L g11888(.A1(new_n11808), .A2(new_n11674), .B(new_n12138), .C(new_n11956), .D(new_n12144), .Y(new_n12145));
  A2O1A1Ixp33_ASAP7_75t_L   g11889(.A1(new_n11674), .A2(new_n11808), .B(new_n12138), .C(new_n11956), .Y(new_n12146));
  INVx1_ASAP7_75t_L         g11890(.A(new_n12144), .Y(new_n12147));
  NOR2xp33_ASAP7_75t_L      g11891(.A(new_n12147), .B(new_n12146), .Y(new_n12148));
  NOR2xp33_ASAP7_75t_L      g11892(.A(new_n12145), .B(new_n12148), .Y(new_n12149));
  INVx1_ASAP7_75t_L         g11893(.A(new_n12149), .Y(new_n12150));
  A2O1A1Ixp33_ASAP7_75t_L   g11894(.A1(new_n11575), .A2(new_n11832), .B(new_n11865), .C(new_n11861), .Y(new_n12151));
  AOI22xp33_ASAP7_75t_L     g11895(.A1(new_n8831), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n9115), .Y(new_n12152));
  OAI221xp5_ASAP7_75t_L     g11896(.A1(new_n10343), .A2(new_n679), .B1(new_n10016), .B2(new_n768), .C(new_n12152), .Y(new_n12153));
  XNOR2x2_ASAP7_75t_L       g11897(.A(\a[56] ), .B(new_n12153), .Y(new_n12154));
  NAND2xp33_ASAP7_75t_L     g11898(.A(new_n11843), .B(new_n11844), .Y(new_n12155));
  A2O1A1Ixp33_ASAP7_75t_L   g11899(.A1(new_n11533), .A2(\b[2] ), .B(new_n11837), .C(new_n11842), .Y(new_n12156));
  NOR2xp33_ASAP7_75t_L      g11900(.A(new_n276), .B(new_n11535), .Y(new_n12157));
  A2O1A1Ixp33_ASAP7_75t_L   g11901(.A1(new_n11533), .A2(\b[3] ), .B(new_n12157), .C(\a[2] ), .Y(new_n12158));
  O2A1O1Ixp33_ASAP7_75t_L   g11902(.A1(new_n11247), .A2(new_n11249), .B(\b[3] ), .C(new_n12157), .Y(new_n12159));
  NAND2xp33_ASAP7_75t_L     g11903(.A(new_n262), .B(new_n12159), .Y(new_n12160));
  NAND2xp33_ASAP7_75t_L     g11904(.A(new_n12158), .B(new_n12160), .Y(new_n12161));
  NOR2xp33_ASAP7_75t_L      g11905(.A(new_n418), .B(new_n10630), .Y(new_n12162));
  AOI221xp5_ASAP7_75t_L     g11906(.A1(\b[4] ), .A2(new_n10939), .B1(\b[5] ), .B2(new_n10632), .C(new_n12162), .Y(new_n12163));
  OAI211xp5_ASAP7_75t_L     g11907(.A1(new_n10629), .A2(new_n390), .B(\a[62] ), .C(new_n12163), .Y(new_n12164));
  INVx1_ASAP7_75t_L         g11908(.A(new_n12164), .Y(new_n12165));
  O2A1O1Ixp33_ASAP7_75t_L   g11909(.A1(new_n10629), .A2(new_n390), .B(new_n12163), .C(\a[62] ), .Y(new_n12166));
  NOR2xp33_ASAP7_75t_L      g11910(.A(new_n12166), .B(new_n12165), .Y(new_n12167));
  NOR2xp33_ASAP7_75t_L      g11911(.A(new_n12161), .B(new_n12167), .Y(new_n12168));
  AOI211xp5_ASAP7_75t_L     g11912(.A1(new_n12160), .A2(new_n12158), .B(new_n12166), .C(new_n12165), .Y(new_n12169));
  AOI211xp5_ASAP7_75t_L     g11913(.A1(new_n12155), .A2(new_n12156), .B(new_n12168), .C(new_n12169), .Y(new_n12170));
  NAND2xp33_ASAP7_75t_L     g11914(.A(new_n12156), .B(new_n12155), .Y(new_n12171));
  NOR2xp33_ASAP7_75t_L      g11915(.A(new_n12169), .B(new_n12168), .Y(new_n12172));
  NOR2xp33_ASAP7_75t_L      g11916(.A(new_n12172), .B(new_n12171), .Y(new_n12173));
  NOR2xp33_ASAP7_75t_L      g11917(.A(new_n12170), .B(new_n12173), .Y(new_n12174));
  AOI22xp33_ASAP7_75t_L     g11918(.A1(new_n9700), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n10027), .Y(new_n12175));
  OAI221xp5_ASAP7_75t_L     g11919(.A1(new_n10024), .A2(new_n488), .B1(new_n9696), .B2(new_n548), .C(new_n12175), .Y(new_n12176));
  XNOR2x2_ASAP7_75t_L       g11920(.A(\a[59] ), .B(new_n12176), .Y(new_n12177));
  XOR2x2_ASAP7_75t_L        g11921(.A(new_n12177), .B(new_n12174), .Y(new_n12178));
  NOR2xp33_ASAP7_75t_L      g11922(.A(new_n11836), .B(new_n11855), .Y(new_n12179));
  O2A1O1Ixp33_ASAP7_75t_L   g11923(.A1(new_n11845), .A2(new_n11846), .B(new_n11849), .C(new_n12179), .Y(new_n12180));
  XNOR2x2_ASAP7_75t_L       g11924(.A(new_n12180), .B(new_n12178), .Y(new_n12181));
  XNOR2x2_ASAP7_75t_L       g11925(.A(new_n12154), .B(new_n12181), .Y(new_n12182));
  XNOR2x2_ASAP7_75t_L       g11926(.A(new_n12151), .B(new_n12182), .Y(new_n12183));
  AOI22xp33_ASAP7_75t_L     g11927(.A1(new_n7960), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n8537), .Y(new_n12184));
  OAI221xp5_ASAP7_75t_L     g11928(.A1(new_n8817), .A2(new_n869), .B1(new_n7957), .B2(new_n950), .C(new_n12184), .Y(new_n12185));
  XNOR2x2_ASAP7_75t_L       g11929(.A(\a[53] ), .B(new_n12185), .Y(new_n12186));
  INVx1_ASAP7_75t_L         g11930(.A(new_n12186), .Y(new_n12187));
  XNOR2x2_ASAP7_75t_L       g11931(.A(new_n12187), .B(new_n12183), .Y(new_n12188));
  NAND3xp33_ASAP7_75t_L     g11932(.A(new_n11874), .B(new_n11875), .C(new_n11872), .Y(new_n12189));
  A2O1A1Ixp33_ASAP7_75t_L   g11933(.A1(new_n11880), .A2(new_n11879), .B(new_n11878), .C(new_n12189), .Y(new_n12190));
  OR2x4_ASAP7_75t_L         g11934(.A(new_n12190), .B(new_n12188), .Y(new_n12191));
  NAND2xp33_ASAP7_75t_L     g11935(.A(new_n12190), .B(new_n12188), .Y(new_n12192));
  AOI22xp33_ASAP7_75t_L     g11936(.A1(new_n7111), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n7391), .Y(new_n12193));
  OAI221xp5_ASAP7_75t_L     g11937(.A1(new_n8558), .A2(new_n1201), .B1(new_n8237), .B2(new_n1320), .C(new_n12193), .Y(new_n12194));
  XNOR2x2_ASAP7_75t_L       g11938(.A(\a[50] ), .B(new_n12194), .Y(new_n12195));
  NAND3xp33_ASAP7_75t_L     g11939(.A(new_n12191), .B(new_n12192), .C(new_n12195), .Y(new_n12196));
  AO21x2_ASAP7_75t_L        g11940(.A1(new_n12192), .A2(new_n12191), .B(new_n12195), .Y(new_n12197));
  AND2x2_ASAP7_75t_L        g11941(.A(new_n12196), .B(new_n12197), .Y(new_n12198));
  NAND2xp33_ASAP7_75t_L     g11942(.A(new_n11882), .B(new_n11896), .Y(new_n12199));
  XOR2x2_ASAP7_75t_L        g11943(.A(new_n12199), .B(new_n12198), .Y(new_n12200));
  AOI22xp33_ASAP7_75t_L     g11944(.A1(new_n6376), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n6648), .Y(new_n12201));
  OAI221xp5_ASAP7_75t_L     g11945(.A1(new_n6646), .A2(new_n1539), .B1(new_n6636), .B2(new_n1662), .C(new_n12201), .Y(new_n12202));
  XNOR2x2_ASAP7_75t_L       g11946(.A(\a[47] ), .B(new_n12202), .Y(new_n12203));
  AND2x2_ASAP7_75t_L        g11947(.A(new_n12203), .B(new_n12200), .Y(new_n12204));
  NOR2xp33_ASAP7_75t_L      g11948(.A(new_n12203), .B(new_n12200), .Y(new_n12205));
  NAND3xp33_ASAP7_75t_L     g11949(.A(new_n11896), .B(new_n11895), .C(new_n11893), .Y(new_n12206));
  A2O1A1Ixp33_ASAP7_75t_L   g11950(.A1(new_n11900), .A2(new_n11901), .B(new_n11899), .C(new_n12206), .Y(new_n12207));
  INVx1_ASAP7_75t_L         g11951(.A(new_n12207), .Y(new_n12208));
  OR3x1_ASAP7_75t_L         g11952(.A(new_n12204), .B(new_n12205), .C(new_n12208), .Y(new_n12209));
  OAI21xp33_ASAP7_75t_L     g11953(.A1(new_n12205), .A2(new_n12204), .B(new_n12208), .Y(new_n12210));
  AOI22xp33_ASAP7_75t_L     g11954(.A1(new_n5624), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n5901), .Y(new_n12211));
  OAI221xp5_ASAP7_75t_L     g11955(.A1(new_n5900), .A2(new_n1909), .B1(new_n5892), .B2(new_n2477), .C(new_n12211), .Y(new_n12212));
  XNOR2x2_ASAP7_75t_L       g11956(.A(\a[44] ), .B(new_n12212), .Y(new_n12213));
  NAND3xp33_ASAP7_75t_L     g11957(.A(new_n12209), .B(new_n12210), .C(new_n12213), .Y(new_n12214));
  AO21x2_ASAP7_75t_L        g11958(.A1(new_n12210), .A2(new_n12209), .B(new_n12213), .Y(new_n12215));
  NAND4xp25_ASAP7_75t_L     g11959(.A(new_n12215), .B(new_n11903), .C(new_n11916), .D(new_n12214), .Y(new_n12216));
  AO22x1_ASAP7_75t_L        g11960(.A1(new_n11903), .A2(new_n11916), .B1(new_n12214), .B2(new_n12215), .Y(new_n12217));
  AOI22xp33_ASAP7_75t_L     g11961(.A1(new_n4920), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n5167), .Y(new_n12218));
  OAI221xp5_ASAP7_75t_L     g11962(.A1(new_n5154), .A2(new_n2348), .B1(new_n5158), .B2(new_n2505), .C(new_n12218), .Y(new_n12219));
  XNOR2x2_ASAP7_75t_L       g11963(.A(\a[41] ), .B(new_n12219), .Y(new_n12220));
  NAND3xp33_ASAP7_75t_L     g11964(.A(new_n12217), .B(new_n12216), .C(new_n12220), .Y(new_n12221));
  AO21x2_ASAP7_75t_L        g11965(.A1(new_n12216), .A2(new_n12217), .B(new_n12220), .Y(new_n12222));
  NAND2xp33_ASAP7_75t_L     g11966(.A(new_n12221), .B(new_n12222), .Y(new_n12223));
  NOR2xp33_ASAP7_75t_L      g11967(.A(new_n11907), .B(new_n11909), .Y(new_n12224));
  NAND2xp33_ASAP7_75t_L     g11968(.A(new_n11913), .B(new_n12224), .Y(new_n12225));
  A2O1A1Ixp33_ASAP7_75t_L   g11969(.A1(new_n11920), .A2(new_n11640), .B(new_n11918), .C(new_n12225), .Y(new_n12226));
  NOR2xp33_ASAP7_75t_L      g11970(.A(new_n12226), .B(new_n12223), .Y(new_n12227));
  INVx1_ASAP7_75t_L         g11971(.A(new_n12224), .Y(new_n12228));
  INVx1_ASAP7_75t_L         g11972(.A(new_n12221), .Y(new_n12229));
  AOI21xp33_ASAP7_75t_L     g11973(.A1(new_n12217), .A2(new_n12216), .B(new_n12220), .Y(new_n12230));
  NOR2xp33_ASAP7_75t_L      g11974(.A(new_n12230), .B(new_n12229), .Y(new_n12231));
  O2A1O1Ixp33_ASAP7_75t_L   g11975(.A1(new_n12228), .A2(new_n11912), .B(new_n11925), .C(new_n12231), .Y(new_n12232));
  AOI22xp33_ASAP7_75t_L     g11976(.A1(new_n4283), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n4512), .Y(new_n12233));
  OAI221xp5_ASAP7_75t_L     g11977(.A1(new_n4277), .A2(new_n2688), .B1(new_n4499), .B2(new_n2990), .C(new_n12233), .Y(new_n12234));
  XNOR2x2_ASAP7_75t_L       g11978(.A(\a[38] ), .B(new_n12234), .Y(new_n12235));
  OAI21xp33_ASAP7_75t_L     g11979(.A1(new_n12227), .A2(new_n12232), .B(new_n12235), .Y(new_n12236));
  NAND3xp33_ASAP7_75t_L     g11980(.A(new_n12231), .B(new_n11925), .C(new_n12225), .Y(new_n12237));
  A2O1A1Ixp33_ASAP7_75t_L   g11981(.A1(new_n11913), .A2(new_n12224), .B(new_n11931), .C(new_n12223), .Y(new_n12238));
  INVx1_ASAP7_75t_L         g11982(.A(new_n12235), .Y(new_n12239));
  NAND3xp33_ASAP7_75t_L     g11983(.A(new_n12237), .B(new_n12238), .C(new_n12239), .Y(new_n12240));
  NAND3xp33_ASAP7_75t_L     g11984(.A(new_n11921), .B(new_n11925), .C(new_n11932), .Y(new_n12241));
  A2O1A1Ixp33_ASAP7_75t_L   g11985(.A1(new_n11933), .A2(new_n11929), .B(new_n11946), .C(new_n12241), .Y(new_n12242));
  NAND3xp33_ASAP7_75t_L     g11986(.A(new_n12236), .B(new_n12240), .C(new_n12242), .Y(new_n12243));
  NAND2xp33_ASAP7_75t_L     g11987(.A(new_n12240), .B(new_n12236), .Y(new_n12244));
  INVx1_ASAP7_75t_L         g11988(.A(new_n12242), .Y(new_n12245));
  NAND2xp33_ASAP7_75t_L     g11989(.A(new_n12245), .B(new_n12244), .Y(new_n12246));
  AOI22xp33_ASAP7_75t_L     g11990(.A1(new_n3633), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n3858), .Y(new_n12247));
  OAI221xp5_ASAP7_75t_L     g11991(.A1(new_n3853), .A2(new_n3207), .B1(new_n3856), .B2(new_n3572), .C(new_n12247), .Y(new_n12248));
  XNOR2x2_ASAP7_75t_L       g11992(.A(\a[35] ), .B(new_n12248), .Y(new_n12249));
  AND3x1_ASAP7_75t_L        g11993(.A(new_n12246), .B(new_n12249), .C(new_n12243), .Y(new_n12250));
  AOI21xp33_ASAP7_75t_L     g11994(.A1(new_n12246), .A2(new_n12243), .B(new_n12249), .Y(new_n12251));
  NOR2xp33_ASAP7_75t_L      g11995(.A(new_n12251), .B(new_n12250), .Y(new_n12252));
  NAND2xp33_ASAP7_75t_L     g11996(.A(\b[35] ), .B(new_n3030), .Y(new_n12253));
  OAI221xp5_ASAP7_75t_L     g11997(.A1(new_n3022), .A2(new_n4216), .B1(new_n3584), .B2(new_n3402), .C(new_n12253), .Y(new_n12254));
  AOI21xp33_ASAP7_75t_L     g11998(.A1(new_n6848), .A2(new_n3021), .B(new_n12254), .Y(new_n12255));
  NAND2xp33_ASAP7_75t_L     g11999(.A(\a[32] ), .B(new_n12255), .Y(new_n12256));
  A2O1A1Ixp33_ASAP7_75t_L   g12000(.A1(new_n6848), .A2(new_n3021), .B(new_n12254), .C(new_n3015), .Y(new_n12257));
  NAND2xp33_ASAP7_75t_L     g12001(.A(new_n12257), .B(new_n12256), .Y(new_n12258));
  AND2x2_ASAP7_75t_L        g12002(.A(new_n11950), .B(new_n11815), .Y(new_n12259));
  O2A1O1Ixp33_ASAP7_75t_L   g12003(.A1(new_n11937), .A2(new_n11941), .B(new_n11944), .C(new_n12259), .Y(new_n12260));
  XNOR2x2_ASAP7_75t_L       g12004(.A(new_n12258), .B(new_n12260), .Y(new_n12261));
  XNOR2x2_ASAP7_75t_L       g12005(.A(new_n12261), .B(new_n12252), .Y(new_n12262));
  NOR2xp33_ASAP7_75t_L      g12006(.A(new_n12150), .B(new_n12262), .Y(new_n12263));
  INVx1_ASAP7_75t_L         g12007(.A(new_n12263), .Y(new_n12264));
  NAND2xp33_ASAP7_75t_L     g12008(.A(new_n12150), .B(new_n12262), .Y(new_n12265));
  NAND4xp25_ASAP7_75t_L     g12009(.A(new_n12264), .B(new_n12135), .C(new_n12137), .D(new_n12265), .Y(new_n12266));
  NAND2xp33_ASAP7_75t_L     g12010(.A(new_n12135), .B(new_n12137), .Y(new_n12267));
  XNOR2x2_ASAP7_75t_L       g12011(.A(new_n12150), .B(new_n12262), .Y(new_n12268));
  NAND2xp33_ASAP7_75t_L     g12012(.A(new_n12267), .B(new_n12268), .Y(new_n12269));
  NAND2xp33_ASAP7_75t_L     g12013(.A(new_n12266), .B(new_n12269), .Y(new_n12270));
  XNOR2x2_ASAP7_75t_L       g12014(.A(new_n12130), .B(new_n12270), .Y(new_n12271));
  OR2x4_ASAP7_75t_L         g12015(.A(new_n12119), .B(new_n12271), .Y(new_n12272));
  NAND2xp33_ASAP7_75t_L     g12016(.A(new_n12119), .B(new_n12271), .Y(new_n12273));
  AND2x2_ASAP7_75t_L        g12017(.A(new_n12273), .B(new_n12272), .Y(new_n12274));
  NAND2xp33_ASAP7_75t_L     g12018(.A(new_n12111), .B(new_n12274), .Y(new_n12275));
  AO21x2_ASAP7_75t_L        g12019(.A1(new_n12273), .A2(new_n12272), .B(new_n12111), .Y(new_n12276));
  NAND2xp33_ASAP7_75t_L     g12020(.A(new_n12275), .B(new_n12276), .Y(new_n12277));
  XOR2x2_ASAP7_75t_L        g12021(.A(new_n12277), .B(new_n12102), .Y(new_n12278));
  NAND3xp33_ASAP7_75t_L     g12022(.A(new_n12089), .B(new_n12090), .C(new_n12278), .Y(new_n12279));
  INVx1_ASAP7_75t_L         g12023(.A(new_n12090), .Y(new_n12280));
  INVx1_ASAP7_75t_L         g12024(.A(new_n12278), .Y(new_n12281));
  OAI21xp33_ASAP7_75t_L     g12025(.A1(new_n12088), .A2(new_n12280), .B(new_n12281), .Y(new_n12282));
  NAND2xp33_ASAP7_75t_L     g12026(.A(new_n12279), .B(new_n12282), .Y(new_n12283));
  AOI22xp33_ASAP7_75t_L     g12027(.A1(new_n444), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n471), .Y(new_n12284));
  OAI221xp5_ASAP7_75t_L     g12028(.A1(new_n468), .A2(new_n9947), .B1(new_n469), .B2(new_n11446), .C(new_n12284), .Y(new_n12285));
  XNOR2x2_ASAP7_75t_L       g12029(.A(\a[8] ), .B(new_n12285), .Y(new_n12286));
  INVx1_ASAP7_75t_L         g12030(.A(new_n12286), .Y(new_n12287));
  NAND3xp33_ASAP7_75t_L     g12031(.A(new_n12036), .B(new_n12028), .C(new_n12287), .Y(new_n12288));
  O2A1O1Ixp33_ASAP7_75t_L   g12032(.A1(new_n12039), .A2(new_n12038), .B(new_n12028), .C(new_n12287), .Y(new_n12289));
  INVx1_ASAP7_75t_L         g12033(.A(new_n12289), .Y(new_n12290));
  NAND3xp33_ASAP7_75t_L     g12034(.A(new_n12283), .B(new_n12288), .C(new_n12290), .Y(new_n12291));
  AO21x2_ASAP7_75t_L        g12035(.A1(new_n12290), .A2(new_n12288), .B(new_n12283), .Y(new_n12292));
  NAND2xp33_ASAP7_75t_L     g12036(.A(new_n12291), .B(new_n12292), .Y(new_n12293));
  AOI22xp33_ASAP7_75t_L     g12037(.A1(new_n344), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n370), .Y(new_n12294));
  A2O1A1Ixp33_ASAP7_75t_L   g12038(.A1(new_n11470), .A2(new_n11473), .B(new_n366), .C(new_n12294), .Y(new_n12295));
  AOI21xp33_ASAP7_75t_L     g12039(.A1(new_n347), .A2(\b[62] ), .B(new_n12295), .Y(new_n12296));
  NAND2xp33_ASAP7_75t_L     g12040(.A(\a[5] ), .B(new_n12296), .Y(new_n12297));
  A2O1A1Ixp33_ASAP7_75t_L   g12041(.A1(\b[62] ), .A2(new_n347), .B(new_n12295), .C(new_n338), .Y(new_n12298));
  NAND2xp33_ASAP7_75t_L     g12042(.A(new_n12298), .B(new_n12297), .Y(new_n12299));
  AOI21xp33_ASAP7_75t_L     g12043(.A1(new_n12046), .A2(new_n12050), .B(new_n12052), .Y(new_n12300));
  NAND2xp33_ASAP7_75t_L     g12044(.A(new_n12299), .B(new_n12300), .Y(new_n12301));
  O2A1O1Ixp33_ASAP7_75t_L   g12045(.A1(new_n12054), .A2(new_n12053), .B(new_n12042), .C(new_n12299), .Y(new_n12302));
  INVx1_ASAP7_75t_L         g12046(.A(new_n12302), .Y(new_n12303));
  NAND2xp33_ASAP7_75t_L     g12047(.A(new_n12301), .B(new_n12303), .Y(new_n12304));
  NOR2xp33_ASAP7_75t_L      g12048(.A(new_n12293), .B(new_n12304), .Y(new_n12305));
  AND2x2_ASAP7_75t_L        g12049(.A(new_n12291), .B(new_n12292), .Y(new_n12306));
  AOI21xp33_ASAP7_75t_L     g12050(.A1(new_n12303), .A2(new_n12301), .B(new_n12306), .Y(new_n12307));
  OAI21xp33_ASAP7_75t_L     g12051(.A1(new_n12305), .A2(new_n12307), .B(new_n12082), .Y(new_n12308));
  NAND3xp33_ASAP7_75t_L     g12052(.A(new_n12306), .B(new_n12301), .C(new_n12303), .Y(new_n12309));
  NAND2xp33_ASAP7_75t_L     g12053(.A(new_n12293), .B(new_n12304), .Y(new_n12310));
  NAND4xp25_ASAP7_75t_L     g12054(.A(new_n12309), .B(new_n12310), .C(new_n12065), .D(new_n12067), .Y(new_n12311));
  NAND2xp33_ASAP7_75t_L     g12055(.A(new_n12311), .B(new_n12308), .Y(new_n12312));
  O2A1O1Ixp33_ASAP7_75t_L   g12056(.A1(new_n12070), .A2(new_n12079), .B(new_n12077), .C(new_n12312), .Y(new_n12313));
  AND2x2_ASAP7_75t_L        g12057(.A(new_n12311), .B(new_n12308), .Y(new_n12314));
  INVx1_ASAP7_75t_L         g12058(.A(new_n11783), .Y(new_n12315));
  A2O1A1Ixp33_ASAP7_75t_L   g12059(.A1(new_n11490), .A2(new_n11493), .B(new_n11491), .C(new_n11788), .Y(new_n12316));
  A2O1A1Ixp33_ASAP7_75t_L   g12060(.A1(new_n12316), .A2(new_n12315), .B(new_n12078), .C(new_n12077), .Y(new_n12317));
  NOR2xp33_ASAP7_75t_L      g12061(.A(new_n12314), .B(new_n12317), .Y(new_n12318));
  NOR2xp33_ASAP7_75t_L      g12062(.A(new_n12313), .B(new_n12318), .Y(\f[66] ));
  INVx1_ASAP7_75t_L         g12063(.A(new_n12311), .Y(new_n12320));
  OA21x2_ASAP7_75t_L        g12064(.A1(new_n12302), .A2(new_n12293), .B(new_n12301), .Y(new_n12321));
  INVx1_ASAP7_75t_L         g12065(.A(new_n11500), .Y(new_n12322));
  NOR2xp33_ASAP7_75t_L      g12066(.A(new_n11172), .B(new_n407), .Y(new_n12323));
  AOI221xp5_ASAP7_75t_L     g12067(.A1(\b[63] ), .A2(new_n347), .B1(new_n341), .B2(new_n12322), .C(new_n12323), .Y(new_n12324));
  XNOR2x2_ASAP7_75t_L       g12068(.A(\a[5] ), .B(new_n12324), .Y(new_n12325));
  A2O1A1O1Ixp25_ASAP7_75t_L g12069(.A1(new_n12282), .A2(new_n12279), .B(new_n12289), .C(new_n12288), .D(new_n12325), .Y(new_n12326));
  A2O1A1Ixp33_ASAP7_75t_L   g12070(.A1(new_n12279), .A2(new_n12282), .B(new_n12289), .C(new_n12288), .Y(new_n12327));
  INVx1_ASAP7_75t_L         g12071(.A(new_n12325), .Y(new_n12328));
  NOR2xp33_ASAP7_75t_L      g12072(.A(new_n12327), .B(new_n12328), .Y(new_n12329));
  NOR2xp33_ASAP7_75t_L      g12073(.A(new_n12326), .B(new_n12329), .Y(new_n12330));
  A2O1A1Ixp33_ASAP7_75t_L   g12074(.A1(new_n11792), .A2(new_n12009), .B(new_n12091), .C(new_n12100), .Y(new_n12331));
  AOI22xp33_ASAP7_75t_L     g12075(.A1(\b[56] ), .A2(new_n651), .B1(\b[58] ), .B2(new_n581), .Y(new_n12332));
  OAI221xp5_ASAP7_75t_L     g12076(.A1(new_n821), .A2(new_n9620), .B1(new_n577), .B2(new_n9925), .C(new_n12332), .Y(new_n12333));
  XNOR2x2_ASAP7_75t_L       g12077(.A(\a[11] ), .B(new_n12333), .Y(new_n12334));
  INVx1_ASAP7_75t_L         g12078(.A(new_n12334), .Y(new_n12335));
  A2O1A1O1Ixp25_ASAP7_75t_L g12079(.A1(new_n12101), .A2(new_n12098), .B(new_n12277), .C(new_n12331), .D(new_n12335), .Y(new_n12336));
  INVx1_ASAP7_75t_L         g12080(.A(new_n12336), .Y(new_n12337));
  A2O1A1Ixp33_ASAP7_75t_L   g12081(.A1(new_n12101), .A2(new_n12098), .B(new_n12277), .C(new_n12331), .Y(new_n12338));
  NOR2xp33_ASAP7_75t_L      g12082(.A(new_n12334), .B(new_n12338), .Y(new_n12339));
  INVx1_ASAP7_75t_L         g12083(.A(new_n12339), .Y(new_n12340));
  AOI22xp33_ASAP7_75t_L     g12084(.A1(new_n811), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n900), .Y(new_n12341));
  OAI221xp5_ASAP7_75t_L     g12085(.A1(new_n904), .A2(new_n8458), .B1(new_n898), .B2(new_n8768), .C(new_n12341), .Y(new_n12342));
  XNOR2x2_ASAP7_75t_L       g12086(.A(\a[14] ), .B(new_n12342), .Y(new_n12343));
  NAND3xp33_ASAP7_75t_L     g12087(.A(new_n12275), .B(new_n12109), .C(new_n12343), .Y(new_n12344));
  INVx1_ASAP7_75t_L         g12088(.A(new_n12343), .Y(new_n12345));
  A2O1A1Ixp33_ASAP7_75t_L   g12089(.A1(new_n12274), .A2(new_n12111), .B(new_n12110), .C(new_n12345), .Y(new_n12346));
  NAND2xp33_ASAP7_75t_L     g12090(.A(new_n12346), .B(new_n12344), .Y(new_n12347));
  AOI22xp33_ASAP7_75t_L     g12091(.A1(new_n1360), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1581), .Y(new_n12348));
  OAI221xp5_ASAP7_75t_L     g12092(.A1(new_n1373), .A2(new_n6830), .B1(new_n1359), .B2(new_n7323), .C(new_n12348), .Y(new_n12349));
  XNOR2x2_ASAP7_75t_L       g12093(.A(\a[20] ), .B(new_n12349), .Y(new_n12350));
  NAND2xp33_ASAP7_75t_L     g12094(.A(new_n12123), .B(new_n12126), .Y(new_n12351));
  OAI211xp5_ASAP7_75t_L     g12095(.A1(new_n12130), .A2(new_n12270), .B(new_n12350), .C(new_n12351), .Y(new_n12352));
  INVx1_ASAP7_75t_L         g12096(.A(new_n12352), .Y(new_n12353));
  O2A1O1Ixp33_ASAP7_75t_L   g12097(.A1(new_n12130), .A2(new_n12270), .B(new_n12351), .C(new_n12350), .Y(new_n12354));
  NOR2xp33_ASAP7_75t_L      g12098(.A(new_n12354), .B(new_n12353), .Y(new_n12355));
  AOI22xp33_ASAP7_75t_L     g12099(.A1(new_n1704), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n1837), .Y(new_n12356));
  OAI221xp5_ASAP7_75t_L     g12100(.A1(new_n1699), .A2(new_n6321), .B1(new_n1827), .B2(new_n6573), .C(new_n12356), .Y(new_n12357));
  XNOR2x2_ASAP7_75t_L       g12101(.A(\a[23] ), .B(new_n12357), .Y(new_n12358));
  INVx1_ASAP7_75t_L         g12102(.A(new_n12358), .Y(new_n12359));
  AOI31xp33_ASAP7_75t_L     g12103(.A1(new_n12264), .A2(new_n12265), .A3(new_n12135), .B(new_n12136), .Y(new_n12360));
  NAND2xp33_ASAP7_75t_L     g12104(.A(new_n12359), .B(new_n12360), .Y(new_n12361));
  O2A1O1Ixp33_ASAP7_75t_L   g12105(.A1(new_n12267), .A2(new_n12268), .B(new_n12137), .C(new_n12359), .Y(new_n12362));
  INVx1_ASAP7_75t_L         g12106(.A(new_n12362), .Y(new_n12363));
  AOI22xp33_ASAP7_75t_L     g12107(.A1(new_n2114), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n2259), .Y(new_n12364));
  OAI221xp5_ASAP7_75t_L     g12108(.A1(new_n2109), .A2(new_n5338), .B1(new_n2257), .B2(new_n6338), .C(new_n12364), .Y(new_n12365));
  XNOR2x2_ASAP7_75t_L       g12109(.A(\a[26] ), .B(new_n12365), .Y(new_n12366));
  INVx1_ASAP7_75t_L         g12110(.A(new_n12366), .Y(new_n12367));
  NOR3xp33_ASAP7_75t_L      g12111(.A(new_n12263), .B(new_n12367), .C(new_n12145), .Y(new_n12368));
  INVx1_ASAP7_75t_L         g12112(.A(new_n12145), .Y(new_n12369));
  O2A1O1Ixp33_ASAP7_75t_L   g12113(.A1(new_n12150), .A2(new_n12262), .B(new_n12369), .C(new_n12366), .Y(new_n12370));
  NOR2xp33_ASAP7_75t_L      g12114(.A(new_n12370), .B(new_n12368), .Y(new_n12371));
  INVx1_ASAP7_75t_L         g12115(.A(new_n4431), .Y(new_n12372));
  NAND2xp33_ASAP7_75t_L     g12116(.A(\b[36] ), .B(new_n3030), .Y(new_n12373));
  OAI221xp5_ASAP7_75t_L     g12117(.A1(new_n3022), .A2(new_n4424), .B1(new_n3804), .B2(new_n3402), .C(new_n12373), .Y(new_n12374));
  AOI21xp33_ASAP7_75t_L     g12118(.A1(new_n12372), .A2(new_n3021), .B(new_n12374), .Y(new_n12375));
  NAND2xp33_ASAP7_75t_L     g12119(.A(\a[32] ), .B(new_n12375), .Y(new_n12376));
  A2O1A1Ixp33_ASAP7_75t_L   g12120(.A1(new_n12372), .A2(new_n3021), .B(new_n12374), .C(new_n3015), .Y(new_n12377));
  NAND2xp33_ASAP7_75t_L     g12121(.A(new_n12377), .B(new_n12376), .Y(new_n12378));
  MAJIxp5_ASAP7_75t_L       g12122(.A(new_n12244), .B(new_n12245), .C(new_n12249), .Y(new_n12379));
  XNOR2x2_ASAP7_75t_L       g12123(.A(new_n12378), .B(new_n12379), .Y(new_n12380));
  AOI22xp33_ASAP7_75t_L     g12124(.A1(new_n3633), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n3858), .Y(new_n12381));
  OAI221xp5_ASAP7_75t_L     g12125(.A1(new_n3853), .A2(new_n3565), .B1(new_n3856), .B2(new_n3591), .C(new_n12381), .Y(new_n12382));
  XNOR2x2_ASAP7_75t_L       g12126(.A(\a[35] ), .B(new_n12382), .Y(new_n12383));
  INVx1_ASAP7_75t_L         g12127(.A(new_n12383), .Y(new_n12384));
  AOI21xp33_ASAP7_75t_L     g12128(.A1(new_n12237), .A2(new_n12239), .B(new_n12232), .Y(new_n12385));
  AOI22xp33_ASAP7_75t_L     g12129(.A1(new_n5624), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n5901), .Y(new_n12386));
  OAI221xp5_ASAP7_75t_L     g12130(.A1(new_n5900), .A2(new_n1929), .B1(new_n5892), .B2(new_n2075), .C(new_n12386), .Y(new_n12387));
  XNOR2x2_ASAP7_75t_L       g12131(.A(\a[44] ), .B(new_n12387), .Y(new_n12388));
  O2A1O1Ixp33_ASAP7_75t_L   g12132(.A1(new_n11887), .A2(new_n11888), .B(new_n11882), .C(new_n12198), .Y(new_n12389));
  AOI22xp33_ASAP7_75t_L     g12133(.A1(\b[5] ), .A2(new_n10939), .B1(\b[7] ), .B2(new_n10938), .Y(new_n12390));
  OAI221xp5_ASAP7_75t_L     g12134(.A1(new_n10937), .A2(new_n418), .B1(new_n10629), .B2(new_n425), .C(new_n12390), .Y(new_n12391));
  XNOR2x2_ASAP7_75t_L       g12135(.A(\a[62] ), .B(new_n12391), .Y(new_n12392));
  NOR2xp33_ASAP7_75t_L      g12136(.A(new_n298), .B(new_n11535), .Y(new_n12393));
  O2A1O1Ixp33_ASAP7_75t_L   g12137(.A1(new_n11247), .A2(new_n11249), .B(\b[4] ), .C(new_n12393), .Y(new_n12394));
  NAND2xp33_ASAP7_75t_L     g12138(.A(\a[2] ), .B(new_n12394), .Y(new_n12395));
  A2O1A1Ixp33_ASAP7_75t_L   g12139(.A1(new_n11533), .A2(\b[4] ), .B(new_n12393), .C(new_n262), .Y(new_n12396));
  AND2x2_ASAP7_75t_L        g12140(.A(new_n12396), .B(new_n12395), .Y(new_n12397));
  XNOR2x2_ASAP7_75t_L       g12141(.A(new_n12397), .B(new_n12392), .Y(new_n12398));
  A2O1A1O1Ixp25_ASAP7_75t_L g12142(.A1(new_n11533), .A2(\b[3] ), .B(new_n12157), .C(\a[2] ), .D(new_n12168), .Y(new_n12399));
  NAND2xp33_ASAP7_75t_L     g12143(.A(new_n12399), .B(new_n12398), .Y(new_n12400));
  O2A1O1Ixp33_ASAP7_75t_L   g12144(.A1(new_n12161), .A2(new_n12167), .B(new_n12158), .C(new_n12398), .Y(new_n12401));
  INVx1_ASAP7_75t_L         g12145(.A(new_n12401), .Y(new_n12402));
  AOI22xp33_ASAP7_75t_L     g12146(.A1(new_n9700), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n10027), .Y(new_n12403));
  OAI221xp5_ASAP7_75t_L     g12147(.A1(new_n10024), .A2(new_n540), .B1(new_n9696), .B2(new_n624), .C(new_n12403), .Y(new_n12404));
  XNOR2x2_ASAP7_75t_L       g12148(.A(\a[59] ), .B(new_n12404), .Y(new_n12405));
  NAND3xp33_ASAP7_75t_L     g12149(.A(new_n12402), .B(new_n12400), .C(new_n12405), .Y(new_n12406));
  AO21x2_ASAP7_75t_L        g12150(.A1(new_n12400), .A2(new_n12402), .B(new_n12405), .Y(new_n12407));
  AND2x2_ASAP7_75t_L        g12151(.A(new_n12406), .B(new_n12407), .Y(new_n12408));
  AND2x2_ASAP7_75t_L        g12152(.A(new_n12177), .B(new_n12174), .Y(new_n12409));
  NOR2xp33_ASAP7_75t_L      g12153(.A(new_n12173), .B(new_n12409), .Y(new_n12410));
  XNOR2x2_ASAP7_75t_L       g12154(.A(new_n12408), .B(new_n12410), .Y(new_n12411));
  AOI22xp33_ASAP7_75t_L     g12155(.A1(new_n8831), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n9115), .Y(new_n12412));
  OAI221xp5_ASAP7_75t_L     g12156(.A1(new_n10343), .A2(new_n760), .B1(new_n10016), .B2(new_n790), .C(new_n12412), .Y(new_n12413));
  XNOR2x2_ASAP7_75t_L       g12157(.A(\a[56] ), .B(new_n12413), .Y(new_n12414));
  INVx1_ASAP7_75t_L         g12158(.A(new_n12414), .Y(new_n12415));
  XNOR2x2_ASAP7_75t_L       g12159(.A(new_n12415), .B(new_n12411), .Y(new_n12416));
  INVx1_ASAP7_75t_L         g12160(.A(new_n12180), .Y(new_n12417));
  MAJx2_ASAP7_75t_L         g12161(.A(new_n12178), .B(new_n12154), .C(new_n12417), .Y(new_n12418));
  XOR2x2_ASAP7_75t_L        g12162(.A(new_n12418), .B(new_n12416), .Y(new_n12419));
  AOI22xp33_ASAP7_75t_L     g12163(.A1(new_n7960), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n8537), .Y(new_n12420));
  OAI221xp5_ASAP7_75t_L     g12164(.A1(new_n8817), .A2(new_n942), .B1(new_n7957), .B2(new_n1035), .C(new_n12420), .Y(new_n12421));
  XNOR2x2_ASAP7_75t_L       g12165(.A(\a[53] ), .B(new_n12421), .Y(new_n12422));
  XNOR2x2_ASAP7_75t_L       g12166(.A(new_n12422), .B(new_n12419), .Y(new_n12423));
  MAJIxp5_ASAP7_75t_L       g12167(.A(new_n12182), .B(new_n12151), .C(new_n12187), .Y(new_n12424));
  INVx1_ASAP7_75t_L         g12168(.A(new_n12424), .Y(new_n12425));
  XNOR2x2_ASAP7_75t_L       g12169(.A(new_n12425), .B(new_n12423), .Y(new_n12426));
  AOI22xp33_ASAP7_75t_L     g12170(.A1(new_n7111), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n7391), .Y(new_n12427));
  OAI221xp5_ASAP7_75t_L     g12171(.A1(new_n8558), .A2(new_n1313), .B1(new_n8237), .B2(new_n1438), .C(new_n12427), .Y(new_n12428));
  XNOR2x2_ASAP7_75t_L       g12172(.A(\a[50] ), .B(new_n12428), .Y(new_n12429));
  INVx1_ASAP7_75t_L         g12173(.A(new_n12429), .Y(new_n12430));
  XNOR2x2_ASAP7_75t_L       g12174(.A(new_n12430), .B(new_n12426), .Y(new_n12431));
  NAND2xp33_ASAP7_75t_L     g12175(.A(new_n12191), .B(new_n12196), .Y(new_n12432));
  XOR2x2_ASAP7_75t_L        g12176(.A(new_n12432), .B(new_n12431), .Y(new_n12433));
  AOI22xp33_ASAP7_75t_L     g12177(.A1(new_n6376), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n6648), .Y(new_n12434));
  OAI221xp5_ASAP7_75t_L     g12178(.A1(new_n6646), .A2(new_n1655), .B1(new_n6636), .B2(new_n1780), .C(new_n12434), .Y(new_n12435));
  XNOR2x2_ASAP7_75t_L       g12179(.A(\a[47] ), .B(new_n12435), .Y(new_n12436));
  INVx1_ASAP7_75t_L         g12180(.A(new_n12436), .Y(new_n12437));
  XNOR2x2_ASAP7_75t_L       g12181(.A(new_n12437), .B(new_n12433), .Y(new_n12438));
  OA21x2_ASAP7_75t_L        g12182(.A1(new_n12389), .A2(new_n12205), .B(new_n12438), .Y(new_n12439));
  NOR3xp33_ASAP7_75t_L      g12183(.A(new_n12438), .B(new_n12205), .C(new_n12389), .Y(new_n12440));
  NOR3xp33_ASAP7_75t_L      g12184(.A(new_n12439), .B(new_n12440), .C(new_n12388), .Y(new_n12441));
  INVx1_ASAP7_75t_L         g12185(.A(new_n12388), .Y(new_n12442));
  NOR2xp33_ASAP7_75t_L      g12186(.A(new_n12440), .B(new_n12439), .Y(new_n12443));
  NOR2xp33_ASAP7_75t_L      g12187(.A(new_n12442), .B(new_n12443), .Y(new_n12444));
  NAND2xp33_ASAP7_75t_L     g12188(.A(new_n12210), .B(new_n12214), .Y(new_n12445));
  OAI21xp33_ASAP7_75t_L     g12189(.A1(new_n12441), .A2(new_n12444), .B(new_n12445), .Y(new_n12446));
  NOR2xp33_ASAP7_75t_L      g12190(.A(new_n12441), .B(new_n12444), .Y(new_n12447));
  NAND3xp33_ASAP7_75t_L     g12191(.A(new_n12447), .B(new_n12214), .C(new_n12210), .Y(new_n12448));
  AOI22xp33_ASAP7_75t_L     g12192(.A1(new_n4920), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n5167), .Y(new_n12449));
  OAI221xp5_ASAP7_75t_L     g12193(.A1(new_n5154), .A2(new_n2497), .B1(new_n5158), .B2(new_n2672), .C(new_n12449), .Y(new_n12450));
  XNOR2x2_ASAP7_75t_L       g12194(.A(\a[41] ), .B(new_n12450), .Y(new_n12451));
  AND3x1_ASAP7_75t_L        g12195(.A(new_n12448), .B(new_n12451), .C(new_n12446), .Y(new_n12452));
  AOI21xp33_ASAP7_75t_L     g12196(.A1(new_n12448), .A2(new_n12446), .B(new_n12451), .Y(new_n12453));
  AND2x2_ASAP7_75t_L        g12197(.A(new_n12216), .B(new_n12221), .Y(new_n12454));
  NOR3xp33_ASAP7_75t_L      g12198(.A(new_n12452), .B(new_n12453), .C(new_n12454), .Y(new_n12455));
  OA21x2_ASAP7_75t_L        g12199(.A1(new_n12453), .A2(new_n12452), .B(new_n12454), .Y(new_n12456));
  AOI22xp33_ASAP7_75t_L     g12200(.A1(new_n4283), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n4512), .Y(new_n12457));
  OAI221xp5_ASAP7_75t_L     g12201(.A1(new_n4277), .A2(new_n2982), .B1(new_n4499), .B2(new_n3187), .C(new_n12457), .Y(new_n12458));
  XNOR2x2_ASAP7_75t_L       g12202(.A(\a[38] ), .B(new_n12458), .Y(new_n12459));
  OAI21xp33_ASAP7_75t_L     g12203(.A1(new_n12455), .A2(new_n12456), .B(new_n12459), .Y(new_n12460));
  OR3x1_ASAP7_75t_L         g12204(.A(new_n12452), .B(new_n12453), .C(new_n12454), .Y(new_n12461));
  OAI21xp33_ASAP7_75t_L     g12205(.A1(new_n12453), .A2(new_n12452), .B(new_n12454), .Y(new_n12462));
  INVx1_ASAP7_75t_L         g12206(.A(new_n12459), .Y(new_n12463));
  NAND3xp33_ASAP7_75t_L     g12207(.A(new_n12461), .B(new_n12462), .C(new_n12463), .Y(new_n12464));
  NAND2xp33_ASAP7_75t_L     g12208(.A(new_n12460), .B(new_n12464), .Y(new_n12465));
  NOR2xp33_ASAP7_75t_L      g12209(.A(new_n12385), .B(new_n12465), .Y(new_n12466));
  INVx1_ASAP7_75t_L         g12210(.A(new_n12385), .Y(new_n12467));
  AOI21xp33_ASAP7_75t_L     g12211(.A1(new_n12461), .A2(new_n12462), .B(new_n12463), .Y(new_n12468));
  NOR3xp33_ASAP7_75t_L      g12212(.A(new_n12456), .B(new_n12459), .C(new_n12455), .Y(new_n12469));
  NOR2xp33_ASAP7_75t_L      g12213(.A(new_n12469), .B(new_n12468), .Y(new_n12470));
  NOR2xp33_ASAP7_75t_L      g12214(.A(new_n12467), .B(new_n12470), .Y(new_n12471));
  OAI21xp33_ASAP7_75t_L     g12215(.A1(new_n12466), .A2(new_n12471), .B(new_n12384), .Y(new_n12472));
  NAND2xp33_ASAP7_75t_L     g12216(.A(new_n12467), .B(new_n12470), .Y(new_n12473));
  NAND2xp33_ASAP7_75t_L     g12217(.A(new_n12385), .B(new_n12465), .Y(new_n12474));
  NAND3xp33_ASAP7_75t_L     g12218(.A(new_n12473), .B(new_n12474), .C(new_n12383), .Y(new_n12475));
  NAND3xp33_ASAP7_75t_L     g12219(.A(new_n12380), .B(new_n12472), .C(new_n12475), .Y(new_n12476));
  AO21x2_ASAP7_75t_L        g12220(.A1(new_n12475), .A2(new_n12472), .B(new_n12380), .Y(new_n12477));
  NAND2xp33_ASAP7_75t_L     g12221(.A(new_n12476), .B(new_n12477), .Y(new_n12478));
  INVx1_ASAP7_75t_L         g12222(.A(new_n12478), .Y(new_n12479));
  NOR2xp33_ASAP7_75t_L      g12223(.A(new_n12261), .B(new_n12252), .Y(new_n12480));
  NAND2xp33_ASAP7_75t_L     g12224(.A(\b[39] ), .B(new_n2553), .Y(new_n12481));
  OAI221xp5_ASAP7_75t_L     g12225(.A1(new_n2545), .A2(new_n4869), .B1(new_n4632), .B2(new_n2747), .C(new_n12481), .Y(new_n12482));
  AOI21xp33_ASAP7_75t_L     g12226(.A1(new_n4876), .A2(new_n2544), .B(new_n12482), .Y(new_n12483));
  NAND2xp33_ASAP7_75t_L     g12227(.A(\a[29] ), .B(new_n12483), .Y(new_n12484));
  A2O1A1Ixp33_ASAP7_75t_L   g12228(.A1(new_n4876), .A2(new_n2544), .B(new_n12482), .C(new_n2538), .Y(new_n12485));
  AND2x2_ASAP7_75t_L        g12229(.A(new_n12485), .B(new_n12484), .Y(new_n12486));
  A2O1A1Ixp33_ASAP7_75t_L   g12230(.A1(new_n12260), .A2(new_n12258), .B(new_n12480), .C(new_n12486), .Y(new_n12487));
  INVx1_ASAP7_75t_L         g12231(.A(new_n12487), .Y(new_n12488));
  AND2x2_ASAP7_75t_L        g12232(.A(new_n12258), .B(new_n12260), .Y(new_n12489));
  NOR3xp33_ASAP7_75t_L      g12233(.A(new_n12480), .B(new_n12489), .C(new_n12486), .Y(new_n12490));
  OAI21xp33_ASAP7_75t_L     g12234(.A1(new_n12490), .A2(new_n12488), .B(new_n12479), .Y(new_n12491));
  INVx1_ASAP7_75t_L         g12235(.A(new_n12490), .Y(new_n12492));
  NAND3xp33_ASAP7_75t_L     g12236(.A(new_n12492), .B(new_n12487), .C(new_n12478), .Y(new_n12493));
  NAND2xp33_ASAP7_75t_L     g12237(.A(new_n12493), .B(new_n12491), .Y(new_n12494));
  XNOR2x2_ASAP7_75t_L       g12238(.A(new_n12494), .B(new_n12371), .Y(new_n12495));
  NAND3xp33_ASAP7_75t_L     g12239(.A(new_n12495), .B(new_n12361), .C(new_n12363), .Y(new_n12496));
  INVx1_ASAP7_75t_L         g12240(.A(new_n12361), .Y(new_n12497));
  NOR3xp33_ASAP7_75t_L      g12241(.A(new_n12494), .B(new_n12370), .C(new_n12368), .Y(new_n12498));
  AOI21xp33_ASAP7_75t_L     g12242(.A1(new_n12493), .A2(new_n12491), .B(new_n12371), .Y(new_n12499));
  OAI22xp33_ASAP7_75t_L     g12243(.A1(new_n12497), .A2(new_n12362), .B1(new_n12499), .B2(new_n12498), .Y(new_n12500));
  NAND3xp33_ASAP7_75t_L     g12244(.A(new_n12355), .B(new_n12496), .C(new_n12500), .Y(new_n12501));
  NAND2xp33_ASAP7_75t_L     g12245(.A(new_n12500), .B(new_n12496), .Y(new_n12502));
  OAI21xp33_ASAP7_75t_L     g12246(.A1(new_n12353), .A2(new_n12354), .B(new_n12502), .Y(new_n12503));
  NAND2xp33_ASAP7_75t_L     g12247(.A(new_n12501), .B(new_n12503), .Y(new_n12504));
  AOI22xp33_ASAP7_75t_L     g12248(.A1(new_n1076), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1253), .Y(new_n12505));
  OAI221xp5_ASAP7_75t_L     g12249(.A1(new_n1154), .A2(new_n7616), .B1(new_n1156), .B2(new_n7906), .C(new_n12505), .Y(new_n12506));
  XNOR2x2_ASAP7_75t_L       g12250(.A(\a[17] ), .B(new_n12506), .Y(new_n12507));
  A2O1A1Ixp33_ASAP7_75t_L   g12251(.A1(new_n12003), .A2(new_n11990), .B(new_n12114), .C(new_n12272), .Y(new_n12508));
  NOR2xp33_ASAP7_75t_L      g12252(.A(new_n12507), .B(new_n12508), .Y(new_n12509));
  INVx1_ASAP7_75t_L         g12253(.A(new_n12507), .Y(new_n12510));
  O2A1O1Ixp33_ASAP7_75t_L   g12254(.A1(new_n12119), .A2(new_n12271), .B(new_n12118), .C(new_n12510), .Y(new_n12511));
  OA21x2_ASAP7_75t_L        g12255(.A1(new_n12511), .A2(new_n12509), .B(new_n12504), .Y(new_n12512));
  NOR3xp33_ASAP7_75t_L      g12256(.A(new_n12509), .B(new_n12511), .C(new_n12504), .Y(new_n12513));
  NOR2xp33_ASAP7_75t_L      g12257(.A(new_n12513), .B(new_n12512), .Y(new_n12514));
  XNOR2x2_ASAP7_75t_L       g12258(.A(new_n12347), .B(new_n12514), .Y(new_n12515));
  NAND3xp33_ASAP7_75t_L     g12259(.A(new_n12515), .B(new_n12340), .C(new_n12337), .Y(new_n12516));
  XOR2x2_ASAP7_75t_L        g12260(.A(new_n12347), .B(new_n12514), .Y(new_n12517));
  OAI21xp33_ASAP7_75t_L     g12261(.A1(new_n12339), .A2(new_n12336), .B(new_n12517), .Y(new_n12518));
  NAND2xp33_ASAP7_75t_L     g12262(.A(new_n12518), .B(new_n12516), .Y(new_n12519));
  NAND2xp33_ASAP7_75t_L     g12263(.A(\b[60] ), .B(new_n447), .Y(new_n12520));
  OAI221xp5_ASAP7_75t_L     g12264(.A1(new_n515), .A2(new_n10847), .B1(new_n9947), .B2(new_n516), .C(new_n12520), .Y(new_n12521));
  AOI21xp33_ASAP7_75t_L     g12265(.A1(new_n11759), .A2(new_n441), .B(new_n12521), .Y(new_n12522));
  NAND2xp33_ASAP7_75t_L     g12266(.A(\a[8] ), .B(new_n12522), .Y(new_n12523));
  A2O1A1Ixp33_ASAP7_75t_L   g12267(.A1(new_n11759), .A2(new_n441), .B(new_n12521), .C(new_n435), .Y(new_n12524));
  NAND2xp33_ASAP7_75t_L     g12268(.A(new_n12524), .B(new_n12523), .Y(new_n12525));
  AOI21xp33_ASAP7_75t_L     g12269(.A1(new_n12278), .A2(new_n12090), .B(new_n12088), .Y(new_n12526));
  NAND2xp33_ASAP7_75t_L     g12270(.A(new_n12525), .B(new_n12526), .Y(new_n12527));
  O2A1O1Ixp33_ASAP7_75t_L   g12271(.A1(new_n12280), .A2(new_n12281), .B(new_n12089), .C(new_n12525), .Y(new_n12528));
  INVx1_ASAP7_75t_L         g12272(.A(new_n12528), .Y(new_n12529));
  NAND3xp33_ASAP7_75t_L     g12273(.A(new_n12529), .B(new_n12519), .C(new_n12527), .Y(new_n12530));
  INVx1_ASAP7_75t_L         g12274(.A(new_n12530), .Y(new_n12531));
  AOI21xp33_ASAP7_75t_L     g12275(.A1(new_n12529), .A2(new_n12527), .B(new_n12519), .Y(new_n12532));
  NOR3xp33_ASAP7_75t_L      g12276(.A(new_n12330), .B(new_n12531), .C(new_n12532), .Y(new_n12533));
  NOR2xp33_ASAP7_75t_L      g12277(.A(new_n12532), .B(new_n12531), .Y(new_n12534));
  NOR3xp33_ASAP7_75t_L      g12278(.A(new_n12534), .B(new_n12329), .C(new_n12326), .Y(new_n12535));
  NOR3xp33_ASAP7_75t_L      g12279(.A(new_n12535), .B(new_n12533), .C(new_n12321), .Y(new_n12536));
  OA21x2_ASAP7_75t_L        g12280(.A1(new_n12533), .A2(new_n12535), .B(new_n12321), .Y(new_n12537));
  NOR2xp33_ASAP7_75t_L      g12281(.A(new_n12536), .B(new_n12537), .Y(new_n12538));
  A2O1A1Ixp33_ASAP7_75t_L   g12282(.A1(new_n12317), .A2(new_n12314), .B(new_n12320), .C(new_n12538), .Y(new_n12539));
  INVx1_ASAP7_75t_L         g12283(.A(new_n12539), .Y(new_n12540));
  A2O1A1Ixp33_ASAP7_75t_L   g12284(.A1(new_n12075), .A2(new_n12077), .B(new_n12312), .C(new_n12311), .Y(new_n12541));
  NOR2xp33_ASAP7_75t_L      g12285(.A(new_n12538), .B(new_n12541), .Y(new_n12542));
  NOR2xp33_ASAP7_75t_L      g12286(.A(new_n12542), .B(new_n12540), .Y(\f[67] ));
  A2O1A1Ixp33_ASAP7_75t_L   g12287(.A1(new_n12030), .A2(new_n12029), .B(new_n12031), .C(new_n12036), .Y(new_n12544));
  O2A1O1Ixp33_ASAP7_75t_L   g12288(.A1(new_n12286), .A2(new_n12544), .B(new_n12291), .C(new_n12328), .Y(new_n12545));
  O2A1O1Ixp33_ASAP7_75t_L   g12289(.A1(new_n12326), .A2(new_n12329), .B(new_n12534), .C(new_n12545), .Y(new_n12546));
  A2O1A1O1Ixp25_ASAP7_75t_L g12290(.A1(new_n12101), .A2(new_n12098), .B(new_n12277), .C(new_n12331), .D(new_n12334), .Y(new_n12547));
  INVx1_ASAP7_75t_L         g12291(.A(new_n12547), .Y(new_n12548));
  NAND2xp33_ASAP7_75t_L     g12292(.A(\b[61] ), .B(new_n447), .Y(new_n12549));
  OAI221xp5_ASAP7_75t_L     g12293(.A1(new_n515), .A2(new_n11172), .B1(new_n10250), .B2(new_n516), .C(new_n12549), .Y(new_n12550));
  AOI21xp33_ASAP7_75t_L     g12294(.A1(new_n11180), .A2(new_n441), .B(new_n12550), .Y(new_n12551));
  NAND2xp33_ASAP7_75t_L     g12295(.A(\a[8] ), .B(new_n12551), .Y(new_n12552));
  A2O1A1Ixp33_ASAP7_75t_L   g12296(.A1(new_n11180), .A2(new_n441), .B(new_n12550), .C(new_n435), .Y(new_n12553));
  NAND2xp33_ASAP7_75t_L     g12297(.A(new_n12553), .B(new_n12552), .Y(new_n12554));
  A2O1A1O1Ixp25_ASAP7_75t_L g12298(.A1(new_n12337), .A2(new_n12340), .B(new_n12517), .C(new_n12548), .D(new_n12554), .Y(new_n12555));
  O2A1O1Ixp33_ASAP7_75t_L   g12299(.A1(new_n12336), .A2(new_n12339), .B(new_n12515), .C(new_n12547), .Y(new_n12556));
  NAND2xp33_ASAP7_75t_L     g12300(.A(new_n12554), .B(new_n12556), .Y(new_n12557));
  INVx1_ASAP7_75t_L         g12301(.A(new_n12557), .Y(new_n12558));
  AOI22xp33_ASAP7_75t_L     g12302(.A1(\b[57] ), .A2(new_n651), .B1(\b[59] ), .B2(new_n581), .Y(new_n12559));
  OAI221xp5_ASAP7_75t_L     g12303(.A1(new_n821), .A2(new_n9920), .B1(new_n577), .B2(new_n11152), .C(new_n12559), .Y(new_n12560));
  XNOR2x2_ASAP7_75t_L       g12304(.A(\a[11] ), .B(new_n12560), .Y(new_n12561));
  OAI311xp33_ASAP7_75t_L    g12305(.A1(new_n12347), .A2(new_n12513), .A3(new_n12512), .B1(new_n12561), .C1(new_n12346), .Y(new_n12562));
  INVx1_ASAP7_75t_L         g12306(.A(new_n12346), .Y(new_n12563));
  INVx1_ASAP7_75t_L         g12307(.A(new_n12561), .Y(new_n12564));
  A2O1A1Ixp33_ASAP7_75t_L   g12308(.A1(new_n12514), .A2(new_n12344), .B(new_n12563), .C(new_n12564), .Y(new_n12565));
  AOI22xp33_ASAP7_75t_L     g12309(.A1(new_n811), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n900), .Y(new_n12566));
  OAI221xp5_ASAP7_75t_L     g12310(.A1(new_n904), .A2(new_n8762), .B1(new_n898), .B2(new_n9331), .C(new_n12566), .Y(new_n12567));
  XNOR2x2_ASAP7_75t_L       g12311(.A(new_n806), .B(new_n12567), .Y(new_n12568));
  INVx1_ASAP7_75t_L         g12312(.A(new_n12568), .Y(new_n12569));
  MAJx2_ASAP7_75t_L         g12313(.A(new_n12504), .B(new_n12510), .C(new_n12508), .Y(new_n12570));
  XNOR2x2_ASAP7_75t_L       g12314(.A(new_n12569), .B(new_n12570), .Y(new_n12571));
  NAND2xp33_ASAP7_75t_L     g12315(.A(\b[52] ), .B(new_n1080), .Y(new_n12572));
  OAI221xp5_ASAP7_75t_L     g12316(.A1(new_n1259), .A2(new_n8165), .B1(new_n7616), .B2(new_n1158), .C(new_n12572), .Y(new_n12573));
  AOI21xp33_ASAP7_75t_L     g12317(.A1(new_n8173), .A2(new_n1073), .B(new_n12573), .Y(new_n12574));
  NAND2xp33_ASAP7_75t_L     g12318(.A(\a[17] ), .B(new_n12574), .Y(new_n12575));
  A2O1A1Ixp33_ASAP7_75t_L   g12319(.A1(new_n8173), .A2(new_n1073), .B(new_n12573), .C(new_n1071), .Y(new_n12576));
  AND2x2_ASAP7_75t_L        g12320(.A(new_n12576), .B(new_n12575), .Y(new_n12577));
  INVx1_ASAP7_75t_L         g12321(.A(new_n12577), .Y(new_n12578));
  AOI31xp33_ASAP7_75t_L     g12322(.A1(new_n12355), .A2(new_n12496), .A3(new_n12500), .B(new_n12353), .Y(new_n12579));
  NAND2xp33_ASAP7_75t_L     g12323(.A(new_n12578), .B(new_n12579), .Y(new_n12580));
  INVx1_ASAP7_75t_L         g12324(.A(new_n12580), .Y(new_n12581));
  O2A1O1Ixp33_ASAP7_75t_L   g12325(.A1(new_n12354), .A2(new_n12502), .B(new_n12352), .C(new_n12578), .Y(new_n12582));
  AOI22xp33_ASAP7_75t_L     g12326(.A1(new_n1360), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1581), .Y(new_n12583));
  INVx1_ASAP7_75t_L         g12327(.A(new_n12583), .Y(new_n12584));
  AOI221xp5_ASAP7_75t_L     g12328(.A1(\b[49] ), .A2(new_n1362), .B1(new_n1365), .B2(new_n7601), .C(new_n12584), .Y(new_n12585));
  XNOR2x2_ASAP7_75t_L       g12329(.A(new_n1356), .B(new_n12585), .Y(new_n12586));
  O2A1O1Ixp33_ASAP7_75t_L   g12330(.A1(new_n12267), .A2(new_n12268), .B(new_n12137), .C(new_n12358), .Y(new_n12587));
  O2A1O1Ixp33_ASAP7_75t_L   g12331(.A1(new_n12497), .A2(new_n12362), .B(new_n12495), .C(new_n12587), .Y(new_n12588));
  XOR2x2_ASAP7_75t_L        g12332(.A(new_n12586), .B(new_n12588), .Y(new_n12589));
  INVx1_ASAP7_75t_L         g12333(.A(new_n12370), .Y(new_n12590));
  AOI22xp33_ASAP7_75t_L     g12334(.A1(new_n1704), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1837), .Y(new_n12591));
  OAI221xp5_ASAP7_75t_L     g12335(.A1(new_n1699), .A2(new_n6568), .B1(new_n1827), .B2(new_n6820), .C(new_n12591), .Y(new_n12592));
  XNOR2x2_ASAP7_75t_L       g12336(.A(\a[23] ), .B(new_n12592), .Y(new_n12593));
  OAI211xp5_ASAP7_75t_L     g12337(.A1(new_n12368), .A2(new_n12494), .B(new_n12593), .C(new_n12590), .Y(new_n12594));
  O2A1O1Ixp33_ASAP7_75t_L   g12338(.A1(new_n12368), .A2(new_n12494), .B(new_n12590), .C(new_n12593), .Y(new_n12595));
  INVx1_ASAP7_75t_L         g12339(.A(new_n12595), .Y(new_n12596));
  NAND2xp33_ASAP7_75t_L     g12340(.A(new_n12378), .B(new_n12379), .Y(new_n12597));
  AOI22xp33_ASAP7_75t_L     g12341(.A1(new_n2552), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n2736), .Y(new_n12598));
  OAI221xp5_ASAP7_75t_L     g12342(.A1(new_n2547), .A2(new_n4869), .B1(new_n2734), .B2(new_n5327), .C(new_n12598), .Y(new_n12599));
  XNOR2x2_ASAP7_75t_L       g12343(.A(\a[29] ), .B(new_n12599), .Y(new_n12600));
  AND3x1_ASAP7_75t_L        g12344(.A(new_n12477), .B(new_n12600), .C(new_n12597), .Y(new_n12601));
  A2O1A1O1Ixp25_ASAP7_75t_L g12345(.A1(new_n12475), .A2(new_n12472), .B(new_n12380), .C(new_n12597), .D(new_n12600), .Y(new_n12602));
  AOI22xp33_ASAP7_75t_L     g12346(.A1(new_n7960), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n8537), .Y(new_n12603));
  OAI221xp5_ASAP7_75t_L     g12347(.A1(new_n8817), .A2(new_n1030), .B1(new_n7957), .B2(new_n1209), .C(new_n12603), .Y(new_n12604));
  XNOR2x2_ASAP7_75t_L       g12348(.A(\a[53] ), .B(new_n12604), .Y(new_n12605));
  INVx1_ASAP7_75t_L         g12349(.A(new_n12605), .Y(new_n12606));
  INVx1_ASAP7_75t_L         g12350(.A(new_n12410), .Y(new_n12607));
  NAND2xp33_ASAP7_75t_L     g12351(.A(new_n12415), .B(new_n12411), .Y(new_n12608));
  AOI22xp33_ASAP7_75t_L     g12352(.A1(\b[6] ), .A2(new_n10939), .B1(\b[8] ), .B2(new_n10938), .Y(new_n12609));
  OAI21xp33_ASAP7_75t_L     g12353(.A1(new_n10629), .A2(new_n494), .B(new_n12609), .Y(new_n12610));
  AOI21xp33_ASAP7_75t_L     g12354(.A1(new_n10632), .A2(\b[7] ), .B(new_n12610), .Y(new_n12611));
  NAND2xp33_ASAP7_75t_L     g12355(.A(\a[62] ), .B(new_n12611), .Y(new_n12612));
  A2O1A1Ixp33_ASAP7_75t_L   g12356(.A1(\b[7] ), .A2(new_n10632), .B(new_n12610), .C(new_n10622), .Y(new_n12613));
  NAND2xp33_ASAP7_75t_L     g12357(.A(new_n12613), .B(new_n12612), .Y(new_n12614));
  NOR2xp33_ASAP7_75t_L      g12358(.A(new_n324), .B(new_n11535), .Y(new_n12615));
  O2A1O1Ixp33_ASAP7_75t_L   g12359(.A1(new_n11247), .A2(new_n11249), .B(\b[5] ), .C(new_n12615), .Y(new_n12616));
  NAND2xp33_ASAP7_75t_L     g12360(.A(\a[2] ), .B(new_n12616), .Y(new_n12617));
  INVx1_ASAP7_75t_L         g12361(.A(new_n12617), .Y(new_n12618));
  INVx1_ASAP7_75t_L         g12362(.A(new_n12615), .Y(new_n12619));
  O2A1O1Ixp33_ASAP7_75t_L   g12363(.A1(new_n354), .A2(new_n11253), .B(new_n12619), .C(\a[2] ), .Y(new_n12620));
  NOR2xp33_ASAP7_75t_L      g12364(.A(new_n12620), .B(new_n12618), .Y(new_n12621));
  INVx1_ASAP7_75t_L         g12365(.A(new_n12621), .Y(new_n12622));
  XNOR2x2_ASAP7_75t_L       g12366(.A(new_n12622), .B(new_n12614), .Y(new_n12623));
  A2O1A1Ixp33_ASAP7_75t_L   g12367(.A1(new_n11533), .A2(\b[4] ), .B(new_n12393), .C(\a[2] ), .Y(new_n12624));
  A2O1A1Ixp33_ASAP7_75t_L   g12368(.A1(new_n12395), .A2(new_n12396), .B(new_n12392), .C(new_n12624), .Y(new_n12625));
  INVx1_ASAP7_75t_L         g12369(.A(new_n12625), .Y(new_n12626));
  NAND2xp33_ASAP7_75t_L     g12370(.A(new_n12626), .B(new_n12623), .Y(new_n12627));
  OR2x4_ASAP7_75t_L         g12371(.A(new_n12626), .B(new_n12623), .Y(new_n12628));
  NAND2xp33_ASAP7_75t_L     g12372(.A(new_n12627), .B(new_n12628), .Y(new_n12629));
  AOI22xp33_ASAP7_75t_L     g12373(.A1(new_n9700), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n10027), .Y(new_n12630));
  OAI221xp5_ASAP7_75t_L     g12374(.A1(new_n10024), .A2(new_n617), .B1(new_n9696), .B2(new_n685), .C(new_n12630), .Y(new_n12631));
  XNOR2x2_ASAP7_75t_L       g12375(.A(\a[59] ), .B(new_n12631), .Y(new_n12632));
  NAND2xp33_ASAP7_75t_L     g12376(.A(new_n12632), .B(new_n12629), .Y(new_n12633));
  NOR2xp33_ASAP7_75t_L      g12377(.A(new_n12632), .B(new_n12629), .Y(new_n12634));
  INVx1_ASAP7_75t_L         g12378(.A(new_n12634), .Y(new_n12635));
  NAND2xp33_ASAP7_75t_L     g12379(.A(new_n12400), .B(new_n12406), .Y(new_n12636));
  INVx1_ASAP7_75t_L         g12380(.A(new_n12636), .Y(new_n12637));
  NAND3xp33_ASAP7_75t_L     g12381(.A(new_n12635), .B(new_n12633), .C(new_n12637), .Y(new_n12638));
  INVx1_ASAP7_75t_L         g12382(.A(new_n12400), .Y(new_n12639));
  NAND2xp33_ASAP7_75t_L     g12383(.A(new_n12633), .B(new_n12635), .Y(new_n12640));
  A2O1A1Ixp33_ASAP7_75t_L   g12384(.A1(new_n12402), .A2(new_n12405), .B(new_n12639), .C(new_n12640), .Y(new_n12641));
  AOI22xp33_ASAP7_75t_L     g12385(.A1(new_n8831), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n9115), .Y(new_n12642));
  OAI221xp5_ASAP7_75t_L     g12386(.A1(new_n10343), .A2(new_n784), .B1(new_n10016), .B2(new_n875), .C(new_n12642), .Y(new_n12643));
  XNOR2x2_ASAP7_75t_L       g12387(.A(\a[56] ), .B(new_n12643), .Y(new_n12644));
  NAND3xp33_ASAP7_75t_L     g12388(.A(new_n12641), .B(new_n12638), .C(new_n12644), .Y(new_n12645));
  AO21x2_ASAP7_75t_L        g12389(.A1(new_n12638), .A2(new_n12641), .B(new_n12644), .Y(new_n12646));
  AND2x2_ASAP7_75t_L        g12390(.A(new_n12645), .B(new_n12646), .Y(new_n12647));
  O2A1O1Ixp33_ASAP7_75t_L   g12391(.A1(new_n12408), .A2(new_n12607), .B(new_n12608), .C(new_n12647), .Y(new_n12648));
  INVx1_ASAP7_75t_L         g12392(.A(new_n12647), .Y(new_n12649));
  A2O1A1Ixp33_ASAP7_75t_L   g12393(.A1(new_n12407), .A2(new_n12406), .B(new_n12607), .C(new_n12608), .Y(new_n12650));
  NOR2xp33_ASAP7_75t_L      g12394(.A(new_n12650), .B(new_n12649), .Y(new_n12651));
  NOR3xp33_ASAP7_75t_L      g12395(.A(new_n12651), .B(new_n12648), .C(new_n12606), .Y(new_n12652));
  XNOR2x2_ASAP7_75t_L       g12396(.A(new_n12647), .B(new_n12650), .Y(new_n12653));
  NOR2xp33_ASAP7_75t_L      g12397(.A(new_n12605), .B(new_n12653), .Y(new_n12654));
  NOR2xp33_ASAP7_75t_L      g12398(.A(new_n12652), .B(new_n12654), .Y(new_n12655));
  NAND2xp33_ASAP7_75t_L     g12399(.A(new_n12418), .B(new_n12416), .Y(new_n12656));
  NAND2xp33_ASAP7_75t_L     g12400(.A(new_n12422), .B(new_n12419), .Y(new_n12657));
  NAND2xp33_ASAP7_75t_L     g12401(.A(new_n12656), .B(new_n12657), .Y(new_n12658));
  XNOR2x2_ASAP7_75t_L       g12402(.A(new_n12658), .B(new_n12655), .Y(new_n12659));
  AOI22xp33_ASAP7_75t_L     g12403(.A1(new_n7111), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n7391), .Y(new_n12660));
  OAI221xp5_ASAP7_75t_L     g12404(.A1(new_n8558), .A2(new_n1432), .B1(new_n8237), .B2(new_n1547), .C(new_n12660), .Y(new_n12661));
  XNOR2x2_ASAP7_75t_L       g12405(.A(\a[50] ), .B(new_n12661), .Y(new_n12662));
  XNOR2x2_ASAP7_75t_L       g12406(.A(new_n12662), .B(new_n12659), .Y(new_n12663));
  MAJIxp5_ASAP7_75t_L       g12407(.A(new_n12423), .B(new_n12425), .C(new_n12430), .Y(new_n12664));
  NOR2xp33_ASAP7_75t_L      g12408(.A(new_n12664), .B(new_n12663), .Y(new_n12665));
  AND2x2_ASAP7_75t_L        g12409(.A(new_n12662), .B(new_n12659), .Y(new_n12666));
  NOR2xp33_ASAP7_75t_L      g12410(.A(new_n12662), .B(new_n12659), .Y(new_n12667));
  NOR2xp33_ASAP7_75t_L      g12411(.A(new_n12667), .B(new_n12666), .Y(new_n12668));
  INVx1_ASAP7_75t_L         g12412(.A(new_n12664), .Y(new_n12669));
  NOR2xp33_ASAP7_75t_L      g12413(.A(new_n12669), .B(new_n12668), .Y(new_n12670));
  NOR2xp33_ASAP7_75t_L      g12414(.A(new_n12665), .B(new_n12670), .Y(new_n12671));
  AOI22xp33_ASAP7_75t_L     g12415(.A1(new_n6376), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n6648), .Y(new_n12672));
  OAI221xp5_ASAP7_75t_L     g12416(.A1(new_n6646), .A2(new_n1774), .B1(new_n6636), .B2(new_n1915), .C(new_n12672), .Y(new_n12673));
  XNOR2x2_ASAP7_75t_L       g12417(.A(\a[47] ), .B(new_n12673), .Y(new_n12674));
  NAND2xp33_ASAP7_75t_L     g12418(.A(new_n12674), .B(new_n12671), .Y(new_n12675));
  INVx1_ASAP7_75t_L         g12419(.A(new_n12674), .Y(new_n12676));
  OAI21xp33_ASAP7_75t_L     g12420(.A1(new_n12665), .A2(new_n12670), .B(new_n12676), .Y(new_n12677));
  NAND2xp33_ASAP7_75t_L     g12421(.A(new_n12677), .B(new_n12675), .Y(new_n12678));
  O2A1O1Ixp33_ASAP7_75t_L   g12422(.A1(new_n12188), .A2(new_n12190), .B(new_n12196), .C(new_n12431), .Y(new_n12679));
  NOR2xp33_ASAP7_75t_L      g12423(.A(new_n12437), .B(new_n12433), .Y(new_n12680));
  NOR2xp33_ASAP7_75t_L      g12424(.A(new_n12679), .B(new_n12680), .Y(new_n12681));
  NOR2xp33_ASAP7_75t_L      g12425(.A(new_n12681), .B(new_n12678), .Y(new_n12682));
  AOI211xp5_ASAP7_75t_L     g12426(.A1(new_n12675), .A2(new_n12677), .B(new_n12680), .C(new_n12679), .Y(new_n12683));
  NOR2xp33_ASAP7_75t_L      g12427(.A(new_n12683), .B(new_n12682), .Y(new_n12684));
  AOI22xp33_ASAP7_75t_L     g12428(.A1(new_n5624), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n5901), .Y(new_n12685));
  OAI221xp5_ASAP7_75t_L     g12429(.A1(new_n5900), .A2(new_n2067), .B1(new_n5892), .B2(new_n2355), .C(new_n12685), .Y(new_n12686));
  XNOR2x2_ASAP7_75t_L       g12430(.A(\a[44] ), .B(new_n12686), .Y(new_n12687));
  XNOR2x2_ASAP7_75t_L       g12431(.A(new_n12687), .B(new_n12684), .Y(new_n12688));
  O2A1O1Ixp33_ASAP7_75t_L   g12432(.A1(new_n12389), .A2(new_n12205), .B(new_n12438), .C(new_n12441), .Y(new_n12689));
  XNOR2x2_ASAP7_75t_L       g12433(.A(new_n12689), .B(new_n12688), .Y(new_n12690));
  AOI22xp33_ASAP7_75t_L     g12434(.A1(new_n4920), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n5167), .Y(new_n12691));
  OAI221xp5_ASAP7_75t_L     g12435(.A1(new_n5154), .A2(new_n2666), .B1(new_n5158), .B2(new_n2695), .C(new_n12691), .Y(new_n12692));
  XNOR2x2_ASAP7_75t_L       g12436(.A(\a[41] ), .B(new_n12692), .Y(new_n12693));
  NAND2xp33_ASAP7_75t_L     g12437(.A(new_n12693), .B(new_n12690), .Y(new_n12694));
  XOR2x2_ASAP7_75t_L        g12438(.A(new_n12687), .B(new_n12684), .Y(new_n12695));
  NAND2xp33_ASAP7_75t_L     g12439(.A(new_n12689), .B(new_n12695), .Y(new_n12696));
  A2O1A1Ixp33_ASAP7_75t_L   g12440(.A1(new_n12443), .A2(new_n12442), .B(new_n12439), .C(new_n12688), .Y(new_n12697));
  NAND2xp33_ASAP7_75t_L     g12441(.A(new_n12696), .B(new_n12697), .Y(new_n12698));
  INVx1_ASAP7_75t_L         g12442(.A(new_n12693), .Y(new_n12699));
  NAND2xp33_ASAP7_75t_L     g12443(.A(new_n12699), .B(new_n12698), .Y(new_n12700));
  NAND2xp33_ASAP7_75t_L     g12444(.A(new_n12694), .B(new_n12700), .Y(new_n12701));
  NAND3xp33_ASAP7_75t_L     g12445(.A(new_n12448), .B(new_n12446), .C(new_n12451), .Y(new_n12702));
  A2O1A1Ixp33_ASAP7_75t_L   g12446(.A1(new_n12214), .A2(new_n12210), .B(new_n12447), .C(new_n12702), .Y(new_n12703));
  INVx1_ASAP7_75t_L         g12447(.A(new_n12703), .Y(new_n12704));
  NOR2xp33_ASAP7_75t_L      g12448(.A(new_n12701), .B(new_n12704), .Y(new_n12705));
  XNOR2x2_ASAP7_75t_L       g12449(.A(new_n12699), .B(new_n12690), .Y(new_n12706));
  NOR2xp33_ASAP7_75t_L      g12450(.A(new_n12703), .B(new_n12706), .Y(new_n12707));
  AOI22xp33_ASAP7_75t_L     g12451(.A1(new_n4283), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n4512), .Y(new_n12708));
  OAI221xp5_ASAP7_75t_L     g12452(.A1(new_n4277), .A2(new_n3180), .B1(new_n4499), .B2(new_n11047), .C(new_n12708), .Y(new_n12709));
  XNOR2x2_ASAP7_75t_L       g12453(.A(\a[38] ), .B(new_n12709), .Y(new_n12710));
  OAI21xp33_ASAP7_75t_L     g12454(.A1(new_n12707), .A2(new_n12705), .B(new_n12710), .Y(new_n12711));
  INVx1_ASAP7_75t_L         g12455(.A(new_n12447), .Y(new_n12712));
  A2O1A1Ixp33_ASAP7_75t_L   g12456(.A1(new_n12445), .A2(new_n12712), .B(new_n12452), .C(new_n12706), .Y(new_n12713));
  NAND2xp33_ASAP7_75t_L     g12457(.A(new_n12701), .B(new_n12704), .Y(new_n12714));
  INVx1_ASAP7_75t_L         g12458(.A(new_n12710), .Y(new_n12715));
  NAND3xp33_ASAP7_75t_L     g12459(.A(new_n12713), .B(new_n12714), .C(new_n12715), .Y(new_n12716));
  NAND2xp33_ASAP7_75t_L     g12460(.A(new_n12462), .B(new_n12464), .Y(new_n12717));
  NAND3xp33_ASAP7_75t_L     g12461(.A(new_n12716), .B(new_n12711), .C(new_n12717), .Y(new_n12718));
  AO21x2_ASAP7_75t_L        g12462(.A1(new_n12711), .A2(new_n12716), .B(new_n12717), .Y(new_n12719));
  AOI22xp33_ASAP7_75t_L     g12463(.A1(new_n3633), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n3858), .Y(new_n12720));
  OAI221xp5_ASAP7_75t_L     g12464(.A1(new_n3853), .A2(new_n3584), .B1(new_n3856), .B2(new_n10137), .C(new_n12720), .Y(new_n12721));
  XNOR2x2_ASAP7_75t_L       g12465(.A(\a[35] ), .B(new_n12721), .Y(new_n12722));
  NAND3xp33_ASAP7_75t_L     g12466(.A(new_n12719), .B(new_n12718), .C(new_n12722), .Y(new_n12723));
  AND3x1_ASAP7_75t_L        g12467(.A(new_n12716), .B(new_n12711), .C(new_n12717), .Y(new_n12724));
  AOI21xp33_ASAP7_75t_L     g12468(.A1(new_n12716), .A2(new_n12711), .B(new_n12717), .Y(new_n12725));
  INVx1_ASAP7_75t_L         g12469(.A(new_n12722), .Y(new_n12726));
  OAI21xp33_ASAP7_75t_L     g12470(.A1(new_n12725), .A2(new_n12724), .B(new_n12726), .Y(new_n12727));
  NAND2xp33_ASAP7_75t_L     g12471(.A(new_n12723), .B(new_n12727), .Y(new_n12728));
  NOR2xp33_ASAP7_75t_L      g12472(.A(new_n4632), .B(new_n3022), .Y(new_n12729));
  AOI221xp5_ASAP7_75t_L     g12473(.A1(\b[36] ), .A2(new_n3258), .B1(\b[37] ), .B2(new_n3030), .C(new_n12729), .Y(new_n12730));
  OAI211xp5_ASAP7_75t_L     g12474(.A1(new_n3256), .A2(new_n4641), .B(\a[32] ), .C(new_n12730), .Y(new_n12731));
  O2A1O1Ixp33_ASAP7_75t_L   g12475(.A1(new_n3256), .A2(new_n4641), .B(new_n12730), .C(\a[32] ), .Y(new_n12732));
  INVx1_ASAP7_75t_L         g12476(.A(new_n12732), .Y(new_n12733));
  AND2x2_ASAP7_75t_L        g12477(.A(new_n12731), .B(new_n12733), .Y(new_n12734));
  INVx1_ASAP7_75t_L         g12478(.A(new_n12734), .Y(new_n12735));
  MAJIxp5_ASAP7_75t_L       g12479(.A(new_n12465), .B(new_n12383), .C(new_n12385), .Y(new_n12736));
  NAND2xp33_ASAP7_75t_L     g12480(.A(new_n12735), .B(new_n12736), .Y(new_n12737));
  A2O1A1Ixp33_ASAP7_75t_L   g12481(.A1(new_n12473), .A2(new_n12383), .B(new_n12471), .C(new_n12734), .Y(new_n12738));
  NAND2xp33_ASAP7_75t_L     g12482(.A(new_n12737), .B(new_n12738), .Y(new_n12739));
  NAND2xp33_ASAP7_75t_L     g12483(.A(new_n12739), .B(new_n12728), .Y(new_n12740));
  NAND4xp25_ASAP7_75t_L     g12484(.A(new_n12727), .B(new_n12723), .C(new_n12737), .D(new_n12738), .Y(new_n12741));
  NAND2xp33_ASAP7_75t_L     g12485(.A(new_n12741), .B(new_n12740), .Y(new_n12742));
  NOR3xp33_ASAP7_75t_L      g12486(.A(new_n12742), .B(new_n12602), .C(new_n12601), .Y(new_n12743));
  OA21x2_ASAP7_75t_L        g12487(.A1(new_n12602), .A2(new_n12601), .B(new_n12742), .Y(new_n12744));
  NOR2xp33_ASAP7_75t_L      g12488(.A(new_n12743), .B(new_n12744), .Y(new_n12745));
  NOR2xp33_ASAP7_75t_L      g12489(.A(new_n12489), .B(new_n12480), .Y(new_n12746));
  MAJIxp5_ASAP7_75t_L       g12490(.A(new_n12478), .B(new_n12486), .C(new_n12746), .Y(new_n12747));
  INVx1_ASAP7_75t_L         g12491(.A(new_n5835), .Y(new_n12748));
  NAND2xp33_ASAP7_75t_L     g12492(.A(\b[43] ), .B(new_n2115), .Y(new_n12749));
  OAI221xp5_ASAP7_75t_L     g12493(.A1(new_n2107), .A2(new_n5829), .B1(new_n5338), .B2(new_n2269), .C(new_n12749), .Y(new_n12750));
  AOI21xp33_ASAP7_75t_L     g12494(.A1(new_n12748), .A2(new_n2106), .B(new_n12750), .Y(new_n12751));
  NAND2xp33_ASAP7_75t_L     g12495(.A(\a[26] ), .B(new_n12751), .Y(new_n12752));
  A2O1A1Ixp33_ASAP7_75t_L   g12496(.A1(new_n12748), .A2(new_n2106), .B(new_n12750), .C(new_n2100), .Y(new_n12753));
  NAND2xp33_ASAP7_75t_L     g12497(.A(new_n12753), .B(new_n12752), .Y(new_n12754));
  XNOR2x2_ASAP7_75t_L       g12498(.A(new_n12754), .B(new_n12747), .Y(new_n12755));
  NOR2xp33_ASAP7_75t_L      g12499(.A(new_n12745), .B(new_n12755), .Y(new_n12756));
  AND2x2_ASAP7_75t_L        g12500(.A(new_n12745), .B(new_n12755), .Y(new_n12757));
  NOR2xp33_ASAP7_75t_L      g12501(.A(new_n12756), .B(new_n12757), .Y(new_n12758));
  NAND3xp33_ASAP7_75t_L     g12502(.A(new_n12758), .B(new_n12596), .C(new_n12594), .Y(new_n12759));
  AO21x2_ASAP7_75t_L        g12503(.A1(new_n12594), .A2(new_n12596), .B(new_n12758), .Y(new_n12760));
  NAND2xp33_ASAP7_75t_L     g12504(.A(new_n12759), .B(new_n12760), .Y(new_n12761));
  XNOR2x2_ASAP7_75t_L       g12505(.A(new_n12761), .B(new_n12589), .Y(new_n12762));
  NOR3xp33_ASAP7_75t_L      g12506(.A(new_n12762), .B(new_n12581), .C(new_n12582), .Y(new_n12763));
  INVx1_ASAP7_75t_L         g12507(.A(new_n12582), .Y(new_n12764));
  XOR2x2_ASAP7_75t_L        g12508(.A(new_n12761), .B(new_n12589), .Y(new_n12765));
  AOI21xp33_ASAP7_75t_L     g12509(.A1(new_n12764), .A2(new_n12580), .B(new_n12765), .Y(new_n12766));
  NOR2xp33_ASAP7_75t_L      g12510(.A(new_n12766), .B(new_n12763), .Y(new_n12767));
  XNOR2x2_ASAP7_75t_L       g12511(.A(new_n12767), .B(new_n12571), .Y(new_n12768));
  NAND3xp33_ASAP7_75t_L     g12512(.A(new_n12768), .B(new_n12565), .C(new_n12562), .Y(new_n12769));
  AO21x2_ASAP7_75t_L        g12513(.A1(new_n12562), .A2(new_n12565), .B(new_n12768), .Y(new_n12770));
  AND2x2_ASAP7_75t_L        g12514(.A(new_n12769), .B(new_n12770), .Y(new_n12771));
  OAI21xp33_ASAP7_75t_L     g12515(.A1(new_n12555), .A2(new_n12558), .B(new_n12771), .Y(new_n12772));
  INVx1_ASAP7_75t_L         g12516(.A(new_n12555), .Y(new_n12773));
  NAND2xp33_ASAP7_75t_L     g12517(.A(new_n12769), .B(new_n12770), .Y(new_n12774));
  NAND3xp33_ASAP7_75t_L     g12518(.A(new_n12774), .B(new_n12557), .C(new_n12773), .Y(new_n12775));
  INVx1_ASAP7_75t_L         g12519(.A(new_n12527), .Y(new_n12776));
  A2O1A1Ixp33_ASAP7_75t_L   g12520(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n341), .Y(new_n12777));
  A2O1A1Ixp33_ASAP7_75t_L   g12521(.A1(new_n12777), .A2(new_n407), .B(new_n11468), .C(\a[5] ), .Y(new_n12778));
  O2A1O1Ixp33_ASAP7_75t_L   g12522(.A1(new_n366), .A2(new_n12060), .B(new_n407), .C(new_n11468), .Y(new_n12779));
  NAND2xp33_ASAP7_75t_L     g12523(.A(new_n338), .B(new_n12779), .Y(new_n12780));
  AND2x2_ASAP7_75t_L        g12524(.A(new_n12780), .B(new_n12778), .Y(new_n12781));
  INVx1_ASAP7_75t_L         g12525(.A(new_n12781), .Y(new_n12782));
  A2O1A1Ixp33_ASAP7_75t_L   g12526(.A1(new_n12529), .A2(new_n12519), .B(new_n12776), .C(new_n12782), .Y(new_n12783));
  NAND3xp33_ASAP7_75t_L     g12527(.A(new_n12530), .B(new_n12527), .C(new_n12781), .Y(new_n12784));
  NAND4xp25_ASAP7_75t_L     g12528(.A(new_n12772), .B(new_n12784), .C(new_n12783), .D(new_n12775), .Y(new_n12785));
  NAND2xp33_ASAP7_75t_L     g12529(.A(new_n12775), .B(new_n12772), .Y(new_n12786));
  NAND2xp33_ASAP7_75t_L     g12530(.A(new_n12783), .B(new_n12784), .Y(new_n12787));
  NAND2xp33_ASAP7_75t_L     g12531(.A(new_n12787), .B(new_n12786), .Y(new_n12788));
  NAND2xp33_ASAP7_75t_L     g12532(.A(new_n12785), .B(new_n12788), .Y(new_n12789));
  XOR2x2_ASAP7_75t_L        g12533(.A(new_n12546), .B(new_n12789), .Y(new_n12790));
  A2O1A1Ixp33_ASAP7_75t_L   g12534(.A1(new_n12541), .A2(new_n12538), .B(new_n12536), .C(new_n12790), .Y(new_n12791));
  INVx1_ASAP7_75t_L         g12535(.A(new_n12791), .Y(new_n12792));
  INVx1_ASAP7_75t_L         g12536(.A(new_n12313), .Y(new_n12793));
  INVx1_ASAP7_75t_L         g12537(.A(new_n12536), .Y(new_n12794));
  A2O1A1Ixp33_ASAP7_75t_L   g12538(.A1(new_n12793), .A2(new_n12311), .B(new_n12537), .C(new_n12794), .Y(new_n12795));
  NOR2xp33_ASAP7_75t_L      g12539(.A(new_n12790), .B(new_n12795), .Y(new_n12796));
  NOR2xp33_ASAP7_75t_L      g12540(.A(new_n12792), .B(new_n12796), .Y(\f[68] ));
  INVx1_ASAP7_75t_L         g12541(.A(new_n12789), .Y(new_n12798));
  A2O1A1Ixp33_ASAP7_75t_L   g12542(.A1(new_n12325), .A2(new_n12327), .B(new_n12533), .C(new_n12798), .Y(new_n12799));
  INVx1_ASAP7_75t_L         g12543(.A(new_n12799), .Y(new_n12800));
  INVx1_ASAP7_75t_L         g12544(.A(new_n12554), .Y(new_n12801));
  A2O1A1O1Ixp25_ASAP7_75t_L g12545(.A1(new_n12337), .A2(new_n12340), .B(new_n12517), .C(new_n12548), .D(new_n12801), .Y(new_n12802));
  INVx1_ASAP7_75t_L         g12546(.A(new_n12802), .Y(new_n12803));
  AOI22xp33_ASAP7_75t_L     g12547(.A1(new_n444), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n471), .Y(new_n12804));
  A2O1A1Ixp33_ASAP7_75t_L   g12548(.A1(new_n11470), .A2(new_n11473), .B(new_n469), .C(new_n12804), .Y(new_n12805));
  AOI21xp33_ASAP7_75t_L     g12549(.A1(new_n447), .A2(\b[62] ), .B(new_n12805), .Y(new_n12806));
  NAND2xp33_ASAP7_75t_L     g12550(.A(\a[8] ), .B(new_n12806), .Y(new_n12807));
  A2O1A1Ixp33_ASAP7_75t_L   g12551(.A1(\b[62] ), .A2(new_n447), .B(new_n12805), .C(new_n435), .Y(new_n12808));
  NAND2xp33_ASAP7_75t_L     g12552(.A(new_n12808), .B(new_n12807), .Y(new_n12809));
  A2O1A1O1Ixp25_ASAP7_75t_L g12553(.A1(new_n12557), .A2(new_n12773), .B(new_n12774), .C(new_n12803), .D(new_n12809), .Y(new_n12810));
  A2O1A1Ixp33_ASAP7_75t_L   g12554(.A1(new_n12557), .A2(new_n12773), .B(new_n12774), .C(new_n12803), .Y(new_n12811));
  AOI21xp33_ASAP7_75t_L     g12555(.A1(new_n12808), .A2(new_n12807), .B(new_n12811), .Y(new_n12812));
  NOR2xp33_ASAP7_75t_L      g12556(.A(new_n12810), .B(new_n12812), .Y(new_n12813));
  AOI22xp33_ASAP7_75t_L     g12557(.A1(\b[58] ), .A2(new_n651), .B1(\b[60] ), .B2(new_n581), .Y(new_n12814));
  OAI221xp5_ASAP7_75t_L     g12558(.A1(new_n821), .A2(new_n9947), .B1(new_n577), .B2(new_n11446), .C(new_n12814), .Y(new_n12815));
  XNOR2x2_ASAP7_75t_L       g12559(.A(\a[11] ), .B(new_n12815), .Y(new_n12816));
  INVx1_ASAP7_75t_L         g12560(.A(new_n12816), .Y(new_n12817));
  NAND2xp33_ASAP7_75t_L     g12561(.A(new_n12565), .B(new_n12769), .Y(new_n12818));
  XNOR2x2_ASAP7_75t_L       g12562(.A(new_n12817), .B(new_n12818), .Y(new_n12819));
  O2A1O1Ixp33_ASAP7_75t_L   g12563(.A1(new_n12119), .A2(new_n12271), .B(new_n12118), .C(new_n12507), .Y(new_n12820));
  O2A1O1Ixp33_ASAP7_75t_L   g12564(.A1(new_n12511), .A2(new_n12509), .B(new_n12504), .C(new_n12820), .Y(new_n12821));
  NAND2xp33_ASAP7_75t_L     g12565(.A(new_n12568), .B(new_n12821), .Y(new_n12822));
  A2O1A1Ixp33_ASAP7_75t_L   g12566(.A1(new_n12508), .A2(new_n12510), .B(new_n12512), .C(new_n12569), .Y(new_n12823));
  AOI22xp33_ASAP7_75t_L     g12567(.A1(new_n811), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n900), .Y(new_n12824));
  OAI221xp5_ASAP7_75t_L     g12568(.A1(new_n904), .A2(new_n9323), .B1(new_n898), .B2(new_n9627), .C(new_n12824), .Y(new_n12825));
  XNOR2x2_ASAP7_75t_L       g12569(.A(\a[14] ), .B(new_n12825), .Y(new_n12826));
  A2O1A1Ixp33_ASAP7_75t_L   g12570(.A1(new_n12508), .A2(new_n12510), .B(new_n12512), .C(new_n12568), .Y(new_n12827));
  A2O1A1O1Ixp25_ASAP7_75t_L g12571(.A1(new_n12823), .A2(new_n12822), .B(new_n12767), .C(new_n12827), .D(new_n12826), .Y(new_n12828));
  INVx1_ASAP7_75t_L         g12572(.A(new_n12828), .Y(new_n12829));
  INVx1_ASAP7_75t_L         g12573(.A(new_n12827), .Y(new_n12830));
  O2A1O1Ixp33_ASAP7_75t_L   g12574(.A1(new_n12763), .A2(new_n12766), .B(new_n12571), .C(new_n12830), .Y(new_n12831));
  NAND2xp33_ASAP7_75t_L     g12575(.A(new_n12826), .B(new_n12831), .Y(new_n12832));
  AOI22xp33_ASAP7_75t_L     g12576(.A1(new_n1704), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1837), .Y(new_n12833));
  OAI221xp5_ASAP7_75t_L     g12577(.A1(new_n1699), .A2(new_n6812), .B1(new_n1827), .B2(new_n6837), .C(new_n12833), .Y(new_n12834));
  XNOR2x2_ASAP7_75t_L       g12578(.A(\a[23] ), .B(new_n12834), .Y(new_n12835));
  AOI21xp33_ASAP7_75t_L     g12579(.A1(new_n12758), .A2(new_n12594), .B(new_n12595), .Y(new_n12836));
  NAND2xp33_ASAP7_75t_L     g12580(.A(new_n12835), .B(new_n12836), .Y(new_n12837));
  INVx1_ASAP7_75t_L         g12581(.A(new_n12835), .Y(new_n12838));
  A2O1A1Ixp33_ASAP7_75t_L   g12582(.A1(new_n12758), .A2(new_n12594), .B(new_n12595), .C(new_n12838), .Y(new_n12839));
  AOI22xp33_ASAP7_75t_L     g12583(.A1(new_n2114), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n2259), .Y(new_n12840));
  OAI221xp5_ASAP7_75t_L     g12584(.A1(new_n2109), .A2(new_n5829), .B1(new_n2257), .B2(new_n6329), .C(new_n12840), .Y(new_n12841));
  XNOR2x2_ASAP7_75t_L       g12585(.A(\a[26] ), .B(new_n12841), .Y(new_n12842));
  A2O1A1Ixp33_ASAP7_75t_L   g12586(.A1(new_n12754), .A2(new_n12747), .B(new_n12756), .C(new_n12842), .Y(new_n12843));
  INVx1_ASAP7_75t_L         g12587(.A(new_n12843), .Y(new_n12844));
  AOI211xp5_ASAP7_75t_L     g12588(.A1(new_n12754), .A2(new_n12747), .B(new_n12842), .C(new_n12756), .Y(new_n12845));
  AOI22xp33_ASAP7_75t_L     g12589(.A1(new_n2552), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n2736), .Y(new_n12846));
  OAI221xp5_ASAP7_75t_L     g12590(.A1(new_n2547), .A2(new_n5321), .B1(new_n2734), .B2(new_n5346), .C(new_n12846), .Y(new_n12847));
  XNOR2x2_ASAP7_75t_L       g12591(.A(\a[29] ), .B(new_n12847), .Y(new_n12848));
  OAI21xp33_ASAP7_75t_L     g12592(.A1(new_n12601), .A2(new_n12743), .B(new_n12848), .Y(new_n12849));
  OR3x1_ASAP7_75t_L         g12593(.A(new_n12743), .B(new_n12601), .C(new_n12848), .Y(new_n12850));
  NAND2xp33_ASAP7_75t_L     g12594(.A(new_n12849), .B(new_n12850), .Y(new_n12851));
  AOI22xp33_ASAP7_75t_L     g12595(.A1(new_n3633), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n3858), .Y(new_n12852));
  OAI221xp5_ASAP7_75t_L     g12596(.A1(new_n3853), .A2(new_n3804), .B1(new_n3856), .B2(new_n4223), .C(new_n12852), .Y(new_n12853));
  XNOR2x2_ASAP7_75t_L       g12597(.A(\a[35] ), .B(new_n12853), .Y(new_n12854));
  INVx1_ASAP7_75t_L         g12598(.A(new_n12854), .Y(new_n12855));
  A2O1A1Ixp33_ASAP7_75t_L   g12599(.A1(new_n12700), .A2(new_n12694), .B(new_n12703), .C(new_n12716), .Y(new_n12856));
  AOI22xp33_ASAP7_75t_L     g12600(.A1(new_n4283), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n4512), .Y(new_n12857));
  OAI221xp5_ASAP7_75t_L     g12601(.A1(new_n4277), .A2(new_n3207), .B1(new_n4499), .B2(new_n3572), .C(new_n12857), .Y(new_n12858));
  XNOR2x2_ASAP7_75t_L       g12602(.A(\a[38] ), .B(new_n12858), .Y(new_n12859));
  INVx1_ASAP7_75t_L         g12603(.A(new_n12859), .Y(new_n12860));
  AOI22xp33_ASAP7_75t_L     g12604(.A1(new_n6376), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n6648), .Y(new_n12861));
  OAI221xp5_ASAP7_75t_L     g12605(.A1(new_n6646), .A2(new_n1909), .B1(new_n6636), .B2(new_n2477), .C(new_n12861), .Y(new_n12862));
  XNOR2x2_ASAP7_75t_L       g12606(.A(\a[47] ), .B(new_n12862), .Y(new_n12863));
  INVx1_ASAP7_75t_L         g12607(.A(new_n12658), .Y(new_n12864));
  O2A1O1Ixp33_ASAP7_75t_L   g12608(.A1(new_n12652), .A2(new_n12654), .B(new_n12864), .C(new_n12667), .Y(new_n12865));
  INVx1_ASAP7_75t_L         g12609(.A(new_n12865), .Y(new_n12866));
  AOI22xp33_ASAP7_75t_L     g12610(.A1(new_n8831), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n9115), .Y(new_n12867));
  OAI221xp5_ASAP7_75t_L     g12611(.A1(new_n10343), .A2(new_n869), .B1(new_n10016), .B2(new_n950), .C(new_n12867), .Y(new_n12868));
  XNOR2x2_ASAP7_75t_L       g12612(.A(\a[56] ), .B(new_n12868), .Y(new_n12869));
  INVx1_ASAP7_75t_L         g12613(.A(new_n12869), .Y(new_n12870));
  AOI22xp33_ASAP7_75t_L     g12614(.A1(new_n9700), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n10027), .Y(new_n12871));
  OAI221xp5_ASAP7_75t_L     g12615(.A1(new_n10024), .A2(new_n679), .B1(new_n9696), .B2(new_n768), .C(new_n12871), .Y(new_n12872));
  XNOR2x2_ASAP7_75t_L       g12616(.A(\a[59] ), .B(new_n12872), .Y(new_n12873));
  O2A1O1Ixp33_ASAP7_75t_L   g12617(.A1(new_n354), .A2(new_n11253), .B(new_n12619), .C(new_n262), .Y(new_n12874));
  O2A1O1Ixp33_ASAP7_75t_L   g12618(.A1(new_n12618), .A2(new_n12620), .B(new_n12614), .C(new_n12874), .Y(new_n12875));
  NOR2xp33_ASAP7_75t_L      g12619(.A(new_n354), .B(new_n11535), .Y(new_n12876));
  INVx1_ASAP7_75t_L         g12620(.A(new_n12876), .Y(new_n12877));
  XNOR2x2_ASAP7_75t_L       g12621(.A(\a[5] ), .B(\a[2] ), .Y(new_n12878));
  O2A1O1Ixp33_ASAP7_75t_L   g12622(.A1(new_n418), .A2(new_n11253), .B(new_n12877), .C(new_n12878), .Y(new_n12879));
  INVx1_ASAP7_75t_L         g12623(.A(new_n12879), .Y(new_n12880));
  O2A1O1Ixp33_ASAP7_75t_L   g12624(.A1(new_n11247), .A2(new_n11249), .B(\b[6] ), .C(new_n12876), .Y(new_n12881));
  NAND2xp33_ASAP7_75t_L     g12625(.A(new_n12878), .B(new_n12881), .Y(new_n12882));
  AND2x2_ASAP7_75t_L        g12626(.A(new_n12882), .B(new_n12880), .Y(new_n12883));
  INVx1_ASAP7_75t_L         g12627(.A(new_n12883), .Y(new_n12884));
  NAND2xp33_ASAP7_75t_L     g12628(.A(new_n12884), .B(new_n12875), .Y(new_n12885));
  INVx1_ASAP7_75t_L         g12629(.A(new_n12874), .Y(new_n12886));
  A2O1A1O1Ixp25_ASAP7_75t_L g12630(.A1(new_n12613), .A2(new_n12612), .B(new_n12621), .C(new_n12886), .D(new_n12884), .Y(new_n12887));
  INVx1_ASAP7_75t_L         g12631(.A(new_n12887), .Y(new_n12888));
  AOI22xp33_ASAP7_75t_L     g12632(.A1(\b[7] ), .A2(new_n10939), .B1(\b[9] ), .B2(new_n10938), .Y(new_n12889));
  OAI221xp5_ASAP7_75t_L     g12633(.A1(new_n10937), .A2(new_n488), .B1(new_n10629), .B2(new_n548), .C(new_n12889), .Y(new_n12890));
  XNOR2x2_ASAP7_75t_L       g12634(.A(\a[62] ), .B(new_n12890), .Y(new_n12891));
  INVx1_ASAP7_75t_L         g12635(.A(new_n12891), .Y(new_n12892));
  AOI21xp33_ASAP7_75t_L     g12636(.A1(new_n12885), .A2(new_n12888), .B(new_n12892), .Y(new_n12893));
  NAND2xp33_ASAP7_75t_L     g12637(.A(new_n12888), .B(new_n12885), .Y(new_n12894));
  NOR2xp33_ASAP7_75t_L      g12638(.A(new_n12891), .B(new_n12894), .Y(new_n12895));
  NOR2xp33_ASAP7_75t_L      g12639(.A(new_n12893), .B(new_n12895), .Y(new_n12896));
  XNOR2x2_ASAP7_75t_L       g12640(.A(new_n12873), .B(new_n12896), .Y(new_n12897));
  INVx1_ASAP7_75t_L         g12641(.A(new_n12897), .Y(new_n12898));
  O2A1O1Ixp33_ASAP7_75t_L   g12642(.A1(new_n12623), .A2(new_n12626), .B(new_n12635), .C(new_n12898), .Y(new_n12899));
  AND2x2_ASAP7_75t_L        g12643(.A(new_n12628), .B(new_n12635), .Y(new_n12900));
  AND2x2_ASAP7_75t_L        g12644(.A(new_n12900), .B(new_n12898), .Y(new_n12901));
  NOR2xp33_ASAP7_75t_L      g12645(.A(new_n12899), .B(new_n12901), .Y(new_n12902));
  XNOR2x2_ASAP7_75t_L       g12646(.A(new_n12870), .B(new_n12902), .Y(new_n12903));
  A2O1A1Ixp33_ASAP7_75t_L   g12647(.A1(new_n12635), .A2(new_n12633), .B(new_n12637), .C(new_n12645), .Y(new_n12904));
  XOR2x2_ASAP7_75t_L        g12648(.A(new_n12904), .B(new_n12903), .Y(new_n12905));
  AOI22xp33_ASAP7_75t_L     g12649(.A1(new_n7960), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n8537), .Y(new_n12906));
  OAI221xp5_ASAP7_75t_L     g12650(.A1(new_n8817), .A2(new_n1201), .B1(new_n7957), .B2(new_n1320), .C(new_n12906), .Y(new_n12907));
  XNOR2x2_ASAP7_75t_L       g12651(.A(\a[53] ), .B(new_n12907), .Y(new_n12908));
  INVx1_ASAP7_75t_L         g12652(.A(new_n12908), .Y(new_n12909));
  XNOR2x2_ASAP7_75t_L       g12653(.A(new_n12909), .B(new_n12905), .Y(new_n12910));
  A2O1A1Ixp33_ASAP7_75t_L   g12654(.A1(new_n12653), .A2(new_n12605), .B(new_n12651), .C(new_n12910), .Y(new_n12911));
  AND2x2_ASAP7_75t_L        g12655(.A(new_n12908), .B(new_n12905), .Y(new_n12912));
  NOR2xp33_ASAP7_75t_L      g12656(.A(new_n12908), .B(new_n12905), .Y(new_n12913));
  NOR2xp33_ASAP7_75t_L      g12657(.A(new_n12651), .B(new_n12652), .Y(new_n12914));
  OAI21xp33_ASAP7_75t_L     g12658(.A1(new_n12913), .A2(new_n12912), .B(new_n12914), .Y(new_n12915));
  NAND2xp33_ASAP7_75t_L     g12659(.A(new_n12915), .B(new_n12911), .Y(new_n12916));
  AOI22xp33_ASAP7_75t_L     g12660(.A1(new_n7111), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n7391), .Y(new_n12917));
  OAI221xp5_ASAP7_75t_L     g12661(.A1(new_n8558), .A2(new_n1539), .B1(new_n8237), .B2(new_n1662), .C(new_n12917), .Y(new_n12918));
  XNOR2x2_ASAP7_75t_L       g12662(.A(\a[50] ), .B(new_n12918), .Y(new_n12919));
  INVx1_ASAP7_75t_L         g12663(.A(new_n12919), .Y(new_n12920));
  XNOR2x2_ASAP7_75t_L       g12664(.A(new_n12920), .B(new_n12916), .Y(new_n12921));
  AND2x2_ASAP7_75t_L        g12665(.A(new_n12921), .B(new_n12866), .Y(new_n12922));
  NOR2xp33_ASAP7_75t_L      g12666(.A(new_n12921), .B(new_n12866), .Y(new_n12923));
  OR3x1_ASAP7_75t_L         g12667(.A(new_n12922), .B(new_n12863), .C(new_n12923), .Y(new_n12924));
  OAI21xp33_ASAP7_75t_L     g12668(.A1(new_n12923), .A2(new_n12922), .B(new_n12863), .Y(new_n12925));
  NAND2xp33_ASAP7_75t_L     g12669(.A(new_n12925), .B(new_n12924), .Y(new_n12926));
  A2O1A1Ixp33_ASAP7_75t_L   g12670(.A1(new_n12671), .A2(new_n12674), .B(new_n12670), .C(new_n12926), .Y(new_n12927));
  INVx1_ASAP7_75t_L         g12671(.A(new_n12670), .Y(new_n12928));
  NAND4xp25_ASAP7_75t_L     g12672(.A(new_n12924), .B(new_n12928), .C(new_n12675), .D(new_n12925), .Y(new_n12929));
  NAND2xp33_ASAP7_75t_L     g12673(.A(new_n12929), .B(new_n12927), .Y(new_n12930));
  AOI22xp33_ASAP7_75t_L     g12674(.A1(new_n5624), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n5901), .Y(new_n12931));
  OAI221xp5_ASAP7_75t_L     g12675(.A1(new_n5900), .A2(new_n2348), .B1(new_n5892), .B2(new_n2505), .C(new_n12931), .Y(new_n12932));
  XNOR2x2_ASAP7_75t_L       g12676(.A(\a[44] ), .B(new_n12932), .Y(new_n12933));
  XOR2x2_ASAP7_75t_L        g12677(.A(new_n12933), .B(new_n12930), .Y(new_n12934));
  AOI21xp33_ASAP7_75t_L     g12678(.A1(new_n12684), .A2(new_n12687), .B(new_n12682), .Y(new_n12935));
  XNOR2x2_ASAP7_75t_L       g12679(.A(new_n12935), .B(new_n12934), .Y(new_n12936));
  AOI22xp33_ASAP7_75t_L     g12680(.A1(new_n4920), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n5167), .Y(new_n12937));
  OAI221xp5_ASAP7_75t_L     g12681(.A1(new_n5154), .A2(new_n2688), .B1(new_n5158), .B2(new_n2990), .C(new_n12937), .Y(new_n12938));
  XNOR2x2_ASAP7_75t_L       g12682(.A(\a[41] ), .B(new_n12938), .Y(new_n12939));
  XNOR2x2_ASAP7_75t_L       g12683(.A(new_n12939), .B(new_n12936), .Y(new_n12940));
  NAND2xp33_ASAP7_75t_L     g12684(.A(new_n12696), .B(new_n12694), .Y(new_n12941));
  XNOR2x2_ASAP7_75t_L       g12685(.A(new_n12941), .B(new_n12940), .Y(new_n12942));
  NOR2xp33_ASAP7_75t_L      g12686(.A(new_n12860), .B(new_n12942), .Y(new_n12943));
  NAND2xp33_ASAP7_75t_L     g12687(.A(new_n12860), .B(new_n12942), .Y(new_n12944));
  INVx1_ASAP7_75t_L         g12688(.A(new_n12944), .Y(new_n12945));
  OAI21xp33_ASAP7_75t_L     g12689(.A1(new_n12943), .A2(new_n12945), .B(new_n12856), .Y(new_n12946));
  INVx1_ASAP7_75t_L         g12690(.A(new_n12856), .Y(new_n12947));
  INVx1_ASAP7_75t_L         g12691(.A(new_n12943), .Y(new_n12948));
  NAND3xp33_ASAP7_75t_L     g12692(.A(new_n12948), .B(new_n12944), .C(new_n12947), .Y(new_n12949));
  NAND3xp33_ASAP7_75t_L     g12693(.A(new_n12946), .B(new_n12949), .C(new_n12855), .Y(new_n12950));
  AO21x2_ASAP7_75t_L        g12694(.A1(new_n12949), .A2(new_n12946), .B(new_n12855), .Y(new_n12951));
  AOI21xp33_ASAP7_75t_L     g12695(.A1(new_n12718), .A2(new_n12722), .B(new_n12725), .Y(new_n12952));
  AO21x2_ASAP7_75t_L        g12696(.A1(new_n12950), .A2(new_n12951), .B(new_n12952), .Y(new_n12953));
  NAND3xp33_ASAP7_75t_L     g12697(.A(new_n12951), .B(new_n12950), .C(new_n12952), .Y(new_n12954));
  AOI22xp33_ASAP7_75t_L     g12698(.A1(new_n3029), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n3258), .Y(new_n12955));
  OAI221xp5_ASAP7_75t_L     g12699(.A1(new_n3024), .A2(new_n4632), .B1(new_n3256), .B2(new_n4858), .C(new_n12955), .Y(new_n12956));
  XNOR2x2_ASAP7_75t_L       g12700(.A(\a[32] ), .B(new_n12956), .Y(new_n12957));
  A2O1A1Ixp33_ASAP7_75t_L   g12701(.A1(new_n12475), .A2(new_n12474), .B(new_n12735), .C(new_n12741), .Y(new_n12958));
  NAND2xp33_ASAP7_75t_L     g12702(.A(new_n12957), .B(new_n12958), .Y(new_n12959));
  NOR2xp33_ASAP7_75t_L      g12703(.A(new_n12957), .B(new_n12958), .Y(new_n12960));
  INVx1_ASAP7_75t_L         g12704(.A(new_n12960), .Y(new_n12961));
  NAND4xp25_ASAP7_75t_L     g12705(.A(new_n12961), .B(new_n12953), .C(new_n12954), .D(new_n12959), .Y(new_n12962));
  AO22x1_ASAP7_75t_L        g12706(.A1(new_n12953), .A2(new_n12954), .B1(new_n12959), .B2(new_n12961), .Y(new_n12963));
  NAND2xp33_ASAP7_75t_L     g12707(.A(new_n12962), .B(new_n12963), .Y(new_n12964));
  XNOR2x2_ASAP7_75t_L       g12708(.A(new_n12964), .B(new_n12851), .Y(new_n12965));
  OA21x2_ASAP7_75t_L        g12709(.A1(new_n12845), .A2(new_n12844), .B(new_n12965), .Y(new_n12966));
  NOR3xp33_ASAP7_75t_L      g12710(.A(new_n12844), .B(new_n12965), .C(new_n12845), .Y(new_n12967));
  NOR2xp33_ASAP7_75t_L      g12711(.A(new_n12967), .B(new_n12966), .Y(new_n12968));
  AND3x1_ASAP7_75t_L        g12712(.A(new_n12968), .B(new_n12839), .C(new_n12837), .Y(new_n12969));
  AOI21xp33_ASAP7_75t_L     g12713(.A1(new_n12839), .A2(new_n12837), .B(new_n12968), .Y(new_n12970));
  AOI22xp33_ASAP7_75t_L     g12714(.A1(new_n1360), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1581), .Y(new_n12971));
  OAI221xp5_ASAP7_75t_L     g12715(.A1(new_n1373), .A2(new_n7593), .B1(new_n1359), .B2(new_n7623), .C(new_n12971), .Y(new_n12972));
  XNOR2x2_ASAP7_75t_L       g12716(.A(\a[20] ), .B(new_n12972), .Y(new_n12973));
  NAND3xp33_ASAP7_75t_L     g12717(.A(new_n12589), .B(new_n12759), .C(new_n12760), .Y(new_n12974));
  O2A1O1Ixp33_ASAP7_75t_L   g12718(.A1(new_n12588), .A2(new_n12586), .B(new_n12974), .C(new_n12973), .Y(new_n12975));
  INVx1_ASAP7_75t_L         g12719(.A(new_n12973), .Y(new_n12976));
  MAJIxp5_ASAP7_75t_L       g12720(.A(new_n12761), .B(new_n12586), .C(new_n12588), .Y(new_n12977));
  NOR2xp33_ASAP7_75t_L      g12721(.A(new_n12976), .B(new_n12977), .Y(new_n12978));
  OAI22xp33_ASAP7_75t_L     g12722(.A1(new_n12975), .A2(new_n12978), .B1(new_n12969), .B2(new_n12970), .Y(new_n12979));
  NOR4xp25_ASAP7_75t_L      g12723(.A(new_n12975), .B(new_n12978), .C(new_n12969), .D(new_n12970), .Y(new_n12980));
  INVx1_ASAP7_75t_L         g12724(.A(new_n12980), .Y(new_n12981));
  NAND2xp33_ASAP7_75t_L     g12725(.A(new_n12979), .B(new_n12981), .Y(new_n12982));
  AOI22xp33_ASAP7_75t_L     g12726(.A1(new_n1076), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1253), .Y(new_n12983));
  OAI221xp5_ASAP7_75t_L     g12727(.A1(new_n1154), .A2(new_n8165), .B1(new_n1156), .B2(new_n8465), .C(new_n12983), .Y(new_n12984));
  XNOR2x2_ASAP7_75t_L       g12728(.A(\a[17] ), .B(new_n12984), .Y(new_n12985));
  NOR3xp33_ASAP7_75t_L      g12729(.A(new_n12763), .B(new_n12985), .C(new_n12582), .Y(new_n12986));
  INVx1_ASAP7_75t_L         g12730(.A(new_n12986), .Y(new_n12987));
  A2O1A1Ixp33_ASAP7_75t_L   g12731(.A1(new_n12765), .A2(new_n12580), .B(new_n12582), .C(new_n12985), .Y(new_n12988));
  NAND3xp33_ASAP7_75t_L     g12732(.A(new_n12982), .B(new_n12987), .C(new_n12988), .Y(new_n12989));
  NOR2xp33_ASAP7_75t_L      g12733(.A(new_n12970), .B(new_n12969), .Y(new_n12990));
  NOR2xp33_ASAP7_75t_L      g12734(.A(new_n12978), .B(new_n12975), .Y(new_n12991));
  NOR2xp33_ASAP7_75t_L      g12735(.A(new_n12990), .B(new_n12991), .Y(new_n12992));
  NOR2xp33_ASAP7_75t_L      g12736(.A(new_n12980), .B(new_n12992), .Y(new_n12993));
  INVx1_ASAP7_75t_L         g12737(.A(new_n12988), .Y(new_n12994));
  OAI21xp33_ASAP7_75t_L     g12738(.A1(new_n12994), .A2(new_n12986), .B(new_n12993), .Y(new_n12995));
  NAND4xp25_ASAP7_75t_L     g12739(.A(new_n12832), .B(new_n12989), .C(new_n12995), .D(new_n12829), .Y(new_n12996));
  INVx1_ASAP7_75t_L         g12740(.A(new_n12826), .Y(new_n12997));
  A2O1A1Ixp33_ASAP7_75t_L   g12741(.A1(new_n12823), .A2(new_n12822), .B(new_n12767), .C(new_n12827), .Y(new_n12998));
  NOR2xp33_ASAP7_75t_L      g12742(.A(new_n12997), .B(new_n12998), .Y(new_n12999));
  NAND2xp33_ASAP7_75t_L     g12743(.A(new_n12995), .B(new_n12989), .Y(new_n13000));
  OAI21xp33_ASAP7_75t_L     g12744(.A1(new_n12828), .A2(new_n12999), .B(new_n13000), .Y(new_n13001));
  AND2x2_ASAP7_75t_L        g12745(.A(new_n12996), .B(new_n13001), .Y(new_n13002));
  XNOR2x2_ASAP7_75t_L       g12746(.A(new_n13002), .B(new_n12819), .Y(new_n13003));
  XOR2x2_ASAP7_75t_L        g12747(.A(new_n12813), .B(new_n13003), .Y(new_n13004));
  O2A1O1Ixp33_ASAP7_75t_L   g12748(.A1(new_n12786), .A2(new_n12787), .B(new_n12783), .C(new_n13004), .Y(new_n13005));
  A2O1A1Ixp33_ASAP7_75t_L   g12749(.A1(new_n12530), .A2(new_n12527), .B(new_n12781), .C(new_n12785), .Y(new_n13006));
  XNOR2x2_ASAP7_75t_L       g12750(.A(new_n12813), .B(new_n13003), .Y(new_n13007));
  NOR2xp33_ASAP7_75t_L      g12751(.A(new_n13006), .B(new_n13007), .Y(new_n13008));
  NOR2xp33_ASAP7_75t_L      g12752(.A(new_n13008), .B(new_n13005), .Y(new_n13009));
  A2O1A1Ixp33_ASAP7_75t_L   g12753(.A1(new_n12795), .A2(new_n12790), .B(new_n12800), .C(new_n13009), .Y(new_n13010));
  INVx1_ASAP7_75t_L         g12754(.A(new_n13010), .Y(new_n13011));
  NOR3xp33_ASAP7_75t_L      g12755(.A(new_n12798), .B(new_n12545), .C(new_n12533), .Y(new_n13012));
  A2O1A1Ixp33_ASAP7_75t_L   g12756(.A1(new_n12539), .A2(new_n12794), .B(new_n13012), .C(new_n12799), .Y(new_n13013));
  NOR2xp33_ASAP7_75t_L      g12757(.A(new_n13009), .B(new_n13013), .Y(new_n13014));
  NOR2xp33_ASAP7_75t_L      g12758(.A(new_n13014), .B(new_n13011), .Y(\f[69] ));
  AOI22xp33_ASAP7_75t_L     g12759(.A1(new_n471), .A2(\b[62] ), .B1(new_n441), .B2(new_n12322), .Y(new_n13016));
  OA211x2_ASAP7_75t_L       g12760(.A1(new_n468), .A2(new_n11468), .B(new_n13016), .C(\a[8] ), .Y(new_n13017));
  O2A1O1Ixp33_ASAP7_75t_L   g12761(.A1(new_n11468), .A2(new_n468), .B(new_n13016), .C(\a[8] ), .Y(new_n13018));
  NOR2xp33_ASAP7_75t_L      g12762(.A(new_n13018), .B(new_n13017), .Y(new_n13019));
  MAJIxp5_ASAP7_75t_L       g12763(.A(new_n13002), .B(new_n12817), .C(new_n12818), .Y(new_n13020));
  XNOR2x2_ASAP7_75t_L       g12764(.A(new_n13019), .B(new_n13020), .Y(new_n13021));
  AOI22xp33_ASAP7_75t_L     g12765(.A1(\b[59] ), .A2(new_n651), .B1(\b[61] ), .B2(new_n581), .Y(new_n13022));
  OAI221xp5_ASAP7_75t_L     g12766(.A1(new_n821), .A2(new_n10250), .B1(new_n577), .B2(new_n10855), .C(new_n13022), .Y(new_n13023));
  XNOR2x2_ASAP7_75t_L       g12767(.A(\a[11] ), .B(new_n13023), .Y(new_n13024));
  AND3x1_ASAP7_75t_L        g12768(.A(new_n12996), .B(new_n13024), .C(new_n12829), .Y(new_n13025));
  O2A1O1Ixp33_ASAP7_75t_L   g12769(.A1(new_n12999), .A2(new_n13000), .B(new_n12829), .C(new_n13024), .Y(new_n13026));
  NOR2xp33_ASAP7_75t_L      g12770(.A(new_n13026), .B(new_n13025), .Y(new_n13027));
  AOI22xp33_ASAP7_75t_L     g12771(.A1(new_n811), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n900), .Y(new_n13028));
  OAI221xp5_ASAP7_75t_L     g12772(.A1(new_n904), .A2(new_n9620), .B1(new_n898), .B2(new_n9925), .C(new_n13028), .Y(new_n13029));
  XNOR2x2_ASAP7_75t_L       g12773(.A(\a[14] ), .B(new_n13029), .Y(new_n13030));
  A2O1A1O1Ixp25_ASAP7_75t_L g12774(.A1(new_n12981), .A2(new_n12979), .B(new_n12994), .C(new_n12987), .D(new_n13030), .Y(new_n13031));
  INVx1_ASAP7_75t_L         g12775(.A(new_n13031), .Y(new_n13032));
  O2A1O1Ixp33_ASAP7_75t_L   g12776(.A1(new_n12980), .A2(new_n12992), .B(new_n12988), .C(new_n12986), .Y(new_n13033));
  NAND2xp33_ASAP7_75t_L     g12777(.A(new_n13030), .B(new_n13033), .Y(new_n13034));
  AND2x2_ASAP7_75t_L        g12778(.A(new_n13034), .B(new_n13032), .Y(new_n13035));
  AOI22xp33_ASAP7_75t_L     g12779(.A1(new_n1076), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1253), .Y(new_n13036));
  OAI221xp5_ASAP7_75t_L     g12780(.A1(new_n1154), .A2(new_n8458), .B1(new_n1156), .B2(new_n8768), .C(new_n13036), .Y(new_n13037));
  XNOR2x2_ASAP7_75t_L       g12781(.A(\a[17] ), .B(new_n13037), .Y(new_n13038));
  A2O1A1Ixp33_ASAP7_75t_L   g12782(.A1(new_n12991), .A2(new_n12990), .B(new_n12978), .C(new_n13038), .Y(new_n13039));
  INVx1_ASAP7_75t_L         g12783(.A(new_n13039), .Y(new_n13040));
  NOR3xp33_ASAP7_75t_L      g12784(.A(new_n12980), .B(new_n13038), .C(new_n12978), .Y(new_n13041));
  AOI22xp33_ASAP7_75t_L     g12785(.A1(new_n1360), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1581), .Y(new_n13042));
  OAI221xp5_ASAP7_75t_L     g12786(.A1(new_n1373), .A2(new_n7616), .B1(new_n1359), .B2(new_n7906), .C(new_n13042), .Y(new_n13043));
  XNOR2x2_ASAP7_75t_L       g12787(.A(new_n1356), .B(new_n13043), .Y(new_n13044));
  MAJIxp5_ASAP7_75t_L       g12788(.A(new_n12968), .B(new_n12835), .C(new_n12836), .Y(new_n13045));
  XNOR2x2_ASAP7_75t_L       g12789(.A(new_n13044), .B(new_n13045), .Y(new_n13046));
  AOI22xp33_ASAP7_75t_L     g12790(.A1(new_n1704), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1837), .Y(new_n13047));
  OAI221xp5_ASAP7_75t_L     g12791(.A1(new_n1699), .A2(new_n6830), .B1(new_n1827), .B2(new_n7323), .C(new_n13047), .Y(new_n13048));
  XNOR2x2_ASAP7_75t_L       g12792(.A(\a[23] ), .B(new_n13048), .Y(new_n13049));
  INVx1_ASAP7_75t_L         g12793(.A(new_n12845), .Y(new_n13050));
  INVx1_ASAP7_75t_L         g12794(.A(new_n12842), .Y(new_n13051));
  A2O1A1Ixp33_ASAP7_75t_L   g12795(.A1(new_n12754), .A2(new_n12747), .B(new_n12756), .C(new_n13051), .Y(new_n13052));
  A2O1A1Ixp33_ASAP7_75t_L   g12796(.A1(new_n13050), .A2(new_n12843), .B(new_n12965), .C(new_n13052), .Y(new_n13053));
  XNOR2x2_ASAP7_75t_L       g12797(.A(new_n13049), .B(new_n13053), .Y(new_n13054));
  AOI22xp33_ASAP7_75t_L     g12798(.A1(new_n2114), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n2259), .Y(new_n13055));
  OAI221xp5_ASAP7_75t_L     g12799(.A1(new_n2109), .A2(new_n6321), .B1(new_n2257), .B2(new_n6573), .C(new_n13055), .Y(new_n13056));
  XNOR2x2_ASAP7_75t_L       g12800(.A(\a[26] ), .B(new_n13056), .Y(new_n13057));
  O2A1O1Ixp33_ASAP7_75t_L   g12801(.A1(new_n12964), .A2(new_n12851), .B(new_n12850), .C(new_n13057), .Y(new_n13058));
  INVx1_ASAP7_75t_L         g12802(.A(new_n13058), .Y(new_n13059));
  OAI211xp5_ASAP7_75t_L     g12803(.A1(new_n12964), .A2(new_n12851), .B(new_n12850), .C(new_n13057), .Y(new_n13060));
  AOI22xp33_ASAP7_75t_L     g12804(.A1(new_n2552), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n2736), .Y(new_n13061));
  OAI221xp5_ASAP7_75t_L     g12805(.A1(new_n2547), .A2(new_n5338), .B1(new_n2734), .B2(new_n6338), .C(new_n13061), .Y(new_n13062));
  XNOR2x2_ASAP7_75t_L       g12806(.A(\a[29] ), .B(new_n13062), .Y(new_n13063));
  INVx1_ASAP7_75t_L         g12807(.A(new_n13063), .Y(new_n13064));
  AND3x1_ASAP7_75t_L        g12808(.A(new_n12962), .B(new_n13064), .C(new_n12961), .Y(new_n13065));
  O2A1O1Ixp33_ASAP7_75t_L   g12809(.A1(new_n12957), .A2(new_n12958), .B(new_n12962), .C(new_n13064), .Y(new_n13066));
  NOR2xp33_ASAP7_75t_L      g12810(.A(new_n13066), .B(new_n13065), .Y(new_n13067));
  AOI22xp33_ASAP7_75t_L     g12811(.A1(new_n3029), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n3258), .Y(new_n13068));
  OAI221xp5_ASAP7_75t_L     g12812(.A1(new_n3024), .A2(new_n4848), .B1(new_n3256), .B2(new_n11686), .C(new_n13068), .Y(new_n13069));
  XNOR2x2_ASAP7_75t_L       g12813(.A(\a[32] ), .B(new_n13069), .Y(new_n13070));
  AND3x1_ASAP7_75t_L        g12814(.A(new_n12946), .B(new_n12949), .C(new_n12855), .Y(new_n13071));
  AOI21xp33_ASAP7_75t_L     g12815(.A1(new_n12951), .A2(new_n12952), .B(new_n13071), .Y(new_n13072));
  NAND2xp33_ASAP7_75t_L     g12816(.A(new_n13070), .B(new_n13072), .Y(new_n13073));
  INVx1_ASAP7_75t_L         g12817(.A(new_n13070), .Y(new_n13074));
  A2O1A1Ixp33_ASAP7_75t_L   g12818(.A1(new_n12951), .A2(new_n12952), .B(new_n13071), .C(new_n13074), .Y(new_n13075));
  NAND2xp33_ASAP7_75t_L     g12819(.A(new_n13075), .B(new_n13073), .Y(new_n13076));
  NAND2xp33_ASAP7_75t_L     g12820(.A(\b[35] ), .B(new_n3858), .Y(new_n13077));
  OAI221xp5_ASAP7_75t_L     g12821(.A1(new_n4061), .A2(new_n4424), .B1(new_n3856), .B2(new_n4431), .C(new_n13077), .Y(new_n13078));
  AOI21xp33_ASAP7_75t_L     g12822(.A1(new_n3639), .A2(\b[36] ), .B(new_n13078), .Y(new_n13079));
  NAND2xp33_ASAP7_75t_L     g12823(.A(\a[35] ), .B(new_n13079), .Y(new_n13080));
  A2O1A1Ixp33_ASAP7_75t_L   g12824(.A1(\b[36] ), .A2(new_n3639), .B(new_n13078), .C(new_n3628), .Y(new_n13081));
  NAND2xp33_ASAP7_75t_L     g12825(.A(new_n13081), .B(new_n13080), .Y(new_n13082));
  INVx1_ASAP7_75t_L         g12826(.A(new_n13082), .Y(new_n13083));
  INVx1_ASAP7_75t_L         g12827(.A(new_n12942), .Y(new_n13084));
  NAND2xp33_ASAP7_75t_L     g12828(.A(new_n12860), .B(new_n13084), .Y(new_n13085));
  A2O1A1Ixp33_ASAP7_75t_L   g12829(.A1(new_n12948), .A2(new_n12944), .B(new_n12947), .C(new_n13085), .Y(new_n13086));
  AOI22xp33_ASAP7_75t_L     g12830(.A1(new_n4283), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n4512), .Y(new_n13087));
  OAI221xp5_ASAP7_75t_L     g12831(.A1(new_n4277), .A2(new_n3565), .B1(new_n4499), .B2(new_n3591), .C(new_n13087), .Y(new_n13088));
  XNOR2x2_ASAP7_75t_L       g12832(.A(\a[38] ), .B(new_n13088), .Y(new_n13089));
  NAND2xp33_ASAP7_75t_L     g12833(.A(new_n12935), .B(new_n12934), .Y(new_n13090));
  NOR2xp33_ASAP7_75t_L      g12834(.A(new_n418), .B(new_n11535), .Y(new_n13091));
  O2A1O1Ixp33_ASAP7_75t_L   g12835(.A1(new_n11247), .A2(new_n11249), .B(\b[7] ), .C(new_n13091), .Y(new_n13092));
  INVx1_ASAP7_75t_L         g12836(.A(new_n13092), .Y(new_n13093));
  O2A1O1Ixp33_ASAP7_75t_L   g12837(.A1(\a[2] ), .A2(\a[5] ), .B(new_n12880), .C(new_n13093), .Y(new_n13094));
  INVx1_ASAP7_75t_L         g12838(.A(new_n13094), .Y(new_n13095));
  AOI21xp33_ASAP7_75t_L     g12839(.A1(new_n338), .A2(new_n262), .B(new_n12879), .Y(new_n13096));
  A2O1A1Ixp33_ASAP7_75t_L   g12840(.A1(\b[7] ), .A2(new_n11533), .B(new_n13091), .C(new_n13096), .Y(new_n13097));
  NAND2xp33_ASAP7_75t_L     g12841(.A(new_n13097), .B(new_n13095), .Y(new_n13098));
  NAND2xp33_ASAP7_75t_L     g12842(.A(\b[9] ), .B(new_n10632), .Y(new_n13099));
  OAI221xp5_ASAP7_75t_L     g12843(.A1(new_n10630), .A2(new_n617), .B1(new_n488), .B2(new_n11257), .C(new_n13099), .Y(new_n13100));
  AOI21xp33_ASAP7_75t_L     g12844(.A1(new_n2143), .A2(new_n11256), .B(new_n13100), .Y(new_n13101));
  NAND2xp33_ASAP7_75t_L     g12845(.A(\a[62] ), .B(new_n13101), .Y(new_n13102));
  A2O1A1Ixp33_ASAP7_75t_L   g12846(.A1(new_n2143), .A2(new_n11256), .B(new_n13100), .C(new_n10622), .Y(new_n13103));
  AO21x2_ASAP7_75t_L        g12847(.A1(new_n13103), .A2(new_n13102), .B(new_n13098), .Y(new_n13104));
  NAND3xp33_ASAP7_75t_L     g12848(.A(new_n13102), .B(new_n13098), .C(new_n13103), .Y(new_n13105));
  AND2x2_ASAP7_75t_L        g12849(.A(new_n13105), .B(new_n13104), .Y(new_n13106));
  INVx1_ASAP7_75t_L         g12850(.A(new_n13106), .Y(new_n13107));
  O2A1O1Ixp33_ASAP7_75t_L   g12851(.A1(new_n12891), .A2(new_n12894), .B(new_n12888), .C(new_n13107), .Y(new_n13108));
  INVx1_ASAP7_75t_L         g12852(.A(new_n13108), .Y(new_n13109));
  A2O1A1O1Ixp25_ASAP7_75t_L g12853(.A1(new_n12622), .A2(new_n12614), .B(new_n12874), .C(new_n12883), .D(new_n12895), .Y(new_n13110));
  NAND2xp33_ASAP7_75t_L     g12854(.A(new_n13107), .B(new_n13110), .Y(new_n13111));
  AOI22xp33_ASAP7_75t_L     g12855(.A1(new_n9700), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n10027), .Y(new_n13112));
  OAI221xp5_ASAP7_75t_L     g12856(.A1(new_n10024), .A2(new_n760), .B1(new_n9696), .B2(new_n790), .C(new_n13112), .Y(new_n13113));
  XNOR2x2_ASAP7_75t_L       g12857(.A(\a[59] ), .B(new_n13113), .Y(new_n13114));
  NAND3xp33_ASAP7_75t_L     g12858(.A(new_n13111), .B(new_n13109), .C(new_n13114), .Y(new_n13115));
  AO21x2_ASAP7_75t_L        g12859(.A1(new_n13109), .A2(new_n13111), .B(new_n13114), .Y(new_n13116));
  NAND2xp33_ASAP7_75t_L     g12860(.A(new_n13115), .B(new_n13116), .Y(new_n13117));
  INVx1_ASAP7_75t_L         g12861(.A(new_n13117), .Y(new_n13118));
  INVx1_ASAP7_75t_L         g12862(.A(new_n12873), .Y(new_n13119));
  NAND2xp33_ASAP7_75t_L     g12863(.A(new_n13119), .B(new_n12896), .Y(new_n13120));
  OAI211xp5_ASAP7_75t_L     g12864(.A1(new_n12898), .A2(new_n12900), .B(new_n13118), .C(new_n13120), .Y(new_n13121));
  INVx1_ASAP7_75t_L         g12865(.A(new_n13121), .Y(new_n13122));
  O2A1O1Ixp33_ASAP7_75t_L   g12866(.A1(new_n12898), .A2(new_n12900), .B(new_n13120), .C(new_n13118), .Y(new_n13123));
  NOR2xp33_ASAP7_75t_L      g12867(.A(new_n13123), .B(new_n13122), .Y(new_n13124));
  AOI22xp33_ASAP7_75t_L     g12868(.A1(new_n8831), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n9115), .Y(new_n13125));
  OAI221xp5_ASAP7_75t_L     g12869(.A1(new_n10343), .A2(new_n942), .B1(new_n10016), .B2(new_n1035), .C(new_n13125), .Y(new_n13126));
  XNOR2x2_ASAP7_75t_L       g12870(.A(\a[56] ), .B(new_n13126), .Y(new_n13127));
  NAND2xp33_ASAP7_75t_L     g12871(.A(new_n13127), .B(new_n13124), .Y(new_n13128));
  A2O1A1Ixp33_ASAP7_75t_L   g12872(.A1(new_n12896), .A2(new_n13119), .B(new_n12899), .C(new_n13117), .Y(new_n13129));
  AO21x2_ASAP7_75t_L        g12873(.A1(new_n13129), .A2(new_n13121), .B(new_n13127), .Y(new_n13130));
  NAND2xp33_ASAP7_75t_L     g12874(.A(new_n13130), .B(new_n13128), .Y(new_n13131));
  INVx1_ASAP7_75t_L         g12875(.A(new_n13131), .Y(new_n13132));
  NOR2xp33_ASAP7_75t_L      g12876(.A(new_n12904), .B(new_n12903), .Y(new_n13133));
  AOI21xp33_ASAP7_75t_L     g12877(.A1(new_n12902), .A2(new_n12870), .B(new_n13133), .Y(new_n13134));
  NAND2xp33_ASAP7_75t_L     g12878(.A(new_n13134), .B(new_n13132), .Y(new_n13135));
  A2O1A1Ixp33_ASAP7_75t_L   g12879(.A1(new_n12902), .A2(new_n12870), .B(new_n13133), .C(new_n13131), .Y(new_n13136));
  AOI22xp33_ASAP7_75t_L     g12880(.A1(new_n7960), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n8537), .Y(new_n13137));
  OAI221xp5_ASAP7_75t_L     g12881(.A1(new_n8817), .A2(new_n1313), .B1(new_n7957), .B2(new_n1438), .C(new_n13137), .Y(new_n13138));
  XNOR2x2_ASAP7_75t_L       g12882(.A(\a[53] ), .B(new_n13138), .Y(new_n13139));
  AND3x1_ASAP7_75t_L        g12883(.A(new_n13135), .B(new_n13139), .C(new_n13136), .Y(new_n13140));
  AOI21xp33_ASAP7_75t_L     g12884(.A1(new_n13136), .A2(new_n13135), .B(new_n13139), .Y(new_n13141));
  NOR2xp33_ASAP7_75t_L      g12885(.A(new_n13141), .B(new_n13140), .Y(new_n13142));
  NAND2xp33_ASAP7_75t_L     g12886(.A(new_n12909), .B(new_n12905), .Y(new_n13143));
  NAND2xp33_ASAP7_75t_L     g12887(.A(new_n13143), .B(new_n12915), .Y(new_n13144));
  XNOR2x2_ASAP7_75t_L       g12888(.A(new_n13144), .B(new_n13142), .Y(new_n13145));
  AOI22xp33_ASAP7_75t_L     g12889(.A1(new_n7111), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n7391), .Y(new_n13146));
  OAI221xp5_ASAP7_75t_L     g12890(.A1(new_n8558), .A2(new_n1655), .B1(new_n8237), .B2(new_n1780), .C(new_n13146), .Y(new_n13147));
  XNOR2x2_ASAP7_75t_L       g12891(.A(\a[50] ), .B(new_n13147), .Y(new_n13148));
  XOR2x2_ASAP7_75t_L        g12892(.A(new_n13148), .B(new_n13145), .Y(new_n13149));
  AOI31xp33_ASAP7_75t_L     g12893(.A1(new_n12915), .A2(new_n12911), .A3(new_n12920), .B(new_n12922), .Y(new_n13150));
  XOR2x2_ASAP7_75t_L        g12894(.A(new_n13149), .B(new_n13150), .Y(new_n13151));
  AOI22xp33_ASAP7_75t_L     g12895(.A1(new_n6376), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n6648), .Y(new_n13152));
  OAI221xp5_ASAP7_75t_L     g12896(.A1(new_n6646), .A2(new_n1929), .B1(new_n6636), .B2(new_n2075), .C(new_n13152), .Y(new_n13153));
  XNOR2x2_ASAP7_75t_L       g12897(.A(\a[47] ), .B(new_n13153), .Y(new_n13154));
  XNOR2x2_ASAP7_75t_L       g12898(.A(new_n13154), .B(new_n13151), .Y(new_n13155));
  NAND2xp33_ASAP7_75t_L     g12899(.A(new_n12924), .B(new_n12929), .Y(new_n13156));
  XNOR2x2_ASAP7_75t_L       g12900(.A(new_n13156), .B(new_n13155), .Y(new_n13157));
  AOI22xp33_ASAP7_75t_L     g12901(.A1(new_n5624), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n5901), .Y(new_n13158));
  OAI221xp5_ASAP7_75t_L     g12902(.A1(new_n5900), .A2(new_n2497), .B1(new_n5892), .B2(new_n2672), .C(new_n13158), .Y(new_n13159));
  XNOR2x2_ASAP7_75t_L       g12903(.A(\a[44] ), .B(new_n13159), .Y(new_n13160));
  XNOR2x2_ASAP7_75t_L       g12904(.A(new_n13160), .B(new_n13157), .Y(new_n13161));
  OAI211xp5_ASAP7_75t_L     g12905(.A1(new_n12930), .A2(new_n12933), .B(new_n13161), .C(new_n13090), .Y(new_n13162));
  INVx1_ASAP7_75t_L         g12906(.A(new_n13160), .Y(new_n13163));
  XNOR2x2_ASAP7_75t_L       g12907(.A(new_n13163), .B(new_n13157), .Y(new_n13164));
  OAI21xp33_ASAP7_75t_L     g12908(.A1(new_n12930), .A2(new_n12933), .B(new_n13090), .Y(new_n13165));
  NAND2xp33_ASAP7_75t_L     g12909(.A(new_n13165), .B(new_n13164), .Y(new_n13166));
  AOI22xp33_ASAP7_75t_L     g12910(.A1(new_n4920), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n5167), .Y(new_n13167));
  OAI221xp5_ASAP7_75t_L     g12911(.A1(new_n5154), .A2(new_n2982), .B1(new_n5158), .B2(new_n3187), .C(new_n13167), .Y(new_n13168));
  XNOR2x2_ASAP7_75t_L       g12912(.A(\a[41] ), .B(new_n13168), .Y(new_n13169));
  INVx1_ASAP7_75t_L         g12913(.A(new_n13169), .Y(new_n13170));
  AO21x2_ASAP7_75t_L        g12914(.A1(new_n13166), .A2(new_n13162), .B(new_n13170), .Y(new_n13171));
  NAND3xp33_ASAP7_75t_L     g12915(.A(new_n13162), .B(new_n13166), .C(new_n13170), .Y(new_n13172));
  NAND2xp33_ASAP7_75t_L     g12916(.A(new_n13172), .B(new_n13171), .Y(new_n13173));
  MAJx2_ASAP7_75t_L         g12917(.A(new_n12941), .B(new_n12939), .C(new_n12936), .Y(new_n13174));
  XNOR2x2_ASAP7_75t_L       g12918(.A(new_n13174), .B(new_n13173), .Y(new_n13175));
  NOR2xp33_ASAP7_75t_L      g12919(.A(new_n13089), .B(new_n13175), .Y(new_n13176));
  INVx1_ASAP7_75t_L         g12920(.A(new_n13089), .Y(new_n13177));
  INVx1_ASAP7_75t_L         g12921(.A(new_n13175), .Y(new_n13178));
  NOR2xp33_ASAP7_75t_L      g12922(.A(new_n13177), .B(new_n13178), .Y(new_n13179));
  NOR2xp33_ASAP7_75t_L      g12923(.A(new_n13176), .B(new_n13179), .Y(new_n13180));
  NAND2xp33_ASAP7_75t_L     g12924(.A(new_n13086), .B(new_n13180), .Y(new_n13181));
  OAI211xp5_ASAP7_75t_L     g12925(.A1(new_n13176), .A2(new_n13179), .B(new_n13085), .C(new_n12946), .Y(new_n13182));
  AO21x2_ASAP7_75t_L        g12926(.A1(new_n13182), .A2(new_n13181), .B(new_n13083), .Y(new_n13183));
  NAND3xp33_ASAP7_75t_L     g12927(.A(new_n13181), .B(new_n13083), .C(new_n13182), .Y(new_n13184));
  NAND2xp33_ASAP7_75t_L     g12928(.A(new_n13184), .B(new_n13183), .Y(new_n13185));
  XNOR2x2_ASAP7_75t_L       g12929(.A(new_n13076), .B(new_n13185), .Y(new_n13186));
  XNOR2x2_ASAP7_75t_L       g12930(.A(new_n13067), .B(new_n13186), .Y(new_n13187));
  NAND3xp33_ASAP7_75t_L     g12931(.A(new_n13187), .B(new_n13060), .C(new_n13059), .Y(new_n13188));
  AO21x2_ASAP7_75t_L        g12932(.A1(new_n13059), .A2(new_n13060), .B(new_n13187), .Y(new_n13189));
  NAND2xp33_ASAP7_75t_L     g12933(.A(new_n13188), .B(new_n13189), .Y(new_n13190));
  XNOR2x2_ASAP7_75t_L       g12934(.A(new_n13054), .B(new_n13190), .Y(new_n13191));
  NOR2xp33_ASAP7_75t_L      g12935(.A(new_n13191), .B(new_n13046), .Y(new_n13192));
  AND2x2_ASAP7_75t_L        g12936(.A(new_n13191), .B(new_n13046), .Y(new_n13193));
  NOR2xp33_ASAP7_75t_L      g12937(.A(new_n13192), .B(new_n13193), .Y(new_n13194));
  NOR3xp33_ASAP7_75t_L      g12938(.A(new_n13194), .B(new_n13041), .C(new_n13040), .Y(new_n13195));
  INVx1_ASAP7_75t_L         g12939(.A(new_n13041), .Y(new_n13196));
  XNOR2x2_ASAP7_75t_L       g12940(.A(new_n13191), .B(new_n13046), .Y(new_n13197));
  AOI21xp33_ASAP7_75t_L     g12941(.A1(new_n13196), .A2(new_n13039), .B(new_n13197), .Y(new_n13198));
  NOR2xp33_ASAP7_75t_L      g12942(.A(new_n13198), .B(new_n13195), .Y(new_n13199));
  XOR2x2_ASAP7_75t_L        g12943(.A(new_n13199), .B(new_n13035), .Y(new_n13200));
  NAND2xp33_ASAP7_75t_L     g12944(.A(new_n13027), .B(new_n13200), .Y(new_n13201));
  OR2x4_ASAP7_75t_L         g12945(.A(new_n13027), .B(new_n13200), .Y(new_n13202));
  AO21x2_ASAP7_75t_L        g12946(.A1(new_n13202), .A2(new_n13201), .B(new_n13021), .Y(new_n13203));
  NAND3xp33_ASAP7_75t_L     g12947(.A(new_n13021), .B(new_n13202), .C(new_n13201), .Y(new_n13204));
  AND2x2_ASAP7_75t_L        g12948(.A(new_n12808), .B(new_n12807), .Y(new_n13205));
  A2O1A1O1Ixp25_ASAP7_75t_L g12949(.A1(new_n12557), .A2(new_n12773), .B(new_n12774), .C(new_n12803), .D(new_n13205), .Y(new_n13206));
  O2A1O1Ixp33_ASAP7_75t_L   g12950(.A1(new_n12810), .A2(new_n12812), .B(new_n13003), .C(new_n13206), .Y(new_n13207));
  AOI21xp33_ASAP7_75t_L     g12951(.A1(new_n13203), .A2(new_n13204), .B(new_n13207), .Y(new_n13208));
  AND3x1_ASAP7_75t_L        g12952(.A(new_n13203), .B(new_n13207), .C(new_n13204), .Y(new_n13209));
  NOR2xp33_ASAP7_75t_L      g12953(.A(new_n13208), .B(new_n13209), .Y(new_n13210));
  A2O1A1Ixp33_ASAP7_75t_L   g12954(.A1(new_n13013), .A2(new_n13009), .B(new_n13005), .C(new_n13210), .Y(new_n13211));
  INVx1_ASAP7_75t_L         g12955(.A(new_n13211), .Y(new_n13212));
  INVx1_ASAP7_75t_L         g12956(.A(new_n13005), .Y(new_n13213));
  A2O1A1Ixp33_ASAP7_75t_L   g12957(.A1(new_n12791), .A2(new_n12799), .B(new_n13008), .C(new_n13213), .Y(new_n13214));
  NOR2xp33_ASAP7_75t_L      g12958(.A(new_n13210), .B(new_n13214), .Y(new_n13215));
  NOR2xp33_ASAP7_75t_L      g12959(.A(new_n13215), .B(new_n13212), .Y(\f[70] ));
  NAND2xp33_ASAP7_75t_L     g12960(.A(new_n13199), .B(new_n13035), .Y(new_n13217));
  A2O1A1Ixp33_ASAP7_75t_L   g12961(.A1(new_n12989), .A2(new_n12987), .B(new_n13030), .C(new_n13217), .Y(new_n13218));
  NAND2xp33_ASAP7_75t_L     g12962(.A(\b[61] ), .B(new_n584), .Y(new_n13219));
  OAI221xp5_ASAP7_75t_L     g12963(.A1(new_n580), .A2(new_n11172), .B1(new_n10250), .B2(new_n706), .C(new_n13219), .Y(new_n13220));
  AOI21xp33_ASAP7_75t_L     g12964(.A1(new_n11180), .A2(new_n578), .B(new_n13220), .Y(new_n13221));
  NAND2xp33_ASAP7_75t_L     g12965(.A(\a[11] ), .B(new_n13221), .Y(new_n13222));
  A2O1A1Ixp33_ASAP7_75t_L   g12966(.A1(new_n11180), .A2(new_n578), .B(new_n13220), .C(new_n574), .Y(new_n13223));
  NAND2xp33_ASAP7_75t_L     g12967(.A(new_n13223), .B(new_n13222), .Y(new_n13224));
  XOR2x2_ASAP7_75t_L        g12968(.A(new_n13224), .B(new_n13218), .Y(new_n13225));
  NOR2xp33_ASAP7_75t_L      g12969(.A(new_n13044), .B(new_n13045), .Y(new_n13226));
  AOI22xp33_ASAP7_75t_L     g12970(.A1(new_n1076), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1253), .Y(new_n13227));
  OAI221xp5_ASAP7_75t_L     g12971(.A1(new_n1154), .A2(new_n8762), .B1(new_n1156), .B2(new_n9331), .C(new_n13227), .Y(new_n13228));
  XNOR2x2_ASAP7_75t_L       g12972(.A(\a[17] ), .B(new_n13228), .Y(new_n13229));
  OAI21xp33_ASAP7_75t_L     g12973(.A1(new_n13226), .A2(new_n13192), .B(new_n13229), .Y(new_n13230));
  OR3x1_ASAP7_75t_L         g12974(.A(new_n13192), .B(new_n13226), .C(new_n13229), .Y(new_n13231));
  NAND2xp33_ASAP7_75t_L     g12975(.A(new_n13230), .B(new_n13231), .Y(new_n13232));
  AOI22xp33_ASAP7_75t_L     g12976(.A1(new_n1704), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1837), .Y(new_n13233));
  OAI221xp5_ASAP7_75t_L     g12977(.A1(new_n1699), .A2(new_n7317), .B1(new_n1827), .B2(new_n7602), .C(new_n13233), .Y(new_n13234));
  XNOR2x2_ASAP7_75t_L       g12978(.A(\a[23] ), .B(new_n13234), .Y(new_n13235));
  AND3x1_ASAP7_75t_L        g12979(.A(new_n13188), .B(new_n13235), .C(new_n13059), .Y(new_n13236));
  AOI21xp33_ASAP7_75t_L     g12980(.A1(new_n13187), .A2(new_n13060), .B(new_n13058), .Y(new_n13237));
  NOR2xp33_ASAP7_75t_L      g12981(.A(new_n13235), .B(new_n13237), .Y(new_n13238));
  AOI22xp33_ASAP7_75t_L     g12982(.A1(new_n2114), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n2259), .Y(new_n13239));
  OAI221xp5_ASAP7_75t_L     g12983(.A1(new_n2109), .A2(new_n6568), .B1(new_n2257), .B2(new_n6820), .C(new_n13239), .Y(new_n13240));
  XNOR2x2_ASAP7_75t_L       g12984(.A(\a[26] ), .B(new_n13240), .Y(new_n13241));
  O2A1O1Ixp33_ASAP7_75t_L   g12985(.A1(new_n12957), .A2(new_n12958), .B(new_n12962), .C(new_n13063), .Y(new_n13242));
  O2A1O1Ixp33_ASAP7_75t_L   g12986(.A1(new_n13065), .A2(new_n13066), .B(new_n13186), .C(new_n13242), .Y(new_n13243));
  XNOR2x2_ASAP7_75t_L       g12987(.A(new_n13241), .B(new_n13243), .Y(new_n13244));
  NOR2xp33_ASAP7_75t_L      g12988(.A(new_n13070), .B(new_n13072), .Y(new_n13245));
  NOR2xp33_ASAP7_75t_L      g12989(.A(new_n5829), .B(new_n2545), .Y(new_n13246));
  AOI221xp5_ASAP7_75t_L     g12990(.A1(\b[42] ), .A2(new_n2736), .B1(\b[43] ), .B2(new_n2553), .C(new_n13246), .Y(new_n13247));
  OA211x2_ASAP7_75t_L       g12991(.A1(new_n2734), .A2(new_n5835), .B(new_n13247), .C(\a[29] ), .Y(new_n13248));
  O2A1O1Ixp33_ASAP7_75t_L   g12992(.A1(new_n2734), .A2(new_n5835), .B(new_n13247), .C(\a[29] ), .Y(new_n13249));
  NOR2xp33_ASAP7_75t_L      g12993(.A(new_n13249), .B(new_n13248), .Y(new_n13250));
  A2O1A1Ixp33_ASAP7_75t_L   g12994(.A1(new_n13185), .A2(new_n13073), .B(new_n13245), .C(new_n13250), .Y(new_n13251));
  AOI21xp33_ASAP7_75t_L     g12995(.A1(new_n13185), .A2(new_n13073), .B(new_n13245), .Y(new_n13252));
  OAI21xp33_ASAP7_75t_L     g12996(.A1(new_n13248), .A2(new_n13249), .B(new_n13252), .Y(new_n13253));
  NAND2xp33_ASAP7_75t_L     g12997(.A(new_n13251), .B(new_n13253), .Y(new_n13254));
  AOI22xp33_ASAP7_75t_L     g12998(.A1(new_n3029), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n3258), .Y(new_n13255));
  OAI221xp5_ASAP7_75t_L     g12999(.A1(new_n3024), .A2(new_n4869), .B1(new_n3256), .B2(new_n5327), .C(new_n13255), .Y(new_n13256));
  XNOR2x2_ASAP7_75t_L       g13000(.A(\a[32] ), .B(new_n13256), .Y(new_n13257));
  MAJIxp5_ASAP7_75t_L       g13001(.A(new_n13180), .B(new_n13082), .C(new_n13086), .Y(new_n13258));
  XNOR2x2_ASAP7_75t_L       g13002(.A(new_n13257), .B(new_n13258), .Y(new_n13259));
  NAND2xp33_ASAP7_75t_L     g13003(.A(new_n13149), .B(new_n13150), .Y(new_n13260));
  INVx1_ASAP7_75t_L         g13004(.A(new_n13260), .Y(new_n13261));
  AOI22xp33_ASAP7_75t_L     g13005(.A1(new_n7111), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n7391), .Y(new_n13262));
  OAI221xp5_ASAP7_75t_L     g13006(.A1(new_n8558), .A2(new_n1774), .B1(new_n8237), .B2(new_n1915), .C(new_n13262), .Y(new_n13263));
  XNOR2x2_ASAP7_75t_L       g13007(.A(\a[50] ), .B(new_n13263), .Y(new_n13264));
  INVx1_ASAP7_75t_L         g13008(.A(new_n13264), .Y(new_n13265));
  A2O1A1Ixp33_ASAP7_75t_L   g13009(.A1(new_n12635), .A2(new_n12628), .B(new_n12898), .C(new_n13120), .Y(new_n13266));
  INVx1_ASAP7_75t_L         g13010(.A(new_n13110), .Y(new_n13267));
  AOI22xp33_ASAP7_75t_L     g13011(.A1(new_n9700), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n10027), .Y(new_n13268));
  OAI221xp5_ASAP7_75t_L     g13012(.A1(new_n10024), .A2(new_n784), .B1(new_n9696), .B2(new_n875), .C(new_n13268), .Y(new_n13269));
  XNOR2x2_ASAP7_75t_L       g13013(.A(\a[59] ), .B(new_n13269), .Y(new_n13270));
  AOI22xp33_ASAP7_75t_L     g13014(.A1(\b[9] ), .A2(new_n10939), .B1(\b[11] ), .B2(new_n10938), .Y(new_n13271));
  OAI221xp5_ASAP7_75t_L     g13015(.A1(new_n10937), .A2(new_n617), .B1(new_n10629), .B2(new_n685), .C(new_n13271), .Y(new_n13272));
  XNOR2x2_ASAP7_75t_L       g13016(.A(\a[62] ), .B(new_n13272), .Y(new_n13273));
  A2O1A1Ixp33_ASAP7_75t_L   g13017(.A1(new_n13102), .A2(new_n13103), .B(new_n13098), .C(new_n13095), .Y(new_n13274));
  NOR2xp33_ASAP7_75t_L      g13018(.A(new_n420), .B(new_n11535), .Y(new_n13275));
  INVx1_ASAP7_75t_L         g13019(.A(new_n13275), .Y(new_n13276));
  O2A1O1Ixp33_ASAP7_75t_L   g13020(.A1(new_n11253), .A2(new_n488), .B(new_n13276), .C(new_n13093), .Y(new_n13277));
  O2A1O1Ixp33_ASAP7_75t_L   g13021(.A1(new_n11247), .A2(new_n11249), .B(\b[8] ), .C(new_n13275), .Y(new_n13278));
  A2O1A1Ixp33_ASAP7_75t_L   g13022(.A1(new_n11533), .A2(\b[7] ), .B(new_n13091), .C(new_n13278), .Y(new_n13279));
  INVx1_ASAP7_75t_L         g13023(.A(new_n13279), .Y(new_n13280));
  NOR3xp33_ASAP7_75t_L      g13024(.A(new_n13274), .B(new_n13277), .C(new_n13280), .Y(new_n13281));
  NOR2xp33_ASAP7_75t_L      g13025(.A(new_n13280), .B(new_n13277), .Y(new_n13282));
  A2O1A1O1Ixp25_ASAP7_75t_L g13026(.A1(new_n13103), .A2(new_n13102), .B(new_n13098), .C(new_n13095), .D(new_n13282), .Y(new_n13283));
  NOR2xp33_ASAP7_75t_L      g13027(.A(new_n13283), .B(new_n13281), .Y(new_n13284));
  NOR2xp33_ASAP7_75t_L      g13028(.A(new_n13273), .B(new_n13284), .Y(new_n13285));
  INVx1_ASAP7_75t_L         g13029(.A(new_n13285), .Y(new_n13286));
  NAND2xp33_ASAP7_75t_L     g13030(.A(new_n13273), .B(new_n13284), .Y(new_n13287));
  NAND2xp33_ASAP7_75t_L     g13031(.A(new_n13287), .B(new_n13286), .Y(new_n13288));
  NOR2xp33_ASAP7_75t_L      g13032(.A(new_n13270), .B(new_n13288), .Y(new_n13289));
  INVx1_ASAP7_75t_L         g13033(.A(new_n13270), .Y(new_n13290));
  AOI21xp33_ASAP7_75t_L     g13034(.A1(new_n13287), .A2(new_n13286), .B(new_n13290), .Y(new_n13291));
  NOR2xp33_ASAP7_75t_L      g13035(.A(new_n13291), .B(new_n13289), .Y(new_n13292));
  O2A1O1Ixp33_ASAP7_75t_L   g13036(.A1(new_n13267), .A2(new_n13106), .B(new_n13115), .C(new_n13292), .Y(new_n13293));
  INVx1_ASAP7_75t_L         g13037(.A(new_n13293), .Y(new_n13294));
  NAND3xp33_ASAP7_75t_L     g13038(.A(new_n13292), .B(new_n13115), .C(new_n13111), .Y(new_n13295));
  AOI22xp33_ASAP7_75t_L     g13039(.A1(new_n8831), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n9115), .Y(new_n13296));
  OAI221xp5_ASAP7_75t_L     g13040(.A1(new_n10343), .A2(new_n1030), .B1(new_n10016), .B2(new_n1209), .C(new_n13296), .Y(new_n13297));
  XNOR2x2_ASAP7_75t_L       g13041(.A(\a[56] ), .B(new_n13297), .Y(new_n13298));
  NAND3xp33_ASAP7_75t_L     g13042(.A(new_n13294), .B(new_n13295), .C(new_n13298), .Y(new_n13299));
  AO21x2_ASAP7_75t_L        g13043(.A1(new_n13295), .A2(new_n13294), .B(new_n13298), .Y(new_n13300));
  NAND2xp33_ASAP7_75t_L     g13044(.A(new_n13299), .B(new_n13300), .Y(new_n13301));
  O2A1O1Ixp33_ASAP7_75t_L   g13045(.A1(new_n13117), .A2(new_n13266), .B(new_n13128), .C(new_n13301), .Y(new_n13302));
  INVx1_ASAP7_75t_L         g13046(.A(new_n13302), .Y(new_n13303));
  NAND3xp33_ASAP7_75t_L     g13047(.A(new_n13128), .B(new_n13121), .C(new_n13301), .Y(new_n13304));
  NAND2xp33_ASAP7_75t_L     g13048(.A(new_n13304), .B(new_n13303), .Y(new_n13305));
  AOI22xp33_ASAP7_75t_L     g13049(.A1(new_n7960), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n8537), .Y(new_n13306));
  OAI221xp5_ASAP7_75t_L     g13050(.A1(new_n8817), .A2(new_n1432), .B1(new_n7957), .B2(new_n1547), .C(new_n13306), .Y(new_n13307));
  XNOR2x2_ASAP7_75t_L       g13051(.A(\a[53] ), .B(new_n13307), .Y(new_n13308));
  XOR2x2_ASAP7_75t_L        g13052(.A(new_n13308), .B(new_n13305), .Y(new_n13309));
  INVx1_ASAP7_75t_L         g13053(.A(new_n13135), .Y(new_n13310));
  AO21x2_ASAP7_75t_L        g13054(.A1(new_n13139), .A2(new_n13136), .B(new_n13310), .Y(new_n13311));
  XNOR2x2_ASAP7_75t_L       g13055(.A(new_n13311), .B(new_n13309), .Y(new_n13312));
  NAND2xp33_ASAP7_75t_L     g13056(.A(new_n13265), .B(new_n13312), .Y(new_n13313));
  INVx1_ASAP7_75t_L         g13057(.A(new_n13312), .Y(new_n13314));
  NAND2xp33_ASAP7_75t_L     g13058(.A(new_n13264), .B(new_n13314), .Y(new_n13315));
  NAND2xp33_ASAP7_75t_L     g13059(.A(new_n13313), .B(new_n13315), .Y(new_n13316));
  NAND2xp33_ASAP7_75t_L     g13060(.A(new_n13148), .B(new_n13145), .Y(new_n13317));
  OAI31xp33_ASAP7_75t_L     g13061(.A1(new_n13140), .A2(new_n13144), .A3(new_n13141), .B(new_n13317), .Y(new_n13318));
  XNOR2x2_ASAP7_75t_L       g13062(.A(new_n13318), .B(new_n13316), .Y(new_n13319));
  AOI22xp33_ASAP7_75t_L     g13063(.A1(new_n6376), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n6648), .Y(new_n13320));
  OAI221xp5_ASAP7_75t_L     g13064(.A1(new_n6646), .A2(new_n2067), .B1(new_n6636), .B2(new_n2355), .C(new_n13320), .Y(new_n13321));
  XNOR2x2_ASAP7_75t_L       g13065(.A(\a[47] ), .B(new_n13321), .Y(new_n13322));
  XNOR2x2_ASAP7_75t_L       g13066(.A(new_n13322), .B(new_n13319), .Y(new_n13323));
  A2O1A1Ixp33_ASAP7_75t_L   g13067(.A1(new_n13151), .A2(new_n13154), .B(new_n13261), .C(new_n13323), .Y(new_n13324));
  NAND2xp33_ASAP7_75t_L     g13068(.A(new_n13154), .B(new_n13151), .Y(new_n13325));
  INVx1_ASAP7_75t_L         g13069(.A(new_n13325), .Y(new_n13326));
  OR3x1_ASAP7_75t_L         g13070(.A(new_n13323), .B(new_n13261), .C(new_n13326), .Y(new_n13327));
  AOI22xp33_ASAP7_75t_L     g13071(.A1(new_n5624), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n5901), .Y(new_n13328));
  OAI221xp5_ASAP7_75t_L     g13072(.A1(new_n5900), .A2(new_n2666), .B1(new_n5892), .B2(new_n2695), .C(new_n13328), .Y(new_n13329));
  XNOR2x2_ASAP7_75t_L       g13073(.A(\a[44] ), .B(new_n13329), .Y(new_n13330));
  NAND3xp33_ASAP7_75t_L     g13074(.A(new_n13327), .B(new_n13324), .C(new_n13330), .Y(new_n13331));
  AO21x2_ASAP7_75t_L        g13075(.A1(new_n13324), .A2(new_n13327), .B(new_n13330), .Y(new_n13332));
  NAND2xp33_ASAP7_75t_L     g13076(.A(new_n13331), .B(new_n13332), .Y(new_n13333));
  MAJx2_ASAP7_75t_L         g13077(.A(new_n13155), .B(new_n13156), .C(new_n13163), .Y(new_n13334));
  XOR2x2_ASAP7_75t_L        g13078(.A(new_n13334), .B(new_n13333), .Y(new_n13335));
  AOI22xp33_ASAP7_75t_L     g13079(.A1(new_n4920), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n5167), .Y(new_n13336));
  OAI221xp5_ASAP7_75t_L     g13080(.A1(new_n5154), .A2(new_n3180), .B1(new_n5158), .B2(new_n11047), .C(new_n13336), .Y(new_n13337));
  XNOR2x2_ASAP7_75t_L       g13081(.A(\a[41] ), .B(new_n13337), .Y(new_n13338));
  INVx1_ASAP7_75t_L         g13082(.A(new_n13338), .Y(new_n13339));
  XNOR2x2_ASAP7_75t_L       g13083(.A(new_n13339), .B(new_n13335), .Y(new_n13340));
  AO21x2_ASAP7_75t_L        g13084(.A1(new_n13166), .A2(new_n13172), .B(new_n13340), .Y(new_n13341));
  NAND3xp33_ASAP7_75t_L     g13085(.A(new_n13340), .B(new_n13172), .C(new_n13166), .Y(new_n13342));
  AOI22xp33_ASAP7_75t_L     g13086(.A1(new_n4283), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n4512), .Y(new_n13343));
  OAI221xp5_ASAP7_75t_L     g13087(.A1(new_n4277), .A2(new_n3584), .B1(new_n4499), .B2(new_n10137), .C(new_n13343), .Y(new_n13344));
  XNOR2x2_ASAP7_75t_L       g13088(.A(\a[38] ), .B(new_n13344), .Y(new_n13345));
  NAND3xp33_ASAP7_75t_L     g13089(.A(new_n13341), .B(new_n13342), .C(new_n13345), .Y(new_n13346));
  AO21x2_ASAP7_75t_L        g13090(.A1(new_n13342), .A2(new_n13341), .B(new_n13345), .Y(new_n13347));
  NOR2xp33_ASAP7_75t_L      g13091(.A(new_n13174), .B(new_n13173), .Y(new_n13348));
  NOR2xp33_ASAP7_75t_L      g13092(.A(new_n13348), .B(new_n13176), .Y(new_n13349));
  NAND3xp33_ASAP7_75t_L     g13093(.A(new_n13349), .B(new_n13347), .C(new_n13346), .Y(new_n13350));
  NAND2xp33_ASAP7_75t_L     g13094(.A(new_n13346), .B(new_n13347), .Y(new_n13351));
  A2O1A1Ixp33_ASAP7_75t_L   g13095(.A1(new_n13178), .A2(new_n13177), .B(new_n13348), .C(new_n13351), .Y(new_n13352));
  NAND2xp33_ASAP7_75t_L     g13096(.A(new_n13352), .B(new_n13350), .Y(new_n13353));
  AOI22xp33_ASAP7_75t_L     g13097(.A1(new_n3633), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n3858), .Y(new_n13354));
  OAI221xp5_ASAP7_75t_L     g13098(.A1(new_n3853), .A2(new_n4424), .B1(new_n3856), .B2(new_n4641), .C(new_n13354), .Y(new_n13355));
  XNOR2x2_ASAP7_75t_L       g13099(.A(\a[35] ), .B(new_n13355), .Y(new_n13356));
  XNOR2x2_ASAP7_75t_L       g13100(.A(new_n13356), .B(new_n13353), .Y(new_n13357));
  XNOR2x2_ASAP7_75t_L       g13101(.A(new_n13259), .B(new_n13357), .Y(new_n13358));
  XOR2x2_ASAP7_75t_L        g13102(.A(new_n13358), .B(new_n13254), .Y(new_n13359));
  XNOR2x2_ASAP7_75t_L       g13103(.A(new_n13359), .B(new_n13244), .Y(new_n13360));
  OAI21xp33_ASAP7_75t_L     g13104(.A1(new_n13238), .A2(new_n13236), .B(new_n13360), .Y(new_n13361));
  OR3x1_ASAP7_75t_L         g13105(.A(new_n13360), .B(new_n13236), .C(new_n13238), .Y(new_n13362));
  AND2x2_ASAP7_75t_L        g13106(.A(new_n13361), .B(new_n13362), .Y(new_n13363));
  INVx1_ASAP7_75t_L         g13107(.A(new_n13190), .Y(new_n13364));
  A2O1A1O1Ixp25_ASAP7_75t_L g13108(.A1(new_n12843), .A2(new_n13050), .B(new_n12965), .C(new_n13052), .D(new_n13049), .Y(new_n13365));
  AOI21xp33_ASAP7_75t_L     g13109(.A1(new_n13364), .A2(new_n13054), .B(new_n13365), .Y(new_n13366));
  NAND2xp33_ASAP7_75t_L     g13110(.A(\b[52] ), .B(new_n1362), .Y(new_n13367));
  OAI221xp5_ASAP7_75t_L     g13111(.A1(new_n1372), .A2(new_n8165), .B1(new_n7616), .B2(new_n1483), .C(new_n13367), .Y(new_n13368));
  AOI21xp33_ASAP7_75t_L     g13112(.A1(new_n8173), .A2(new_n1365), .B(new_n13368), .Y(new_n13369));
  NAND2xp33_ASAP7_75t_L     g13113(.A(\a[20] ), .B(new_n13369), .Y(new_n13370));
  A2O1A1Ixp33_ASAP7_75t_L   g13114(.A1(new_n8173), .A2(new_n1365), .B(new_n13368), .C(new_n1356), .Y(new_n13371));
  NAND2xp33_ASAP7_75t_L     g13115(.A(new_n13371), .B(new_n13370), .Y(new_n13372));
  XNOR2x2_ASAP7_75t_L       g13116(.A(new_n13372), .B(new_n13366), .Y(new_n13373));
  XOR2x2_ASAP7_75t_L        g13117(.A(new_n13363), .B(new_n13373), .Y(new_n13374));
  OR2x4_ASAP7_75t_L         g13118(.A(new_n13232), .B(new_n13374), .Y(new_n13375));
  NAND2xp33_ASAP7_75t_L     g13119(.A(new_n13232), .B(new_n13374), .Y(new_n13376));
  NAND2xp33_ASAP7_75t_L     g13120(.A(new_n13376), .B(new_n13375), .Y(new_n13377));
  AOI22xp33_ASAP7_75t_L     g13121(.A1(new_n811), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n900), .Y(new_n13378));
  OAI221xp5_ASAP7_75t_L     g13122(.A1(new_n904), .A2(new_n9920), .B1(new_n898), .B2(new_n11152), .C(new_n13378), .Y(new_n13379));
  XNOR2x2_ASAP7_75t_L       g13123(.A(\a[14] ), .B(new_n13379), .Y(new_n13380));
  NOR3xp33_ASAP7_75t_L      g13124(.A(new_n13195), .B(new_n13380), .C(new_n13041), .Y(new_n13381));
  INVx1_ASAP7_75t_L         g13125(.A(new_n13380), .Y(new_n13382));
  O2A1O1Ixp33_ASAP7_75t_L   g13126(.A1(new_n13040), .A2(new_n13194), .B(new_n13196), .C(new_n13382), .Y(new_n13383));
  NOR2xp33_ASAP7_75t_L      g13127(.A(new_n13383), .B(new_n13381), .Y(new_n13384));
  XNOR2x2_ASAP7_75t_L       g13128(.A(new_n13384), .B(new_n13377), .Y(new_n13385));
  NAND2xp33_ASAP7_75t_L     g13129(.A(new_n13385), .B(new_n13225), .Y(new_n13386));
  O2A1O1Ixp33_ASAP7_75t_L   g13130(.A1(new_n13033), .A2(new_n13030), .B(new_n13217), .C(new_n13224), .Y(new_n13387));
  AOI21xp33_ASAP7_75t_L     g13131(.A1(new_n13223), .A2(new_n13222), .B(new_n13218), .Y(new_n13388));
  NOR2xp33_ASAP7_75t_L      g13132(.A(new_n13387), .B(new_n13388), .Y(new_n13389));
  XOR2x2_ASAP7_75t_L        g13133(.A(new_n13384), .B(new_n13377), .Y(new_n13390));
  NAND2xp33_ASAP7_75t_L     g13134(.A(new_n13390), .B(new_n13389), .Y(new_n13391));
  NAND2xp33_ASAP7_75t_L     g13135(.A(new_n13386), .B(new_n13391), .Y(new_n13392));
  A2O1A1Ixp33_ASAP7_75t_L   g13136(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n441), .Y(new_n13393));
  A2O1A1Ixp33_ASAP7_75t_L   g13137(.A1(new_n13393), .A2(new_n516), .B(new_n11468), .C(\a[8] ), .Y(new_n13394));
  O2A1O1Ixp33_ASAP7_75t_L   g13138(.A1(new_n469), .A2(new_n12060), .B(new_n516), .C(new_n11468), .Y(new_n13395));
  NAND2xp33_ASAP7_75t_L     g13139(.A(new_n435), .B(new_n13395), .Y(new_n13396));
  AND2x2_ASAP7_75t_L        g13140(.A(new_n13396), .B(new_n13394), .Y(new_n13397));
  A2O1A1O1Ixp25_ASAP7_75t_L g13141(.A1(new_n12996), .A2(new_n12829), .B(new_n13024), .C(new_n13201), .D(new_n13397), .Y(new_n13398));
  A2O1A1Ixp33_ASAP7_75t_L   g13142(.A1(new_n12996), .A2(new_n12829), .B(new_n13024), .C(new_n13201), .Y(new_n13399));
  INVx1_ASAP7_75t_L         g13143(.A(new_n13397), .Y(new_n13400));
  NOR2xp33_ASAP7_75t_L      g13144(.A(new_n13400), .B(new_n13399), .Y(new_n13401));
  NOR3xp33_ASAP7_75t_L      g13145(.A(new_n13392), .B(new_n13398), .C(new_n13401), .Y(new_n13402));
  INVx1_ASAP7_75t_L         g13146(.A(new_n13398), .Y(new_n13403));
  INVx1_ASAP7_75t_L         g13147(.A(new_n13401), .Y(new_n13404));
  AOI22xp33_ASAP7_75t_L     g13148(.A1(new_n13386), .A2(new_n13391), .B1(new_n13403), .B2(new_n13404), .Y(new_n13405));
  NAND2xp33_ASAP7_75t_L     g13149(.A(new_n13019), .B(new_n13020), .Y(new_n13406));
  A2O1A1Ixp33_ASAP7_75t_L   g13150(.A1(new_n13202), .A2(new_n13201), .B(new_n13021), .C(new_n13406), .Y(new_n13407));
  NOR3xp33_ASAP7_75t_L      g13151(.A(new_n13402), .B(new_n13405), .C(new_n13407), .Y(new_n13408));
  NAND4xp25_ASAP7_75t_L     g13152(.A(new_n13404), .B(new_n13386), .C(new_n13391), .D(new_n13403), .Y(new_n13409));
  OAI21xp33_ASAP7_75t_L     g13153(.A1(new_n13398), .A2(new_n13401), .B(new_n13392), .Y(new_n13410));
  AOI22xp33_ASAP7_75t_L     g13154(.A1(new_n13406), .A2(new_n13203), .B1(new_n13409), .B2(new_n13410), .Y(new_n13411));
  NOR2xp33_ASAP7_75t_L      g13155(.A(new_n13411), .B(new_n13408), .Y(new_n13412));
  A2O1A1Ixp33_ASAP7_75t_L   g13156(.A1(new_n13214), .A2(new_n13210), .B(new_n13208), .C(new_n13412), .Y(new_n13413));
  INVx1_ASAP7_75t_L         g13157(.A(new_n13413), .Y(new_n13414));
  A2O1A1Ixp33_ASAP7_75t_L   g13158(.A1(new_n13204), .A2(new_n13203), .B(new_n13207), .C(new_n13211), .Y(new_n13415));
  NOR2xp33_ASAP7_75t_L      g13159(.A(new_n13412), .B(new_n13415), .Y(new_n13416));
  NOR2xp33_ASAP7_75t_L      g13160(.A(new_n13414), .B(new_n13416), .Y(\f[71] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13161(.A1(new_n13199), .A2(new_n13034), .B(new_n13031), .C(new_n13224), .Y(new_n13418));
  AOI22xp33_ASAP7_75t_L     g13162(.A1(\b[61] ), .A2(new_n651), .B1(\b[63] ), .B2(new_n581), .Y(new_n13419));
  A2O1A1Ixp33_ASAP7_75t_L   g13163(.A1(new_n11470), .A2(new_n11473), .B(new_n577), .C(new_n13419), .Y(new_n13420));
  AOI21xp33_ASAP7_75t_L     g13164(.A1(new_n584), .A2(\b[62] ), .B(new_n13420), .Y(new_n13421));
  NAND2xp33_ASAP7_75t_L     g13165(.A(\a[11] ), .B(new_n13421), .Y(new_n13422));
  A2O1A1Ixp33_ASAP7_75t_L   g13166(.A1(\b[62] ), .A2(new_n584), .B(new_n13420), .C(new_n574), .Y(new_n13423));
  AND2x2_ASAP7_75t_L        g13167(.A(new_n13423), .B(new_n13422), .Y(new_n13424));
  INVx1_ASAP7_75t_L         g13168(.A(new_n13424), .Y(new_n13425));
  O2A1O1Ixp33_ASAP7_75t_L   g13169(.A1(new_n13390), .A2(new_n13389), .B(new_n13418), .C(new_n13425), .Y(new_n13426));
  NAND3xp33_ASAP7_75t_L     g13170(.A(new_n13386), .B(new_n13418), .C(new_n13425), .Y(new_n13427));
  INVx1_ASAP7_75t_L         g13171(.A(new_n13427), .Y(new_n13428));
  A2O1A1Ixp33_ASAP7_75t_L   g13172(.A1(new_n13197), .A2(new_n13039), .B(new_n13041), .C(new_n13382), .Y(new_n13429));
  A2O1A1Ixp33_ASAP7_75t_L   g13173(.A1(new_n13375), .A2(new_n13376), .B(new_n13384), .C(new_n13429), .Y(new_n13430));
  AOI22xp33_ASAP7_75t_L     g13174(.A1(new_n811), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n900), .Y(new_n13431));
  OAI221xp5_ASAP7_75t_L     g13175(.A1(new_n904), .A2(new_n9947), .B1(new_n898), .B2(new_n11446), .C(new_n13431), .Y(new_n13432));
  XNOR2x2_ASAP7_75t_L       g13176(.A(\a[14] ), .B(new_n13432), .Y(new_n13433));
  XNOR2x2_ASAP7_75t_L       g13177(.A(new_n13433), .B(new_n13430), .Y(new_n13434));
  AOI22xp33_ASAP7_75t_L     g13178(.A1(new_n1076), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1253), .Y(new_n13435));
  OAI221xp5_ASAP7_75t_L     g13179(.A1(new_n1154), .A2(new_n9323), .B1(new_n1156), .B2(new_n9627), .C(new_n13435), .Y(new_n13436));
  XNOR2x2_ASAP7_75t_L       g13180(.A(\a[17] ), .B(new_n13436), .Y(new_n13437));
  INVx1_ASAP7_75t_L         g13181(.A(new_n13437), .Y(new_n13438));
  O2A1O1Ixp33_ASAP7_75t_L   g13182(.A1(new_n13232), .A2(new_n13374), .B(new_n13230), .C(new_n13438), .Y(new_n13439));
  INVx1_ASAP7_75t_L         g13183(.A(new_n13439), .Y(new_n13440));
  NAND3xp33_ASAP7_75t_L     g13184(.A(new_n13375), .B(new_n13230), .C(new_n13438), .Y(new_n13441));
  NAND2xp33_ASAP7_75t_L     g13185(.A(new_n13440), .B(new_n13441), .Y(new_n13442));
  NAND2xp33_ASAP7_75t_L     g13186(.A(new_n13363), .B(new_n13373), .Y(new_n13443));
  AOI22xp33_ASAP7_75t_L     g13187(.A1(new_n1360), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1581), .Y(new_n13444));
  OAI221xp5_ASAP7_75t_L     g13188(.A1(new_n1373), .A2(new_n8165), .B1(new_n1359), .B2(new_n8465), .C(new_n13444), .Y(new_n13445));
  XNOR2x2_ASAP7_75t_L       g13189(.A(\a[20] ), .B(new_n13445), .Y(new_n13446));
  INVx1_ASAP7_75t_L         g13190(.A(new_n13446), .Y(new_n13447));
  A2O1A1O1Ixp25_ASAP7_75t_L g13191(.A1(new_n13370), .A2(new_n13371), .B(new_n13366), .C(new_n13443), .D(new_n13447), .Y(new_n13448));
  A2O1A1Ixp33_ASAP7_75t_L   g13192(.A1(new_n13370), .A2(new_n13371), .B(new_n13366), .C(new_n13443), .Y(new_n13449));
  NOR2xp33_ASAP7_75t_L      g13193(.A(new_n13446), .B(new_n13449), .Y(new_n13450));
  AOI22xp33_ASAP7_75t_L     g13194(.A1(new_n1704), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1837), .Y(new_n13451));
  OAI221xp5_ASAP7_75t_L     g13195(.A1(new_n1699), .A2(new_n7593), .B1(new_n1827), .B2(new_n7623), .C(new_n13451), .Y(new_n13452));
  XNOR2x2_ASAP7_75t_L       g13196(.A(\a[23] ), .B(new_n13452), .Y(new_n13453));
  INVx1_ASAP7_75t_L         g13197(.A(new_n13453), .Y(new_n13454));
  A2O1A1Ixp33_ASAP7_75t_L   g13198(.A1(new_n13188), .A2(new_n13059), .B(new_n13235), .C(new_n13362), .Y(new_n13455));
  NAND2xp33_ASAP7_75t_L     g13199(.A(new_n13454), .B(new_n13455), .Y(new_n13456));
  OAI211xp5_ASAP7_75t_L     g13200(.A1(new_n13237), .A2(new_n13235), .B(new_n13362), .C(new_n13453), .Y(new_n13457));
  AOI22xp33_ASAP7_75t_L     g13201(.A1(new_n2114), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n2259), .Y(new_n13458));
  OAI221xp5_ASAP7_75t_L     g13202(.A1(new_n2109), .A2(new_n6812), .B1(new_n2257), .B2(new_n6837), .C(new_n13458), .Y(new_n13459));
  XNOR2x2_ASAP7_75t_L       g13203(.A(\a[26] ), .B(new_n13459), .Y(new_n13460));
  MAJIxp5_ASAP7_75t_L       g13204(.A(new_n13359), .B(new_n13241), .C(new_n13243), .Y(new_n13461));
  XNOR2x2_ASAP7_75t_L       g13205(.A(new_n13460), .B(new_n13461), .Y(new_n13462));
  MAJIxp5_ASAP7_75t_L       g13206(.A(new_n13358), .B(new_n13250), .C(new_n13252), .Y(new_n13463));
  AOI22xp33_ASAP7_75t_L     g13207(.A1(new_n2552), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n2736), .Y(new_n13464));
  OAI221xp5_ASAP7_75t_L     g13208(.A1(new_n2547), .A2(new_n5829), .B1(new_n2734), .B2(new_n6329), .C(new_n13464), .Y(new_n13465));
  XNOR2x2_ASAP7_75t_L       g13209(.A(\a[29] ), .B(new_n13465), .Y(new_n13466));
  INVx1_ASAP7_75t_L         g13210(.A(new_n13466), .Y(new_n13467));
  XNOR2x2_ASAP7_75t_L       g13211(.A(new_n13467), .B(new_n13463), .Y(new_n13468));
  MAJx2_ASAP7_75t_L         g13212(.A(new_n13357), .B(new_n13258), .C(new_n13257), .Y(new_n13469));
  AOI22xp33_ASAP7_75t_L     g13213(.A1(new_n3029), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n3258), .Y(new_n13470));
  OAI221xp5_ASAP7_75t_L     g13214(.A1(new_n3024), .A2(new_n5321), .B1(new_n3256), .B2(new_n5346), .C(new_n13470), .Y(new_n13471));
  XNOR2x2_ASAP7_75t_L       g13215(.A(\a[32] ), .B(new_n13471), .Y(new_n13472));
  XOR2x2_ASAP7_75t_L        g13216(.A(new_n13472), .B(new_n13469), .Y(new_n13473));
  AOI22xp33_ASAP7_75t_L     g13217(.A1(new_n4283), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n4512), .Y(new_n13474));
  OAI221xp5_ASAP7_75t_L     g13218(.A1(new_n4277), .A2(new_n3804), .B1(new_n4499), .B2(new_n4223), .C(new_n13474), .Y(new_n13475));
  XNOR2x2_ASAP7_75t_L       g13219(.A(\a[38] ), .B(new_n13475), .Y(new_n13476));
  MAJx2_ASAP7_75t_L         g13220(.A(new_n13333), .B(new_n13334), .C(new_n13339), .Y(new_n13477));
  AOI22xp33_ASAP7_75t_L     g13221(.A1(new_n4920), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n5167), .Y(new_n13478));
  OAI221xp5_ASAP7_75t_L     g13222(.A1(new_n5154), .A2(new_n3207), .B1(new_n5158), .B2(new_n3572), .C(new_n13478), .Y(new_n13479));
  XNOR2x2_ASAP7_75t_L       g13223(.A(\a[41] ), .B(new_n13479), .Y(new_n13480));
  INVx1_ASAP7_75t_L         g13224(.A(new_n13309), .Y(new_n13481));
  AOI22xp33_ASAP7_75t_L     g13225(.A1(new_n7111), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n7391), .Y(new_n13482));
  OAI221xp5_ASAP7_75t_L     g13226(.A1(new_n8558), .A2(new_n1909), .B1(new_n8237), .B2(new_n2477), .C(new_n13482), .Y(new_n13483));
  XNOR2x2_ASAP7_75t_L       g13227(.A(\a[50] ), .B(new_n13483), .Y(new_n13484));
  AOI22xp33_ASAP7_75t_L     g13228(.A1(\b[10] ), .A2(new_n10939), .B1(\b[12] ), .B2(new_n10938), .Y(new_n13485));
  OAI221xp5_ASAP7_75t_L     g13229(.A1(new_n10937), .A2(new_n679), .B1(new_n10629), .B2(new_n768), .C(new_n13485), .Y(new_n13486));
  XNOR2x2_ASAP7_75t_L       g13230(.A(\a[62] ), .B(new_n13486), .Y(new_n13487));
  NOR2xp33_ASAP7_75t_L      g13231(.A(new_n488), .B(new_n11535), .Y(new_n13488));
  O2A1O1Ixp33_ASAP7_75t_L   g13232(.A1(new_n488), .A2(new_n11253), .B(new_n13276), .C(new_n435), .Y(new_n13489));
  AOI211xp5_ASAP7_75t_L     g13233(.A1(new_n11533), .A2(\b[8] ), .B(new_n13275), .C(\a[8] ), .Y(new_n13490));
  NOR2xp33_ASAP7_75t_L      g13234(.A(new_n13490), .B(new_n13489), .Y(new_n13491));
  INVx1_ASAP7_75t_L         g13235(.A(new_n13491), .Y(new_n13492));
  A2O1A1Ixp33_ASAP7_75t_L   g13236(.A1(new_n11533), .A2(\b[9] ), .B(new_n13488), .C(new_n13492), .Y(new_n13493));
  O2A1O1Ixp33_ASAP7_75t_L   g13237(.A1(new_n11247), .A2(new_n11249), .B(\b[9] ), .C(new_n13488), .Y(new_n13494));
  NAND2xp33_ASAP7_75t_L     g13238(.A(new_n13494), .B(new_n13491), .Y(new_n13495));
  AND2x2_ASAP7_75t_L        g13239(.A(new_n13495), .B(new_n13493), .Y(new_n13496));
  A2O1A1O1Ixp25_ASAP7_75t_L g13240(.A1(new_n13103), .A2(new_n13102), .B(new_n13098), .C(new_n13095), .D(new_n13277), .Y(new_n13497));
  A2O1A1Ixp33_ASAP7_75t_L   g13241(.A1(new_n13093), .A2(new_n13278), .B(new_n13497), .C(new_n13496), .Y(new_n13498));
  OR3x1_ASAP7_75t_L         g13242(.A(new_n13497), .B(new_n13280), .C(new_n13496), .Y(new_n13499));
  NAND3xp33_ASAP7_75t_L     g13243(.A(new_n13487), .B(new_n13498), .C(new_n13499), .Y(new_n13500));
  AO21x2_ASAP7_75t_L        g13244(.A1(new_n13499), .A2(new_n13498), .B(new_n13487), .Y(new_n13501));
  NAND2xp33_ASAP7_75t_L     g13245(.A(new_n13500), .B(new_n13501), .Y(new_n13502));
  AOI22xp33_ASAP7_75t_L     g13246(.A1(new_n9700), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n10027), .Y(new_n13503));
  OAI221xp5_ASAP7_75t_L     g13247(.A1(new_n10024), .A2(new_n869), .B1(new_n9696), .B2(new_n950), .C(new_n13503), .Y(new_n13504));
  XNOR2x2_ASAP7_75t_L       g13248(.A(new_n9693), .B(new_n13504), .Y(new_n13505));
  NAND2xp33_ASAP7_75t_L     g13249(.A(new_n13502), .B(new_n13505), .Y(new_n13506));
  OR2x4_ASAP7_75t_L         g13250(.A(new_n13502), .B(new_n13505), .Y(new_n13507));
  OAI211xp5_ASAP7_75t_L     g13251(.A1(new_n13285), .A2(new_n13289), .B(new_n13507), .C(new_n13506), .Y(new_n13508));
  INVx1_ASAP7_75t_L         g13252(.A(new_n13289), .Y(new_n13509));
  NAND2xp33_ASAP7_75t_L     g13253(.A(new_n13506), .B(new_n13507), .Y(new_n13510));
  NAND3xp33_ASAP7_75t_L     g13254(.A(new_n13510), .B(new_n13509), .C(new_n13286), .Y(new_n13511));
  NAND2xp33_ASAP7_75t_L     g13255(.A(new_n13508), .B(new_n13511), .Y(new_n13512));
  AOI22xp33_ASAP7_75t_L     g13256(.A1(new_n8831), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n9115), .Y(new_n13513));
  OAI221xp5_ASAP7_75t_L     g13257(.A1(new_n10343), .A2(new_n1201), .B1(new_n10016), .B2(new_n1320), .C(new_n13513), .Y(new_n13514));
  XNOR2x2_ASAP7_75t_L       g13258(.A(\a[56] ), .B(new_n13514), .Y(new_n13515));
  XOR2x2_ASAP7_75t_L        g13259(.A(new_n13515), .B(new_n13512), .Y(new_n13516));
  AO21x2_ASAP7_75t_L        g13260(.A1(new_n13294), .A2(new_n13299), .B(new_n13516), .Y(new_n13517));
  NAND3xp33_ASAP7_75t_L     g13261(.A(new_n13516), .B(new_n13299), .C(new_n13294), .Y(new_n13518));
  NAND2xp33_ASAP7_75t_L     g13262(.A(new_n13518), .B(new_n13517), .Y(new_n13519));
  AOI22xp33_ASAP7_75t_L     g13263(.A1(new_n7960), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n8537), .Y(new_n13520));
  OAI221xp5_ASAP7_75t_L     g13264(.A1(new_n8817), .A2(new_n1539), .B1(new_n7957), .B2(new_n1662), .C(new_n13520), .Y(new_n13521));
  XNOR2x2_ASAP7_75t_L       g13265(.A(\a[53] ), .B(new_n13521), .Y(new_n13522));
  XNOR2x2_ASAP7_75t_L       g13266(.A(new_n13522), .B(new_n13519), .Y(new_n13523));
  O2A1O1Ixp33_ASAP7_75t_L   g13267(.A1(new_n13302), .A2(new_n13308), .B(new_n13304), .C(new_n13523), .Y(new_n13524));
  OA211x2_ASAP7_75t_L       g13268(.A1(new_n13302), .A2(new_n13308), .B(new_n13523), .C(new_n13304), .Y(new_n13525));
  NOR2xp33_ASAP7_75t_L      g13269(.A(new_n13524), .B(new_n13525), .Y(new_n13526));
  XNOR2x2_ASAP7_75t_L       g13270(.A(new_n13484), .B(new_n13526), .Y(new_n13527));
  O2A1O1Ixp33_ASAP7_75t_L   g13271(.A1(new_n13481), .A2(new_n13311), .B(new_n13313), .C(new_n13527), .Y(new_n13528));
  OR3x1_ASAP7_75t_L         g13272(.A(new_n13481), .B(new_n13310), .C(new_n13140), .Y(new_n13529));
  AND3x1_ASAP7_75t_L        g13273(.A(new_n13527), .B(new_n13313), .C(new_n13529), .Y(new_n13530));
  NOR2xp33_ASAP7_75t_L      g13274(.A(new_n13528), .B(new_n13530), .Y(new_n13531));
  AOI22xp33_ASAP7_75t_L     g13275(.A1(new_n6376), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n6648), .Y(new_n13532));
  OAI221xp5_ASAP7_75t_L     g13276(.A1(new_n6646), .A2(new_n2348), .B1(new_n6636), .B2(new_n2505), .C(new_n13532), .Y(new_n13533));
  XNOR2x2_ASAP7_75t_L       g13277(.A(\a[47] ), .B(new_n13533), .Y(new_n13534));
  XNOR2x2_ASAP7_75t_L       g13278(.A(new_n13534), .B(new_n13531), .Y(new_n13535));
  MAJx2_ASAP7_75t_L         g13279(.A(new_n13316), .B(new_n13318), .C(new_n13322), .Y(new_n13536));
  XNOR2x2_ASAP7_75t_L       g13280(.A(new_n13536), .B(new_n13535), .Y(new_n13537));
  AOI22xp33_ASAP7_75t_L     g13281(.A1(new_n5624), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n5901), .Y(new_n13538));
  OAI221xp5_ASAP7_75t_L     g13282(.A1(new_n5900), .A2(new_n2688), .B1(new_n5892), .B2(new_n2990), .C(new_n13538), .Y(new_n13539));
  XNOR2x2_ASAP7_75t_L       g13283(.A(\a[44] ), .B(new_n13539), .Y(new_n13540));
  XNOR2x2_ASAP7_75t_L       g13284(.A(new_n13540), .B(new_n13537), .Y(new_n13541));
  NAND2xp33_ASAP7_75t_L     g13285(.A(new_n13324), .B(new_n13331), .Y(new_n13542));
  XOR2x2_ASAP7_75t_L        g13286(.A(new_n13541), .B(new_n13542), .Y(new_n13543));
  XNOR2x2_ASAP7_75t_L       g13287(.A(new_n13480), .B(new_n13543), .Y(new_n13544));
  XNOR2x2_ASAP7_75t_L       g13288(.A(new_n13477), .B(new_n13544), .Y(new_n13545));
  XNOR2x2_ASAP7_75t_L       g13289(.A(new_n13476), .B(new_n13545), .Y(new_n13546));
  NAND2xp33_ASAP7_75t_L     g13290(.A(new_n13342), .B(new_n13346), .Y(new_n13547));
  XOR2x2_ASAP7_75t_L        g13291(.A(new_n13547), .B(new_n13546), .Y(new_n13548));
  AOI22xp33_ASAP7_75t_L     g13292(.A1(new_n3633), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n3858), .Y(new_n13549));
  OAI221xp5_ASAP7_75t_L     g13293(.A1(new_n3853), .A2(new_n4632), .B1(new_n3856), .B2(new_n4858), .C(new_n13549), .Y(new_n13550));
  XNOR2x2_ASAP7_75t_L       g13294(.A(\a[35] ), .B(new_n13550), .Y(new_n13551));
  INVx1_ASAP7_75t_L         g13295(.A(new_n13551), .Y(new_n13552));
  XNOR2x2_ASAP7_75t_L       g13296(.A(new_n13552), .B(new_n13548), .Y(new_n13553));
  OAI21xp33_ASAP7_75t_L     g13297(.A1(new_n13356), .A2(new_n13353), .B(new_n13352), .Y(new_n13554));
  XOR2x2_ASAP7_75t_L        g13298(.A(new_n13554), .B(new_n13553), .Y(new_n13555));
  XNOR2x2_ASAP7_75t_L       g13299(.A(new_n13555), .B(new_n13473), .Y(new_n13556));
  XNOR2x2_ASAP7_75t_L       g13300(.A(new_n13468), .B(new_n13556), .Y(new_n13557));
  XNOR2x2_ASAP7_75t_L       g13301(.A(new_n13557), .B(new_n13462), .Y(new_n13558));
  AO21x2_ASAP7_75t_L        g13302(.A1(new_n13457), .A2(new_n13456), .B(new_n13558), .Y(new_n13559));
  NAND3xp33_ASAP7_75t_L     g13303(.A(new_n13456), .B(new_n13457), .C(new_n13558), .Y(new_n13560));
  NAND2xp33_ASAP7_75t_L     g13304(.A(new_n13560), .B(new_n13559), .Y(new_n13561));
  OAI21xp33_ASAP7_75t_L     g13305(.A1(new_n13448), .A2(new_n13450), .B(new_n13561), .Y(new_n13562));
  INVx1_ASAP7_75t_L         g13306(.A(new_n13448), .Y(new_n13563));
  A2O1A1Ixp33_ASAP7_75t_L   g13307(.A1(new_n13364), .A2(new_n13054), .B(new_n13365), .C(new_n13372), .Y(new_n13564));
  AND2x2_ASAP7_75t_L        g13308(.A(new_n13564), .B(new_n13443), .Y(new_n13565));
  NAND2xp33_ASAP7_75t_L     g13309(.A(new_n13447), .B(new_n13565), .Y(new_n13566));
  NAND4xp25_ASAP7_75t_L     g13310(.A(new_n13566), .B(new_n13559), .C(new_n13560), .D(new_n13563), .Y(new_n13567));
  NAND2xp33_ASAP7_75t_L     g13311(.A(new_n13562), .B(new_n13567), .Y(new_n13568));
  XOR2x2_ASAP7_75t_L        g13312(.A(new_n13568), .B(new_n13442), .Y(new_n13569));
  XOR2x2_ASAP7_75t_L        g13313(.A(new_n13434), .B(new_n13569), .Y(new_n13570));
  OAI21xp33_ASAP7_75t_L     g13314(.A1(new_n13426), .A2(new_n13428), .B(new_n13570), .Y(new_n13571));
  INVx1_ASAP7_75t_L         g13315(.A(new_n13426), .Y(new_n13572));
  XNOR2x2_ASAP7_75t_L       g13316(.A(new_n13434), .B(new_n13569), .Y(new_n13573));
  NAND3xp33_ASAP7_75t_L     g13317(.A(new_n13573), .B(new_n13427), .C(new_n13572), .Y(new_n13574));
  OAI211xp5_ASAP7_75t_L     g13318(.A1(new_n13402), .A2(new_n13398), .B(new_n13571), .C(new_n13574), .Y(new_n13575));
  INVx1_ASAP7_75t_L         g13319(.A(new_n13399), .Y(new_n13576));
  A2O1A1Ixp33_ASAP7_75t_L   g13320(.A1(new_n13394), .A2(new_n13396), .B(new_n13576), .C(new_n13409), .Y(new_n13577));
  AO21x2_ASAP7_75t_L        g13321(.A1(new_n13574), .A2(new_n13571), .B(new_n13577), .Y(new_n13578));
  AND2x2_ASAP7_75t_L        g13322(.A(new_n13575), .B(new_n13578), .Y(new_n13579));
  A2O1A1Ixp33_ASAP7_75t_L   g13323(.A1(new_n13415), .A2(new_n13412), .B(new_n13408), .C(new_n13579), .Y(new_n13580));
  INVx1_ASAP7_75t_L         g13324(.A(new_n13580), .Y(new_n13581));
  INVx1_ASAP7_75t_L         g13325(.A(new_n13208), .Y(new_n13582));
  INVx1_ASAP7_75t_L         g13326(.A(new_n13408), .Y(new_n13583));
  A2O1A1Ixp33_ASAP7_75t_L   g13327(.A1(new_n13211), .A2(new_n13582), .B(new_n13411), .C(new_n13583), .Y(new_n13584));
  NOR2xp33_ASAP7_75t_L      g13328(.A(new_n13579), .B(new_n13584), .Y(new_n13585));
  NOR2xp33_ASAP7_75t_L      g13329(.A(new_n13585), .B(new_n13581), .Y(\f[72] ));
  INVx1_ASAP7_75t_L         g13330(.A(new_n13575), .Y(new_n13587));
  O2A1O1Ixp33_ASAP7_75t_L   g13331(.A1(new_n13390), .A2(new_n13389), .B(new_n13418), .C(new_n13424), .Y(new_n13588));
  O2A1O1Ixp33_ASAP7_75t_L   g13332(.A1(new_n13426), .A2(new_n13428), .B(new_n13570), .C(new_n13588), .Y(new_n13589));
  A2O1A1O1Ixp25_ASAP7_75t_L g13333(.A1(new_n13376), .A2(new_n13375), .B(new_n13384), .C(new_n13429), .D(new_n13433), .Y(new_n13590));
  NOR2xp33_ASAP7_75t_L      g13334(.A(new_n577), .B(new_n11500), .Y(new_n13591));
  AOI21xp33_ASAP7_75t_L     g13335(.A1(new_n651), .A2(\b[62] ), .B(new_n13591), .Y(new_n13592));
  OAI211xp5_ASAP7_75t_L     g13336(.A1(new_n11468), .A2(new_n821), .B(new_n13592), .C(\a[11] ), .Y(new_n13593));
  O2A1O1Ixp33_ASAP7_75t_L   g13337(.A1(new_n11468), .A2(new_n821), .B(new_n13592), .C(\a[11] ), .Y(new_n13594));
  INVx1_ASAP7_75t_L         g13338(.A(new_n13594), .Y(new_n13595));
  AND2x2_ASAP7_75t_L        g13339(.A(new_n13593), .B(new_n13595), .Y(new_n13596));
  A2O1A1Ixp33_ASAP7_75t_L   g13340(.A1(new_n13569), .A2(new_n13434), .B(new_n13590), .C(new_n13596), .Y(new_n13597));
  AOI211xp5_ASAP7_75t_L     g13341(.A1(new_n13569), .A2(new_n13434), .B(new_n13590), .C(new_n13596), .Y(new_n13598));
  INVx1_ASAP7_75t_L         g13342(.A(new_n13598), .Y(new_n13599));
  NAND2xp33_ASAP7_75t_L     g13343(.A(\b[59] ), .B(new_n900), .Y(new_n13600));
  OAI221xp5_ASAP7_75t_L     g13344(.A1(new_n977), .A2(new_n10847), .B1(new_n898), .B2(new_n10855), .C(new_n13600), .Y(new_n13601));
  AOI211xp5_ASAP7_75t_L     g13345(.A1(\b[60] ), .A2(new_n815), .B(new_n806), .C(new_n13601), .Y(new_n13602));
  INVx1_ASAP7_75t_L         g13346(.A(new_n13602), .Y(new_n13603));
  A2O1A1Ixp33_ASAP7_75t_L   g13347(.A1(\b[60] ), .A2(new_n815), .B(new_n13601), .C(new_n806), .Y(new_n13604));
  NAND2xp33_ASAP7_75t_L     g13348(.A(new_n13604), .B(new_n13603), .Y(new_n13605));
  OAI211xp5_ASAP7_75t_L     g13349(.A1(new_n13439), .A2(new_n13568), .B(new_n13605), .C(new_n13441), .Y(new_n13606));
  INVx1_ASAP7_75t_L         g13350(.A(new_n13606), .Y(new_n13607));
  O2A1O1Ixp33_ASAP7_75t_L   g13351(.A1(new_n13439), .A2(new_n13568), .B(new_n13441), .C(new_n13605), .Y(new_n13608));
  NAND2xp33_ASAP7_75t_L     g13352(.A(new_n13563), .B(new_n13566), .Y(new_n13609));
  A2O1A1O1Ixp25_ASAP7_75t_L g13353(.A1(new_n13370), .A2(new_n13371), .B(new_n13366), .C(new_n13443), .D(new_n13446), .Y(new_n13610));
  NOR2xp33_ASAP7_75t_L      g13354(.A(new_n9920), .B(new_n1259), .Y(new_n13611));
  AOI221xp5_ASAP7_75t_L     g13355(.A1(\b[57] ), .A2(new_n1080), .B1(\b[56] ), .B2(new_n1253), .C(new_n13611), .Y(new_n13612));
  OAI211xp5_ASAP7_75t_L     g13356(.A1(new_n1156), .A2(new_n9925), .B(\a[17] ), .C(new_n13612), .Y(new_n13613));
  O2A1O1Ixp33_ASAP7_75t_L   g13357(.A1(new_n1156), .A2(new_n9925), .B(new_n13612), .C(\a[17] ), .Y(new_n13614));
  INVx1_ASAP7_75t_L         g13358(.A(new_n13614), .Y(new_n13615));
  AND2x2_ASAP7_75t_L        g13359(.A(new_n13613), .B(new_n13615), .Y(new_n13616));
  A2O1A1Ixp33_ASAP7_75t_L   g13360(.A1(new_n13609), .A2(new_n13561), .B(new_n13610), .C(new_n13616), .Y(new_n13617));
  O2A1O1Ixp33_ASAP7_75t_L   g13361(.A1(new_n13448), .A2(new_n13450), .B(new_n13561), .C(new_n13610), .Y(new_n13618));
  INVx1_ASAP7_75t_L         g13362(.A(new_n13616), .Y(new_n13619));
  NAND2xp33_ASAP7_75t_L     g13363(.A(new_n13619), .B(new_n13618), .Y(new_n13620));
  AOI22xp33_ASAP7_75t_L     g13364(.A1(new_n1360), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1581), .Y(new_n13621));
  OAI221xp5_ASAP7_75t_L     g13365(.A1(new_n1373), .A2(new_n8458), .B1(new_n1359), .B2(new_n8768), .C(new_n13621), .Y(new_n13622));
  XNOR2x2_ASAP7_75t_L       g13366(.A(\a[20] ), .B(new_n13622), .Y(new_n13623));
  OA21x2_ASAP7_75t_L        g13367(.A1(new_n13235), .A2(new_n13237), .B(new_n13362), .Y(new_n13624));
  MAJx2_ASAP7_75t_L         g13368(.A(new_n13558), .B(new_n13453), .C(new_n13624), .Y(new_n13625));
  XNOR2x2_ASAP7_75t_L       g13369(.A(new_n13623), .B(new_n13625), .Y(new_n13626));
  AOI22xp33_ASAP7_75t_L     g13370(.A1(new_n1704), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1837), .Y(new_n13627));
  OAI221xp5_ASAP7_75t_L     g13371(.A1(new_n1699), .A2(new_n7616), .B1(new_n1827), .B2(new_n7906), .C(new_n13627), .Y(new_n13628));
  XNOR2x2_ASAP7_75t_L       g13372(.A(\a[23] ), .B(new_n13628), .Y(new_n13629));
  INVx1_ASAP7_75t_L         g13373(.A(new_n13460), .Y(new_n13630));
  MAJIxp5_ASAP7_75t_L       g13374(.A(new_n13557), .B(new_n13630), .C(new_n13461), .Y(new_n13631));
  XNOR2x2_ASAP7_75t_L       g13375(.A(new_n13629), .B(new_n13631), .Y(new_n13632));
  AOI22xp33_ASAP7_75t_L     g13376(.A1(new_n2114), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n2259), .Y(new_n13633));
  OAI221xp5_ASAP7_75t_L     g13377(.A1(new_n2109), .A2(new_n6830), .B1(new_n2257), .B2(new_n7323), .C(new_n13633), .Y(new_n13634));
  XNOR2x2_ASAP7_75t_L       g13378(.A(\a[26] ), .B(new_n13634), .Y(new_n13635));
  INVx1_ASAP7_75t_L         g13379(.A(new_n13635), .Y(new_n13636));
  MAJIxp5_ASAP7_75t_L       g13380(.A(new_n13556), .B(new_n13463), .C(new_n13467), .Y(new_n13637));
  NAND2xp33_ASAP7_75t_L     g13381(.A(new_n13636), .B(new_n13637), .Y(new_n13638));
  INVx1_ASAP7_75t_L         g13382(.A(new_n13638), .Y(new_n13639));
  NOR2xp33_ASAP7_75t_L      g13383(.A(new_n13636), .B(new_n13637), .Y(new_n13640));
  MAJIxp5_ASAP7_75t_L       g13384(.A(new_n13555), .B(new_n13472), .C(new_n13469), .Y(new_n13641));
  NAND2xp33_ASAP7_75t_L     g13385(.A(\b[45] ), .B(new_n2553), .Y(new_n13642));
  OAI221xp5_ASAP7_75t_L     g13386(.A1(new_n2545), .A2(new_n6568), .B1(new_n5829), .B2(new_n2747), .C(new_n13642), .Y(new_n13643));
  AOI21xp33_ASAP7_75t_L     g13387(.A1(new_n7919), .A2(new_n2544), .B(new_n13643), .Y(new_n13644));
  NAND2xp33_ASAP7_75t_L     g13388(.A(\a[29] ), .B(new_n13644), .Y(new_n13645));
  A2O1A1Ixp33_ASAP7_75t_L   g13389(.A1(new_n7919), .A2(new_n2544), .B(new_n13643), .C(new_n2538), .Y(new_n13646));
  NAND2xp33_ASAP7_75t_L     g13390(.A(new_n13646), .B(new_n13645), .Y(new_n13647));
  XNOR2x2_ASAP7_75t_L       g13391(.A(new_n13647), .B(new_n13641), .Y(new_n13648));
  AOI22xp33_ASAP7_75t_L     g13392(.A1(new_n3029), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n3258), .Y(new_n13649));
  OAI221xp5_ASAP7_75t_L     g13393(.A1(new_n3024), .A2(new_n5338), .B1(new_n3256), .B2(new_n6338), .C(new_n13649), .Y(new_n13650));
  XNOR2x2_ASAP7_75t_L       g13394(.A(\a[32] ), .B(new_n13650), .Y(new_n13651));
  MAJIxp5_ASAP7_75t_L       g13395(.A(new_n13554), .B(new_n13548), .C(new_n13552), .Y(new_n13652));
  NAND2xp33_ASAP7_75t_L     g13396(.A(new_n13651), .B(new_n13652), .Y(new_n13653));
  O2A1O1Ixp33_ASAP7_75t_L   g13397(.A1(new_n13353), .A2(new_n13356), .B(new_n13352), .C(new_n13553), .Y(new_n13654));
  INVx1_ASAP7_75t_L         g13398(.A(new_n13651), .Y(new_n13655));
  A2O1A1Ixp33_ASAP7_75t_L   g13399(.A1(new_n13552), .A2(new_n13548), .B(new_n13654), .C(new_n13655), .Y(new_n13656));
  NAND2xp33_ASAP7_75t_L     g13400(.A(new_n13653), .B(new_n13656), .Y(new_n13657));
  AOI22xp33_ASAP7_75t_L     g13401(.A1(new_n3633), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n3858), .Y(new_n13658));
  OAI221xp5_ASAP7_75t_L     g13402(.A1(new_n3853), .A2(new_n4848), .B1(new_n3856), .B2(new_n11686), .C(new_n13658), .Y(new_n13659));
  XNOR2x2_ASAP7_75t_L       g13403(.A(\a[35] ), .B(new_n13659), .Y(new_n13660));
  MAJIxp5_ASAP7_75t_L       g13404(.A(new_n13547), .B(new_n13476), .C(new_n13545), .Y(new_n13661));
  AOI22xp33_ASAP7_75t_L     g13405(.A1(new_n4283), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n4512), .Y(new_n13662));
  OAI221xp5_ASAP7_75t_L     g13406(.A1(new_n4277), .A2(new_n4216), .B1(new_n4499), .B2(new_n4431), .C(new_n13662), .Y(new_n13663));
  XNOR2x2_ASAP7_75t_L       g13407(.A(\a[38] ), .B(new_n13663), .Y(new_n13664));
  INVx1_ASAP7_75t_L         g13408(.A(new_n13543), .Y(new_n13665));
  NAND2xp33_ASAP7_75t_L     g13409(.A(new_n13477), .B(new_n13544), .Y(new_n13666));
  OAI21xp33_ASAP7_75t_L     g13410(.A1(new_n13480), .A2(new_n13665), .B(new_n13666), .Y(new_n13667));
  AOI22xp33_ASAP7_75t_L     g13411(.A1(new_n4920), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n5167), .Y(new_n13668));
  OAI221xp5_ASAP7_75t_L     g13412(.A1(new_n5154), .A2(new_n3565), .B1(new_n5158), .B2(new_n3591), .C(new_n13668), .Y(new_n13669));
  XNOR2x2_ASAP7_75t_L       g13413(.A(\a[41] ), .B(new_n13669), .Y(new_n13670));
  AOI22xp33_ASAP7_75t_L     g13414(.A1(new_n9700), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n10027), .Y(new_n13671));
  OAI221xp5_ASAP7_75t_L     g13415(.A1(new_n10024), .A2(new_n942), .B1(new_n9696), .B2(new_n1035), .C(new_n13671), .Y(new_n13672));
  XNOR2x2_ASAP7_75t_L       g13416(.A(\a[59] ), .B(new_n13672), .Y(new_n13673));
  AOI22xp33_ASAP7_75t_L     g13417(.A1(\b[11] ), .A2(new_n10939), .B1(\b[13] ), .B2(new_n10938), .Y(new_n13674));
  OAI21xp33_ASAP7_75t_L     g13418(.A1(new_n10629), .A2(new_n790), .B(new_n13674), .Y(new_n13675));
  AOI21xp33_ASAP7_75t_L     g13419(.A1(new_n10632), .A2(\b[12] ), .B(new_n13675), .Y(new_n13676));
  NAND2xp33_ASAP7_75t_L     g13420(.A(\a[62] ), .B(new_n13676), .Y(new_n13677));
  A2O1A1Ixp33_ASAP7_75t_L   g13421(.A1(\b[12] ), .A2(new_n10632), .B(new_n13675), .C(new_n10622), .Y(new_n13678));
  NAND2xp33_ASAP7_75t_L     g13422(.A(new_n13678), .B(new_n13677), .Y(new_n13679));
  NOR2xp33_ASAP7_75t_L      g13423(.A(new_n540), .B(new_n11535), .Y(new_n13680));
  O2A1O1Ixp33_ASAP7_75t_L   g13424(.A1(new_n11247), .A2(new_n11249), .B(\b[10] ), .C(new_n13680), .Y(new_n13681));
  INVx1_ASAP7_75t_L         g13425(.A(new_n13494), .Y(new_n13682));
  O2A1O1Ixp33_ASAP7_75t_L   g13426(.A1(new_n488), .A2(new_n11253), .B(new_n13276), .C(\a[8] ), .Y(new_n13683));
  O2A1O1Ixp33_ASAP7_75t_L   g13427(.A1(new_n13490), .A2(new_n13489), .B(new_n13682), .C(new_n13683), .Y(new_n13684));
  NAND2xp33_ASAP7_75t_L     g13428(.A(new_n13681), .B(new_n13684), .Y(new_n13685));
  INVx1_ASAP7_75t_L         g13429(.A(new_n13681), .Y(new_n13686));
  A2O1A1Ixp33_ASAP7_75t_L   g13430(.A1(new_n13492), .A2(new_n13682), .B(new_n13683), .C(new_n13686), .Y(new_n13687));
  AND2x2_ASAP7_75t_L        g13431(.A(new_n13685), .B(new_n13687), .Y(new_n13688));
  XNOR2x2_ASAP7_75t_L       g13432(.A(new_n13688), .B(new_n13679), .Y(new_n13689));
  NAND3xp33_ASAP7_75t_L     g13433(.A(new_n13689), .B(new_n13500), .C(new_n13499), .Y(new_n13690));
  A2O1A1Ixp33_ASAP7_75t_L   g13434(.A1(new_n13104), .A2(new_n13095), .B(new_n13277), .C(new_n13279), .Y(new_n13691));
  O2A1O1Ixp33_ASAP7_75t_L   g13435(.A1(new_n13496), .A2(new_n13691), .B(new_n13500), .C(new_n13689), .Y(new_n13692));
  INVx1_ASAP7_75t_L         g13436(.A(new_n13692), .Y(new_n13693));
  NAND3xp33_ASAP7_75t_L     g13437(.A(new_n13693), .B(new_n13690), .C(new_n13673), .Y(new_n13694));
  AO21x2_ASAP7_75t_L        g13438(.A1(new_n13690), .A2(new_n13693), .B(new_n13673), .Y(new_n13695));
  NAND4xp25_ASAP7_75t_L     g13439(.A(new_n13695), .B(new_n13506), .C(new_n13508), .D(new_n13694), .Y(new_n13696));
  INVx1_ASAP7_75t_L         g13440(.A(new_n13508), .Y(new_n13697));
  NAND2xp33_ASAP7_75t_L     g13441(.A(new_n13694), .B(new_n13695), .Y(new_n13698));
  A2O1A1Ixp33_ASAP7_75t_L   g13442(.A1(new_n13505), .A2(new_n13502), .B(new_n13697), .C(new_n13698), .Y(new_n13699));
  NAND2xp33_ASAP7_75t_L     g13443(.A(\b[17] ), .B(new_n9115), .Y(new_n13700));
  OAI221xp5_ASAP7_75t_L     g13444(.A1(new_n9113), .A2(new_n1432), .B1(new_n10016), .B2(new_n1438), .C(new_n13700), .Y(new_n13701));
  AOI21xp33_ASAP7_75t_L     g13445(.A1(new_n8835), .A2(\b[18] ), .B(new_n13701), .Y(new_n13702));
  NAND2xp33_ASAP7_75t_L     g13446(.A(\a[56] ), .B(new_n13702), .Y(new_n13703));
  A2O1A1Ixp33_ASAP7_75t_L   g13447(.A1(\b[18] ), .A2(new_n8835), .B(new_n13701), .C(new_n8826), .Y(new_n13704));
  AND2x2_ASAP7_75t_L        g13448(.A(new_n13704), .B(new_n13703), .Y(new_n13705));
  NAND3xp33_ASAP7_75t_L     g13449(.A(new_n13699), .B(new_n13696), .C(new_n13705), .Y(new_n13706));
  AO21x2_ASAP7_75t_L        g13450(.A1(new_n13696), .A2(new_n13699), .B(new_n13705), .Y(new_n13707));
  NAND2xp33_ASAP7_75t_L     g13451(.A(new_n13706), .B(new_n13707), .Y(new_n13708));
  OAI21xp33_ASAP7_75t_L     g13452(.A1(new_n13512), .A2(new_n13515), .B(new_n13518), .Y(new_n13709));
  NOR2xp33_ASAP7_75t_L      g13453(.A(new_n13708), .B(new_n13709), .Y(new_n13710));
  INVx1_ASAP7_75t_L         g13454(.A(new_n13710), .Y(new_n13711));
  NAND2xp33_ASAP7_75t_L     g13455(.A(new_n13708), .B(new_n13709), .Y(new_n13712));
  AOI22xp33_ASAP7_75t_L     g13456(.A1(new_n7960), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n8537), .Y(new_n13713));
  OAI221xp5_ASAP7_75t_L     g13457(.A1(new_n8817), .A2(new_n1655), .B1(new_n7957), .B2(new_n1780), .C(new_n13713), .Y(new_n13714));
  XNOR2x2_ASAP7_75t_L       g13458(.A(\a[53] ), .B(new_n13714), .Y(new_n13715));
  AND3x1_ASAP7_75t_L        g13459(.A(new_n13711), .B(new_n13715), .C(new_n13712), .Y(new_n13716));
  INVx1_ASAP7_75t_L         g13460(.A(new_n13716), .Y(new_n13717));
  AO21x2_ASAP7_75t_L        g13461(.A1(new_n13712), .A2(new_n13711), .B(new_n13715), .Y(new_n13718));
  AND2x2_ASAP7_75t_L        g13462(.A(new_n13718), .B(new_n13717), .Y(new_n13719));
  INVx1_ASAP7_75t_L         g13463(.A(new_n13524), .Y(new_n13720));
  OA21x2_ASAP7_75t_L        g13464(.A1(new_n13519), .A2(new_n13522), .B(new_n13720), .Y(new_n13721));
  AND2x2_ASAP7_75t_L        g13465(.A(new_n13719), .B(new_n13721), .Y(new_n13722));
  INVx1_ASAP7_75t_L         g13466(.A(new_n13722), .Y(new_n13723));
  O2A1O1Ixp33_ASAP7_75t_L   g13467(.A1(new_n13519), .A2(new_n13522), .B(new_n13720), .C(new_n13719), .Y(new_n13724));
  INVx1_ASAP7_75t_L         g13468(.A(new_n13724), .Y(new_n13725));
  AOI22xp33_ASAP7_75t_L     g13469(.A1(new_n7111), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n7391), .Y(new_n13726));
  OAI221xp5_ASAP7_75t_L     g13470(.A1(new_n8558), .A2(new_n1929), .B1(new_n8237), .B2(new_n2075), .C(new_n13726), .Y(new_n13727));
  XNOR2x2_ASAP7_75t_L       g13471(.A(\a[50] ), .B(new_n13727), .Y(new_n13728));
  NAND3xp33_ASAP7_75t_L     g13472(.A(new_n13723), .B(new_n13725), .C(new_n13728), .Y(new_n13729));
  AO21x2_ASAP7_75t_L        g13473(.A1(new_n13725), .A2(new_n13723), .B(new_n13728), .Y(new_n13730));
  INVx1_ASAP7_75t_L         g13474(.A(new_n13529), .Y(new_n13731));
  NOR3xp33_ASAP7_75t_L      g13475(.A(new_n13525), .B(new_n13524), .C(new_n13484), .Y(new_n13732));
  A2O1A1O1Ixp25_ASAP7_75t_L g13476(.A1(new_n13265), .A2(new_n13312), .B(new_n13731), .C(new_n13527), .D(new_n13732), .Y(new_n13733));
  AND3x1_ASAP7_75t_L        g13477(.A(new_n13730), .B(new_n13733), .C(new_n13729), .Y(new_n13734));
  AOI21xp33_ASAP7_75t_L     g13478(.A1(new_n13730), .A2(new_n13729), .B(new_n13733), .Y(new_n13735));
  NOR2xp33_ASAP7_75t_L      g13479(.A(new_n13735), .B(new_n13734), .Y(new_n13736));
  AOI22xp33_ASAP7_75t_L     g13480(.A1(new_n6376), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n6648), .Y(new_n13737));
  OAI221xp5_ASAP7_75t_L     g13481(.A1(new_n6646), .A2(new_n2497), .B1(new_n6636), .B2(new_n2672), .C(new_n13737), .Y(new_n13738));
  XNOR2x2_ASAP7_75t_L       g13482(.A(\a[47] ), .B(new_n13738), .Y(new_n13739));
  XNOR2x2_ASAP7_75t_L       g13483(.A(new_n13739), .B(new_n13736), .Y(new_n13740));
  NOR2xp33_ASAP7_75t_L      g13484(.A(new_n13534), .B(new_n13531), .Y(new_n13741));
  NOR2xp33_ASAP7_75t_L      g13485(.A(new_n13536), .B(new_n13535), .Y(new_n13742));
  NOR2xp33_ASAP7_75t_L      g13486(.A(new_n13741), .B(new_n13742), .Y(new_n13743));
  XOR2x2_ASAP7_75t_L        g13487(.A(new_n13740), .B(new_n13743), .Y(new_n13744));
  AOI22xp33_ASAP7_75t_L     g13488(.A1(new_n5624), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n5901), .Y(new_n13745));
  OAI221xp5_ASAP7_75t_L     g13489(.A1(new_n5900), .A2(new_n2982), .B1(new_n5892), .B2(new_n3187), .C(new_n13745), .Y(new_n13746));
  XNOR2x2_ASAP7_75t_L       g13490(.A(\a[44] ), .B(new_n13746), .Y(new_n13747));
  XNOR2x2_ASAP7_75t_L       g13491(.A(new_n13747), .B(new_n13744), .Y(new_n13748));
  MAJx2_ASAP7_75t_L         g13492(.A(new_n13542), .B(new_n13540), .C(new_n13537), .Y(new_n13749));
  XNOR2x2_ASAP7_75t_L       g13493(.A(new_n13749), .B(new_n13748), .Y(new_n13750));
  XNOR2x2_ASAP7_75t_L       g13494(.A(new_n13670), .B(new_n13750), .Y(new_n13751));
  XNOR2x2_ASAP7_75t_L       g13495(.A(new_n13751), .B(new_n13667), .Y(new_n13752));
  XNOR2x2_ASAP7_75t_L       g13496(.A(new_n13664), .B(new_n13752), .Y(new_n13753));
  XOR2x2_ASAP7_75t_L        g13497(.A(new_n13661), .B(new_n13753), .Y(new_n13754));
  XNOR2x2_ASAP7_75t_L       g13498(.A(new_n13660), .B(new_n13754), .Y(new_n13755));
  XNOR2x2_ASAP7_75t_L       g13499(.A(new_n13755), .B(new_n13657), .Y(new_n13756));
  XNOR2x2_ASAP7_75t_L       g13500(.A(new_n13756), .B(new_n13648), .Y(new_n13757));
  OA21x2_ASAP7_75t_L        g13501(.A1(new_n13640), .A2(new_n13639), .B(new_n13757), .Y(new_n13758));
  NOR3xp33_ASAP7_75t_L      g13502(.A(new_n13639), .B(new_n13640), .C(new_n13757), .Y(new_n13759));
  NOR3xp33_ASAP7_75t_L      g13503(.A(new_n13632), .B(new_n13758), .C(new_n13759), .Y(new_n13760));
  OA21x2_ASAP7_75t_L        g13504(.A1(new_n13758), .A2(new_n13759), .B(new_n13632), .Y(new_n13761));
  NOR2xp33_ASAP7_75t_L      g13505(.A(new_n13760), .B(new_n13761), .Y(new_n13762));
  XNOR2x2_ASAP7_75t_L       g13506(.A(new_n13762), .B(new_n13626), .Y(new_n13763));
  NAND3xp33_ASAP7_75t_L     g13507(.A(new_n13763), .B(new_n13617), .C(new_n13620), .Y(new_n13764));
  O2A1O1Ixp33_ASAP7_75t_L   g13508(.A1(new_n13565), .A2(new_n13446), .B(new_n13562), .C(new_n13619), .Y(new_n13765));
  AOI211xp5_ASAP7_75t_L     g13509(.A1(new_n13609), .A2(new_n13561), .B(new_n13610), .C(new_n13616), .Y(new_n13766));
  INVx1_ASAP7_75t_L         g13510(.A(new_n13457), .Y(new_n13767));
  A2O1A1Ixp33_ASAP7_75t_L   g13511(.A1(new_n13456), .A2(new_n13558), .B(new_n13767), .C(new_n13623), .Y(new_n13768));
  OR2x4_ASAP7_75t_L         g13512(.A(new_n13623), .B(new_n13625), .Y(new_n13769));
  NAND3xp33_ASAP7_75t_L     g13513(.A(new_n13762), .B(new_n13769), .C(new_n13768), .Y(new_n13770));
  OAI21xp33_ASAP7_75t_L     g13514(.A1(new_n13760), .A2(new_n13761), .B(new_n13626), .Y(new_n13771));
  NAND2xp33_ASAP7_75t_L     g13515(.A(new_n13770), .B(new_n13771), .Y(new_n13772));
  OAI21xp33_ASAP7_75t_L     g13516(.A1(new_n13765), .A2(new_n13766), .B(new_n13772), .Y(new_n13773));
  NAND2xp33_ASAP7_75t_L     g13517(.A(new_n13764), .B(new_n13773), .Y(new_n13774));
  OAI21xp33_ASAP7_75t_L     g13518(.A1(new_n13608), .A2(new_n13607), .B(new_n13774), .Y(new_n13775));
  INVx1_ASAP7_75t_L         g13519(.A(new_n13608), .Y(new_n13776));
  AND2x2_ASAP7_75t_L        g13520(.A(new_n13764), .B(new_n13773), .Y(new_n13777));
  NAND3xp33_ASAP7_75t_L     g13521(.A(new_n13777), .B(new_n13776), .C(new_n13606), .Y(new_n13778));
  NAND2xp33_ASAP7_75t_L     g13522(.A(new_n13775), .B(new_n13778), .Y(new_n13779));
  AOI21xp33_ASAP7_75t_L     g13523(.A1(new_n13597), .A2(new_n13599), .B(new_n13779), .Y(new_n13780));
  INVx1_ASAP7_75t_L         g13524(.A(new_n13597), .Y(new_n13781));
  AOI211xp5_ASAP7_75t_L     g13525(.A1(new_n13775), .A2(new_n13778), .B(new_n13598), .C(new_n13781), .Y(new_n13782));
  NOR3xp33_ASAP7_75t_L      g13526(.A(new_n13780), .B(new_n13782), .C(new_n13589), .Y(new_n13783));
  OA21x2_ASAP7_75t_L        g13527(.A1(new_n13782), .A2(new_n13780), .B(new_n13589), .Y(new_n13784));
  NOR2xp33_ASAP7_75t_L      g13528(.A(new_n13783), .B(new_n13784), .Y(new_n13785));
  A2O1A1Ixp33_ASAP7_75t_L   g13529(.A1(new_n13584), .A2(new_n13579), .B(new_n13587), .C(new_n13785), .Y(new_n13786));
  INVx1_ASAP7_75t_L         g13530(.A(new_n13786), .Y(new_n13787));
  NAND2xp33_ASAP7_75t_L     g13531(.A(new_n13575), .B(new_n13578), .Y(new_n13788));
  A2O1A1Ixp33_ASAP7_75t_L   g13532(.A1(new_n13413), .A2(new_n13583), .B(new_n13788), .C(new_n13575), .Y(new_n13789));
  NOR2xp33_ASAP7_75t_L      g13533(.A(new_n13785), .B(new_n13789), .Y(new_n13790));
  NOR2xp33_ASAP7_75t_L      g13534(.A(new_n13790), .B(new_n13787), .Y(\f[73] ));
  INVx1_ASAP7_75t_L         g13535(.A(new_n13596), .Y(new_n13792));
  A2O1A1Ixp33_ASAP7_75t_L   g13536(.A1(new_n13569), .A2(new_n13434), .B(new_n13590), .C(new_n13792), .Y(new_n13793));
  A2O1A1Ixp33_ASAP7_75t_L   g13537(.A1(new_n13599), .A2(new_n13597), .B(new_n13779), .C(new_n13793), .Y(new_n13794));
  O2A1O1Ixp33_ASAP7_75t_L   g13538(.A1(new_n13565), .A2(new_n13446), .B(new_n13562), .C(new_n13616), .Y(new_n13795));
  INVx1_ASAP7_75t_L         g13539(.A(new_n13795), .Y(new_n13796));
  NAND2xp33_ASAP7_75t_L     g13540(.A(\b[61] ), .B(new_n815), .Y(new_n13797));
  OAI221xp5_ASAP7_75t_L     g13541(.A1(new_n977), .A2(new_n11172), .B1(new_n10250), .B2(new_n978), .C(new_n13797), .Y(new_n13798));
  AOI21xp33_ASAP7_75t_L     g13542(.A1(new_n11180), .A2(new_n808), .B(new_n13798), .Y(new_n13799));
  NAND2xp33_ASAP7_75t_L     g13543(.A(\a[14] ), .B(new_n13799), .Y(new_n13800));
  A2O1A1Ixp33_ASAP7_75t_L   g13544(.A1(new_n11180), .A2(new_n808), .B(new_n13798), .C(new_n806), .Y(new_n13801));
  AND2x2_ASAP7_75t_L        g13545(.A(new_n13801), .B(new_n13800), .Y(new_n13802));
  A2O1A1O1Ixp25_ASAP7_75t_L g13546(.A1(new_n13620), .A2(new_n13617), .B(new_n13772), .C(new_n13796), .D(new_n13802), .Y(new_n13803));
  INVx1_ASAP7_75t_L         g13547(.A(new_n13803), .Y(new_n13804));
  O2A1O1Ixp33_ASAP7_75t_L   g13548(.A1(new_n13765), .A2(new_n13766), .B(new_n13763), .C(new_n13795), .Y(new_n13805));
  NAND2xp33_ASAP7_75t_L     g13549(.A(new_n13802), .B(new_n13805), .Y(new_n13806));
  NAND2xp33_ASAP7_75t_L     g13550(.A(new_n13806), .B(new_n13804), .Y(new_n13807));
  AOI22xp33_ASAP7_75t_L     g13551(.A1(new_n1076), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1253), .Y(new_n13808));
  OAI221xp5_ASAP7_75t_L     g13552(.A1(new_n1154), .A2(new_n9920), .B1(new_n1156), .B2(new_n11152), .C(new_n13808), .Y(new_n13809));
  XNOR2x2_ASAP7_75t_L       g13553(.A(\a[17] ), .B(new_n13809), .Y(new_n13810));
  AND2x2_ASAP7_75t_L        g13554(.A(new_n13769), .B(new_n13770), .Y(new_n13811));
  NAND2xp33_ASAP7_75t_L     g13555(.A(new_n13810), .B(new_n13811), .Y(new_n13812));
  AO21x2_ASAP7_75t_L        g13556(.A1(new_n13769), .A2(new_n13770), .B(new_n13810), .Y(new_n13813));
  AOI22xp33_ASAP7_75t_L     g13557(.A1(new_n1360), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1581), .Y(new_n13814));
  OAI221xp5_ASAP7_75t_L     g13558(.A1(new_n1373), .A2(new_n8762), .B1(new_n1359), .B2(new_n9331), .C(new_n13814), .Y(new_n13815));
  XNOR2x2_ASAP7_75t_L       g13559(.A(\a[20] ), .B(new_n13815), .Y(new_n13816));
  NOR2xp33_ASAP7_75t_L      g13560(.A(new_n13629), .B(new_n13631), .Y(new_n13817));
  NOR2xp33_ASAP7_75t_L      g13561(.A(new_n13817), .B(new_n13760), .Y(new_n13818));
  XOR2x2_ASAP7_75t_L        g13562(.A(new_n13816), .B(new_n13818), .Y(new_n13819));
  INVx1_ASAP7_75t_L         g13563(.A(new_n13637), .Y(new_n13820));
  MAJx2_ASAP7_75t_L         g13564(.A(new_n13820), .B(new_n13636), .C(new_n13757), .Y(new_n13821));
  NOR2xp33_ASAP7_75t_L      g13565(.A(new_n8165), .B(new_n1696), .Y(new_n13822));
  AOI221xp5_ASAP7_75t_L     g13566(.A1(\b[51] ), .A2(new_n1837), .B1(\b[52] ), .B2(new_n1706), .C(new_n13822), .Y(new_n13823));
  OAI211xp5_ASAP7_75t_L     g13567(.A1(new_n1827), .A2(new_n8174), .B(\a[23] ), .C(new_n13823), .Y(new_n13824));
  INVx1_ASAP7_75t_L         g13568(.A(new_n13824), .Y(new_n13825));
  O2A1O1Ixp33_ASAP7_75t_L   g13569(.A1(new_n1827), .A2(new_n8174), .B(new_n13823), .C(\a[23] ), .Y(new_n13826));
  NOR2xp33_ASAP7_75t_L      g13570(.A(new_n13826), .B(new_n13825), .Y(new_n13827));
  INVx1_ASAP7_75t_L         g13571(.A(new_n13827), .Y(new_n13828));
  XNOR2x2_ASAP7_75t_L       g13572(.A(new_n13828), .B(new_n13821), .Y(new_n13829));
  MAJIxp5_ASAP7_75t_L       g13573(.A(new_n13756), .B(new_n13641), .C(new_n13647), .Y(new_n13830));
  NAND2xp33_ASAP7_75t_L     g13574(.A(\b[49] ), .B(new_n2115), .Y(new_n13831));
  OAI221xp5_ASAP7_75t_L     g13575(.A1(new_n2107), .A2(new_n7593), .B1(new_n6830), .B2(new_n2269), .C(new_n13831), .Y(new_n13832));
  AOI21xp33_ASAP7_75t_L     g13576(.A1(new_n7601), .A2(new_n2106), .B(new_n13832), .Y(new_n13833));
  NAND2xp33_ASAP7_75t_L     g13577(.A(\a[26] ), .B(new_n13833), .Y(new_n13834));
  A2O1A1Ixp33_ASAP7_75t_L   g13578(.A1(new_n7601), .A2(new_n2106), .B(new_n13832), .C(new_n2100), .Y(new_n13835));
  AND2x2_ASAP7_75t_L        g13579(.A(new_n13835), .B(new_n13834), .Y(new_n13836));
  NOR2xp33_ASAP7_75t_L      g13580(.A(new_n13836), .B(new_n13830), .Y(new_n13837));
  INVx1_ASAP7_75t_L         g13581(.A(new_n13837), .Y(new_n13838));
  NAND2xp33_ASAP7_75t_L     g13582(.A(new_n13836), .B(new_n13830), .Y(new_n13839));
  AND2x2_ASAP7_75t_L        g13583(.A(new_n13839), .B(new_n13838), .Y(new_n13840));
  AOI22xp33_ASAP7_75t_L     g13584(.A1(new_n2552), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n2736), .Y(new_n13841));
  OAI221xp5_ASAP7_75t_L     g13585(.A1(new_n2547), .A2(new_n6568), .B1(new_n2734), .B2(new_n6820), .C(new_n13841), .Y(new_n13842));
  XNOR2x2_ASAP7_75t_L       g13586(.A(\a[29] ), .B(new_n13842), .Y(new_n13843));
  NAND2xp33_ASAP7_75t_L     g13587(.A(new_n13653), .B(new_n13755), .Y(new_n13844));
  AND3x1_ASAP7_75t_L        g13588(.A(new_n13844), .B(new_n13843), .C(new_n13656), .Y(new_n13845));
  O2A1O1Ixp33_ASAP7_75t_L   g13589(.A1(new_n13652), .A2(new_n13651), .B(new_n13844), .C(new_n13843), .Y(new_n13846));
  NAND2xp33_ASAP7_75t_L     g13590(.A(new_n13660), .B(new_n13754), .Y(new_n13847));
  NOR2xp33_ASAP7_75t_L      g13591(.A(new_n5829), .B(new_n3022), .Y(new_n13848));
  AOI221xp5_ASAP7_75t_L     g13592(.A1(\b[42] ), .A2(new_n3258), .B1(\b[43] ), .B2(new_n3030), .C(new_n13848), .Y(new_n13849));
  OAI211xp5_ASAP7_75t_L     g13593(.A1(new_n3256), .A2(new_n5835), .B(\a[32] ), .C(new_n13849), .Y(new_n13850));
  O2A1O1Ixp33_ASAP7_75t_L   g13594(.A1(new_n3256), .A2(new_n5835), .B(new_n13849), .C(\a[32] ), .Y(new_n13851));
  INVx1_ASAP7_75t_L         g13595(.A(new_n13851), .Y(new_n13852));
  AND2x2_ASAP7_75t_L        g13596(.A(new_n13850), .B(new_n13852), .Y(new_n13853));
  INVx1_ASAP7_75t_L         g13597(.A(new_n13853), .Y(new_n13854));
  OA211x2_ASAP7_75t_L       g13598(.A1(new_n13661), .A2(new_n13753), .B(new_n13847), .C(new_n13854), .Y(new_n13855));
  O2A1O1Ixp33_ASAP7_75t_L   g13599(.A1(new_n13661), .A2(new_n13753), .B(new_n13847), .C(new_n13854), .Y(new_n13856));
  NOR2xp33_ASAP7_75t_L      g13600(.A(new_n13856), .B(new_n13855), .Y(new_n13857));
  AOI22xp33_ASAP7_75t_L     g13601(.A1(new_n3633), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n3858), .Y(new_n13858));
  OAI221xp5_ASAP7_75t_L     g13602(.A1(new_n3853), .A2(new_n4869), .B1(new_n3856), .B2(new_n5327), .C(new_n13858), .Y(new_n13859));
  XNOR2x2_ASAP7_75t_L       g13603(.A(\a[35] ), .B(new_n13859), .Y(new_n13860));
  INVx1_ASAP7_75t_L         g13604(.A(new_n13667), .Y(new_n13861));
  MAJIxp5_ASAP7_75t_L       g13605(.A(new_n13861), .B(new_n13664), .C(new_n13751), .Y(new_n13862));
  INVx1_ASAP7_75t_L         g13606(.A(new_n13862), .Y(new_n13863));
  INVx1_ASAP7_75t_L         g13607(.A(new_n13743), .Y(new_n13864));
  NOR2xp33_ASAP7_75t_L      g13608(.A(new_n13747), .B(new_n13744), .Y(new_n13865));
  AOI22xp33_ASAP7_75t_L     g13609(.A1(new_n7111), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n7391), .Y(new_n13866));
  OAI221xp5_ASAP7_75t_L     g13610(.A1(new_n8558), .A2(new_n2067), .B1(new_n8237), .B2(new_n2355), .C(new_n13866), .Y(new_n13867));
  XNOR2x2_ASAP7_75t_L       g13611(.A(\a[50] ), .B(new_n13867), .Y(new_n13868));
  INVx1_ASAP7_75t_L         g13612(.A(new_n13868), .Y(new_n13869));
  AOI22xp33_ASAP7_75t_L     g13613(.A1(new_n7960), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n8537), .Y(new_n13870));
  OAI221xp5_ASAP7_75t_L     g13614(.A1(new_n8817), .A2(new_n1774), .B1(new_n7957), .B2(new_n1915), .C(new_n13870), .Y(new_n13871));
  XNOR2x2_ASAP7_75t_L       g13615(.A(\a[53] ), .B(new_n13871), .Y(new_n13872));
  AOI22xp33_ASAP7_75t_L     g13616(.A1(new_n9700), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n10027), .Y(new_n13873));
  OAI221xp5_ASAP7_75t_L     g13617(.A1(new_n10024), .A2(new_n1030), .B1(new_n9696), .B2(new_n1209), .C(new_n13873), .Y(new_n13874));
  XNOR2x2_ASAP7_75t_L       g13618(.A(\a[59] ), .B(new_n13874), .Y(new_n13875));
  A2O1A1Ixp33_ASAP7_75t_L   g13619(.A1(new_n13492), .A2(new_n13682), .B(new_n13683), .C(new_n13681), .Y(new_n13876));
  A2O1A1Ixp33_ASAP7_75t_L   g13620(.A1(new_n13677), .A2(new_n13678), .B(new_n13688), .C(new_n13876), .Y(new_n13877));
  NOR2xp33_ASAP7_75t_L      g13621(.A(new_n617), .B(new_n11535), .Y(new_n13878));
  O2A1O1Ixp33_ASAP7_75t_L   g13622(.A1(new_n11247), .A2(new_n11249), .B(\b[11] ), .C(new_n13878), .Y(new_n13879));
  NAND2xp33_ASAP7_75t_L     g13623(.A(new_n13879), .B(new_n13681), .Y(new_n13880));
  A2O1A1Ixp33_ASAP7_75t_L   g13624(.A1(\b[11] ), .A2(new_n11533), .B(new_n13878), .C(new_n13686), .Y(new_n13881));
  AND2x2_ASAP7_75t_L        g13625(.A(new_n13880), .B(new_n13881), .Y(new_n13882));
  XNOR2x2_ASAP7_75t_L       g13626(.A(new_n13882), .B(new_n13877), .Y(new_n13883));
  AOI22xp33_ASAP7_75t_L     g13627(.A1(\b[12] ), .A2(new_n10939), .B1(\b[14] ), .B2(new_n10938), .Y(new_n13884));
  OAI221xp5_ASAP7_75t_L     g13628(.A1(new_n10937), .A2(new_n784), .B1(new_n10629), .B2(new_n875), .C(new_n13884), .Y(new_n13885));
  XNOR2x2_ASAP7_75t_L       g13629(.A(\a[62] ), .B(new_n13885), .Y(new_n13886));
  INVx1_ASAP7_75t_L         g13630(.A(new_n13886), .Y(new_n13887));
  NAND2xp33_ASAP7_75t_L     g13631(.A(new_n13887), .B(new_n13883), .Y(new_n13888));
  INVx1_ASAP7_75t_L         g13632(.A(new_n13883), .Y(new_n13889));
  NAND2xp33_ASAP7_75t_L     g13633(.A(new_n13886), .B(new_n13889), .Y(new_n13890));
  NAND3xp33_ASAP7_75t_L     g13634(.A(new_n13890), .B(new_n13875), .C(new_n13888), .Y(new_n13891));
  AO21x2_ASAP7_75t_L        g13635(.A1(new_n13888), .A2(new_n13890), .B(new_n13875), .Y(new_n13892));
  AND2x2_ASAP7_75t_L        g13636(.A(new_n13891), .B(new_n13892), .Y(new_n13893));
  A2O1A1Ixp33_ASAP7_75t_L   g13637(.A1(new_n13690), .A2(new_n13673), .B(new_n13692), .C(new_n13893), .Y(new_n13894));
  A2O1A1Ixp33_ASAP7_75t_L   g13638(.A1(new_n13500), .A2(new_n13499), .B(new_n13689), .C(new_n13694), .Y(new_n13895));
  NOR2xp33_ASAP7_75t_L      g13639(.A(new_n13895), .B(new_n13893), .Y(new_n13896));
  INVx1_ASAP7_75t_L         g13640(.A(new_n13896), .Y(new_n13897));
  NAND2xp33_ASAP7_75t_L     g13641(.A(new_n13894), .B(new_n13897), .Y(new_n13898));
  AOI22xp33_ASAP7_75t_L     g13642(.A1(new_n8831), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n9115), .Y(new_n13899));
  OAI221xp5_ASAP7_75t_L     g13643(.A1(new_n10343), .A2(new_n1432), .B1(new_n10016), .B2(new_n1547), .C(new_n13899), .Y(new_n13900));
  XNOR2x2_ASAP7_75t_L       g13644(.A(\a[56] ), .B(new_n13900), .Y(new_n13901));
  NAND2xp33_ASAP7_75t_L     g13645(.A(new_n13901), .B(new_n13898), .Y(new_n13902));
  NOR2xp33_ASAP7_75t_L      g13646(.A(new_n13901), .B(new_n13898), .Y(new_n13903));
  INVx1_ASAP7_75t_L         g13647(.A(new_n13903), .Y(new_n13904));
  NAND2xp33_ASAP7_75t_L     g13648(.A(new_n13904), .B(new_n13902), .Y(new_n13905));
  NAND2xp33_ASAP7_75t_L     g13649(.A(new_n13696), .B(new_n13706), .Y(new_n13906));
  NOR2xp33_ASAP7_75t_L      g13650(.A(new_n13906), .B(new_n13905), .Y(new_n13907));
  AOI22xp33_ASAP7_75t_L     g13651(.A1(new_n13696), .A2(new_n13706), .B1(new_n13902), .B2(new_n13904), .Y(new_n13908));
  NOR3xp33_ASAP7_75t_L      g13652(.A(new_n13907), .B(new_n13908), .C(new_n13872), .Y(new_n13909));
  INVx1_ASAP7_75t_L         g13653(.A(new_n13909), .Y(new_n13910));
  OAI21xp33_ASAP7_75t_L     g13654(.A1(new_n13908), .A2(new_n13907), .B(new_n13872), .Y(new_n13911));
  NAND2xp33_ASAP7_75t_L     g13655(.A(new_n13911), .B(new_n13910), .Y(new_n13912));
  NOR3xp33_ASAP7_75t_L      g13656(.A(new_n13912), .B(new_n13716), .C(new_n13710), .Y(new_n13913));
  A2O1A1Ixp33_ASAP7_75t_L   g13657(.A1(new_n13712), .A2(new_n13715), .B(new_n13710), .C(new_n13912), .Y(new_n13914));
  INVx1_ASAP7_75t_L         g13658(.A(new_n13914), .Y(new_n13915));
  NOR2xp33_ASAP7_75t_L      g13659(.A(new_n13913), .B(new_n13915), .Y(new_n13916));
  NAND2xp33_ASAP7_75t_L     g13660(.A(new_n13869), .B(new_n13916), .Y(new_n13917));
  OAI21xp33_ASAP7_75t_L     g13661(.A1(new_n13913), .A2(new_n13915), .B(new_n13868), .Y(new_n13918));
  NAND2xp33_ASAP7_75t_L     g13662(.A(new_n13918), .B(new_n13917), .Y(new_n13919));
  AOI21xp33_ASAP7_75t_L     g13663(.A1(new_n13725), .A2(new_n13728), .B(new_n13722), .Y(new_n13920));
  XNOR2x2_ASAP7_75t_L       g13664(.A(new_n13920), .B(new_n13919), .Y(new_n13921));
  AOI22xp33_ASAP7_75t_L     g13665(.A1(new_n6376), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n6648), .Y(new_n13922));
  OAI221xp5_ASAP7_75t_L     g13666(.A1(new_n6646), .A2(new_n2666), .B1(new_n6636), .B2(new_n2695), .C(new_n13922), .Y(new_n13923));
  XNOR2x2_ASAP7_75t_L       g13667(.A(\a[47] ), .B(new_n13923), .Y(new_n13924));
  XOR2x2_ASAP7_75t_L        g13668(.A(new_n13924), .B(new_n13921), .Y(new_n13925));
  AOI21xp33_ASAP7_75t_L     g13669(.A1(new_n13736), .A2(new_n13739), .B(new_n13734), .Y(new_n13926));
  XNOR2x2_ASAP7_75t_L       g13670(.A(new_n13926), .B(new_n13925), .Y(new_n13927));
  AOI22xp33_ASAP7_75t_L     g13671(.A1(new_n5624), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n5901), .Y(new_n13928));
  OAI221xp5_ASAP7_75t_L     g13672(.A1(new_n5900), .A2(new_n3180), .B1(new_n5892), .B2(new_n11047), .C(new_n13928), .Y(new_n13929));
  XNOR2x2_ASAP7_75t_L       g13673(.A(\a[44] ), .B(new_n13929), .Y(new_n13930));
  XNOR2x2_ASAP7_75t_L       g13674(.A(new_n13930), .B(new_n13927), .Y(new_n13931));
  A2O1A1Ixp33_ASAP7_75t_L   g13675(.A1(new_n13864), .A2(new_n13740), .B(new_n13865), .C(new_n13931), .Y(new_n13932));
  AND2x2_ASAP7_75t_L        g13676(.A(new_n13740), .B(new_n13864), .Y(new_n13933));
  OR3x1_ASAP7_75t_L         g13677(.A(new_n13931), .B(new_n13933), .C(new_n13865), .Y(new_n13934));
  AOI22xp33_ASAP7_75t_L     g13678(.A1(new_n4920), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n5167), .Y(new_n13935));
  OAI221xp5_ASAP7_75t_L     g13679(.A1(new_n5154), .A2(new_n3584), .B1(new_n5158), .B2(new_n10137), .C(new_n13935), .Y(new_n13936));
  XNOR2x2_ASAP7_75t_L       g13680(.A(\a[41] ), .B(new_n13936), .Y(new_n13937));
  NAND3xp33_ASAP7_75t_L     g13681(.A(new_n13932), .B(new_n13934), .C(new_n13937), .Y(new_n13938));
  AO21x2_ASAP7_75t_L        g13682(.A1(new_n13932), .A2(new_n13934), .B(new_n13937), .Y(new_n13939));
  NAND2xp33_ASAP7_75t_L     g13683(.A(new_n13938), .B(new_n13939), .Y(new_n13940));
  MAJIxp5_ASAP7_75t_L       g13684(.A(new_n13748), .B(new_n13670), .C(new_n13749), .Y(new_n13941));
  INVx1_ASAP7_75t_L         g13685(.A(new_n13941), .Y(new_n13942));
  XNOR2x2_ASAP7_75t_L       g13686(.A(new_n13942), .B(new_n13940), .Y(new_n13943));
  AOI22xp33_ASAP7_75t_L     g13687(.A1(new_n4283), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n4512), .Y(new_n13944));
  OAI221xp5_ASAP7_75t_L     g13688(.A1(new_n4277), .A2(new_n4424), .B1(new_n4499), .B2(new_n4641), .C(new_n13944), .Y(new_n13945));
  XNOR2x2_ASAP7_75t_L       g13689(.A(\a[38] ), .B(new_n13945), .Y(new_n13946));
  INVx1_ASAP7_75t_L         g13690(.A(new_n13946), .Y(new_n13947));
  XNOR2x2_ASAP7_75t_L       g13691(.A(new_n13947), .B(new_n13943), .Y(new_n13948));
  NOR2xp33_ASAP7_75t_L      g13692(.A(new_n13863), .B(new_n13948), .Y(new_n13949));
  NAND2xp33_ASAP7_75t_L     g13693(.A(new_n13863), .B(new_n13948), .Y(new_n13950));
  INVx1_ASAP7_75t_L         g13694(.A(new_n13950), .Y(new_n13951));
  NOR2xp33_ASAP7_75t_L      g13695(.A(new_n13949), .B(new_n13951), .Y(new_n13952));
  NOR2xp33_ASAP7_75t_L      g13696(.A(new_n13860), .B(new_n13952), .Y(new_n13953));
  AND2x2_ASAP7_75t_L        g13697(.A(new_n13860), .B(new_n13952), .Y(new_n13954));
  NOR2xp33_ASAP7_75t_L      g13698(.A(new_n13953), .B(new_n13954), .Y(new_n13955));
  NAND2xp33_ASAP7_75t_L     g13699(.A(new_n13857), .B(new_n13955), .Y(new_n13956));
  OAI22xp33_ASAP7_75t_L     g13700(.A1(new_n13954), .A2(new_n13953), .B1(new_n13856), .B2(new_n13855), .Y(new_n13957));
  AND2x2_ASAP7_75t_L        g13701(.A(new_n13957), .B(new_n13956), .Y(new_n13958));
  OR3x1_ASAP7_75t_L         g13702(.A(new_n13958), .B(new_n13845), .C(new_n13846), .Y(new_n13959));
  OAI21xp33_ASAP7_75t_L     g13703(.A1(new_n13845), .A2(new_n13846), .B(new_n13958), .Y(new_n13960));
  NAND2xp33_ASAP7_75t_L     g13704(.A(new_n13960), .B(new_n13959), .Y(new_n13961));
  INVx1_ASAP7_75t_L         g13705(.A(new_n13961), .Y(new_n13962));
  NAND2xp33_ASAP7_75t_L     g13706(.A(new_n13962), .B(new_n13840), .Y(new_n13963));
  NAND2xp33_ASAP7_75t_L     g13707(.A(new_n13839), .B(new_n13838), .Y(new_n13964));
  NAND2xp33_ASAP7_75t_L     g13708(.A(new_n13961), .B(new_n13964), .Y(new_n13965));
  NAND2xp33_ASAP7_75t_L     g13709(.A(new_n13965), .B(new_n13963), .Y(new_n13966));
  XNOR2x2_ASAP7_75t_L       g13710(.A(new_n13829), .B(new_n13966), .Y(new_n13967));
  XNOR2x2_ASAP7_75t_L       g13711(.A(new_n13967), .B(new_n13819), .Y(new_n13968));
  NAND3xp33_ASAP7_75t_L     g13712(.A(new_n13968), .B(new_n13813), .C(new_n13812), .Y(new_n13969));
  AO21x2_ASAP7_75t_L        g13713(.A1(new_n13812), .A2(new_n13813), .B(new_n13968), .Y(new_n13970));
  NAND2xp33_ASAP7_75t_L     g13714(.A(new_n13969), .B(new_n13970), .Y(new_n13971));
  INVx1_ASAP7_75t_L         g13715(.A(new_n13971), .Y(new_n13972));
  NOR2xp33_ASAP7_75t_L      g13716(.A(new_n13807), .B(new_n13972), .Y(new_n13973));
  INVx1_ASAP7_75t_L         g13717(.A(new_n13807), .Y(new_n13974));
  NOR2xp33_ASAP7_75t_L      g13718(.A(new_n13971), .B(new_n13974), .Y(new_n13975));
  NAND2xp33_ASAP7_75t_L     g13719(.A(new_n13606), .B(new_n13776), .Y(new_n13976));
  INVx1_ASAP7_75t_L         g13720(.A(new_n13605), .Y(new_n13977));
  O2A1O1Ixp33_ASAP7_75t_L   g13721(.A1(new_n13439), .A2(new_n13568), .B(new_n13441), .C(new_n13977), .Y(new_n13978));
  A2O1A1O1Ixp25_ASAP7_75t_L g13722(.A1(new_n578), .A2(new_n12061), .B(new_n651), .C(\b[63] ), .D(new_n574), .Y(new_n13979));
  A2O1A1O1Ixp25_ASAP7_75t_L g13723(.A1(\b[61] ), .A2(new_n11471), .B(\b[62] ), .C(new_n578), .D(new_n651), .Y(new_n13980));
  NOR3xp33_ASAP7_75t_L      g13724(.A(new_n13980), .B(new_n11468), .C(\a[11] ), .Y(new_n13981));
  NOR2xp33_ASAP7_75t_L      g13725(.A(new_n13979), .B(new_n13981), .Y(new_n13982));
  INVx1_ASAP7_75t_L         g13726(.A(new_n13982), .Y(new_n13983));
  A2O1A1Ixp33_ASAP7_75t_L   g13727(.A1(new_n13976), .A2(new_n13774), .B(new_n13978), .C(new_n13983), .Y(new_n13984));
  O2A1O1Ixp33_ASAP7_75t_L   g13728(.A1(new_n13608), .A2(new_n13607), .B(new_n13774), .C(new_n13978), .Y(new_n13985));
  NAND2xp33_ASAP7_75t_L     g13729(.A(new_n13982), .B(new_n13985), .Y(new_n13986));
  NAND2xp33_ASAP7_75t_L     g13730(.A(new_n13984), .B(new_n13986), .Y(new_n13987));
  NOR3xp33_ASAP7_75t_L      g13731(.A(new_n13973), .B(new_n13975), .C(new_n13987), .Y(new_n13988));
  NAND2xp33_ASAP7_75t_L     g13732(.A(new_n13971), .B(new_n13974), .Y(new_n13989));
  NAND2xp33_ASAP7_75t_L     g13733(.A(new_n13807), .B(new_n13972), .Y(new_n13990));
  AND2x2_ASAP7_75t_L        g13734(.A(new_n13984), .B(new_n13986), .Y(new_n13991));
  AOI21xp33_ASAP7_75t_L     g13735(.A1(new_n13990), .A2(new_n13989), .B(new_n13991), .Y(new_n13992));
  OA21x2_ASAP7_75t_L        g13736(.A1(new_n13988), .A2(new_n13992), .B(new_n13794), .Y(new_n13993));
  NOR3xp33_ASAP7_75t_L      g13737(.A(new_n13992), .B(new_n13988), .C(new_n13794), .Y(new_n13994));
  NOR2xp33_ASAP7_75t_L      g13738(.A(new_n13994), .B(new_n13993), .Y(new_n13995));
  A2O1A1Ixp33_ASAP7_75t_L   g13739(.A1(new_n13789), .A2(new_n13785), .B(new_n13783), .C(new_n13995), .Y(new_n13996));
  INVx1_ASAP7_75t_L         g13740(.A(new_n13996), .Y(new_n13997));
  INVx1_ASAP7_75t_L         g13741(.A(new_n13783), .Y(new_n13998));
  A2O1A1Ixp33_ASAP7_75t_L   g13742(.A1(new_n13580), .A2(new_n13575), .B(new_n13784), .C(new_n13998), .Y(new_n13999));
  NOR2xp33_ASAP7_75t_L      g13743(.A(new_n13995), .B(new_n13999), .Y(new_n14000));
  NOR2xp33_ASAP7_75t_L      g13744(.A(new_n13997), .B(new_n14000), .Y(\f[74] ));
  AOI22xp33_ASAP7_75t_L     g13745(.A1(new_n1076), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1253), .Y(new_n14002));
  OAI221xp5_ASAP7_75t_L     g13746(.A1(new_n1154), .A2(new_n9947), .B1(new_n1156), .B2(new_n11446), .C(new_n14002), .Y(new_n14003));
  XNOR2x2_ASAP7_75t_L       g13747(.A(\a[17] ), .B(new_n14003), .Y(new_n14004));
  INVx1_ASAP7_75t_L         g13748(.A(new_n14004), .Y(new_n14005));
  O2A1O1Ixp33_ASAP7_75t_L   g13749(.A1(new_n13810), .A2(new_n13811), .B(new_n13969), .C(new_n14005), .Y(new_n14006));
  INVx1_ASAP7_75t_L         g13750(.A(new_n13813), .Y(new_n14007));
  AOI21xp33_ASAP7_75t_L     g13751(.A1(new_n13968), .A2(new_n13812), .B(new_n14007), .Y(new_n14008));
  NAND2xp33_ASAP7_75t_L     g13752(.A(new_n14005), .B(new_n14008), .Y(new_n14009));
  INVx1_ASAP7_75t_L         g13753(.A(new_n14009), .Y(new_n14010));
  AOI22xp33_ASAP7_75t_L     g13754(.A1(new_n1360), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1581), .Y(new_n14011));
  OAI221xp5_ASAP7_75t_L     g13755(.A1(new_n1373), .A2(new_n9323), .B1(new_n1359), .B2(new_n9627), .C(new_n14011), .Y(new_n14012));
  XNOR2x2_ASAP7_75t_L       g13756(.A(\a[20] ), .B(new_n14012), .Y(new_n14013));
  MAJIxp5_ASAP7_75t_L       g13757(.A(new_n13967), .B(new_n13816), .C(new_n13818), .Y(new_n14014));
  INVx1_ASAP7_75t_L         g13758(.A(new_n14014), .Y(new_n14015));
  NAND2xp33_ASAP7_75t_L     g13759(.A(new_n14013), .B(new_n14015), .Y(new_n14016));
  INVx1_ASAP7_75t_L         g13760(.A(new_n14013), .Y(new_n14017));
  NAND2xp33_ASAP7_75t_L     g13761(.A(new_n14017), .B(new_n14014), .Y(new_n14018));
  A2O1A1Ixp33_ASAP7_75t_L   g13762(.A1(new_n13820), .A2(new_n13636), .B(new_n13758), .C(new_n13828), .Y(new_n14019));
  OA21x2_ASAP7_75t_L        g13763(.A1(new_n13829), .A2(new_n13966), .B(new_n14019), .Y(new_n14020));
  AOI22xp33_ASAP7_75t_L     g13764(.A1(new_n1704), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1837), .Y(new_n14021));
  OAI221xp5_ASAP7_75t_L     g13765(.A1(new_n1699), .A2(new_n8165), .B1(new_n1827), .B2(new_n8465), .C(new_n14021), .Y(new_n14022));
  XNOR2x2_ASAP7_75t_L       g13766(.A(\a[23] ), .B(new_n14022), .Y(new_n14023));
  XOR2x2_ASAP7_75t_L        g13767(.A(new_n14023), .B(new_n14020), .Y(new_n14024));
  AOI22xp33_ASAP7_75t_L     g13768(.A1(new_n2114), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n2259), .Y(new_n14025));
  OAI221xp5_ASAP7_75t_L     g13769(.A1(new_n2109), .A2(new_n7593), .B1(new_n2257), .B2(new_n7623), .C(new_n14025), .Y(new_n14026));
  XNOR2x2_ASAP7_75t_L       g13770(.A(\a[26] ), .B(new_n14026), .Y(new_n14027));
  AOI21xp33_ASAP7_75t_L     g13771(.A1(new_n13962), .A2(new_n13839), .B(new_n13837), .Y(new_n14028));
  NAND2xp33_ASAP7_75t_L     g13772(.A(new_n14027), .B(new_n14028), .Y(new_n14029));
  O2A1O1Ixp33_ASAP7_75t_L   g13773(.A1(new_n13961), .A2(new_n13964), .B(new_n13838), .C(new_n14027), .Y(new_n14030));
  INVx1_ASAP7_75t_L         g13774(.A(new_n14030), .Y(new_n14031));
  INVx1_ASAP7_75t_L         g13775(.A(new_n13846), .Y(new_n14032));
  AOI22xp33_ASAP7_75t_L     g13776(.A1(new_n2552), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n2736), .Y(new_n14033));
  OAI221xp5_ASAP7_75t_L     g13777(.A1(new_n2547), .A2(new_n6812), .B1(new_n2734), .B2(new_n6837), .C(new_n14033), .Y(new_n14034));
  XNOR2x2_ASAP7_75t_L       g13778(.A(\a[29] ), .B(new_n14034), .Y(new_n14035));
  INVx1_ASAP7_75t_L         g13779(.A(new_n14035), .Y(new_n14036));
  A2O1A1O1Ixp25_ASAP7_75t_L g13780(.A1(new_n13957), .A2(new_n13956), .B(new_n13845), .C(new_n14032), .D(new_n14036), .Y(new_n14037));
  A2O1A1Ixp33_ASAP7_75t_L   g13781(.A1(new_n13956), .A2(new_n13957), .B(new_n13845), .C(new_n14032), .Y(new_n14038));
  NOR2xp33_ASAP7_75t_L      g13782(.A(new_n14035), .B(new_n14038), .Y(new_n14039));
  NOR2xp33_ASAP7_75t_L      g13783(.A(new_n14037), .B(new_n14039), .Y(new_n14040));
  AOI22xp33_ASAP7_75t_L     g13784(.A1(new_n3633), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n3858), .Y(new_n14041));
  OAI221xp5_ASAP7_75t_L     g13785(.A1(new_n3853), .A2(new_n5321), .B1(new_n3856), .B2(new_n5346), .C(new_n14041), .Y(new_n14042));
  XNOR2x2_ASAP7_75t_L       g13786(.A(\a[35] ), .B(new_n14042), .Y(new_n14043));
  NAND2xp33_ASAP7_75t_L     g13787(.A(new_n13947), .B(new_n13943), .Y(new_n14044));
  A2O1A1Ixp33_ASAP7_75t_L   g13788(.A1(new_n13939), .A2(new_n13938), .B(new_n13942), .C(new_n14044), .Y(new_n14045));
  AOI22xp33_ASAP7_75t_L     g13789(.A1(new_n4920), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n5167), .Y(new_n14046));
  OAI221xp5_ASAP7_75t_L     g13790(.A1(new_n5154), .A2(new_n3804), .B1(new_n5158), .B2(new_n4223), .C(new_n14046), .Y(new_n14047));
  XNOR2x2_ASAP7_75t_L       g13791(.A(\a[41] ), .B(new_n14047), .Y(new_n14048));
  INVx1_ASAP7_75t_L         g13792(.A(new_n13926), .Y(new_n14049));
  MAJIxp5_ASAP7_75t_L       g13793(.A(new_n13925), .B(new_n14049), .C(new_n13930), .Y(new_n14050));
  AOI22xp33_ASAP7_75t_L     g13794(.A1(new_n5624), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n5901), .Y(new_n14051));
  OAI221xp5_ASAP7_75t_L     g13795(.A1(new_n5900), .A2(new_n3207), .B1(new_n5892), .B2(new_n3572), .C(new_n14051), .Y(new_n14052));
  XNOR2x2_ASAP7_75t_L       g13796(.A(\a[44] ), .B(new_n14052), .Y(new_n14053));
  AOI21xp33_ASAP7_75t_L     g13797(.A1(new_n13914), .A2(new_n13869), .B(new_n13913), .Y(new_n14054));
  NOR2xp33_ASAP7_75t_L      g13798(.A(new_n13907), .B(new_n13909), .Y(new_n14055));
  AOI22xp33_ASAP7_75t_L     g13799(.A1(new_n7960), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n8537), .Y(new_n14056));
  OAI221xp5_ASAP7_75t_L     g13800(.A1(new_n8817), .A2(new_n1909), .B1(new_n7957), .B2(new_n2477), .C(new_n14056), .Y(new_n14057));
  XNOR2x2_ASAP7_75t_L       g13801(.A(\a[53] ), .B(new_n14057), .Y(new_n14058));
  INVx1_ASAP7_75t_L         g13802(.A(new_n14058), .Y(new_n14059));
  A2O1A1O1Ixp25_ASAP7_75t_L g13803(.A1(new_n13678), .A2(new_n13677), .B(new_n13688), .C(new_n13876), .D(new_n13882), .Y(new_n14060));
  A2O1A1O1Ixp25_ASAP7_75t_L g13804(.A1(new_n11533), .A2(\b[11] ), .B(new_n13878), .C(new_n13681), .D(new_n14060), .Y(new_n14061));
  AOI22xp33_ASAP7_75t_L     g13805(.A1(\b[13] ), .A2(new_n10939), .B1(\b[15] ), .B2(new_n10938), .Y(new_n14062));
  OAI221xp5_ASAP7_75t_L     g13806(.A1(new_n10937), .A2(new_n869), .B1(new_n10629), .B2(new_n950), .C(new_n14062), .Y(new_n14063));
  XNOR2x2_ASAP7_75t_L       g13807(.A(new_n10622), .B(new_n14063), .Y(new_n14064));
  NOR2xp33_ASAP7_75t_L      g13808(.A(new_n679), .B(new_n11535), .Y(new_n14065));
  O2A1O1Ixp33_ASAP7_75t_L   g13809(.A1(new_n11247), .A2(new_n11249), .B(\b[12] ), .C(new_n14065), .Y(new_n14066));
  A2O1A1Ixp33_ASAP7_75t_L   g13810(.A1(new_n11533), .A2(\b[10] ), .B(new_n13680), .C(\a[11] ), .Y(new_n14067));
  NOR2xp33_ASAP7_75t_L      g13811(.A(\a[11] ), .B(new_n13686), .Y(new_n14068));
  INVx1_ASAP7_75t_L         g13812(.A(new_n14068), .Y(new_n14069));
  AOI21xp33_ASAP7_75t_L     g13813(.A1(new_n14069), .A2(new_n14067), .B(new_n14066), .Y(new_n14070));
  AND3x1_ASAP7_75t_L        g13814(.A(new_n14069), .B(new_n14067), .C(new_n14066), .Y(new_n14071));
  NOR2xp33_ASAP7_75t_L      g13815(.A(new_n14070), .B(new_n14071), .Y(new_n14072));
  XNOR2x2_ASAP7_75t_L       g13816(.A(new_n14072), .B(new_n14064), .Y(new_n14073));
  XNOR2x2_ASAP7_75t_L       g13817(.A(new_n14061), .B(new_n14073), .Y(new_n14074));
  AOI22xp33_ASAP7_75t_L     g13818(.A1(new_n9700), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n10027), .Y(new_n14075));
  OAI221xp5_ASAP7_75t_L     g13819(.A1(new_n10024), .A2(new_n1201), .B1(new_n9696), .B2(new_n1320), .C(new_n14075), .Y(new_n14076));
  XNOR2x2_ASAP7_75t_L       g13820(.A(\a[59] ), .B(new_n14076), .Y(new_n14077));
  NOR2xp33_ASAP7_75t_L      g13821(.A(new_n14077), .B(new_n14074), .Y(new_n14078));
  INVx1_ASAP7_75t_L         g13822(.A(new_n14078), .Y(new_n14079));
  NAND2xp33_ASAP7_75t_L     g13823(.A(new_n14077), .B(new_n14074), .Y(new_n14080));
  AND2x2_ASAP7_75t_L        g13824(.A(new_n14080), .B(new_n14079), .Y(new_n14081));
  O2A1O1Ixp33_ASAP7_75t_L   g13825(.A1(new_n13883), .A2(new_n13887), .B(new_n13891), .C(new_n14081), .Y(new_n14082));
  NAND4xp25_ASAP7_75t_L     g13826(.A(new_n14079), .B(new_n13890), .C(new_n13891), .D(new_n14080), .Y(new_n14083));
  INVx1_ASAP7_75t_L         g13827(.A(new_n14083), .Y(new_n14084));
  NOR2xp33_ASAP7_75t_L      g13828(.A(new_n14084), .B(new_n14082), .Y(new_n14085));
  AOI22xp33_ASAP7_75t_L     g13829(.A1(new_n8831), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n9115), .Y(new_n14086));
  OAI221xp5_ASAP7_75t_L     g13830(.A1(new_n10343), .A2(new_n1539), .B1(new_n10016), .B2(new_n1662), .C(new_n14086), .Y(new_n14087));
  XNOR2x2_ASAP7_75t_L       g13831(.A(\a[56] ), .B(new_n14087), .Y(new_n14088));
  INVx1_ASAP7_75t_L         g13832(.A(new_n14088), .Y(new_n14089));
  XNOR2x2_ASAP7_75t_L       g13833(.A(new_n14089), .B(new_n14085), .Y(new_n14090));
  NOR2xp33_ASAP7_75t_L      g13834(.A(new_n13896), .B(new_n13903), .Y(new_n14091));
  XOR2x2_ASAP7_75t_L        g13835(.A(new_n14091), .B(new_n14090), .Y(new_n14092));
  XNOR2x2_ASAP7_75t_L       g13836(.A(new_n14059), .B(new_n14092), .Y(new_n14093));
  XNOR2x2_ASAP7_75t_L       g13837(.A(new_n14055), .B(new_n14093), .Y(new_n14094));
  AOI22xp33_ASAP7_75t_L     g13838(.A1(new_n7111), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n7391), .Y(new_n14095));
  OAI221xp5_ASAP7_75t_L     g13839(.A1(new_n8558), .A2(new_n2348), .B1(new_n8237), .B2(new_n2505), .C(new_n14095), .Y(new_n14096));
  XNOR2x2_ASAP7_75t_L       g13840(.A(\a[50] ), .B(new_n14096), .Y(new_n14097));
  XNOR2x2_ASAP7_75t_L       g13841(.A(new_n14097), .B(new_n14094), .Y(new_n14098));
  XOR2x2_ASAP7_75t_L        g13842(.A(new_n14054), .B(new_n14098), .Y(new_n14099));
  AOI22xp33_ASAP7_75t_L     g13843(.A1(new_n6376), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n6648), .Y(new_n14100));
  OAI221xp5_ASAP7_75t_L     g13844(.A1(new_n6646), .A2(new_n2688), .B1(new_n6636), .B2(new_n2990), .C(new_n14100), .Y(new_n14101));
  XNOR2x2_ASAP7_75t_L       g13845(.A(\a[47] ), .B(new_n14101), .Y(new_n14102));
  INVx1_ASAP7_75t_L         g13846(.A(new_n14102), .Y(new_n14103));
  XNOR2x2_ASAP7_75t_L       g13847(.A(new_n14103), .B(new_n14099), .Y(new_n14104));
  NAND2xp33_ASAP7_75t_L     g13848(.A(new_n13924), .B(new_n13921), .Y(new_n14105));
  A2O1A1Ixp33_ASAP7_75t_L   g13849(.A1(new_n13918), .A2(new_n13917), .B(new_n13920), .C(new_n14105), .Y(new_n14106));
  XOR2x2_ASAP7_75t_L        g13850(.A(new_n14104), .B(new_n14106), .Y(new_n14107));
  XNOR2x2_ASAP7_75t_L       g13851(.A(new_n14053), .B(new_n14107), .Y(new_n14108));
  XNOR2x2_ASAP7_75t_L       g13852(.A(new_n14050), .B(new_n14108), .Y(new_n14109));
  XNOR2x2_ASAP7_75t_L       g13853(.A(new_n14048), .B(new_n14109), .Y(new_n14110));
  NAND2xp33_ASAP7_75t_L     g13854(.A(new_n13934), .B(new_n13938), .Y(new_n14111));
  XNOR2x2_ASAP7_75t_L       g13855(.A(new_n14111), .B(new_n14110), .Y(new_n14112));
  AOI22xp33_ASAP7_75t_L     g13856(.A1(new_n4283), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n4512), .Y(new_n14113));
  OAI221xp5_ASAP7_75t_L     g13857(.A1(new_n4277), .A2(new_n4632), .B1(new_n4499), .B2(new_n4858), .C(new_n14113), .Y(new_n14114));
  XNOR2x2_ASAP7_75t_L       g13858(.A(\a[38] ), .B(new_n14114), .Y(new_n14115));
  XOR2x2_ASAP7_75t_L        g13859(.A(new_n14115), .B(new_n14112), .Y(new_n14116));
  XNOR2x2_ASAP7_75t_L       g13860(.A(new_n14045), .B(new_n14116), .Y(new_n14117));
  XNOR2x2_ASAP7_75t_L       g13861(.A(new_n14043), .B(new_n14117), .Y(new_n14118));
  A2O1A1Ixp33_ASAP7_75t_L   g13862(.A1(new_n13952), .A2(new_n13860), .B(new_n13951), .C(new_n14118), .Y(new_n14119));
  OR3x1_ASAP7_75t_L         g13863(.A(new_n14118), .B(new_n13954), .C(new_n13951), .Y(new_n14120));
  NAND2xp33_ASAP7_75t_L     g13864(.A(new_n14119), .B(new_n14120), .Y(new_n14121));
  AOI22xp33_ASAP7_75t_L     g13865(.A1(new_n3029), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n3258), .Y(new_n14122));
  OAI221xp5_ASAP7_75t_L     g13866(.A1(new_n3024), .A2(new_n5829), .B1(new_n3256), .B2(new_n6329), .C(new_n14122), .Y(new_n14123));
  XNOR2x2_ASAP7_75t_L       g13867(.A(\a[32] ), .B(new_n14123), .Y(new_n14124));
  AO21x2_ASAP7_75t_L        g13868(.A1(new_n13857), .A2(new_n13955), .B(new_n13856), .Y(new_n14125));
  XNOR2x2_ASAP7_75t_L       g13869(.A(new_n14124), .B(new_n14125), .Y(new_n14126));
  XNOR2x2_ASAP7_75t_L       g13870(.A(new_n14121), .B(new_n14126), .Y(new_n14127));
  XOR2x2_ASAP7_75t_L        g13871(.A(new_n14040), .B(new_n14127), .Y(new_n14128));
  AND3x1_ASAP7_75t_L        g13872(.A(new_n14029), .B(new_n14128), .C(new_n14031), .Y(new_n14129));
  AOI21xp33_ASAP7_75t_L     g13873(.A1(new_n14029), .A2(new_n14031), .B(new_n14128), .Y(new_n14130));
  NOR2xp33_ASAP7_75t_L      g13874(.A(new_n14129), .B(new_n14130), .Y(new_n14131));
  XOR2x2_ASAP7_75t_L        g13875(.A(new_n14131), .B(new_n14024), .Y(new_n14132));
  NAND3xp33_ASAP7_75t_L     g13876(.A(new_n14132), .B(new_n14018), .C(new_n14016), .Y(new_n14133));
  AO21x2_ASAP7_75t_L        g13877(.A1(new_n14016), .A2(new_n14018), .B(new_n14132), .Y(new_n14134));
  NAND2xp33_ASAP7_75t_L     g13878(.A(new_n14133), .B(new_n14134), .Y(new_n14135));
  INVx1_ASAP7_75t_L         g13879(.A(new_n14135), .Y(new_n14136));
  OAI21xp33_ASAP7_75t_L     g13880(.A1(new_n14006), .A2(new_n14010), .B(new_n14136), .Y(new_n14137));
  INVx1_ASAP7_75t_L         g13881(.A(new_n14137), .Y(new_n14138));
  NOR3xp33_ASAP7_75t_L      g13882(.A(new_n14136), .B(new_n14010), .C(new_n14006), .Y(new_n14139));
  NOR2xp33_ASAP7_75t_L      g13883(.A(new_n14139), .B(new_n14138), .Y(new_n14140));
  AOI22xp33_ASAP7_75t_L     g13884(.A1(new_n811), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n900), .Y(new_n14141));
  A2O1A1Ixp33_ASAP7_75t_L   g13885(.A1(new_n11470), .A2(new_n11473), .B(new_n898), .C(new_n14141), .Y(new_n14142));
  AOI21xp33_ASAP7_75t_L     g13886(.A1(new_n815), .A2(\b[62] ), .B(new_n14142), .Y(new_n14143));
  NAND2xp33_ASAP7_75t_L     g13887(.A(\a[14] ), .B(new_n14143), .Y(new_n14144));
  A2O1A1Ixp33_ASAP7_75t_L   g13888(.A1(\b[62] ), .A2(new_n815), .B(new_n14142), .C(new_n806), .Y(new_n14145));
  AND2x2_ASAP7_75t_L        g13889(.A(new_n14145), .B(new_n14144), .Y(new_n14146));
  A2O1A1Ixp33_ASAP7_75t_L   g13890(.A1(new_n13970), .A2(new_n13969), .B(new_n13803), .C(new_n13806), .Y(new_n14147));
  NOR2xp33_ASAP7_75t_L      g13891(.A(new_n14146), .B(new_n14147), .Y(new_n14148));
  INVx1_ASAP7_75t_L         g13892(.A(new_n14148), .Y(new_n14149));
  INVx1_ASAP7_75t_L         g13893(.A(new_n14146), .Y(new_n14150));
  A2O1A1O1Ixp25_ASAP7_75t_L g13894(.A1(new_n13969), .A2(new_n13970), .B(new_n13803), .C(new_n13806), .D(new_n14150), .Y(new_n14151));
  INVx1_ASAP7_75t_L         g13895(.A(new_n14151), .Y(new_n14152));
  NAND3xp33_ASAP7_75t_L     g13896(.A(new_n14140), .B(new_n14149), .C(new_n14152), .Y(new_n14153));
  OR3x1_ASAP7_75t_L         g13897(.A(new_n14136), .B(new_n14010), .C(new_n14006), .Y(new_n14154));
  NAND2xp33_ASAP7_75t_L     g13898(.A(new_n14137), .B(new_n14154), .Y(new_n14155));
  OAI21xp33_ASAP7_75t_L     g13899(.A1(new_n14148), .A2(new_n14151), .B(new_n14155), .Y(new_n14156));
  OAI31xp33_ASAP7_75t_L     g13900(.A1(new_n13973), .A2(new_n13975), .A3(new_n13987), .B(new_n13986), .Y(new_n14157));
  INVx1_ASAP7_75t_L         g13901(.A(new_n14157), .Y(new_n14158));
  NAND3xp33_ASAP7_75t_L     g13902(.A(new_n14153), .B(new_n14156), .C(new_n14158), .Y(new_n14159));
  NOR3xp33_ASAP7_75t_L      g13903(.A(new_n14155), .B(new_n14148), .C(new_n14151), .Y(new_n14160));
  AOI21xp33_ASAP7_75t_L     g13904(.A1(new_n14152), .A2(new_n14149), .B(new_n14140), .Y(new_n14161));
  OAI21xp33_ASAP7_75t_L     g13905(.A1(new_n14160), .A2(new_n14161), .B(new_n14157), .Y(new_n14162));
  AND2x2_ASAP7_75t_L        g13906(.A(new_n14159), .B(new_n14162), .Y(new_n14163));
  A2O1A1Ixp33_ASAP7_75t_L   g13907(.A1(new_n13999), .A2(new_n13995), .B(new_n13993), .C(new_n14163), .Y(new_n14164));
  INVx1_ASAP7_75t_L         g13908(.A(new_n14164), .Y(new_n14165));
  INVx1_ASAP7_75t_L         g13909(.A(new_n13993), .Y(new_n14166));
  A2O1A1Ixp33_ASAP7_75t_L   g13910(.A1(new_n13786), .A2(new_n13998), .B(new_n13994), .C(new_n14166), .Y(new_n14167));
  NOR2xp33_ASAP7_75t_L      g13911(.A(new_n14163), .B(new_n14167), .Y(new_n14168));
  NOR2xp33_ASAP7_75t_L      g13912(.A(new_n14168), .B(new_n14165), .Y(\f[75] ));
  INVx1_ASAP7_75t_L         g13913(.A(new_n14159), .Y(new_n14170));
  AOI21xp33_ASAP7_75t_L     g13914(.A1(new_n14140), .A2(new_n14152), .B(new_n14148), .Y(new_n14171));
  MAJIxp5_ASAP7_75t_L       g13915(.A(new_n14135), .B(new_n14008), .C(new_n14004), .Y(new_n14172));
  NOR2xp33_ASAP7_75t_L      g13916(.A(new_n898), .B(new_n11500), .Y(new_n14173));
  AOI21xp33_ASAP7_75t_L     g13917(.A1(new_n900), .A2(\b[62] ), .B(new_n14173), .Y(new_n14174));
  OAI211xp5_ASAP7_75t_L     g13918(.A1(new_n11468), .A2(new_n904), .B(new_n14174), .C(\a[14] ), .Y(new_n14175));
  O2A1O1Ixp33_ASAP7_75t_L   g13919(.A1(new_n11468), .A2(new_n904), .B(new_n14174), .C(\a[14] ), .Y(new_n14176));
  INVx1_ASAP7_75t_L         g13920(.A(new_n14176), .Y(new_n14177));
  AND2x2_ASAP7_75t_L        g13921(.A(new_n14175), .B(new_n14177), .Y(new_n14178));
  INVx1_ASAP7_75t_L         g13922(.A(new_n14178), .Y(new_n14179));
  XNOR2x2_ASAP7_75t_L       g13923(.A(new_n14179), .B(new_n14172), .Y(new_n14180));
  AOI22xp33_ASAP7_75t_L     g13924(.A1(new_n1076), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1253), .Y(new_n14181));
  OAI221xp5_ASAP7_75t_L     g13925(.A1(new_n1154), .A2(new_n10250), .B1(new_n1156), .B2(new_n10855), .C(new_n14181), .Y(new_n14182));
  XNOR2x2_ASAP7_75t_L       g13926(.A(\a[17] ), .B(new_n14182), .Y(new_n14183));
  NAND2xp33_ASAP7_75t_L     g13927(.A(new_n14018), .B(new_n14133), .Y(new_n14184));
  XNOR2x2_ASAP7_75t_L       g13928(.A(new_n14183), .B(new_n14184), .Y(new_n14185));
  O2A1O1Ixp33_ASAP7_75t_L   g13929(.A1(new_n13829), .A2(new_n13966), .B(new_n14019), .C(new_n14023), .Y(new_n14186));
  NOR2xp33_ASAP7_75t_L      g13930(.A(new_n9920), .B(new_n1372), .Y(new_n14187));
  AOI221xp5_ASAP7_75t_L     g13931(.A1(\b[56] ), .A2(new_n1581), .B1(\b[57] ), .B2(new_n1362), .C(new_n14187), .Y(new_n14188));
  OAI211xp5_ASAP7_75t_L     g13932(.A1(new_n1359), .A2(new_n9925), .B(\a[20] ), .C(new_n14188), .Y(new_n14189));
  O2A1O1Ixp33_ASAP7_75t_L   g13933(.A1(new_n1359), .A2(new_n9925), .B(new_n14188), .C(\a[20] ), .Y(new_n14190));
  INVx1_ASAP7_75t_L         g13934(.A(new_n14190), .Y(new_n14191));
  AND2x2_ASAP7_75t_L        g13935(.A(new_n14189), .B(new_n14191), .Y(new_n14192));
  A2O1A1Ixp33_ASAP7_75t_L   g13936(.A1(new_n14024), .A2(new_n14131), .B(new_n14186), .C(new_n14192), .Y(new_n14193));
  AO21x2_ASAP7_75t_L        g13937(.A1(new_n14131), .A2(new_n14024), .B(new_n14186), .Y(new_n14194));
  AO21x2_ASAP7_75t_L        g13938(.A1(new_n14191), .A2(new_n14189), .B(new_n14194), .Y(new_n14195));
  NAND2xp33_ASAP7_75t_L     g13939(.A(new_n14193), .B(new_n14195), .Y(new_n14196));
  AOI22xp33_ASAP7_75t_L     g13940(.A1(new_n1704), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1837), .Y(new_n14197));
  OAI221xp5_ASAP7_75t_L     g13941(.A1(new_n1699), .A2(new_n8458), .B1(new_n1827), .B2(new_n8768), .C(new_n14197), .Y(new_n14198));
  XNOR2x2_ASAP7_75t_L       g13942(.A(\a[23] ), .B(new_n14198), .Y(new_n14199));
  INVx1_ASAP7_75t_L         g13943(.A(new_n14199), .Y(new_n14200));
  AOI21xp33_ASAP7_75t_L     g13944(.A1(new_n14029), .A2(new_n14128), .B(new_n14030), .Y(new_n14201));
  NAND2xp33_ASAP7_75t_L     g13945(.A(new_n14200), .B(new_n14201), .Y(new_n14202));
  A2O1A1Ixp33_ASAP7_75t_L   g13946(.A1(new_n14029), .A2(new_n14128), .B(new_n14030), .C(new_n14199), .Y(new_n14203));
  AOI22xp33_ASAP7_75t_L     g13947(.A1(new_n2552), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n2736), .Y(new_n14204));
  OAI221xp5_ASAP7_75t_L     g13948(.A1(new_n2547), .A2(new_n6830), .B1(new_n2734), .B2(new_n7323), .C(new_n14204), .Y(new_n14205));
  XNOR2x2_ASAP7_75t_L       g13949(.A(\a[29] ), .B(new_n14205), .Y(new_n14206));
  MAJIxp5_ASAP7_75t_L       g13950(.A(new_n14121), .B(new_n14124), .C(new_n14125), .Y(new_n14207));
  NOR2xp33_ASAP7_75t_L      g13951(.A(new_n14206), .B(new_n14207), .Y(new_n14208));
  INVx1_ASAP7_75t_L         g13952(.A(new_n14208), .Y(new_n14209));
  NAND2xp33_ASAP7_75t_L     g13953(.A(new_n14206), .B(new_n14207), .Y(new_n14210));
  NAND2xp33_ASAP7_75t_L     g13954(.A(new_n14045), .B(new_n14116), .Y(new_n14211));
  OAI21xp33_ASAP7_75t_L     g13955(.A1(new_n14112), .A2(new_n14115), .B(new_n14211), .Y(new_n14212));
  AOI22xp33_ASAP7_75t_L     g13956(.A1(new_n4283), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n4512), .Y(new_n14213));
  OAI221xp5_ASAP7_75t_L     g13957(.A1(new_n4277), .A2(new_n4848), .B1(new_n4499), .B2(new_n11686), .C(new_n14213), .Y(new_n14214));
  XNOR2x2_ASAP7_75t_L       g13958(.A(\a[38] ), .B(new_n14214), .Y(new_n14215));
  MAJx2_ASAP7_75t_L         g13959(.A(new_n14111), .B(new_n14109), .C(new_n14048), .Y(new_n14216));
  AOI22xp33_ASAP7_75t_L     g13960(.A1(new_n4920), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n5167), .Y(new_n14217));
  OAI221xp5_ASAP7_75t_L     g13961(.A1(new_n5154), .A2(new_n4216), .B1(new_n5158), .B2(new_n4431), .C(new_n14217), .Y(new_n14218));
  XNOR2x2_ASAP7_75t_L       g13962(.A(\a[41] ), .B(new_n14218), .Y(new_n14219));
  INVx1_ASAP7_75t_L         g13963(.A(new_n14219), .Y(new_n14220));
  INVx1_ASAP7_75t_L         g13964(.A(new_n14107), .Y(new_n14221));
  NAND2xp33_ASAP7_75t_L     g13965(.A(new_n14050), .B(new_n14108), .Y(new_n14222));
  OAI21xp33_ASAP7_75t_L     g13966(.A1(new_n14053), .A2(new_n14221), .B(new_n14222), .Y(new_n14223));
  AOI22xp33_ASAP7_75t_L     g13967(.A1(new_n5624), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n5901), .Y(new_n14224));
  OAI221xp5_ASAP7_75t_L     g13968(.A1(new_n5900), .A2(new_n3565), .B1(new_n5892), .B2(new_n3591), .C(new_n14224), .Y(new_n14225));
  XNOR2x2_ASAP7_75t_L       g13969(.A(\a[44] ), .B(new_n14225), .Y(new_n14226));
  INVx1_ASAP7_75t_L         g13970(.A(new_n14226), .Y(new_n14227));
  AOI22xp33_ASAP7_75t_L     g13971(.A1(new_n6376), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n6648), .Y(new_n14228));
  OAI221xp5_ASAP7_75t_L     g13972(.A1(new_n6646), .A2(new_n2982), .B1(new_n6636), .B2(new_n3187), .C(new_n14228), .Y(new_n14229));
  XNOR2x2_ASAP7_75t_L       g13973(.A(\a[47] ), .B(new_n14229), .Y(new_n14230));
  NOR2xp33_ASAP7_75t_L      g13974(.A(new_n14097), .B(new_n14094), .Y(new_n14231));
  NAND2xp33_ASAP7_75t_L     g13975(.A(new_n14097), .B(new_n14094), .Y(new_n14232));
  A2O1A1O1Ixp25_ASAP7_75t_L g13976(.A1(new_n13869), .A2(new_n13916), .B(new_n13913), .C(new_n14232), .D(new_n14231), .Y(new_n14233));
  NOR2xp33_ASAP7_75t_L      g13977(.A(new_n760), .B(new_n11535), .Y(new_n14234));
  O2A1O1Ixp33_ASAP7_75t_L   g13978(.A1(new_n11247), .A2(new_n11249), .B(\b[13] ), .C(new_n14234), .Y(new_n14235));
  A2O1A1Ixp33_ASAP7_75t_L   g13979(.A1(new_n11533), .A2(\b[10] ), .B(new_n13680), .C(new_n574), .Y(new_n14236));
  A2O1A1Ixp33_ASAP7_75t_L   g13980(.A1(new_n14069), .A2(new_n14067), .B(new_n14066), .C(new_n14236), .Y(new_n14237));
  INVx1_ASAP7_75t_L         g13981(.A(new_n14237), .Y(new_n14238));
  NAND2xp33_ASAP7_75t_L     g13982(.A(new_n14235), .B(new_n14238), .Y(new_n14239));
  A2O1A1Ixp33_ASAP7_75t_L   g13983(.A1(new_n11533), .A2(\b[13] ), .B(new_n14234), .C(new_n14237), .Y(new_n14240));
  AND2x2_ASAP7_75t_L        g13984(.A(new_n14240), .B(new_n14239), .Y(new_n14241));
  AOI22xp33_ASAP7_75t_L     g13985(.A1(\b[14] ), .A2(new_n10939), .B1(\b[16] ), .B2(new_n10938), .Y(new_n14242));
  OAI221xp5_ASAP7_75t_L     g13986(.A1(new_n10937), .A2(new_n942), .B1(new_n10629), .B2(new_n1035), .C(new_n14242), .Y(new_n14243));
  XNOR2x2_ASAP7_75t_L       g13987(.A(\a[62] ), .B(new_n14243), .Y(new_n14244));
  XOR2x2_ASAP7_75t_L        g13988(.A(new_n14241), .B(new_n14244), .Y(new_n14245));
  AND2x2_ASAP7_75t_L        g13989(.A(new_n14072), .B(new_n14064), .Y(new_n14246));
  INVx1_ASAP7_75t_L         g13990(.A(new_n13877), .Y(new_n14247));
  A2O1A1Ixp33_ASAP7_75t_L   g13991(.A1(\b[11] ), .A2(new_n11533), .B(new_n13878), .C(new_n13681), .Y(new_n14248));
  O2A1O1Ixp33_ASAP7_75t_L   g13992(.A1(new_n14247), .A2(new_n13882), .B(new_n14248), .C(new_n14073), .Y(new_n14249));
  OR3x1_ASAP7_75t_L         g13993(.A(new_n14249), .B(new_n14245), .C(new_n14246), .Y(new_n14250));
  A2O1A1Ixp33_ASAP7_75t_L   g13994(.A1(new_n14064), .A2(new_n14072), .B(new_n14249), .C(new_n14245), .Y(new_n14251));
  NAND2xp33_ASAP7_75t_L     g13995(.A(new_n14251), .B(new_n14250), .Y(new_n14252));
  NAND2xp33_ASAP7_75t_L     g13996(.A(\b[17] ), .B(new_n10027), .Y(new_n14253));
  OAI221xp5_ASAP7_75t_L     g13997(.A1(new_n9699), .A2(new_n1432), .B1(new_n9696), .B2(new_n1438), .C(new_n14253), .Y(new_n14254));
  AOI21xp33_ASAP7_75t_L     g13998(.A1(new_n9703), .A2(\b[18] ), .B(new_n14254), .Y(new_n14255));
  NAND2xp33_ASAP7_75t_L     g13999(.A(\a[59] ), .B(new_n14255), .Y(new_n14256));
  A2O1A1Ixp33_ASAP7_75t_L   g14000(.A1(\b[18] ), .A2(new_n9703), .B(new_n14254), .C(new_n9693), .Y(new_n14257));
  NAND2xp33_ASAP7_75t_L     g14001(.A(new_n14257), .B(new_n14256), .Y(new_n14258));
  NOR2xp33_ASAP7_75t_L      g14002(.A(new_n14258), .B(new_n14252), .Y(new_n14259));
  INVx1_ASAP7_75t_L         g14003(.A(new_n14259), .Y(new_n14260));
  NAND2xp33_ASAP7_75t_L     g14004(.A(new_n14258), .B(new_n14252), .Y(new_n14261));
  NAND2xp33_ASAP7_75t_L     g14005(.A(new_n14261), .B(new_n14260), .Y(new_n14262));
  NAND2xp33_ASAP7_75t_L     g14006(.A(new_n14079), .B(new_n14083), .Y(new_n14263));
  NOR2xp33_ASAP7_75t_L      g14007(.A(new_n14263), .B(new_n14262), .Y(new_n14264));
  INVx1_ASAP7_75t_L         g14008(.A(new_n14262), .Y(new_n14265));
  O2A1O1Ixp33_ASAP7_75t_L   g14009(.A1(new_n14074), .A2(new_n14077), .B(new_n14083), .C(new_n14265), .Y(new_n14266));
  NOR2xp33_ASAP7_75t_L      g14010(.A(new_n14264), .B(new_n14266), .Y(new_n14267));
  AOI22xp33_ASAP7_75t_L     g14011(.A1(new_n8831), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n9115), .Y(new_n14268));
  OAI221xp5_ASAP7_75t_L     g14012(.A1(new_n10343), .A2(new_n1655), .B1(new_n10016), .B2(new_n1780), .C(new_n14268), .Y(new_n14269));
  XNOR2x2_ASAP7_75t_L       g14013(.A(\a[56] ), .B(new_n14269), .Y(new_n14270));
  NAND2xp33_ASAP7_75t_L     g14014(.A(new_n14270), .B(new_n14267), .Y(new_n14271));
  INVx1_ASAP7_75t_L         g14015(.A(new_n14270), .Y(new_n14272));
  OAI21xp33_ASAP7_75t_L     g14016(.A1(new_n14266), .A2(new_n14264), .B(new_n14272), .Y(new_n14273));
  O2A1O1Ixp33_ASAP7_75t_L   g14017(.A1(new_n13898), .A2(new_n13901), .B(new_n13897), .C(new_n14090), .Y(new_n14274));
  AOI21xp33_ASAP7_75t_L     g14018(.A1(new_n14089), .A2(new_n14085), .B(new_n14274), .Y(new_n14275));
  NAND3xp33_ASAP7_75t_L     g14019(.A(new_n14275), .B(new_n14273), .C(new_n14271), .Y(new_n14276));
  NAND2xp33_ASAP7_75t_L     g14020(.A(new_n14273), .B(new_n14271), .Y(new_n14277));
  A2O1A1Ixp33_ASAP7_75t_L   g14021(.A1(new_n14089), .A2(new_n14085), .B(new_n14274), .C(new_n14277), .Y(new_n14278));
  NAND2xp33_ASAP7_75t_L     g14022(.A(new_n14278), .B(new_n14276), .Y(new_n14279));
  AOI22xp33_ASAP7_75t_L     g14023(.A1(new_n7960), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n8537), .Y(new_n14280));
  OAI221xp5_ASAP7_75t_L     g14024(.A1(new_n8817), .A2(new_n1929), .B1(new_n7957), .B2(new_n2075), .C(new_n14280), .Y(new_n14281));
  XNOR2x2_ASAP7_75t_L       g14025(.A(\a[53] ), .B(new_n14281), .Y(new_n14282));
  XNOR2x2_ASAP7_75t_L       g14026(.A(new_n14282), .B(new_n14279), .Y(new_n14283));
  INVx1_ASAP7_75t_L         g14027(.A(new_n13907), .Y(new_n14284));
  NAND2xp33_ASAP7_75t_L     g14028(.A(new_n14059), .B(new_n14092), .Y(new_n14285));
  A2O1A1Ixp33_ASAP7_75t_L   g14029(.A1(new_n13910), .A2(new_n14284), .B(new_n14093), .C(new_n14285), .Y(new_n14286));
  XNOR2x2_ASAP7_75t_L       g14030(.A(new_n14286), .B(new_n14283), .Y(new_n14287));
  AOI22xp33_ASAP7_75t_L     g14031(.A1(new_n7111), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n7391), .Y(new_n14288));
  OAI221xp5_ASAP7_75t_L     g14032(.A1(new_n8558), .A2(new_n2497), .B1(new_n8237), .B2(new_n2672), .C(new_n14288), .Y(new_n14289));
  XNOR2x2_ASAP7_75t_L       g14033(.A(\a[50] ), .B(new_n14289), .Y(new_n14290));
  INVx1_ASAP7_75t_L         g14034(.A(new_n14290), .Y(new_n14291));
  XNOR2x2_ASAP7_75t_L       g14035(.A(new_n14291), .B(new_n14287), .Y(new_n14292));
  XOR2x2_ASAP7_75t_L        g14036(.A(new_n14233), .B(new_n14292), .Y(new_n14293));
  XNOR2x2_ASAP7_75t_L       g14037(.A(new_n14230), .B(new_n14293), .Y(new_n14294));
  NOR2xp33_ASAP7_75t_L      g14038(.A(new_n14104), .B(new_n14106), .Y(new_n14295));
  AOI21xp33_ASAP7_75t_L     g14039(.A1(new_n14103), .A2(new_n14099), .B(new_n14295), .Y(new_n14296));
  XNOR2x2_ASAP7_75t_L       g14040(.A(new_n14294), .B(new_n14296), .Y(new_n14297));
  XNOR2x2_ASAP7_75t_L       g14041(.A(new_n14227), .B(new_n14297), .Y(new_n14298));
  XNOR2x2_ASAP7_75t_L       g14042(.A(new_n14223), .B(new_n14298), .Y(new_n14299));
  XNOR2x2_ASAP7_75t_L       g14043(.A(new_n14220), .B(new_n14299), .Y(new_n14300));
  XOR2x2_ASAP7_75t_L        g14044(.A(new_n14216), .B(new_n14300), .Y(new_n14301));
  XNOR2x2_ASAP7_75t_L       g14045(.A(new_n14215), .B(new_n14301), .Y(new_n14302));
  XNOR2x2_ASAP7_75t_L       g14046(.A(new_n14212), .B(new_n14302), .Y(new_n14303));
  AOI22xp33_ASAP7_75t_L     g14047(.A1(new_n3633), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n3858), .Y(new_n14304));
  OAI221xp5_ASAP7_75t_L     g14048(.A1(new_n3853), .A2(new_n5338), .B1(new_n3856), .B2(new_n6338), .C(new_n14304), .Y(new_n14305));
  XNOR2x2_ASAP7_75t_L       g14049(.A(new_n3628), .B(new_n14305), .Y(new_n14306));
  NOR2xp33_ASAP7_75t_L      g14050(.A(new_n14306), .B(new_n14303), .Y(new_n14307));
  AND2x2_ASAP7_75t_L        g14051(.A(new_n14306), .B(new_n14303), .Y(new_n14308));
  NOR2xp33_ASAP7_75t_L      g14052(.A(new_n14307), .B(new_n14308), .Y(new_n14309));
  OA21x2_ASAP7_75t_L        g14053(.A1(new_n14043), .A2(new_n14117), .B(new_n14120), .Y(new_n14310));
  NOR2xp33_ASAP7_75t_L      g14054(.A(new_n6568), .B(new_n3022), .Y(new_n14311));
  AOI221xp5_ASAP7_75t_L     g14055(.A1(\b[44] ), .A2(new_n3258), .B1(\b[45] ), .B2(new_n3030), .C(new_n14311), .Y(new_n14312));
  OA211x2_ASAP7_75t_L       g14056(.A1(new_n3256), .A2(new_n6573), .B(new_n14312), .C(\a[32] ), .Y(new_n14313));
  O2A1O1Ixp33_ASAP7_75t_L   g14057(.A1(new_n3256), .A2(new_n6573), .B(new_n14312), .C(\a[32] ), .Y(new_n14314));
  NOR2xp33_ASAP7_75t_L      g14058(.A(new_n14314), .B(new_n14313), .Y(new_n14315));
  XNOR2x2_ASAP7_75t_L       g14059(.A(new_n14315), .B(new_n14310), .Y(new_n14316));
  XOR2x2_ASAP7_75t_L        g14060(.A(new_n14309), .B(new_n14316), .Y(new_n14317));
  AOI21xp33_ASAP7_75t_L     g14061(.A1(new_n14209), .A2(new_n14210), .B(new_n14317), .Y(new_n14318));
  AND3x1_ASAP7_75t_L        g14062(.A(new_n14317), .B(new_n14210), .C(new_n14209), .Y(new_n14319));
  NOR2xp33_ASAP7_75t_L      g14063(.A(new_n14040), .B(new_n14127), .Y(new_n14320));
  INVx1_ASAP7_75t_L         g14064(.A(new_n7906), .Y(new_n14321));
  NAND2xp33_ASAP7_75t_L     g14065(.A(\b[51] ), .B(new_n2115), .Y(new_n14322));
  OAI221xp5_ASAP7_75t_L     g14066(.A1(new_n2107), .A2(new_n7900), .B1(new_n7593), .B2(new_n2269), .C(new_n14322), .Y(new_n14323));
  AOI21xp33_ASAP7_75t_L     g14067(.A1(new_n14321), .A2(new_n2106), .B(new_n14323), .Y(new_n14324));
  NAND2xp33_ASAP7_75t_L     g14068(.A(\a[26] ), .B(new_n14324), .Y(new_n14325));
  A2O1A1Ixp33_ASAP7_75t_L   g14069(.A1(new_n14321), .A2(new_n2106), .B(new_n14323), .C(new_n2100), .Y(new_n14326));
  AND2x2_ASAP7_75t_L        g14070(.A(new_n14326), .B(new_n14325), .Y(new_n14327));
  INVx1_ASAP7_75t_L         g14071(.A(new_n14327), .Y(new_n14328));
  A2O1A1Ixp33_ASAP7_75t_L   g14072(.A1(new_n14036), .A2(new_n14038), .B(new_n14320), .C(new_n14328), .Y(new_n14329));
  NAND2xp33_ASAP7_75t_L     g14073(.A(new_n14036), .B(new_n14038), .Y(new_n14330));
  OAI211xp5_ASAP7_75t_L     g14074(.A1(new_n14040), .A2(new_n14127), .B(new_n14330), .C(new_n14327), .Y(new_n14331));
  NAND2xp33_ASAP7_75t_L     g14075(.A(new_n14331), .B(new_n14329), .Y(new_n14332));
  OAI21xp33_ASAP7_75t_L     g14076(.A1(new_n14318), .A2(new_n14319), .B(new_n14332), .Y(new_n14333));
  OR3x1_ASAP7_75t_L         g14077(.A(new_n14332), .B(new_n14318), .C(new_n14319), .Y(new_n14334));
  NAND2xp33_ASAP7_75t_L     g14078(.A(new_n14333), .B(new_n14334), .Y(new_n14335));
  INVx1_ASAP7_75t_L         g14079(.A(new_n14335), .Y(new_n14336));
  AOI21xp33_ASAP7_75t_L     g14080(.A1(new_n14203), .A2(new_n14202), .B(new_n14336), .Y(new_n14337));
  INVx1_ASAP7_75t_L         g14081(.A(new_n14202), .Y(new_n14338));
  INVx1_ASAP7_75t_L         g14082(.A(new_n14203), .Y(new_n14339));
  NOR3xp33_ASAP7_75t_L      g14083(.A(new_n14335), .B(new_n14339), .C(new_n14338), .Y(new_n14340));
  NOR2xp33_ASAP7_75t_L      g14084(.A(new_n14340), .B(new_n14337), .Y(new_n14341));
  XNOR2x2_ASAP7_75t_L       g14085(.A(new_n14341), .B(new_n14196), .Y(new_n14342));
  XOR2x2_ASAP7_75t_L        g14086(.A(new_n14342), .B(new_n14185), .Y(new_n14343));
  NOR2xp33_ASAP7_75t_L      g14087(.A(new_n14180), .B(new_n14343), .Y(new_n14344));
  XNOR2x2_ASAP7_75t_L       g14088(.A(new_n14178), .B(new_n14172), .Y(new_n14345));
  XNOR2x2_ASAP7_75t_L       g14089(.A(new_n14342), .B(new_n14185), .Y(new_n14346));
  NOR2xp33_ASAP7_75t_L      g14090(.A(new_n14345), .B(new_n14346), .Y(new_n14347));
  NOR3xp33_ASAP7_75t_L      g14091(.A(new_n14171), .B(new_n14344), .C(new_n14347), .Y(new_n14348));
  OA21x2_ASAP7_75t_L        g14092(.A1(new_n14347), .A2(new_n14344), .B(new_n14171), .Y(new_n14349));
  NOR2xp33_ASAP7_75t_L      g14093(.A(new_n14348), .B(new_n14349), .Y(new_n14350));
  A2O1A1Ixp33_ASAP7_75t_L   g14094(.A1(new_n14167), .A2(new_n14163), .B(new_n14170), .C(new_n14350), .Y(new_n14351));
  INVx1_ASAP7_75t_L         g14095(.A(new_n14351), .Y(new_n14352));
  NAND2xp33_ASAP7_75t_L     g14096(.A(new_n14159), .B(new_n14162), .Y(new_n14353));
  A2O1A1Ixp33_ASAP7_75t_L   g14097(.A1(new_n13996), .A2(new_n14166), .B(new_n14353), .C(new_n14159), .Y(new_n14354));
  NOR2xp33_ASAP7_75t_L      g14098(.A(new_n14350), .B(new_n14354), .Y(new_n14355));
  NOR2xp33_ASAP7_75t_L      g14099(.A(new_n14355), .B(new_n14352), .Y(\f[76] ));
  O2A1O1Ixp33_ASAP7_75t_L   g14100(.A1(new_n13810), .A2(new_n13811), .B(new_n13969), .C(new_n14004), .Y(new_n14357));
  O2A1O1Ixp33_ASAP7_75t_L   g14101(.A1(new_n14138), .A2(new_n14357), .B(new_n14179), .C(new_n14344), .Y(new_n14358));
  INVx1_ASAP7_75t_L         g14102(.A(new_n14192), .Y(new_n14359));
  MAJIxp5_ASAP7_75t_L       g14103(.A(new_n14341), .B(new_n14194), .C(new_n14359), .Y(new_n14360));
  NAND2xp33_ASAP7_75t_L     g14104(.A(\b[61] ), .B(new_n1080), .Y(new_n14361));
  OAI221xp5_ASAP7_75t_L     g14105(.A1(new_n1259), .A2(new_n11172), .B1(new_n10250), .B2(new_n1158), .C(new_n14361), .Y(new_n14362));
  AOI21xp33_ASAP7_75t_L     g14106(.A1(new_n11180), .A2(new_n1073), .B(new_n14362), .Y(new_n14363));
  NAND2xp33_ASAP7_75t_L     g14107(.A(\a[17] ), .B(new_n14363), .Y(new_n14364));
  A2O1A1Ixp33_ASAP7_75t_L   g14108(.A1(new_n11180), .A2(new_n1073), .B(new_n14362), .C(new_n1071), .Y(new_n14365));
  NAND2xp33_ASAP7_75t_L     g14109(.A(new_n14365), .B(new_n14364), .Y(new_n14366));
  XOR2x2_ASAP7_75t_L        g14110(.A(new_n14366), .B(new_n14360), .Y(new_n14367));
  AOI22xp33_ASAP7_75t_L     g14111(.A1(new_n1360), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1581), .Y(new_n14368));
  OAI221xp5_ASAP7_75t_L     g14112(.A1(new_n1373), .A2(new_n9920), .B1(new_n1359), .B2(new_n11152), .C(new_n14368), .Y(new_n14369));
  XNOR2x2_ASAP7_75t_L       g14113(.A(\a[20] ), .B(new_n14369), .Y(new_n14370));
  A2O1A1Ixp33_ASAP7_75t_L   g14114(.A1(new_n14029), .A2(new_n14128), .B(new_n14030), .C(new_n14200), .Y(new_n14371));
  INVx1_ASAP7_75t_L         g14115(.A(new_n14371), .Y(new_n14372));
  O2A1O1Ixp33_ASAP7_75t_L   g14116(.A1(new_n14338), .A2(new_n14339), .B(new_n14335), .C(new_n14372), .Y(new_n14373));
  NAND2xp33_ASAP7_75t_L     g14117(.A(new_n14370), .B(new_n14373), .Y(new_n14374));
  A2O1A1O1Ixp25_ASAP7_75t_L g14118(.A1(new_n14203), .A2(new_n14202), .B(new_n14336), .C(new_n14371), .D(new_n14370), .Y(new_n14375));
  INVx1_ASAP7_75t_L         g14119(.A(new_n14375), .Y(new_n14376));
  AND2x2_ASAP7_75t_L        g14120(.A(new_n14374), .B(new_n14376), .Y(new_n14377));
  AOI22xp33_ASAP7_75t_L     g14121(.A1(new_n1704), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1837), .Y(new_n14378));
  OAI221xp5_ASAP7_75t_L     g14122(.A1(new_n1699), .A2(new_n8762), .B1(new_n1827), .B2(new_n9331), .C(new_n14378), .Y(new_n14379));
  XNOR2x2_ASAP7_75t_L       g14123(.A(\a[23] ), .B(new_n14379), .Y(new_n14380));
  NAND2xp33_ASAP7_75t_L     g14124(.A(new_n14331), .B(new_n14334), .Y(new_n14381));
  NAND2xp33_ASAP7_75t_L     g14125(.A(new_n14380), .B(new_n14381), .Y(new_n14382));
  NOR2xp33_ASAP7_75t_L      g14126(.A(new_n14380), .B(new_n14381), .Y(new_n14383));
  INVx1_ASAP7_75t_L         g14127(.A(new_n14383), .Y(new_n14384));
  AOI22xp33_ASAP7_75t_L     g14128(.A1(new_n2114), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n2259), .Y(new_n14385));
  OAI221xp5_ASAP7_75t_L     g14129(.A1(new_n2109), .A2(new_n7900), .B1(new_n2257), .B2(new_n8174), .C(new_n14385), .Y(new_n14386));
  XNOR2x2_ASAP7_75t_L       g14130(.A(new_n2100), .B(new_n14386), .Y(new_n14387));
  INVx1_ASAP7_75t_L         g14131(.A(new_n14317), .Y(new_n14388));
  INVx1_ASAP7_75t_L         g14132(.A(new_n14206), .Y(new_n14389));
  NAND2xp33_ASAP7_75t_L     g14133(.A(new_n14389), .B(new_n14207), .Y(new_n14390));
  A2O1A1Ixp33_ASAP7_75t_L   g14134(.A1(new_n14210), .A2(new_n14209), .B(new_n14388), .C(new_n14390), .Y(new_n14391));
  NOR2xp33_ASAP7_75t_L      g14135(.A(new_n14387), .B(new_n14391), .Y(new_n14392));
  NAND2xp33_ASAP7_75t_L     g14136(.A(new_n14387), .B(new_n14391), .Y(new_n14393));
  INVx1_ASAP7_75t_L         g14137(.A(new_n14393), .Y(new_n14394));
  NOR2xp33_ASAP7_75t_L      g14138(.A(new_n14392), .B(new_n14394), .Y(new_n14395));
  NAND2xp33_ASAP7_75t_L     g14139(.A(\b[46] ), .B(new_n3030), .Y(new_n14396));
  OAI221xp5_ASAP7_75t_L     g14140(.A1(new_n3022), .A2(new_n6812), .B1(new_n6321), .B2(new_n3402), .C(new_n14396), .Y(new_n14397));
  AOI21xp33_ASAP7_75t_L     g14141(.A1(new_n8186), .A2(new_n3021), .B(new_n14397), .Y(new_n14398));
  NAND2xp33_ASAP7_75t_L     g14142(.A(\a[32] ), .B(new_n14398), .Y(new_n14399));
  A2O1A1Ixp33_ASAP7_75t_L   g14143(.A1(new_n8186), .A2(new_n3021), .B(new_n14397), .C(new_n3015), .Y(new_n14400));
  NAND2xp33_ASAP7_75t_L     g14144(.A(new_n14400), .B(new_n14399), .Y(new_n14401));
  NOR2xp33_ASAP7_75t_L      g14145(.A(new_n14212), .B(new_n14302), .Y(new_n14402));
  NOR2xp33_ASAP7_75t_L      g14146(.A(new_n14402), .B(new_n14307), .Y(new_n14403));
  XNOR2x2_ASAP7_75t_L       g14147(.A(new_n14401), .B(new_n14403), .Y(new_n14404));
  AOI22xp33_ASAP7_75t_L     g14148(.A1(new_n3633), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n3858), .Y(new_n14405));
  OAI221xp5_ASAP7_75t_L     g14149(.A1(new_n3853), .A2(new_n5805), .B1(new_n3856), .B2(new_n5835), .C(new_n14405), .Y(new_n14406));
  XNOR2x2_ASAP7_75t_L       g14150(.A(\a[35] ), .B(new_n14406), .Y(new_n14407));
  MAJx2_ASAP7_75t_L         g14151(.A(new_n14300), .B(new_n14216), .C(new_n14215), .Y(new_n14408));
  AOI22xp33_ASAP7_75t_L     g14152(.A1(new_n4283), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n4512), .Y(new_n14409));
  OAI221xp5_ASAP7_75t_L     g14153(.A1(new_n4277), .A2(new_n4869), .B1(new_n4499), .B2(new_n5327), .C(new_n14409), .Y(new_n14410));
  XNOR2x2_ASAP7_75t_L       g14154(.A(new_n4268), .B(new_n14410), .Y(new_n14411));
  O2A1O1Ixp33_ASAP7_75t_L   g14155(.A1(new_n14053), .A2(new_n14221), .B(new_n14222), .C(new_n14298), .Y(new_n14412));
  AO21x2_ASAP7_75t_L        g14156(.A1(new_n14220), .A2(new_n14299), .B(new_n14412), .Y(new_n14413));
  MAJIxp5_ASAP7_75t_L       g14157(.A(new_n14292), .B(new_n14230), .C(new_n14233), .Y(new_n14414));
  AOI22xp33_ASAP7_75t_L     g14158(.A1(new_n6376), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n6648), .Y(new_n14415));
  OAI221xp5_ASAP7_75t_L     g14159(.A1(new_n6646), .A2(new_n3180), .B1(new_n6636), .B2(new_n11047), .C(new_n14415), .Y(new_n14416));
  XNOR2x2_ASAP7_75t_L       g14160(.A(\a[47] ), .B(new_n14416), .Y(new_n14417));
  AOI22xp33_ASAP7_75t_L     g14161(.A1(new_n7960), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n8537), .Y(new_n14418));
  OAI221xp5_ASAP7_75t_L     g14162(.A1(new_n8817), .A2(new_n2067), .B1(new_n7957), .B2(new_n2355), .C(new_n14418), .Y(new_n14419));
  XNOR2x2_ASAP7_75t_L       g14163(.A(\a[53] ), .B(new_n14419), .Y(new_n14420));
  A2O1A1Ixp33_ASAP7_75t_L   g14164(.A1(new_n13686), .A2(new_n574), .B(new_n14070), .C(new_n14235), .Y(new_n14421));
  NOR2xp33_ASAP7_75t_L      g14165(.A(new_n784), .B(new_n11535), .Y(new_n14422));
  A2O1A1Ixp33_ASAP7_75t_L   g14166(.A1(\b[14] ), .A2(new_n11533), .B(new_n14422), .C(new_n14235), .Y(new_n14423));
  O2A1O1Ixp33_ASAP7_75t_L   g14167(.A1(new_n11247), .A2(new_n11249), .B(\b[14] ), .C(new_n14422), .Y(new_n14424));
  A2O1A1Ixp33_ASAP7_75t_L   g14168(.A1(new_n11533), .A2(\b[13] ), .B(new_n14234), .C(new_n14424), .Y(new_n14425));
  NAND2xp33_ASAP7_75t_L     g14169(.A(new_n14425), .B(new_n14423), .Y(new_n14426));
  INVx1_ASAP7_75t_L         g14170(.A(new_n14426), .Y(new_n14427));
  NOR2xp33_ASAP7_75t_L      g14171(.A(new_n1201), .B(new_n10630), .Y(new_n14428));
  AOI221xp5_ASAP7_75t_L     g14172(.A1(\b[15] ), .A2(new_n10939), .B1(\b[16] ), .B2(new_n10632), .C(new_n14428), .Y(new_n14429));
  OA211x2_ASAP7_75t_L       g14173(.A1(new_n10629), .A2(new_n1209), .B(\a[62] ), .C(new_n14429), .Y(new_n14430));
  O2A1O1Ixp33_ASAP7_75t_L   g14174(.A1(new_n10629), .A2(new_n1209), .B(new_n14429), .C(\a[62] ), .Y(new_n14431));
  OR2x4_ASAP7_75t_L         g14175(.A(new_n14431), .B(new_n14430), .Y(new_n14432));
  AND2x2_ASAP7_75t_L        g14176(.A(new_n14427), .B(new_n14432), .Y(new_n14433));
  INVx1_ASAP7_75t_L         g14177(.A(new_n14433), .Y(new_n14434));
  OR3x1_ASAP7_75t_L         g14178(.A(new_n14430), .B(new_n14431), .C(new_n14427), .Y(new_n14435));
  NAND2xp33_ASAP7_75t_L     g14179(.A(new_n14435), .B(new_n14434), .Y(new_n14436));
  O2A1O1Ixp33_ASAP7_75t_L   g14180(.A1(new_n14241), .A2(new_n14244), .B(new_n14421), .C(new_n14436), .Y(new_n14437));
  INVx1_ASAP7_75t_L         g14181(.A(new_n14437), .Y(new_n14438));
  A2O1A1Ixp33_ASAP7_75t_L   g14182(.A1(new_n14240), .A2(new_n14239), .B(new_n14244), .C(new_n14421), .Y(new_n14439));
  INVx1_ASAP7_75t_L         g14183(.A(new_n14436), .Y(new_n14440));
  NOR2xp33_ASAP7_75t_L      g14184(.A(new_n14439), .B(new_n14440), .Y(new_n14441));
  INVx1_ASAP7_75t_L         g14185(.A(new_n14441), .Y(new_n14442));
  AOI22xp33_ASAP7_75t_L     g14186(.A1(new_n9700), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n10027), .Y(new_n14443));
  OAI221xp5_ASAP7_75t_L     g14187(.A1(new_n10024), .A2(new_n1432), .B1(new_n9696), .B2(new_n1547), .C(new_n14443), .Y(new_n14444));
  XNOR2x2_ASAP7_75t_L       g14188(.A(\a[59] ), .B(new_n14444), .Y(new_n14445));
  NAND3xp33_ASAP7_75t_L     g14189(.A(new_n14442), .B(new_n14438), .C(new_n14445), .Y(new_n14446));
  AO21x2_ASAP7_75t_L        g14190(.A1(new_n14438), .A2(new_n14442), .B(new_n14445), .Y(new_n14447));
  NAND2xp33_ASAP7_75t_L     g14191(.A(new_n14446), .B(new_n14447), .Y(new_n14448));
  O2A1O1Ixp33_ASAP7_75t_L   g14192(.A1(new_n14252), .A2(new_n14258), .B(new_n14250), .C(new_n14448), .Y(new_n14449));
  AND2x2_ASAP7_75t_L        g14193(.A(new_n14446), .B(new_n14447), .Y(new_n14450));
  NAND2xp33_ASAP7_75t_L     g14194(.A(new_n14250), .B(new_n14260), .Y(new_n14451));
  NOR2xp33_ASAP7_75t_L      g14195(.A(new_n14451), .B(new_n14450), .Y(new_n14452));
  AOI22xp33_ASAP7_75t_L     g14196(.A1(new_n8831), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n9115), .Y(new_n14453));
  OAI221xp5_ASAP7_75t_L     g14197(.A1(new_n10343), .A2(new_n1774), .B1(new_n10016), .B2(new_n1915), .C(new_n14453), .Y(new_n14454));
  XNOR2x2_ASAP7_75t_L       g14198(.A(\a[56] ), .B(new_n14454), .Y(new_n14455));
  OAI21xp33_ASAP7_75t_L     g14199(.A1(new_n14449), .A2(new_n14452), .B(new_n14455), .Y(new_n14456));
  NOR2xp33_ASAP7_75t_L      g14200(.A(new_n14449), .B(new_n14452), .Y(new_n14457));
  INVx1_ASAP7_75t_L         g14201(.A(new_n14455), .Y(new_n14458));
  NAND2xp33_ASAP7_75t_L     g14202(.A(new_n14458), .B(new_n14457), .Y(new_n14459));
  NAND2xp33_ASAP7_75t_L     g14203(.A(new_n14456), .B(new_n14459), .Y(new_n14460));
  OAI21xp33_ASAP7_75t_L     g14204(.A1(new_n14262), .A2(new_n14263), .B(new_n14271), .Y(new_n14461));
  NOR2xp33_ASAP7_75t_L      g14205(.A(new_n14461), .B(new_n14460), .Y(new_n14462));
  AND2x2_ASAP7_75t_L        g14206(.A(new_n14461), .B(new_n14460), .Y(new_n14463));
  NOR3xp33_ASAP7_75t_L      g14207(.A(new_n14463), .B(new_n14462), .C(new_n14420), .Y(new_n14464));
  INVx1_ASAP7_75t_L         g14208(.A(new_n14464), .Y(new_n14465));
  OAI21xp33_ASAP7_75t_L     g14209(.A1(new_n14462), .A2(new_n14463), .B(new_n14420), .Y(new_n14466));
  NAND2xp33_ASAP7_75t_L     g14210(.A(new_n14466), .B(new_n14465), .Y(new_n14467));
  NAND3xp33_ASAP7_75t_L     g14211(.A(new_n14276), .B(new_n14278), .C(new_n14282), .Y(new_n14468));
  NAND2xp33_ASAP7_75t_L     g14212(.A(new_n14276), .B(new_n14468), .Y(new_n14469));
  NOR2xp33_ASAP7_75t_L      g14213(.A(new_n14469), .B(new_n14467), .Y(new_n14470));
  INVx1_ASAP7_75t_L         g14214(.A(new_n14282), .Y(new_n14471));
  INVx1_ASAP7_75t_L         g14215(.A(new_n14466), .Y(new_n14472));
  NOR2xp33_ASAP7_75t_L      g14216(.A(new_n14464), .B(new_n14472), .Y(new_n14473));
  O2A1O1Ixp33_ASAP7_75t_L   g14217(.A1(new_n14279), .A2(new_n14471), .B(new_n14276), .C(new_n14473), .Y(new_n14474));
  NOR2xp33_ASAP7_75t_L      g14218(.A(new_n14470), .B(new_n14474), .Y(new_n14475));
  AOI22xp33_ASAP7_75t_L     g14219(.A1(new_n7111), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n7391), .Y(new_n14476));
  OAI221xp5_ASAP7_75t_L     g14220(.A1(new_n8558), .A2(new_n2666), .B1(new_n8237), .B2(new_n2695), .C(new_n14476), .Y(new_n14477));
  XNOR2x2_ASAP7_75t_L       g14221(.A(\a[50] ), .B(new_n14477), .Y(new_n14478));
  NAND2xp33_ASAP7_75t_L     g14222(.A(new_n14478), .B(new_n14475), .Y(new_n14479));
  XNOR2x2_ASAP7_75t_L       g14223(.A(new_n14469), .B(new_n14467), .Y(new_n14480));
  INVx1_ASAP7_75t_L         g14224(.A(new_n14478), .Y(new_n14481));
  NAND2xp33_ASAP7_75t_L     g14225(.A(new_n14481), .B(new_n14480), .Y(new_n14482));
  NAND2xp33_ASAP7_75t_L     g14226(.A(new_n14482), .B(new_n14479), .Y(new_n14483));
  NAND2xp33_ASAP7_75t_L     g14227(.A(new_n14471), .B(new_n14279), .Y(new_n14484));
  INVx1_ASAP7_75t_L         g14228(.A(new_n14286), .Y(new_n14485));
  NAND2xp33_ASAP7_75t_L     g14229(.A(new_n14291), .B(new_n14287), .Y(new_n14486));
  A2O1A1Ixp33_ASAP7_75t_L   g14230(.A1(new_n14484), .A2(new_n14468), .B(new_n14485), .C(new_n14486), .Y(new_n14487));
  XOR2x2_ASAP7_75t_L        g14231(.A(new_n14487), .B(new_n14483), .Y(new_n14488));
  XNOR2x2_ASAP7_75t_L       g14232(.A(new_n14417), .B(new_n14488), .Y(new_n14489));
  OR2x4_ASAP7_75t_L         g14233(.A(new_n14414), .B(new_n14489), .Y(new_n14490));
  NAND2xp33_ASAP7_75t_L     g14234(.A(new_n14414), .B(new_n14489), .Y(new_n14491));
  AOI22xp33_ASAP7_75t_L     g14235(.A1(new_n5624), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n5901), .Y(new_n14492));
  OAI221xp5_ASAP7_75t_L     g14236(.A1(new_n5900), .A2(new_n3584), .B1(new_n5892), .B2(new_n10137), .C(new_n14492), .Y(new_n14493));
  XNOR2x2_ASAP7_75t_L       g14237(.A(\a[44] ), .B(new_n14493), .Y(new_n14494));
  NAND3xp33_ASAP7_75t_L     g14238(.A(new_n14490), .B(new_n14491), .C(new_n14494), .Y(new_n14495));
  AO21x2_ASAP7_75t_L        g14239(.A1(new_n14491), .A2(new_n14490), .B(new_n14494), .Y(new_n14496));
  NAND2xp33_ASAP7_75t_L     g14240(.A(new_n14495), .B(new_n14496), .Y(new_n14497));
  A2O1A1Ixp33_ASAP7_75t_L   g14241(.A1(new_n14103), .A2(new_n14099), .B(new_n14295), .C(new_n14294), .Y(new_n14498));
  NAND2xp33_ASAP7_75t_L     g14242(.A(new_n14227), .B(new_n14297), .Y(new_n14499));
  NAND2xp33_ASAP7_75t_L     g14243(.A(new_n14498), .B(new_n14499), .Y(new_n14500));
  XOR2x2_ASAP7_75t_L        g14244(.A(new_n14500), .B(new_n14497), .Y(new_n14501));
  INVx1_ASAP7_75t_L         g14245(.A(new_n14501), .Y(new_n14502));
  AOI22xp33_ASAP7_75t_L     g14246(.A1(new_n4920), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n5167), .Y(new_n14503));
  OAI221xp5_ASAP7_75t_L     g14247(.A1(new_n5154), .A2(new_n4424), .B1(new_n5158), .B2(new_n4641), .C(new_n14503), .Y(new_n14504));
  XNOR2x2_ASAP7_75t_L       g14248(.A(\a[41] ), .B(new_n14504), .Y(new_n14505));
  NAND2xp33_ASAP7_75t_L     g14249(.A(new_n14505), .B(new_n14502), .Y(new_n14506));
  INVx1_ASAP7_75t_L         g14250(.A(new_n14505), .Y(new_n14507));
  NAND2xp33_ASAP7_75t_L     g14251(.A(new_n14507), .B(new_n14501), .Y(new_n14508));
  NAND3xp33_ASAP7_75t_L     g14252(.A(new_n14506), .B(new_n14413), .C(new_n14508), .Y(new_n14509));
  AO21x2_ASAP7_75t_L        g14253(.A1(new_n14508), .A2(new_n14506), .B(new_n14413), .Y(new_n14510));
  NAND3xp33_ASAP7_75t_L     g14254(.A(new_n14510), .B(new_n14509), .C(new_n14411), .Y(new_n14511));
  AO21x2_ASAP7_75t_L        g14255(.A1(new_n14509), .A2(new_n14510), .B(new_n14411), .Y(new_n14512));
  NAND2xp33_ASAP7_75t_L     g14256(.A(new_n14511), .B(new_n14512), .Y(new_n14513));
  XOR2x2_ASAP7_75t_L        g14257(.A(new_n14408), .B(new_n14513), .Y(new_n14514));
  XNOR2x2_ASAP7_75t_L       g14258(.A(new_n14407), .B(new_n14514), .Y(new_n14515));
  XNOR2x2_ASAP7_75t_L       g14259(.A(new_n14515), .B(new_n14404), .Y(new_n14516));
  MAJIxp5_ASAP7_75t_L       g14260(.A(new_n14310), .B(new_n14315), .C(new_n14309), .Y(new_n14517));
  NAND2xp33_ASAP7_75t_L     g14261(.A(\b[49] ), .B(new_n2553), .Y(new_n14518));
  OAI221xp5_ASAP7_75t_L     g14262(.A1(new_n2545), .A2(new_n7593), .B1(new_n6830), .B2(new_n2747), .C(new_n14518), .Y(new_n14519));
  AOI21xp33_ASAP7_75t_L     g14263(.A1(new_n7601), .A2(new_n2544), .B(new_n14519), .Y(new_n14520));
  NAND2xp33_ASAP7_75t_L     g14264(.A(\a[29] ), .B(new_n14520), .Y(new_n14521));
  A2O1A1Ixp33_ASAP7_75t_L   g14265(.A1(new_n7601), .A2(new_n2544), .B(new_n14519), .C(new_n2538), .Y(new_n14522));
  NAND2xp33_ASAP7_75t_L     g14266(.A(new_n14522), .B(new_n14521), .Y(new_n14523));
  NAND2xp33_ASAP7_75t_L     g14267(.A(new_n14523), .B(new_n14517), .Y(new_n14524));
  OR2x4_ASAP7_75t_L         g14268(.A(new_n14523), .B(new_n14517), .Y(new_n14525));
  NAND2xp33_ASAP7_75t_L     g14269(.A(new_n14524), .B(new_n14525), .Y(new_n14526));
  NAND2xp33_ASAP7_75t_L     g14270(.A(new_n14516), .B(new_n14526), .Y(new_n14527));
  OR2x4_ASAP7_75t_L         g14271(.A(new_n14516), .B(new_n14526), .Y(new_n14528));
  NAND2xp33_ASAP7_75t_L     g14272(.A(new_n14527), .B(new_n14528), .Y(new_n14529));
  XOR2x2_ASAP7_75t_L        g14273(.A(new_n14529), .B(new_n14395), .Y(new_n14530));
  NAND3xp33_ASAP7_75t_L     g14274(.A(new_n14384), .B(new_n14382), .C(new_n14530), .Y(new_n14531));
  AO21x2_ASAP7_75t_L        g14275(.A1(new_n14382), .A2(new_n14384), .B(new_n14530), .Y(new_n14532));
  AND3x1_ASAP7_75t_L        g14276(.A(new_n14377), .B(new_n14532), .C(new_n14531), .Y(new_n14533));
  AND2x2_ASAP7_75t_L        g14277(.A(new_n14531), .B(new_n14532), .Y(new_n14534));
  NOR2xp33_ASAP7_75t_L      g14278(.A(new_n14377), .B(new_n14534), .Y(new_n14535));
  OR3x1_ASAP7_75t_L         g14279(.A(new_n14367), .B(new_n14533), .C(new_n14535), .Y(new_n14536));
  OAI21xp33_ASAP7_75t_L     g14280(.A1(new_n14533), .A2(new_n14535), .B(new_n14367), .Y(new_n14537));
  NAND2xp33_ASAP7_75t_L     g14281(.A(new_n14537), .B(new_n14536), .Y(new_n14538));
  INVx1_ASAP7_75t_L         g14282(.A(new_n14184), .Y(new_n14539));
  MAJIxp5_ASAP7_75t_L       g14283(.A(new_n14342), .B(new_n14183), .C(new_n14539), .Y(new_n14540));
  A2O1A1Ixp33_ASAP7_75t_L   g14284(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n808), .Y(new_n14541));
  A2O1A1Ixp33_ASAP7_75t_L   g14285(.A1(new_n14541), .A2(new_n978), .B(new_n11468), .C(\a[14] ), .Y(new_n14542));
  O2A1O1Ixp33_ASAP7_75t_L   g14286(.A1(new_n898), .A2(new_n12060), .B(new_n978), .C(new_n11468), .Y(new_n14543));
  NAND2xp33_ASAP7_75t_L     g14287(.A(new_n806), .B(new_n14543), .Y(new_n14544));
  AND2x2_ASAP7_75t_L        g14288(.A(new_n14544), .B(new_n14542), .Y(new_n14545));
  INVx1_ASAP7_75t_L         g14289(.A(new_n14545), .Y(new_n14546));
  XNOR2x2_ASAP7_75t_L       g14290(.A(new_n14546), .B(new_n14540), .Y(new_n14547));
  NOR2xp33_ASAP7_75t_L      g14291(.A(new_n14538), .B(new_n14547), .Y(new_n14548));
  INVx1_ASAP7_75t_L         g14292(.A(new_n14538), .Y(new_n14549));
  AND2x2_ASAP7_75t_L        g14293(.A(new_n14546), .B(new_n14540), .Y(new_n14550));
  NOR2xp33_ASAP7_75t_L      g14294(.A(new_n14546), .B(new_n14540), .Y(new_n14551));
  NOR2xp33_ASAP7_75t_L      g14295(.A(new_n14551), .B(new_n14550), .Y(new_n14552));
  NOR2xp33_ASAP7_75t_L      g14296(.A(new_n14552), .B(new_n14549), .Y(new_n14553));
  NOR3xp33_ASAP7_75t_L      g14297(.A(new_n14553), .B(new_n14548), .C(new_n14358), .Y(new_n14554));
  INVx1_ASAP7_75t_L         g14298(.A(new_n14357), .Y(new_n14555));
  NAND2xp33_ASAP7_75t_L     g14299(.A(new_n14345), .B(new_n14346), .Y(new_n14556));
  A2O1A1Ixp33_ASAP7_75t_L   g14300(.A1(new_n14555), .A2(new_n14137), .B(new_n14178), .C(new_n14556), .Y(new_n14557));
  NAND2xp33_ASAP7_75t_L     g14301(.A(new_n14552), .B(new_n14549), .Y(new_n14558));
  NAND2xp33_ASAP7_75t_L     g14302(.A(new_n14538), .B(new_n14547), .Y(new_n14559));
  AOI21xp33_ASAP7_75t_L     g14303(.A1(new_n14558), .A2(new_n14559), .B(new_n14557), .Y(new_n14560));
  NOR2xp33_ASAP7_75t_L      g14304(.A(new_n14560), .B(new_n14554), .Y(new_n14561));
  A2O1A1Ixp33_ASAP7_75t_L   g14305(.A1(new_n14354), .A2(new_n14350), .B(new_n14348), .C(new_n14561), .Y(new_n14562));
  INVx1_ASAP7_75t_L         g14306(.A(new_n14562), .Y(new_n14563));
  INVx1_ASAP7_75t_L         g14307(.A(new_n14348), .Y(new_n14564));
  A2O1A1Ixp33_ASAP7_75t_L   g14308(.A1(new_n14164), .A2(new_n14159), .B(new_n14349), .C(new_n14564), .Y(new_n14565));
  NOR2xp33_ASAP7_75t_L      g14309(.A(new_n14561), .B(new_n14565), .Y(new_n14566));
  NOR2xp33_ASAP7_75t_L      g14310(.A(new_n14563), .B(new_n14566), .Y(\f[77] ));
  NOR2xp33_ASAP7_75t_L      g14311(.A(new_n14550), .B(new_n14548), .Y(new_n14568));
  AOI22xp33_ASAP7_75t_L     g14312(.A1(new_n1076), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1253), .Y(new_n14569));
  A2O1A1Ixp33_ASAP7_75t_L   g14313(.A1(new_n11470), .A2(new_n11473), .B(new_n1156), .C(new_n14569), .Y(new_n14570));
  AOI21xp33_ASAP7_75t_L     g14314(.A1(new_n1080), .A2(\b[62] ), .B(new_n14570), .Y(new_n14571));
  NAND2xp33_ASAP7_75t_L     g14315(.A(\a[17] ), .B(new_n14571), .Y(new_n14572));
  A2O1A1Ixp33_ASAP7_75t_L   g14316(.A1(\b[62] ), .A2(new_n1080), .B(new_n14570), .C(new_n1071), .Y(new_n14573));
  AND2x2_ASAP7_75t_L        g14317(.A(new_n14573), .B(new_n14572), .Y(new_n14574));
  INVx1_ASAP7_75t_L         g14318(.A(new_n14574), .Y(new_n14575));
  A2O1A1O1Ixp25_ASAP7_75t_L g14319(.A1(new_n14364), .A2(new_n14365), .B(new_n14360), .C(new_n14536), .D(new_n14575), .Y(new_n14576));
  INVx1_ASAP7_75t_L         g14320(.A(new_n14576), .Y(new_n14577));
  A2O1A1Ixp33_ASAP7_75t_L   g14321(.A1(new_n14364), .A2(new_n14365), .B(new_n14360), .C(new_n14536), .Y(new_n14578));
  NOR2xp33_ASAP7_75t_L      g14322(.A(new_n14574), .B(new_n14578), .Y(new_n14579));
  INVx1_ASAP7_75t_L         g14323(.A(new_n14579), .Y(new_n14580));
  AOI22xp33_ASAP7_75t_L     g14324(.A1(new_n1360), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1581), .Y(new_n14581));
  OAI221xp5_ASAP7_75t_L     g14325(.A1(new_n1373), .A2(new_n9947), .B1(new_n1359), .B2(new_n11446), .C(new_n14581), .Y(new_n14582));
  XNOR2x2_ASAP7_75t_L       g14326(.A(\a[20] ), .B(new_n14582), .Y(new_n14583));
  INVx1_ASAP7_75t_L         g14327(.A(new_n14583), .Y(new_n14584));
  NOR3xp33_ASAP7_75t_L      g14328(.A(new_n14533), .B(new_n14584), .C(new_n14375), .Y(new_n14585));
  INVx1_ASAP7_75t_L         g14329(.A(new_n14585), .Y(new_n14586));
  A2O1A1Ixp33_ASAP7_75t_L   g14330(.A1(new_n14534), .A2(new_n14374), .B(new_n14375), .C(new_n14584), .Y(new_n14587));
  AOI22xp33_ASAP7_75t_L     g14331(.A1(new_n1704), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1837), .Y(new_n14588));
  OAI221xp5_ASAP7_75t_L     g14332(.A1(new_n1699), .A2(new_n9323), .B1(new_n1827), .B2(new_n9627), .C(new_n14588), .Y(new_n14589));
  XNOR2x2_ASAP7_75t_L       g14333(.A(\a[23] ), .B(new_n14589), .Y(new_n14590));
  A2O1A1Ixp33_ASAP7_75t_L   g14334(.A1(new_n14530), .A2(new_n14382), .B(new_n14383), .C(new_n14590), .Y(new_n14591));
  INVx1_ASAP7_75t_L         g14335(.A(new_n14591), .Y(new_n14592));
  INVx1_ASAP7_75t_L         g14336(.A(new_n14531), .Y(new_n14593));
  NOR3xp33_ASAP7_75t_L      g14337(.A(new_n14593), .B(new_n14590), .C(new_n14383), .Y(new_n14594));
  AOI22xp33_ASAP7_75t_L     g14338(.A1(new_n2114), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n2259), .Y(new_n14595));
  OAI221xp5_ASAP7_75t_L     g14339(.A1(new_n2109), .A2(new_n8165), .B1(new_n2257), .B2(new_n8465), .C(new_n14595), .Y(new_n14596));
  XNOR2x2_ASAP7_75t_L       g14340(.A(\a[26] ), .B(new_n14596), .Y(new_n14597));
  A2O1A1Ixp33_ASAP7_75t_L   g14341(.A1(new_n14527), .A2(new_n14528), .B(new_n14392), .C(new_n14393), .Y(new_n14598));
  XOR2x2_ASAP7_75t_L        g14342(.A(new_n14597), .B(new_n14598), .Y(new_n14599));
  AOI22xp33_ASAP7_75t_L     g14343(.A1(new_n2552), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n2736), .Y(new_n14600));
  OAI221xp5_ASAP7_75t_L     g14344(.A1(new_n2547), .A2(new_n7593), .B1(new_n2734), .B2(new_n7623), .C(new_n14600), .Y(new_n14601));
  XNOR2x2_ASAP7_75t_L       g14345(.A(\a[29] ), .B(new_n14601), .Y(new_n14602));
  INVx1_ASAP7_75t_L         g14346(.A(new_n14602), .Y(new_n14603));
  O2A1O1Ixp33_ASAP7_75t_L   g14347(.A1(new_n14516), .A2(new_n14526), .B(new_n14525), .C(new_n14603), .Y(new_n14604));
  AND3x1_ASAP7_75t_L        g14348(.A(new_n14528), .B(new_n14603), .C(new_n14525), .Y(new_n14605));
  NOR2xp33_ASAP7_75t_L      g14349(.A(new_n14604), .B(new_n14605), .Y(new_n14606));
  NAND2xp33_ASAP7_75t_L     g14350(.A(new_n14509), .B(new_n14511), .Y(new_n14607));
  AOI22xp33_ASAP7_75t_L     g14351(.A1(new_n4283), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n4512), .Y(new_n14608));
  OAI221xp5_ASAP7_75t_L     g14352(.A1(new_n4277), .A2(new_n5321), .B1(new_n4499), .B2(new_n5346), .C(new_n14608), .Y(new_n14609));
  XNOR2x2_ASAP7_75t_L       g14353(.A(\a[38] ), .B(new_n14609), .Y(new_n14610));
  INVx1_ASAP7_75t_L         g14354(.A(new_n14497), .Y(new_n14611));
  A2O1A1Ixp33_ASAP7_75t_L   g14355(.A1(new_n14499), .A2(new_n14498), .B(new_n14611), .C(new_n14508), .Y(new_n14612));
  AOI22xp33_ASAP7_75t_L     g14356(.A1(new_n5624), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n5901), .Y(new_n14613));
  OAI221xp5_ASAP7_75t_L     g14357(.A1(new_n5900), .A2(new_n3804), .B1(new_n5892), .B2(new_n4223), .C(new_n14613), .Y(new_n14614));
  XNOR2x2_ASAP7_75t_L       g14358(.A(\a[44] ), .B(new_n14614), .Y(new_n14615));
  INVx1_ASAP7_75t_L         g14359(.A(new_n14615), .Y(new_n14616));
  AOI22xp33_ASAP7_75t_L     g14360(.A1(new_n7960), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n8537), .Y(new_n14617));
  OAI221xp5_ASAP7_75t_L     g14361(.A1(new_n8817), .A2(new_n2348), .B1(new_n7957), .B2(new_n2505), .C(new_n14617), .Y(new_n14618));
  XNOR2x2_ASAP7_75t_L       g14362(.A(\a[53] ), .B(new_n14618), .Y(new_n14619));
  A2O1A1Ixp33_ASAP7_75t_L   g14363(.A1(new_n14447), .A2(new_n14446), .B(new_n14451), .C(new_n14459), .Y(new_n14620));
  AOI22xp33_ASAP7_75t_L     g14364(.A1(\b[16] ), .A2(new_n10939), .B1(\b[18] ), .B2(new_n10938), .Y(new_n14621));
  OAI221xp5_ASAP7_75t_L     g14365(.A1(new_n10937), .A2(new_n1201), .B1(new_n10629), .B2(new_n1320), .C(new_n14621), .Y(new_n14622));
  XNOR2x2_ASAP7_75t_L       g14366(.A(\a[62] ), .B(new_n14622), .Y(new_n14623));
  NOR2xp33_ASAP7_75t_L      g14367(.A(new_n869), .B(new_n11535), .Y(new_n14624));
  AOI211xp5_ASAP7_75t_L     g14368(.A1(new_n11533), .A2(\b[15] ), .B(new_n14624), .C(\a[14] ), .Y(new_n14625));
  INVx1_ASAP7_75t_L         g14369(.A(new_n14625), .Y(new_n14626));
  A2O1A1Ixp33_ASAP7_75t_L   g14370(.A1(new_n11533), .A2(\b[15] ), .B(new_n14624), .C(\a[14] ), .Y(new_n14627));
  NAND2xp33_ASAP7_75t_L     g14371(.A(new_n14627), .B(new_n14626), .Y(new_n14628));
  A2O1A1Ixp33_ASAP7_75t_L   g14372(.A1(new_n11533), .A2(\b[13] ), .B(new_n14234), .C(new_n14628), .Y(new_n14629));
  INVx1_ASAP7_75t_L         g14373(.A(new_n14629), .Y(new_n14630));
  AND3x1_ASAP7_75t_L        g14374(.A(new_n14626), .B(new_n14627), .C(new_n14235), .Y(new_n14631));
  NOR2xp33_ASAP7_75t_L      g14375(.A(new_n14631), .B(new_n14630), .Y(new_n14632));
  XNOR2x2_ASAP7_75t_L       g14376(.A(new_n14632), .B(new_n14623), .Y(new_n14633));
  A2O1A1O1Ixp25_ASAP7_75t_L g14377(.A1(new_n11533), .A2(\b[14] ), .B(new_n14422), .C(new_n14235), .D(new_n14433), .Y(new_n14634));
  XOR2x2_ASAP7_75t_L        g14378(.A(new_n14634), .B(new_n14633), .Y(new_n14635));
  AOI22xp33_ASAP7_75t_L     g14379(.A1(new_n9700), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n10027), .Y(new_n14636));
  OAI221xp5_ASAP7_75t_L     g14380(.A1(new_n10024), .A2(new_n1539), .B1(new_n9696), .B2(new_n1662), .C(new_n14636), .Y(new_n14637));
  XNOR2x2_ASAP7_75t_L       g14381(.A(\a[59] ), .B(new_n14637), .Y(new_n14638));
  XOR2x2_ASAP7_75t_L        g14382(.A(new_n14638), .B(new_n14635), .Y(new_n14639));
  AO21x2_ASAP7_75t_L        g14383(.A1(new_n14442), .A2(new_n14446), .B(new_n14639), .Y(new_n14640));
  NAND3xp33_ASAP7_75t_L     g14384(.A(new_n14639), .B(new_n14446), .C(new_n14442), .Y(new_n14641));
  NAND2xp33_ASAP7_75t_L     g14385(.A(new_n14641), .B(new_n14640), .Y(new_n14642));
  AOI22xp33_ASAP7_75t_L     g14386(.A1(new_n8831), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n9115), .Y(new_n14643));
  OAI221xp5_ASAP7_75t_L     g14387(.A1(new_n10343), .A2(new_n1909), .B1(new_n10016), .B2(new_n2477), .C(new_n14643), .Y(new_n14644));
  XNOR2x2_ASAP7_75t_L       g14388(.A(\a[56] ), .B(new_n14644), .Y(new_n14645));
  NOR2xp33_ASAP7_75t_L      g14389(.A(new_n14645), .B(new_n14642), .Y(new_n14646));
  INVx1_ASAP7_75t_L         g14390(.A(new_n14646), .Y(new_n14647));
  NAND2xp33_ASAP7_75t_L     g14391(.A(new_n14645), .B(new_n14642), .Y(new_n14648));
  AOI21xp33_ASAP7_75t_L     g14392(.A1(new_n14648), .A2(new_n14647), .B(new_n14620), .Y(new_n14649));
  NAND2xp33_ASAP7_75t_L     g14393(.A(new_n14648), .B(new_n14647), .Y(new_n14650));
  O2A1O1Ixp33_ASAP7_75t_L   g14394(.A1(new_n14450), .A2(new_n14451), .B(new_n14459), .C(new_n14650), .Y(new_n14651));
  NOR2xp33_ASAP7_75t_L      g14395(.A(new_n14649), .B(new_n14651), .Y(new_n14652));
  XNOR2x2_ASAP7_75t_L       g14396(.A(new_n14619), .B(new_n14652), .Y(new_n14653));
  NOR2xp33_ASAP7_75t_L      g14397(.A(new_n14462), .B(new_n14464), .Y(new_n14654));
  XNOR2x2_ASAP7_75t_L       g14398(.A(new_n14654), .B(new_n14653), .Y(new_n14655));
  AOI22xp33_ASAP7_75t_L     g14399(.A1(new_n7111), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n7391), .Y(new_n14656));
  OAI221xp5_ASAP7_75t_L     g14400(.A1(new_n8558), .A2(new_n2688), .B1(new_n8237), .B2(new_n2990), .C(new_n14656), .Y(new_n14657));
  XNOR2x2_ASAP7_75t_L       g14401(.A(\a[50] ), .B(new_n14657), .Y(new_n14658));
  INVx1_ASAP7_75t_L         g14402(.A(new_n14658), .Y(new_n14659));
  XNOR2x2_ASAP7_75t_L       g14403(.A(new_n14659), .B(new_n14655), .Y(new_n14660));
  NOR2xp33_ASAP7_75t_L      g14404(.A(new_n14481), .B(new_n14480), .Y(new_n14661));
  O2A1O1Ixp33_ASAP7_75t_L   g14405(.A1(new_n14464), .A2(new_n14472), .B(new_n14469), .C(new_n14661), .Y(new_n14662));
  XOR2x2_ASAP7_75t_L        g14406(.A(new_n14662), .B(new_n14660), .Y(new_n14663));
  AOI22xp33_ASAP7_75t_L     g14407(.A1(new_n6376), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n6648), .Y(new_n14664));
  OAI221xp5_ASAP7_75t_L     g14408(.A1(new_n6646), .A2(new_n3207), .B1(new_n6636), .B2(new_n3572), .C(new_n14664), .Y(new_n14665));
  XNOR2x2_ASAP7_75t_L       g14409(.A(\a[47] ), .B(new_n14665), .Y(new_n14666));
  XNOR2x2_ASAP7_75t_L       g14410(.A(new_n14666), .B(new_n14663), .Y(new_n14667));
  NOR2xp33_ASAP7_75t_L      g14411(.A(new_n14487), .B(new_n14483), .Y(new_n14668));
  INVx1_ASAP7_75t_L         g14412(.A(new_n14417), .Y(new_n14669));
  INVx1_ASAP7_75t_L         g14413(.A(new_n14483), .Y(new_n14670));
  O2A1O1Ixp33_ASAP7_75t_L   g14414(.A1(new_n14283), .A2(new_n14485), .B(new_n14486), .C(new_n14670), .Y(new_n14671));
  NOR3xp33_ASAP7_75t_L      g14415(.A(new_n14671), .B(new_n14668), .C(new_n14669), .Y(new_n14672));
  NOR2xp33_ASAP7_75t_L      g14416(.A(new_n14668), .B(new_n14672), .Y(new_n14673));
  XNOR2x2_ASAP7_75t_L       g14417(.A(new_n14667), .B(new_n14673), .Y(new_n14674));
  XNOR2x2_ASAP7_75t_L       g14418(.A(new_n14616), .B(new_n14674), .Y(new_n14675));
  NAND2xp33_ASAP7_75t_L     g14419(.A(new_n14490), .B(new_n14495), .Y(new_n14676));
  XNOR2x2_ASAP7_75t_L       g14420(.A(new_n14676), .B(new_n14675), .Y(new_n14677));
  AOI22xp33_ASAP7_75t_L     g14421(.A1(new_n4920), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n5167), .Y(new_n14678));
  OAI221xp5_ASAP7_75t_L     g14422(.A1(new_n5154), .A2(new_n4632), .B1(new_n5158), .B2(new_n4858), .C(new_n14678), .Y(new_n14679));
  XNOR2x2_ASAP7_75t_L       g14423(.A(\a[41] ), .B(new_n14679), .Y(new_n14680));
  XOR2x2_ASAP7_75t_L        g14424(.A(new_n14680), .B(new_n14677), .Y(new_n14681));
  XNOR2x2_ASAP7_75t_L       g14425(.A(new_n14612), .B(new_n14681), .Y(new_n14682));
  OR2x4_ASAP7_75t_L         g14426(.A(new_n14610), .B(new_n14682), .Y(new_n14683));
  NAND2xp33_ASAP7_75t_L     g14427(.A(new_n14610), .B(new_n14682), .Y(new_n14684));
  NAND2xp33_ASAP7_75t_L     g14428(.A(new_n14684), .B(new_n14683), .Y(new_n14685));
  XOR2x2_ASAP7_75t_L        g14429(.A(new_n14607), .B(new_n14685), .Y(new_n14686));
  AOI22xp33_ASAP7_75t_L     g14430(.A1(new_n3633), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n3858), .Y(new_n14687));
  OAI221xp5_ASAP7_75t_L     g14431(.A1(new_n3853), .A2(new_n5829), .B1(new_n3856), .B2(new_n6329), .C(new_n14687), .Y(new_n14688));
  XNOR2x2_ASAP7_75t_L       g14432(.A(\a[35] ), .B(new_n14688), .Y(new_n14689));
  XOR2x2_ASAP7_75t_L        g14433(.A(new_n14689), .B(new_n14686), .Y(new_n14690));
  MAJx2_ASAP7_75t_L         g14434(.A(new_n14513), .B(new_n14408), .C(new_n14407), .Y(new_n14691));
  XNOR2x2_ASAP7_75t_L       g14435(.A(new_n14691), .B(new_n14690), .Y(new_n14692));
  AOI22xp33_ASAP7_75t_L     g14436(.A1(new_n3029), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n3258), .Y(new_n14693));
  OAI221xp5_ASAP7_75t_L     g14437(.A1(new_n3024), .A2(new_n6812), .B1(new_n3256), .B2(new_n6837), .C(new_n14693), .Y(new_n14694));
  XNOR2x2_ASAP7_75t_L       g14438(.A(\a[32] ), .B(new_n14694), .Y(new_n14695));
  INVx1_ASAP7_75t_L         g14439(.A(new_n14695), .Y(new_n14696));
  MAJx2_ASAP7_75t_L         g14440(.A(new_n14515), .B(new_n14403), .C(new_n14401), .Y(new_n14697));
  XNOR2x2_ASAP7_75t_L       g14441(.A(new_n14696), .B(new_n14697), .Y(new_n14698));
  XNOR2x2_ASAP7_75t_L       g14442(.A(new_n14692), .B(new_n14698), .Y(new_n14699));
  XNOR2x2_ASAP7_75t_L       g14443(.A(new_n14699), .B(new_n14606), .Y(new_n14700));
  NOR2xp33_ASAP7_75t_L      g14444(.A(new_n14700), .B(new_n14599), .Y(new_n14701));
  AND2x2_ASAP7_75t_L        g14445(.A(new_n14700), .B(new_n14599), .Y(new_n14702));
  NOR2xp33_ASAP7_75t_L      g14446(.A(new_n14701), .B(new_n14702), .Y(new_n14703));
  INVx1_ASAP7_75t_L         g14447(.A(new_n14703), .Y(new_n14704));
  OA21x2_ASAP7_75t_L        g14448(.A1(new_n14592), .A2(new_n14594), .B(new_n14704), .Y(new_n14705));
  NOR3xp33_ASAP7_75t_L      g14449(.A(new_n14594), .B(new_n14704), .C(new_n14592), .Y(new_n14706));
  NOR2xp33_ASAP7_75t_L      g14450(.A(new_n14706), .B(new_n14705), .Y(new_n14707));
  INVx1_ASAP7_75t_L         g14451(.A(new_n14707), .Y(new_n14708));
  NAND3xp33_ASAP7_75t_L     g14452(.A(new_n14708), .B(new_n14586), .C(new_n14587), .Y(new_n14709));
  INVx1_ASAP7_75t_L         g14453(.A(new_n14587), .Y(new_n14710));
  OAI21xp33_ASAP7_75t_L     g14454(.A1(new_n14710), .A2(new_n14585), .B(new_n14707), .Y(new_n14711));
  NAND2xp33_ASAP7_75t_L     g14455(.A(new_n14711), .B(new_n14709), .Y(new_n14712));
  AOI21xp33_ASAP7_75t_L     g14456(.A1(new_n14580), .A2(new_n14577), .B(new_n14712), .Y(new_n14713));
  AND2x2_ASAP7_75t_L        g14457(.A(new_n14711), .B(new_n14709), .Y(new_n14714));
  NOR3xp33_ASAP7_75t_L      g14458(.A(new_n14714), .B(new_n14579), .C(new_n14576), .Y(new_n14715));
  OAI21xp33_ASAP7_75t_L     g14459(.A1(new_n14715), .A2(new_n14713), .B(new_n14568), .Y(new_n14716));
  OAI21xp33_ASAP7_75t_L     g14460(.A1(new_n14579), .A2(new_n14576), .B(new_n14714), .Y(new_n14717));
  NAND3xp33_ASAP7_75t_L     g14461(.A(new_n14580), .B(new_n14712), .C(new_n14577), .Y(new_n14718));
  OAI211xp5_ASAP7_75t_L     g14462(.A1(new_n14548), .A2(new_n14550), .B(new_n14717), .C(new_n14718), .Y(new_n14719));
  AND2x2_ASAP7_75t_L        g14463(.A(new_n14716), .B(new_n14719), .Y(new_n14720));
  A2O1A1Ixp33_ASAP7_75t_L   g14464(.A1(new_n14565), .A2(new_n14561), .B(new_n14554), .C(new_n14720), .Y(new_n14721));
  INVx1_ASAP7_75t_L         g14465(.A(new_n14721), .Y(new_n14722));
  INVx1_ASAP7_75t_L         g14466(.A(new_n14554), .Y(new_n14723));
  A2O1A1Ixp33_ASAP7_75t_L   g14467(.A1(new_n14351), .A2(new_n14564), .B(new_n14560), .C(new_n14723), .Y(new_n14724));
  NOR2xp33_ASAP7_75t_L      g14468(.A(new_n14720), .B(new_n14724), .Y(new_n14725));
  NOR2xp33_ASAP7_75t_L      g14469(.A(new_n14725), .B(new_n14722), .Y(\f[78] ));
  INVx1_ASAP7_75t_L         g14470(.A(new_n14719), .Y(new_n14727));
  OAI22xp33_ASAP7_75t_L     g14471(.A1(new_n11500), .A2(new_n1156), .B1(new_n11172), .B2(new_n1158), .Y(new_n14728));
  AOI21xp33_ASAP7_75t_L     g14472(.A1(new_n1080), .A2(\b[63] ), .B(new_n14728), .Y(new_n14729));
  NAND2xp33_ASAP7_75t_L     g14473(.A(\a[17] ), .B(new_n14729), .Y(new_n14730));
  A2O1A1Ixp33_ASAP7_75t_L   g14474(.A1(\b[63] ), .A2(new_n1080), .B(new_n14728), .C(new_n1071), .Y(new_n14731));
  NAND2xp33_ASAP7_75t_L     g14475(.A(new_n14731), .B(new_n14730), .Y(new_n14732));
  INVx1_ASAP7_75t_L         g14476(.A(new_n14732), .Y(new_n14733));
  O2A1O1Ixp33_ASAP7_75t_L   g14477(.A1(new_n14585), .A2(new_n14707), .B(new_n14587), .C(new_n14733), .Y(new_n14734));
  INVx1_ASAP7_75t_L         g14478(.A(new_n14734), .Y(new_n14735));
  O2A1O1Ixp33_ASAP7_75t_L   g14479(.A1(new_n14705), .A2(new_n14706), .B(new_n14586), .C(new_n14710), .Y(new_n14736));
  NAND2xp33_ASAP7_75t_L     g14480(.A(new_n14733), .B(new_n14736), .Y(new_n14737));
  AOI22xp33_ASAP7_75t_L     g14481(.A1(new_n1360), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1581), .Y(new_n14738));
  OAI221xp5_ASAP7_75t_L     g14482(.A1(new_n1373), .A2(new_n10250), .B1(new_n1359), .B2(new_n10855), .C(new_n14738), .Y(new_n14739));
  XNOR2x2_ASAP7_75t_L       g14483(.A(\a[20] ), .B(new_n14739), .Y(new_n14740));
  NOR2xp33_ASAP7_75t_L      g14484(.A(new_n14383), .B(new_n14593), .Y(new_n14741));
  MAJIxp5_ASAP7_75t_L       g14485(.A(new_n14741), .B(new_n14590), .C(new_n14704), .Y(new_n14742));
  INVx1_ASAP7_75t_L         g14486(.A(new_n14742), .Y(new_n14743));
  NAND2xp33_ASAP7_75t_L     g14487(.A(new_n14740), .B(new_n14743), .Y(new_n14744));
  INVx1_ASAP7_75t_L         g14488(.A(new_n14740), .Y(new_n14745));
  NAND2xp33_ASAP7_75t_L     g14489(.A(new_n14745), .B(new_n14742), .Y(new_n14746));
  A2O1A1O1Ixp25_ASAP7_75t_L g14490(.A1(new_n14527), .A2(new_n14528), .B(new_n14392), .C(new_n14393), .D(new_n14597), .Y(new_n14747));
  NOR2xp33_ASAP7_75t_L      g14491(.A(new_n14747), .B(new_n14701), .Y(new_n14748));
  AOI22xp33_ASAP7_75t_L     g14492(.A1(new_n1704), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n1837), .Y(new_n14749));
  OAI221xp5_ASAP7_75t_L     g14493(.A1(new_n1699), .A2(new_n9620), .B1(new_n1827), .B2(new_n9925), .C(new_n14749), .Y(new_n14750));
  XNOR2x2_ASAP7_75t_L       g14494(.A(\a[23] ), .B(new_n14750), .Y(new_n14751));
  NOR2xp33_ASAP7_75t_L      g14495(.A(new_n14751), .B(new_n14748), .Y(new_n14752));
  INVx1_ASAP7_75t_L         g14496(.A(new_n14752), .Y(new_n14753));
  NAND2xp33_ASAP7_75t_L     g14497(.A(new_n14751), .B(new_n14748), .Y(new_n14754));
  AOI22xp33_ASAP7_75t_L     g14498(.A1(new_n2114), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n2259), .Y(new_n14755));
  OAI221xp5_ASAP7_75t_L     g14499(.A1(new_n2109), .A2(new_n8458), .B1(new_n2257), .B2(new_n8768), .C(new_n14755), .Y(new_n14756));
  XNOR2x2_ASAP7_75t_L       g14500(.A(\a[26] ), .B(new_n14756), .Y(new_n14757));
  AOI21xp33_ASAP7_75t_L     g14501(.A1(new_n14606), .A2(new_n14699), .B(new_n14605), .Y(new_n14758));
  XNOR2x2_ASAP7_75t_L       g14502(.A(new_n14757), .B(new_n14758), .Y(new_n14759));
  AOI22xp33_ASAP7_75t_L     g14503(.A1(new_n2552), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n2736), .Y(new_n14760));
  OAI221xp5_ASAP7_75t_L     g14504(.A1(new_n2547), .A2(new_n7616), .B1(new_n2734), .B2(new_n7906), .C(new_n14760), .Y(new_n14761));
  XNOR2x2_ASAP7_75t_L       g14505(.A(\a[29] ), .B(new_n14761), .Y(new_n14762));
  INVx1_ASAP7_75t_L         g14506(.A(new_n14762), .Y(new_n14763));
  MAJx2_ASAP7_75t_L         g14507(.A(new_n14692), .B(new_n14696), .C(new_n14697), .Y(new_n14764));
  XNOR2x2_ASAP7_75t_L       g14508(.A(new_n14763), .B(new_n14764), .Y(new_n14765));
  INVx1_ASAP7_75t_L         g14509(.A(new_n14765), .Y(new_n14766));
  AOI22xp33_ASAP7_75t_L     g14510(.A1(new_n3029), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n3258), .Y(new_n14767));
  OAI221xp5_ASAP7_75t_L     g14511(.A1(new_n3024), .A2(new_n6830), .B1(new_n3256), .B2(new_n7323), .C(new_n14767), .Y(new_n14768));
  XNOR2x2_ASAP7_75t_L       g14512(.A(\a[32] ), .B(new_n14768), .Y(new_n14769));
  MAJIxp5_ASAP7_75t_L       g14513(.A(new_n14686), .B(new_n14689), .C(new_n14691), .Y(new_n14770));
  XNOR2x2_ASAP7_75t_L       g14514(.A(new_n14769), .B(new_n14770), .Y(new_n14771));
  INVx1_ASAP7_75t_L         g14515(.A(new_n14771), .Y(new_n14772));
  NOR2xp33_ASAP7_75t_L      g14516(.A(new_n14680), .B(new_n14677), .Y(new_n14773));
  AOI22xp33_ASAP7_75t_L     g14517(.A1(new_n4920), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n5167), .Y(new_n14774));
  OAI221xp5_ASAP7_75t_L     g14518(.A1(new_n5154), .A2(new_n4848), .B1(new_n5158), .B2(new_n11686), .C(new_n14774), .Y(new_n14775));
  XNOR2x2_ASAP7_75t_L       g14519(.A(\a[41] ), .B(new_n14775), .Y(new_n14776));
  INVx1_ASAP7_75t_L         g14520(.A(new_n14776), .Y(new_n14777));
  NOR2xp33_ASAP7_75t_L      g14521(.A(new_n14676), .B(new_n14675), .Y(new_n14778));
  AOI21xp33_ASAP7_75t_L     g14522(.A1(new_n14674), .A2(new_n14616), .B(new_n14778), .Y(new_n14779));
  AOI22xp33_ASAP7_75t_L     g14523(.A1(new_n5624), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n5901), .Y(new_n14780));
  OAI221xp5_ASAP7_75t_L     g14524(.A1(new_n5900), .A2(new_n4216), .B1(new_n5892), .B2(new_n4431), .C(new_n14780), .Y(new_n14781));
  XNOR2x2_ASAP7_75t_L       g14525(.A(\a[44] ), .B(new_n14781), .Y(new_n14782));
  INVx1_ASAP7_75t_L         g14526(.A(new_n14663), .Y(new_n14783));
  INVx1_ASAP7_75t_L         g14527(.A(new_n14666), .Y(new_n14784));
  NOR3xp33_ASAP7_75t_L      g14528(.A(new_n14667), .B(new_n14672), .C(new_n14668), .Y(new_n14785));
  AOI21xp33_ASAP7_75t_L     g14529(.A1(new_n14784), .A2(new_n14783), .B(new_n14785), .Y(new_n14786));
  INVx1_ASAP7_75t_L         g14530(.A(new_n14651), .Y(new_n14787));
  INVx1_ASAP7_75t_L         g14531(.A(new_n11247), .Y(new_n14788));
  INVx1_ASAP7_75t_L         g14532(.A(new_n11249), .Y(new_n14789));
  INVx1_ASAP7_75t_L         g14533(.A(new_n14422), .Y(new_n14790));
  A2O1A1Ixp33_ASAP7_75t_L   g14534(.A1(new_n14788), .A2(new_n14789), .B(new_n869), .C(new_n14790), .Y(new_n14791));
  A2O1A1Ixp33_ASAP7_75t_L   g14535(.A1(new_n14791), .A2(new_n14235), .B(new_n14433), .C(new_n14633), .Y(new_n14792));
  OAI31xp33_ASAP7_75t_L     g14536(.A1(new_n14623), .A2(new_n14631), .A3(new_n14630), .B(new_n14792), .Y(new_n14793));
  NOR2xp33_ASAP7_75t_L      g14537(.A(new_n942), .B(new_n11535), .Y(new_n14794));
  A2O1A1O1Ixp25_ASAP7_75t_L g14538(.A1(new_n11533), .A2(\b[15] ), .B(new_n14624), .C(new_n806), .D(new_n14630), .Y(new_n14795));
  A2O1A1Ixp33_ASAP7_75t_L   g14539(.A1(new_n11533), .A2(\b[16] ), .B(new_n14794), .C(new_n14795), .Y(new_n14796));
  O2A1O1Ixp33_ASAP7_75t_L   g14540(.A1(new_n11247), .A2(new_n11249), .B(\b[16] ), .C(new_n14794), .Y(new_n14797));
  INVx1_ASAP7_75t_L         g14541(.A(new_n14797), .Y(new_n14798));
  A2O1A1Ixp33_ASAP7_75t_L   g14542(.A1(new_n11533), .A2(\b[15] ), .B(new_n14624), .C(new_n806), .Y(new_n14799));
  A2O1A1O1Ixp25_ASAP7_75t_L g14543(.A1(new_n14627), .A2(new_n14626), .B(new_n14235), .C(new_n14799), .D(new_n14798), .Y(new_n14800));
  INVx1_ASAP7_75t_L         g14544(.A(new_n14800), .Y(new_n14801));
  NAND2xp33_ASAP7_75t_L     g14545(.A(new_n14801), .B(new_n14796), .Y(new_n14802));
  NOR2xp33_ASAP7_75t_L      g14546(.A(new_n1432), .B(new_n10630), .Y(new_n14803));
  AOI221xp5_ASAP7_75t_L     g14547(.A1(\b[17] ), .A2(new_n10939), .B1(\b[18] ), .B2(new_n10632), .C(new_n14803), .Y(new_n14804));
  OAI211xp5_ASAP7_75t_L     g14548(.A1(new_n10629), .A2(new_n1438), .B(\a[62] ), .C(new_n14804), .Y(new_n14805));
  O2A1O1Ixp33_ASAP7_75t_L   g14549(.A1(new_n10629), .A2(new_n1438), .B(new_n14804), .C(\a[62] ), .Y(new_n14806));
  INVx1_ASAP7_75t_L         g14550(.A(new_n14806), .Y(new_n14807));
  AO21x2_ASAP7_75t_L        g14551(.A1(new_n14805), .A2(new_n14807), .B(new_n14802), .Y(new_n14808));
  NAND3xp33_ASAP7_75t_L     g14552(.A(new_n14807), .B(new_n14805), .C(new_n14802), .Y(new_n14809));
  NAND2xp33_ASAP7_75t_L     g14553(.A(new_n14809), .B(new_n14808), .Y(new_n14810));
  INVx1_ASAP7_75t_L         g14554(.A(new_n14810), .Y(new_n14811));
  NAND2xp33_ASAP7_75t_L     g14555(.A(new_n14811), .B(new_n14793), .Y(new_n14812));
  NOR2xp33_ASAP7_75t_L      g14556(.A(new_n14811), .B(new_n14793), .Y(new_n14813));
  INVx1_ASAP7_75t_L         g14557(.A(new_n14813), .Y(new_n14814));
  AOI22xp33_ASAP7_75t_L     g14558(.A1(new_n9700), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n10027), .Y(new_n14815));
  OAI221xp5_ASAP7_75t_L     g14559(.A1(new_n10024), .A2(new_n1655), .B1(new_n9696), .B2(new_n1780), .C(new_n14815), .Y(new_n14816));
  XNOR2x2_ASAP7_75t_L       g14560(.A(\a[59] ), .B(new_n14816), .Y(new_n14817));
  AND3x1_ASAP7_75t_L        g14561(.A(new_n14814), .B(new_n14817), .C(new_n14812), .Y(new_n14818));
  INVx1_ASAP7_75t_L         g14562(.A(new_n14818), .Y(new_n14819));
  AO21x2_ASAP7_75t_L        g14563(.A1(new_n14812), .A2(new_n14814), .B(new_n14817), .Y(new_n14820));
  NAND2xp33_ASAP7_75t_L     g14564(.A(new_n14820), .B(new_n14819), .Y(new_n14821));
  OAI21xp33_ASAP7_75t_L     g14565(.A1(new_n14635), .A2(new_n14638), .B(new_n14641), .Y(new_n14822));
  OR2x4_ASAP7_75t_L         g14566(.A(new_n14822), .B(new_n14821), .Y(new_n14823));
  NAND2xp33_ASAP7_75t_L     g14567(.A(new_n14822), .B(new_n14821), .Y(new_n14824));
  NAND2xp33_ASAP7_75t_L     g14568(.A(\b[23] ), .B(new_n9115), .Y(new_n14825));
  OAI221xp5_ASAP7_75t_L     g14569(.A1(new_n9113), .A2(new_n2067), .B1(new_n10016), .B2(new_n2075), .C(new_n14825), .Y(new_n14826));
  AOI21xp33_ASAP7_75t_L     g14570(.A1(new_n8835), .A2(\b[24] ), .B(new_n14826), .Y(new_n14827));
  NAND2xp33_ASAP7_75t_L     g14571(.A(\a[56] ), .B(new_n14827), .Y(new_n14828));
  A2O1A1Ixp33_ASAP7_75t_L   g14572(.A1(\b[24] ), .A2(new_n8835), .B(new_n14826), .C(new_n8826), .Y(new_n14829));
  NAND4xp25_ASAP7_75t_L     g14573(.A(new_n14823), .B(new_n14829), .C(new_n14828), .D(new_n14824), .Y(new_n14830));
  NAND2xp33_ASAP7_75t_L     g14574(.A(new_n14824), .B(new_n14823), .Y(new_n14831));
  NAND2xp33_ASAP7_75t_L     g14575(.A(new_n14829), .B(new_n14828), .Y(new_n14832));
  NAND2xp33_ASAP7_75t_L     g14576(.A(new_n14832), .B(new_n14831), .Y(new_n14833));
  NAND2xp33_ASAP7_75t_L     g14577(.A(new_n14830), .B(new_n14833), .Y(new_n14834));
  O2A1O1Ixp33_ASAP7_75t_L   g14578(.A1(new_n14642), .A2(new_n14645), .B(new_n14787), .C(new_n14834), .Y(new_n14835));
  INVx1_ASAP7_75t_L         g14579(.A(new_n14834), .Y(new_n14836));
  NOR3xp33_ASAP7_75t_L      g14580(.A(new_n14836), .B(new_n14651), .C(new_n14646), .Y(new_n14837));
  NOR2xp33_ASAP7_75t_L      g14581(.A(new_n14835), .B(new_n14837), .Y(new_n14838));
  NAND2xp33_ASAP7_75t_L     g14582(.A(\b[26] ), .B(new_n8537), .Y(new_n14839));
  OAI221xp5_ASAP7_75t_L     g14583(.A1(new_n8243), .A2(new_n2666), .B1(new_n7957), .B2(new_n2672), .C(new_n14839), .Y(new_n14840));
  AOI21xp33_ASAP7_75t_L     g14584(.A1(new_n7963), .A2(\b[27] ), .B(new_n14840), .Y(new_n14841));
  NAND2xp33_ASAP7_75t_L     g14585(.A(\a[53] ), .B(new_n14841), .Y(new_n14842));
  A2O1A1Ixp33_ASAP7_75t_L   g14586(.A1(\b[27] ), .A2(new_n7963), .B(new_n14840), .C(new_n7954), .Y(new_n14843));
  AND2x2_ASAP7_75t_L        g14587(.A(new_n14843), .B(new_n14842), .Y(new_n14844));
  NAND2xp33_ASAP7_75t_L     g14588(.A(new_n14844), .B(new_n14838), .Y(new_n14845));
  INVx1_ASAP7_75t_L         g14589(.A(new_n14844), .Y(new_n14846));
  OAI21xp33_ASAP7_75t_L     g14590(.A1(new_n14835), .A2(new_n14837), .B(new_n14846), .Y(new_n14847));
  OAI21xp33_ASAP7_75t_L     g14591(.A1(new_n14462), .A2(new_n14464), .B(new_n14653), .Y(new_n14848));
  INVx1_ASAP7_75t_L         g14592(.A(new_n14619), .Y(new_n14849));
  NAND2xp33_ASAP7_75t_L     g14593(.A(new_n14849), .B(new_n14652), .Y(new_n14850));
  NAND2xp33_ASAP7_75t_L     g14594(.A(new_n14850), .B(new_n14848), .Y(new_n14851));
  NAND3xp33_ASAP7_75t_L     g14595(.A(new_n14845), .B(new_n14847), .C(new_n14851), .Y(new_n14852));
  AO21x2_ASAP7_75t_L        g14596(.A1(new_n14847), .A2(new_n14845), .B(new_n14851), .Y(new_n14853));
  NAND2xp33_ASAP7_75t_L     g14597(.A(new_n14852), .B(new_n14853), .Y(new_n14854));
  NAND2xp33_ASAP7_75t_L     g14598(.A(\b[29] ), .B(new_n7391), .Y(new_n14855));
  OAI221xp5_ASAP7_75t_L     g14599(.A1(new_n7389), .A2(new_n3180), .B1(new_n8237), .B2(new_n3187), .C(new_n14855), .Y(new_n14856));
  AOI21xp33_ASAP7_75t_L     g14600(.A1(new_n7115), .A2(\b[30] ), .B(new_n14856), .Y(new_n14857));
  NAND2xp33_ASAP7_75t_L     g14601(.A(\a[50] ), .B(new_n14857), .Y(new_n14858));
  A2O1A1Ixp33_ASAP7_75t_L   g14602(.A1(\b[30] ), .A2(new_n7115), .B(new_n14856), .C(new_n7106), .Y(new_n14859));
  NAND2xp33_ASAP7_75t_L     g14603(.A(new_n14859), .B(new_n14858), .Y(new_n14860));
  XNOR2x2_ASAP7_75t_L       g14604(.A(new_n14860), .B(new_n14854), .Y(new_n14861));
  INVx1_ASAP7_75t_L         g14605(.A(new_n14662), .Y(new_n14862));
  NOR2xp33_ASAP7_75t_L      g14606(.A(new_n14660), .B(new_n14862), .Y(new_n14863));
  AOI21xp33_ASAP7_75t_L     g14607(.A1(new_n14659), .A2(new_n14655), .B(new_n14863), .Y(new_n14864));
  XNOR2x2_ASAP7_75t_L       g14608(.A(new_n14861), .B(new_n14864), .Y(new_n14865));
  AOI22xp33_ASAP7_75t_L     g14609(.A1(new_n6376), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n6648), .Y(new_n14866));
  OAI221xp5_ASAP7_75t_L     g14610(.A1(new_n6646), .A2(new_n3565), .B1(new_n6636), .B2(new_n3591), .C(new_n14866), .Y(new_n14867));
  XNOR2x2_ASAP7_75t_L       g14611(.A(\a[47] ), .B(new_n14867), .Y(new_n14868));
  XNOR2x2_ASAP7_75t_L       g14612(.A(new_n14868), .B(new_n14865), .Y(new_n14869));
  XNOR2x2_ASAP7_75t_L       g14613(.A(new_n14786), .B(new_n14869), .Y(new_n14870));
  XNOR2x2_ASAP7_75t_L       g14614(.A(new_n14782), .B(new_n14870), .Y(new_n14871));
  XNOR2x2_ASAP7_75t_L       g14615(.A(new_n14779), .B(new_n14871), .Y(new_n14872));
  AND2x2_ASAP7_75t_L        g14616(.A(new_n14777), .B(new_n14872), .Y(new_n14873));
  NOR2xp33_ASAP7_75t_L      g14617(.A(new_n14777), .B(new_n14872), .Y(new_n14874));
  NOR2xp33_ASAP7_75t_L      g14618(.A(new_n14874), .B(new_n14873), .Y(new_n14875));
  A2O1A1Ixp33_ASAP7_75t_L   g14619(.A1(new_n14681), .A2(new_n14612), .B(new_n14773), .C(new_n14875), .Y(new_n14876));
  INVx1_ASAP7_75t_L         g14620(.A(new_n14294), .Y(new_n14877));
  O2A1O1Ixp33_ASAP7_75t_L   g14621(.A1(new_n14877), .A2(new_n14296), .B(new_n14499), .C(new_n14611), .Y(new_n14878));
  A2O1A1O1Ixp25_ASAP7_75t_L g14622(.A1(new_n14501), .A2(new_n14507), .B(new_n14878), .C(new_n14681), .D(new_n14773), .Y(new_n14879));
  OAI21xp33_ASAP7_75t_L     g14623(.A1(new_n14874), .A2(new_n14873), .B(new_n14879), .Y(new_n14880));
  NAND2xp33_ASAP7_75t_L     g14624(.A(new_n14880), .B(new_n14876), .Y(new_n14881));
  NAND2xp33_ASAP7_75t_L     g14625(.A(\b[41] ), .B(new_n4512), .Y(new_n14882));
  OAI221xp5_ASAP7_75t_L     g14626(.A1(new_n4275), .A2(new_n5805), .B1(new_n4499), .B2(new_n6338), .C(new_n14882), .Y(new_n14883));
  AOI21xp33_ASAP7_75t_L     g14627(.A1(new_n4285), .A2(\b[42] ), .B(new_n14883), .Y(new_n14884));
  NAND2xp33_ASAP7_75t_L     g14628(.A(\a[38] ), .B(new_n14884), .Y(new_n14885));
  A2O1A1Ixp33_ASAP7_75t_L   g14629(.A1(\b[42] ), .A2(new_n4285), .B(new_n14883), .C(new_n4268), .Y(new_n14886));
  NAND2xp33_ASAP7_75t_L     g14630(.A(new_n14886), .B(new_n14885), .Y(new_n14887));
  XNOR2x2_ASAP7_75t_L       g14631(.A(new_n14887), .B(new_n14881), .Y(new_n14888));
  A2O1A1Ixp33_ASAP7_75t_L   g14632(.A1(new_n14509), .A2(new_n14511), .B(new_n14685), .C(new_n14683), .Y(new_n14889));
  XNOR2x2_ASAP7_75t_L       g14633(.A(new_n14889), .B(new_n14888), .Y(new_n14890));
  AOI22xp33_ASAP7_75t_L     g14634(.A1(new_n3633), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n3858), .Y(new_n14891));
  OAI221xp5_ASAP7_75t_L     g14635(.A1(new_n3853), .A2(new_n6321), .B1(new_n3856), .B2(new_n6573), .C(new_n14891), .Y(new_n14892));
  XNOR2x2_ASAP7_75t_L       g14636(.A(\a[35] ), .B(new_n14892), .Y(new_n14893));
  INVx1_ASAP7_75t_L         g14637(.A(new_n14893), .Y(new_n14894));
  OR2x4_ASAP7_75t_L         g14638(.A(new_n14894), .B(new_n14890), .Y(new_n14895));
  NAND2xp33_ASAP7_75t_L     g14639(.A(new_n14894), .B(new_n14890), .Y(new_n14896));
  NAND2xp33_ASAP7_75t_L     g14640(.A(new_n14896), .B(new_n14895), .Y(new_n14897));
  XNOR2x2_ASAP7_75t_L       g14641(.A(new_n14772), .B(new_n14897), .Y(new_n14898));
  AND2x2_ASAP7_75t_L        g14642(.A(new_n14898), .B(new_n14766), .Y(new_n14899));
  NOR2xp33_ASAP7_75t_L      g14643(.A(new_n14898), .B(new_n14766), .Y(new_n14900));
  NOR2xp33_ASAP7_75t_L      g14644(.A(new_n14900), .B(new_n14899), .Y(new_n14901));
  INVx1_ASAP7_75t_L         g14645(.A(new_n14901), .Y(new_n14902));
  NOR2xp33_ASAP7_75t_L      g14646(.A(new_n14902), .B(new_n14759), .Y(new_n14903));
  AND2x2_ASAP7_75t_L        g14647(.A(new_n14902), .B(new_n14759), .Y(new_n14904));
  NOR2xp33_ASAP7_75t_L      g14648(.A(new_n14903), .B(new_n14904), .Y(new_n14905));
  NAND3xp33_ASAP7_75t_L     g14649(.A(new_n14753), .B(new_n14754), .C(new_n14905), .Y(new_n14906));
  AO21x2_ASAP7_75t_L        g14650(.A1(new_n14754), .A2(new_n14753), .B(new_n14905), .Y(new_n14907));
  AND2x2_ASAP7_75t_L        g14651(.A(new_n14906), .B(new_n14907), .Y(new_n14908));
  AND3x1_ASAP7_75t_L        g14652(.A(new_n14908), .B(new_n14744), .C(new_n14746), .Y(new_n14909));
  AOI21xp33_ASAP7_75t_L     g14653(.A1(new_n14744), .A2(new_n14746), .B(new_n14908), .Y(new_n14910));
  NOR2xp33_ASAP7_75t_L      g14654(.A(new_n14910), .B(new_n14909), .Y(new_n14911));
  INVx1_ASAP7_75t_L         g14655(.A(new_n14911), .Y(new_n14912));
  NAND3xp33_ASAP7_75t_L     g14656(.A(new_n14912), .B(new_n14735), .C(new_n14737), .Y(new_n14913));
  NAND2xp33_ASAP7_75t_L     g14657(.A(new_n14735), .B(new_n14737), .Y(new_n14914));
  NAND2xp33_ASAP7_75t_L     g14658(.A(new_n14911), .B(new_n14914), .Y(new_n14915));
  A2O1A1O1Ixp25_ASAP7_75t_L g14659(.A1(new_n14364), .A2(new_n14365), .B(new_n14360), .C(new_n14536), .D(new_n14574), .Y(new_n14916));
  O2A1O1Ixp33_ASAP7_75t_L   g14660(.A1(new_n14576), .A2(new_n14579), .B(new_n14714), .C(new_n14916), .Y(new_n14917));
  AND3x1_ASAP7_75t_L        g14661(.A(new_n14913), .B(new_n14915), .C(new_n14917), .Y(new_n14918));
  AOI21xp33_ASAP7_75t_L     g14662(.A1(new_n14913), .A2(new_n14915), .B(new_n14917), .Y(new_n14919));
  NOR2xp33_ASAP7_75t_L      g14663(.A(new_n14919), .B(new_n14918), .Y(new_n14920));
  A2O1A1Ixp33_ASAP7_75t_L   g14664(.A1(new_n14724), .A2(new_n14720), .B(new_n14727), .C(new_n14920), .Y(new_n14921));
  INVx1_ASAP7_75t_L         g14665(.A(new_n14921), .Y(new_n14922));
  NAND2xp33_ASAP7_75t_L     g14666(.A(new_n14716), .B(new_n14719), .Y(new_n14923));
  A2O1A1Ixp33_ASAP7_75t_L   g14667(.A1(new_n14562), .A2(new_n14723), .B(new_n14923), .C(new_n14719), .Y(new_n14924));
  NOR2xp33_ASAP7_75t_L      g14668(.A(new_n14920), .B(new_n14924), .Y(new_n14925));
  NOR2xp33_ASAP7_75t_L      g14669(.A(new_n14925), .B(new_n14922), .Y(\f[79] ));
  AOI22xp33_ASAP7_75t_L     g14670(.A1(new_n1360), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n1581), .Y(new_n14927));
  OAI221xp5_ASAP7_75t_L     g14671(.A1(new_n1373), .A2(new_n10847), .B1(new_n1359), .B2(new_n12047), .C(new_n14927), .Y(new_n14928));
  XNOR2x2_ASAP7_75t_L       g14672(.A(\a[20] ), .B(new_n14928), .Y(new_n14929));
  INVx1_ASAP7_75t_L         g14673(.A(new_n14929), .Y(new_n14930));
  NAND2xp33_ASAP7_75t_L     g14674(.A(new_n14753), .B(new_n14906), .Y(new_n14931));
  NOR2xp33_ASAP7_75t_L      g14675(.A(new_n14930), .B(new_n14931), .Y(new_n14932));
  A2O1A1Ixp33_ASAP7_75t_L   g14676(.A1(new_n14754), .A2(new_n14905), .B(new_n14752), .C(new_n14930), .Y(new_n14933));
  INVx1_ASAP7_75t_L         g14677(.A(new_n14933), .Y(new_n14934));
  AOI22xp33_ASAP7_75t_L     g14678(.A1(new_n1704), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1837), .Y(new_n14935));
  OAI221xp5_ASAP7_75t_L     g14679(.A1(new_n1699), .A2(new_n9920), .B1(new_n1827), .B2(new_n11152), .C(new_n14935), .Y(new_n14936));
  XNOR2x2_ASAP7_75t_L       g14680(.A(\a[23] ), .B(new_n14936), .Y(new_n14937));
  MAJIxp5_ASAP7_75t_L       g14681(.A(new_n14902), .B(new_n14757), .C(new_n14758), .Y(new_n14938));
  XNOR2x2_ASAP7_75t_L       g14682(.A(new_n14937), .B(new_n14938), .Y(new_n14939));
  AOI22xp33_ASAP7_75t_L     g14683(.A1(new_n2114), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n2259), .Y(new_n14940));
  OAI221xp5_ASAP7_75t_L     g14684(.A1(new_n2109), .A2(new_n8762), .B1(new_n2257), .B2(new_n9331), .C(new_n14940), .Y(new_n14941));
  XNOR2x2_ASAP7_75t_L       g14685(.A(\a[26] ), .B(new_n14941), .Y(new_n14942));
  AOI21xp33_ASAP7_75t_L     g14686(.A1(new_n14764), .A2(new_n14763), .B(new_n14899), .Y(new_n14943));
  AND2x2_ASAP7_75t_L        g14687(.A(new_n14942), .B(new_n14943), .Y(new_n14944));
  NOR2xp33_ASAP7_75t_L      g14688(.A(new_n14942), .B(new_n14943), .Y(new_n14945));
  NOR2xp33_ASAP7_75t_L      g14689(.A(new_n14945), .B(new_n14944), .Y(new_n14946));
  AOI22xp33_ASAP7_75t_L     g14690(.A1(new_n2552), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n2736), .Y(new_n14947));
  OAI221xp5_ASAP7_75t_L     g14691(.A1(new_n2547), .A2(new_n7900), .B1(new_n2734), .B2(new_n8174), .C(new_n14947), .Y(new_n14948));
  NOR2xp33_ASAP7_75t_L      g14692(.A(new_n2538), .B(new_n14948), .Y(new_n14949));
  AND2x2_ASAP7_75t_L        g14693(.A(new_n2538), .B(new_n14948), .Y(new_n14950));
  NOR2xp33_ASAP7_75t_L      g14694(.A(new_n14949), .B(new_n14950), .Y(new_n14951));
  INVx1_ASAP7_75t_L         g14695(.A(new_n14769), .Y(new_n14952));
  NAND2xp33_ASAP7_75t_L     g14696(.A(new_n14952), .B(new_n14770), .Y(new_n14953));
  A2O1A1Ixp33_ASAP7_75t_L   g14697(.A1(new_n14895), .A2(new_n14896), .B(new_n14772), .C(new_n14953), .Y(new_n14954));
  NOR2xp33_ASAP7_75t_L      g14698(.A(new_n14951), .B(new_n14954), .Y(new_n14955));
  INVx1_ASAP7_75t_L         g14699(.A(new_n14951), .Y(new_n14956));
  A2O1A1O1Ixp25_ASAP7_75t_L g14700(.A1(new_n14896), .A2(new_n14895), .B(new_n14772), .C(new_n14953), .D(new_n14956), .Y(new_n14957));
  NOR2xp33_ASAP7_75t_L      g14701(.A(new_n14957), .B(new_n14955), .Y(new_n14958));
  AOI22xp33_ASAP7_75t_L     g14702(.A1(new_n3029), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n3258), .Y(new_n14959));
  OAI221xp5_ASAP7_75t_L     g14703(.A1(new_n3024), .A2(new_n7317), .B1(new_n3256), .B2(new_n7602), .C(new_n14959), .Y(new_n14960));
  XNOR2x2_ASAP7_75t_L       g14704(.A(\a[32] ), .B(new_n14960), .Y(new_n14961));
  MAJx2_ASAP7_75t_L         g14705(.A(new_n14888), .B(new_n14889), .C(new_n14894), .Y(new_n14962));
  INVx1_ASAP7_75t_L         g14706(.A(new_n14962), .Y(new_n14963));
  AND2x2_ASAP7_75t_L        g14707(.A(new_n14961), .B(new_n14963), .Y(new_n14964));
  NOR2xp33_ASAP7_75t_L      g14708(.A(new_n14961), .B(new_n14963), .Y(new_n14965));
  NOR2xp33_ASAP7_75t_L      g14709(.A(new_n14965), .B(new_n14964), .Y(new_n14966));
  AOI22xp33_ASAP7_75t_L     g14710(.A1(new_n4283), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n4512), .Y(new_n14967));
  OAI221xp5_ASAP7_75t_L     g14711(.A1(new_n4277), .A2(new_n5805), .B1(new_n4499), .B2(new_n5835), .C(new_n14967), .Y(new_n14968));
  XNOR2x2_ASAP7_75t_L       g14712(.A(\a[38] ), .B(new_n14968), .Y(new_n14969));
  INVx1_ASAP7_75t_L         g14713(.A(new_n14969), .Y(new_n14970));
  A2O1A1O1Ixp25_ASAP7_75t_L g14714(.A1(new_n14674), .A2(new_n14616), .B(new_n14778), .C(new_n14871), .D(new_n14873), .Y(new_n14971));
  AOI22xp33_ASAP7_75t_L     g14715(.A1(new_n4920), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n5167), .Y(new_n14972));
  OAI221xp5_ASAP7_75t_L     g14716(.A1(new_n5154), .A2(new_n4869), .B1(new_n5158), .B2(new_n5327), .C(new_n14972), .Y(new_n14973));
  XNOR2x2_ASAP7_75t_L       g14717(.A(\a[41] ), .B(new_n14973), .Y(new_n14974));
  INVx1_ASAP7_75t_L         g14718(.A(new_n14974), .Y(new_n14975));
  A2O1A1Ixp33_ASAP7_75t_L   g14719(.A1(new_n14784), .A2(new_n14783), .B(new_n14785), .C(new_n14869), .Y(new_n14976));
  INVx1_ASAP7_75t_L         g14720(.A(new_n14870), .Y(new_n14977));
  OAI21xp33_ASAP7_75t_L     g14721(.A1(new_n14782), .A2(new_n14977), .B(new_n14976), .Y(new_n14978));
  AOI22xp33_ASAP7_75t_L     g14722(.A1(new_n5624), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n5901), .Y(new_n14979));
  OAI221xp5_ASAP7_75t_L     g14723(.A1(new_n5900), .A2(new_n4424), .B1(new_n5892), .B2(new_n4641), .C(new_n14979), .Y(new_n14980));
  XNOR2x2_ASAP7_75t_L       g14724(.A(\a[44] ), .B(new_n14980), .Y(new_n14981));
  INVx1_ASAP7_75t_L         g14725(.A(new_n14981), .Y(new_n14982));
  A2O1A1Ixp33_ASAP7_75t_L   g14726(.A1(new_n14659), .A2(new_n14655), .B(new_n14863), .C(new_n14861), .Y(new_n14983));
  INVx1_ASAP7_75t_L         g14727(.A(new_n14865), .Y(new_n14984));
  INVx1_ASAP7_75t_L         g14728(.A(new_n14852), .Y(new_n14985));
  AOI22xp33_ASAP7_75t_L     g14729(.A1(new_n7111), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n7391), .Y(new_n14986));
  OAI221xp5_ASAP7_75t_L     g14730(.A1(new_n8558), .A2(new_n3180), .B1(new_n8237), .B2(new_n11047), .C(new_n14986), .Y(new_n14987));
  XNOR2x2_ASAP7_75t_L       g14731(.A(\a[50] ), .B(new_n14987), .Y(new_n14988));
  AOI22xp33_ASAP7_75t_L     g14732(.A1(new_n8831), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n9115), .Y(new_n14989));
  OAI221xp5_ASAP7_75t_L     g14733(.A1(new_n10343), .A2(new_n2067), .B1(new_n10016), .B2(new_n2355), .C(new_n14989), .Y(new_n14990));
  XNOR2x2_ASAP7_75t_L       g14734(.A(\a[56] ), .B(new_n14990), .Y(new_n14991));
  A2O1A1Ixp33_ASAP7_75t_L   g14735(.A1(new_n14807), .A2(new_n14805), .B(new_n14802), .C(new_n14801), .Y(new_n14992));
  AOI22xp33_ASAP7_75t_L     g14736(.A1(\b[18] ), .A2(new_n10939), .B1(\b[20] ), .B2(new_n10938), .Y(new_n14993));
  OAI221xp5_ASAP7_75t_L     g14737(.A1(new_n10937), .A2(new_n1432), .B1(new_n10629), .B2(new_n1547), .C(new_n14993), .Y(new_n14994));
  XNOR2x2_ASAP7_75t_L       g14738(.A(\a[62] ), .B(new_n14994), .Y(new_n14995));
  NOR2xp33_ASAP7_75t_L      g14739(.A(new_n1030), .B(new_n11535), .Y(new_n14996));
  A2O1A1Ixp33_ASAP7_75t_L   g14740(.A1(\b[17] ), .A2(new_n11533), .B(new_n14996), .C(new_n14797), .Y(new_n14997));
  O2A1O1Ixp33_ASAP7_75t_L   g14741(.A1(new_n11247), .A2(new_n11249), .B(\b[17] ), .C(new_n14996), .Y(new_n14998));
  A2O1A1Ixp33_ASAP7_75t_L   g14742(.A1(new_n11533), .A2(\b[16] ), .B(new_n14794), .C(new_n14998), .Y(new_n14999));
  AND2x2_ASAP7_75t_L        g14743(.A(new_n14997), .B(new_n14999), .Y(new_n15000));
  XOR2x2_ASAP7_75t_L        g14744(.A(new_n15000), .B(new_n14995), .Y(new_n15001));
  XOR2x2_ASAP7_75t_L        g14745(.A(new_n14992), .B(new_n15001), .Y(new_n15002));
  AOI22xp33_ASAP7_75t_L     g14746(.A1(new_n9700), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n10027), .Y(new_n15003));
  OAI221xp5_ASAP7_75t_L     g14747(.A1(new_n10024), .A2(new_n1774), .B1(new_n9696), .B2(new_n1915), .C(new_n15003), .Y(new_n15004));
  XNOR2x2_ASAP7_75t_L       g14748(.A(\a[59] ), .B(new_n15004), .Y(new_n15005));
  NAND2xp33_ASAP7_75t_L     g14749(.A(new_n15005), .B(new_n15002), .Y(new_n15006));
  NOR2xp33_ASAP7_75t_L      g14750(.A(new_n15005), .B(new_n15002), .Y(new_n15007));
  INVx1_ASAP7_75t_L         g14751(.A(new_n15007), .Y(new_n15008));
  NAND2xp33_ASAP7_75t_L     g14752(.A(new_n15006), .B(new_n15008), .Y(new_n15009));
  INVx1_ASAP7_75t_L         g14753(.A(new_n15009), .Y(new_n15010));
  NOR2xp33_ASAP7_75t_L      g14754(.A(new_n14813), .B(new_n14818), .Y(new_n15011));
  NAND2xp33_ASAP7_75t_L     g14755(.A(new_n15011), .B(new_n15010), .Y(new_n15012));
  INVx1_ASAP7_75t_L         g14756(.A(new_n15012), .Y(new_n15013));
  O2A1O1Ixp33_ASAP7_75t_L   g14757(.A1(new_n14793), .A2(new_n14811), .B(new_n14819), .C(new_n15010), .Y(new_n15014));
  NOR3xp33_ASAP7_75t_L      g14758(.A(new_n15013), .B(new_n15014), .C(new_n14991), .Y(new_n15015));
  INVx1_ASAP7_75t_L         g14759(.A(new_n14991), .Y(new_n15016));
  A2O1A1Ixp33_ASAP7_75t_L   g14760(.A1(new_n14817), .A2(new_n14812), .B(new_n14813), .C(new_n15009), .Y(new_n15017));
  AOI21xp33_ASAP7_75t_L     g14761(.A1(new_n15012), .A2(new_n15017), .B(new_n15016), .Y(new_n15018));
  NAND2xp33_ASAP7_75t_L     g14762(.A(new_n14823), .B(new_n14830), .Y(new_n15019));
  NOR3xp33_ASAP7_75t_L      g14763(.A(new_n15019), .B(new_n15018), .C(new_n15015), .Y(new_n15020));
  NOR2xp33_ASAP7_75t_L      g14764(.A(new_n15018), .B(new_n15015), .Y(new_n15021));
  O2A1O1Ixp33_ASAP7_75t_L   g14765(.A1(new_n14831), .A2(new_n14832), .B(new_n14823), .C(new_n15021), .Y(new_n15022));
  NOR2xp33_ASAP7_75t_L      g14766(.A(new_n15020), .B(new_n15022), .Y(new_n15023));
  AOI22xp33_ASAP7_75t_L     g14767(.A1(new_n7960), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n8537), .Y(new_n15024));
  OAI221xp5_ASAP7_75t_L     g14768(.A1(new_n8817), .A2(new_n2666), .B1(new_n7957), .B2(new_n2695), .C(new_n15024), .Y(new_n15025));
  XNOR2x2_ASAP7_75t_L       g14769(.A(\a[53] ), .B(new_n15025), .Y(new_n15026));
  XNOR2x2_ASAP7_75t_L       g14770(.A(new_n15026), .B(new_n15023), .Y(new_n15027));
  O2A1O1Ixp33_ASAP7_75t_L   g14771(.A1(new_n14642), .A2(new_n14645), .B(new_n14787), .C(new_n14836), .Y(new_n15028));
  O2A1O1Ixp33_ASAP7_75t_L   g14772(.A1(new_n14835), .A2(new_n14837), .B(new_n14846), .C(new_n15028), .Y(new_n15029));
  INVx1_ASAP7_75t_L         g14773(.A(new_n15029), .Y(new_n15030));
  NAND2xp33_ASAP7_75t_L     g14774(.A(new_n15027), .B(new_n15030), .Y(new_n15031));
  NOR2xp33_ASAP7_75t_L      g14775(.A(new_n15027), .B(new_n15030), .Y(new_n15032));
  INVx1_ASAP7_75t_L         g14776(.A(new_n15032), .Y(new_n15033));
  NAND3xp33_ASAP7_75t_L     g14777(.A(new_n15033), .B(new_n15031), .C(new_n14988), .Y(new_n15034));
  AO21x2_ASAP7_75t_L        g14778(.A1(new_n15031), .A2(new_n15033), .B(new_n14988), .Y(new_n15035));
  NAND2xp33_ASAP7_75t_L     g14779(.A(new_n15034), .B(new_n15035), .Y(new_n15036));
  O2A1O1Ixp33_ASAP7_75t_L   g14780(.A1(new_n14985), .A2(new_n14860), .B(new_n14853), .C(new_n15036), .Y(new_n15037));
  INVx1_ASAP7_75t_L         g14781(.A(new_n15037), .Y(new_n15038));
  OAI21xp33_ASAP7_75t_L     g14782(.A1(new_n14860), .A2(new_n14985), .B(new_n14853), .Y(new_n15039));
  INVx1_ASAP7_75t_L         g14783(.A(new_n15039), .Y(new_n15040));
  NAND2xp33_ASAP7_75t_L     g14784(.A(new_n15040), .B(new_n15036), .Y(new_n15041));
  AOI22xp33_ASAP7_75t_L     g14785(.A1(new_n6376), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n6648), .Y(new_n15042));
  OAI221xp5_ASAP7_75t_L     g14786(.A1(new_n6646), .A2(new_n3584), .B1(new_n6636), .B2(new_n10137), .C(new_n15042), .Y(new_n15043));
  XNOR2x2_ASAP7_75t_L       g14787(.A(\a[47] ), .B(new_n15043), .Y(new_n15044));
  AND3x1_ASAP7_75t_L        g14788(.A(new_n15038), .B(new_n15044), .C(new_n15041), .Y(new_n15045));
  AOI21xp33_ASAP7_75t_L     g14789(.A1(new_n15038), .A2(new_n15041), .B(new_n15044), .Y(new_n15046));
  NOR2xp33_ASAP7_75t_L      g14790(.A(new_n15045), .B(new_n15046), .Y(new_n15047));
  O2A1O1Ixp33_ASAP7_75t_L   g14791(.A1(new_n14984), .A2(new_n14868), .B(new_n14983), .C(new_n15047), .Y(new_n15048));
  OAI21xp33_ASAP7_75t_L     g14792(.A1(new_n14868), .A2(new_n14984), .B(new_n14983), .Y(new_n15049));
  NOR3xp33_ASAP7_75t_L      g14793(.A(new_n15049), .B(new_n15046), .C(new_n15045), .Y(new_n15050));
  NOR2xp33_ASAP7_75t_L      g14794(.A(new_n15050), .B(new_n15048), .Y(new_n15051));
  XNOR2x2_ASAP7_75t_L       g14795(.A(new_n14982), .B(new_n15051), .Y(new_n15052));
  XNOR2x2_ASAP7_75t_L       g14796(.A(new_n14978), .B(new_n15052), .Y(new_n15053));
  XNOR2x2_ASAP7_75t_L       g14797(.A(new_n14975), .B(new_n15053), .Y(new_n15054));
  XOR2x2_ASAP7_75t_L        g14798(.A(new_n15054), .B(new_n14971), .Y(new_n15055));
  NAND2xp33_ASAP7_75t_L     g14799(.A(new_n14970), .B(new_n15055), .Y(new_n15056));
  INVx1_ASAP7_75t_L         g14800(.A(new_n15056), .Y(new_n15057));
  NOR2xp33_ASAP7_75t_L      g14801(.A(new_n14970), .B(new_n15055), .Y(new_n15058));
  OR2x4_ASAP7_75t_L         g14802(.A(new_n15058), .B(new_n15057), .Y(new_n15059));
  NOR2xp33_ASAP7_75t_L      g14803(.A(new_n14887), .B(new_n14881), .Y(new_n15060));
  O2A1O1Ixp33_ASAP7_75t_L   g14804(.A1(new_n14873), .A2(new_n14874), .B(new_n14879), .C(new_n15060), .Y(new_n15061));
  XNOR2x2_ASAP7_75t_L       g14805(.A(new_n15061), .B(new_n15059), .Y(new_n15062));
  AOI22xp33_ASAP7_75t_L     g14806(.A1(new_n3633), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n3858), .Y(new_n15063));
  OAI221xp5_ASAP7_75t_L     g14807(.A1(new_n3853), .A2(new_n6568), .B1(new_n3856), .B2(new_n6820), .C(new_n15063), .Y(new_n15064));
  XNOR2x2_ASAP7_75t_L       g14808(.A(\a[35] ), .B(new_n15064), .Y(new_n15065));
  XNOR2x2_ASAP7_75t_L       g14809(.A(new_n15065), .B(new_n15062), .Y(new_n15066));
  XNOR2x2_ASAP7_75t_L       g14810(.A(new_n14966), .B(new_n15066), .Y(new_n15067));
  NOR2xp33_ASAP7_75t_L      g14811(.A(new_n14958), .B(new_n15067), .Y(new_n15068));
  AND2x2_ASAP7_75t_L        g14812(.A(new_n14958), .B(new_n15067), .Y(new_n15069));
  NOR2xp33_ASAP7_75t_L      g14813(.A(new_n15068), .B(new_n15069), .Y(new_n15070));
  NAND2xp33_ASAP7_75t_L     g14814(.A(new_n15070), .B(new_n14946), .Y(new_n15071));
  OAI22xp33_ASAP7_75t_L     g14815(.A1(new_n14944), .A2(new_n14945), .B1(new_n15069), .B2(new_n15068), .Y(new_n15072));
  NAND2xp33_ASAP7_75t_L     g14816(.A(new_n15072), .B(new_n15071), .Y(new_n15073));
  XOR2x2_ASAP7_75t_L        g14817(.A(new_n14939), .B(new_n15073), .Y(new_n15074));
  OAI21xp33_ASAP7_75t_L     g14818(.A1(new_n14934), .A2(new_n14932), .B(new_n15074), .Y(new_n15075));
  NOR2xp33_ASAP7_75t_L      g14819(.A(new_n14934), .B(new_n14932), .Y(new_n15076));
  INVx1_ASAP7_75t_L         g14820(.A(new_n15074), .Y(new_n15077));
  NAND2xp33_ASAP7_75t_L     g14821(.A(new_n15077), .B(new_n15076), .Y(new_n15078));
  INVx1_ASAP7_75t_L         g14822(.A(new_n14746), .Y(new_n15079));
  A2O1A1Ixp33_ASAP7_75t_L   g14823(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n1073), .Y(new_n15080));
  A2O1A1Ixp33_ASAP7_75t_L   g14824(.A1(new_n15080), .A2(new_n1158), .B(new_n11468), .C(\a[17] ), .Y(new_n15081));
  O2A1O1Ixp33_ASAP7_75t_L   g14825(.A1(new_n1156), .A2(new_n12060), .B(new_n1158), .C(new_n11468), .Y(new_n15082));
  NAND2xp33_ASAP7_75t_L     g14826(.A(new_n1071), .B(new_n15082), .Y(new_n15083));
  AND2x2_ASAP7_75t_L        g14827(.A(new_n15083), .B(new_n15081), .Y(new_n15084));
  INVx1_ASAP7_75t_L         g14828(.A(new_n15084), .Y(new_n15085));
  A2O1A1Ixp33_ASAP7_75t_L   g14829(.A1(new_n14908), .A2(new_n14744), .B(new_n15079), .C(new_n15085), .Y(new_n15086));
  INVx1_ASAP7_75t_L         g14830(.A(new_n14909), .Y(new_n15087));
  NAND3xp33_ASAP7_75t_L     g14831(.A(new_n15087), .B(new_n14746), .C(new_n15084), .Y(new_n15088));
  NAND4xp25_ASAP7_75t_L     g14832(.A(new_n15088), .B(new_n15075), .C(new_n15078), .D(new_n15086), .Y(new_n15089));
  INVx1_ASAP7_75t_L         g14833(.A(new_n15089), .Y(new_n15090));
  AOI22xp33_ASAP7_75t_L     g14834(.A1(new_n15075), .A2(new_n15078), .B1(new_n15086), .B2(new_n15088), .Y(new_n15091));
  INVx1_ASAP7_75t_L         g14835(.A(new_n14910), .Y(new_n15092));
  A2O1A1Ixp33_ASAP7_75t_L   g14836(.A1(new_n15087), .A2(new_n15092), .B(new_n14734), .C(new_n14737), .Y(new_n15093));
  NOR3xp33_ASAP7_75t_L      g14837(.A(new_n15090), .B(new_n15093), .C(new_n15091), .Y(new_n15094));
  OA21x2_ASAP7_75t_L        g14838(.A1(new_n15091), .A2(new_n15090), .B(new_n15093), .Y(new_n15095));
  NOR2xp33_ASAP7_75t_L      g14839(.A(new_n15094), .B(new_n15095), .Y(new_n15096));
  A2O1A1Ixp33_ASAP7_75t_L   g14840(.A1(new_n14924), .A2(new_n14920), .B(new_n14919), .C(new_n15096), .Y(new_n15097));
  INVx1_ASAP7_75t_L         g14841(.A(new_n15097), .Y(new_n15098));
  INVx1_ASAP7_75t_L         g14842(.A(new_n14919), .Y(new_n15099));
  A2O1A1Ixp33_ASAP7_75t_L   g14843(.A1(new_n14721), .A2(new_n14719), .B(new_n14918), .C(new_n15099), .Y(new_n15100));
  NOR2xp33_ASAP7_75t_L      g14844(.A(new_n15096), .B(new_n15100), .Y(new_n15101));
  NOR2xp33_ASAP7_75t_L      g14845(.A(new_n15098), .B(new_n15101), .Y(\f[80] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14846(.A1(new_n15087), .A2(new_n14746), .B(new_n15084), .C(new_n15089), .Y(new_n15103));
  INVx1_ASAP7_75t_L         g14847(.A(new_n15103), .Y(new_n15104));
  AOI22xp33_ASAP7_75t_L     g14848(.A1(new_n1360), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1581), .Y(new_n15105));
  A2O1A1Ixp33_ASAP7_75t_L   g14849(.A1(new_n11470), .A2(new_n11473), .B(new_n1359), .C(new_n15105), .Y(new_n15106));
  AOI21xp33_ASAP7_75t_L     g14850(.A1(new_n1362), .A2(\b[62] ), .B(new_n15106), .Y(new_n15107));
  NAND2xp33_ASAP7_75t_L     g14851(.A(\a[20] ), .B(new_n15107), .Y(new_n15108));
  A2O1A1Ixp33_ASAP7_75t_L   g14852(.A1(\b[62] ), .A2(new_n1362), .B(new_n15106), .C(new_n1356), .Y(new_n15109));
  AND2x2_ASAP7_75t_L        g14853(.A(new_n15109), .B(new_n15108), .Y(new_n15110));
  INVx1_ASAP7_75t_L         g14854(.A(new_n15110), .Y(new_n15111));
  O2A1O1Ixp33_ASAP7_75t_L   g14855(.A1(new_n15074), .A2(new_n14932), .B(new_n14933), .C(new_n15111), .Y(new_n15112));
  A2O1A1Ixp33_ASAP7_75t_L   g14856(.A1(new_n14906), .A2(new_n14753), .B(new_n14929), .C(new_n15078), .Y(new_n15113));
  NOR2xp33_ASAP7_75t_L      g14857(.A(new_n15110), .B(new_n15113), .Y(new_n15114));
  AOI22xp33_ASAP7_75t_L     g14858(.A1(new_n1704), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1837), .Y(new_n15115));
  OAI221xp5_ASAP7_75t_L     g14859(.A1(new_n1699), .A2(new_n9947), .B1(new_n1827), .B2(new_n11446), .C(new_n15115), .Y(new_n15116));
  XNOR2x2_ASAP7_75t_L       g14860(.A(\a[23] ), .B(new_n15116), .Y(new_n15117));
  INVx1_ASAP7_75t_L         g14861(.A(new_n15117), .Y(new_n15118));
  INVx1_ASAP7_75t_L         g14862(.A(new_n14938), .Y(new_n15119));
  MAJIxp5_ASAP7_75t_L       g14863(.A(new_n15073), .B(new_n14937), .C(new_n15119), .Y(new_n15120));
  OR2x4_ASAP7_75t_L         g14864(.A(new_n15118), .B(new_n15120), .Y(new_n15121));
  NAND2xp33_ASAP7_75t_L     g14865(.A(new_n15118), .B(new_n15120), .Y(new_n15122));
  NAND2xp33_ASAP7_75t_L     g14866(.A(new_n15122), .B(new_n15121), .Y(new_n15123));
  AOI22xp33_ASAP7_75t_L     g14867(.A1(new_n2552), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n2736), .Y(new_n15124));
  OAI221xp5_ASAP7_75t_L     g14868(.A1(new_n2547), .A2(new_n8165), .B1(new_n2734), .B2(new_n8465), .C(new_n15124), .Y(new_n15125));
  XNOR2x2_ASAP7_75t_L       g14869(.A(\a[29] ), .B(new_n15125), .Y(new_n15126));
  INVx1_ASAP7_75t_L         g14870(.A(new_n15126), .Y(new_n15127));
  A2O1A1O1Ixp25_ASAP7_75t_L g14871(.A1(new_n14896), .A2(new_n14895), .B(new_n14772), .C(new_n14953), .D(new_n14951), .Y(new_n15128));
  OR3x1_ASAP7_75t_L         g14872(.A(new_n15068), .B(new_n15127), .C(new_n15128), .Y(new_n15129));
  A2O1A1Ixp33_ASAP7_75t_L   g14873(.A1(new_n14954), .A2(new_n14956), .B(new_n15068), .C(new_n15127), .Y(new_n15130));
  INVx1_ASAP7_75t_L         g14874(.A(new_n15059), .Y(new_n15131));
  O2A1O1Ixp33_ASAP7_75t_L   g14875(.A1(new_n14881), .A2(new_n14887), .B(new_n14880), .C(new_n15131), .Y(new_n15132));
  O2A1O1Ixp33_ASAP7_75t_L   g14876(.A1(new_n14782), .A2(new_n14977), .B(new_n14976), .C(new_n15052), .Y(new_n15133));
  AOI21xp33_ASAP7_75t_L     g14877(.A1(new_n15053), .A2(new_n14975), .B(new_n15133), .Y(new_n15134));
  INVx1_ASAP7_75t_L         g14878(.A(new_n15134), .Y(new_n15135));
  AOI22xp33_ASAP7_75t_L     g14879(.A1(new_n4920), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n5167), .Y(new_n15136));
  OAI221xp5_ASAP7_75t_L     g14880(.A1(new_n5154), .A2(new_n5321), .B1(new_n5158), .B2(new_n5346), .C(new_n15136), .Y(new_n15137));
  XNOR2x2_ASAP7_75t_L       g14881(.A(\a[41] ), .B(new_n15137), .Y(new_n15138));
  INVx1_ASAP7_75t_L         g14882(.A(new_n15048), .Y(new_n15139));
  INVx1_ASAP7_75t_L         g14883(.A(new_n15001), .Y(new_n15140));
  AOI22xp33_ASAP7_75t_L     g14884(.A1(new_n9700), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n10027), .Y(new_n15141));
  OAI221xp5_ASAP7_75t_L     g14885(.A1(new_n10024), .A2(new_n1909), .B1(new_n9696), .B2(new_n2477), .C(new_n15141), .Y(new_n15142));
  XNOR2x2_ASAP7_75t_L       g14886(.A(\a[59] ), .B(new_n15142), .Y(new_n15143));
  AOI22xp33_ASAP7_75t_L     g14887(.A1(\b[19] ), .A2(new_n10939), .B1(\b[21] ), .B2(new_n10938), .Y(new_n15144));
  OAI221xp5_ASAP7_75t_L     g14888(.A1(new_n10937), .A2(new_n1539), .B1(new_n10629), .B2(new_n1662), .C(new_n15144), .Y(new_n15145));
  XNOR2x2_ASAP7_75t_L       g14889(.A(\a[62] ), .B(new_n15145), .Y(new_n15146));
  INVx1_ASAP7_75t_L         g14890(.A(new_n14998), .Y(new_n15147));
  NOR2xp33_ASAP7_75t_L      g14891(.A(new_n1201), .B(new_n11535), .Y(new_n15148));
  A2O1A1Ixp33_ASAP7_75t_L   g14892(.A1(new_n11533), .A2(\b[18] ), .B(new_n15148), .C(new_n1071), .Y(new_n15149));
  O2A1O1Ixp33_ASAP7_75t_L   g14893(.A1(new_n11247), .A2(new_n11249), .B(\b[18] ), .C(new_n15148), .Y(new_n15150));
  NAND2xp33_ASAP7_75t_L     g14894(.A(\a[17] ), .B(new_n15150), .Y(new_n15151));
  NAND2xp33_ASAP7_75t_L     g14895(.A(new_n15149), .B(new_n15151), .Y(new_n15152));
  XNOR2x2_ASAP7_75t_L       g14896(.A(new_n15147), .B(new_n15152), .Y(new_n15153));
  INVx1_ASAP7_75t_L         g14897(.A(new_n15153), .Y(new_n15154));
  XNOR2x2_ASAP7_75t_L       g14898(.A(new_n15154), .B(new_n15146), .Y(new_n15155));
  INVx1_ASAP7_75t_L         g14899(.A(new_n15155), .Y(new_n15156));
  A2O1A1O1Ixp25_ASAP7_75t_L g14900(.A1(\b[17] ), .A2(new_n11533), .B(new_n14996), .C(new_n14797), .D(new_n14995), .Y(new_n15157));
  A2O1A1Ixp33_ASAP7_75t_L   g14901(.A1(new_n14798), .A2(new_n14998), .B(new_n15157), .C(new_n15156), .Y(new_n15158));
  A2O1A1O1Ixp25_ASAP7_75t_L g14902(.A1(new_n11533), .A2(\b[16] ), .B(new_n14794), .C(new_n14998), .D(new_n15157), .Y(new_n15159));
  NAND2xp33_ASAP7_75t_L     g14903(.A(new_n15159), .B(new_n15155), .Y(new_n15160));
  AND2x2_ASAP7_75t_L        g14904(.A(new_n15160), .B(new_n15158), .Y(new_n15161));
  INVx1_ASAP7_75t_L         g14905(.A(new_n15161), .Y(new_n15162));
  NAND2xp33_ASAP7_75t_L     g14906(.A(new_n15143), .B(new_n15162), .Y(new_n15163));
  INVx1_ASAP7_75t_L         g14907(.A(new_n15143), .Y(new_n15164));
  NAND2xp33_ASAP7_75t_L     g14908(.A(new_n15164), .B(new_n15161), .Y(new_n15165));
  AND2x2_ASAP7_75t_L        g14909(.A(new_n15165), .B(new_n15163), .Y(new_n15166));
  A2O1A1Ixp33_ASAP7_75t_L   g14910(.A1(new_n15140), .A2(new_n14992), .B(new_n15007), .C(new_n15166), .Y(new_n15167));
  A2O1A1Ixp33_ASAP7_75t_L   g14911(.A1(new_n14808), .A2(new_n14801), .B(new_n15001), .C(new_n15008), .Y(new_n15168));
  AO21x2_ASAP7_75t_L        g14912(.A1(new_n15165), .A2(new_n15163), .B(new_n15168), .Y(new_n15169));
  NAND2xp33_ASAP7_75t_L     g14913(.A(new_n15169), .B(new_n15167), .Y(new_n15170));
  AOI22xp33_ASAP7_75t_L     g14914(.A1(new_n8831), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n9115), .Y(new_n15171));
  OAI221xp5_ASAP7_75t_L     g14915(.A1(new_n10343), .A2(new_n2348), .B1(new_n10016), .B2(new_n2505), .C(new_n15171), .Y(new_n15172));
  XNOR2x2_ASAP7_75t_L       g14916(.A(\a[56] ), .B(new_n15172), .Y(new_n15173));
  XNOR2x2_ASAP7_75t_L       g14917(.A(new_n15173), .B(new_n15170), .Y(new_n15174));
  INVx1_ASAP7_75t_L         g14918(.A(new_n15174), .Y(new_n15175));
  NOR3xp33_ASAP7_75t_L      g14919(.A(new_n15175), .B(new_n15015), .C(new_n15013), .Y(new_n15176));
  O2A1O1Ixp33_ASAP7_75t_L   g14920(.A1(new_n14991), .A2(new_n15014), .B(new_n15012), .C(new_n15174), .Y(new_n15177));
  NOR2xp33_ASAP7_75t_L      g14921(.A(new_n15177), .B(new_n15176), .Y(new_n15178));
  AOI22xp33_ASAP7_75t_L     g14922(.A1(new_n7960), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n8537), .Y(new_n15179));
  OAI221xp5_ASAP7_75t_L     g14923(.A1(new_n8817), .A2(new_n2688), .B1(new_n7957), .B2(new_n2990), .C(new_n15179), .Y(new_n15180));
  XNOR2x2_ASAP7_75t_L       g14924(.A(\a[53] ), .B(new_n15180), .Y(new_n15181));
  INVx1_ASAP7_75t_L         g14925(.A(new_n15181), .Y(new_n15182));
  XNOR2x2_ASAP7_75t_L       g14926(.A(new_n15182), .B(new_n15178), .Y(new_n15183));
  A2O1A1Ixp33_ASAP7_75t_L   g14927(.A1(new_n15023), .A2(new_n15026), .B(new_n15022), .C(new_n15183), .Y(new_n15184));
  NAND2xp33_ASAP7_75t_L     g14928(.A(new_n15026), .B(new_n15023), .Y(new_n15185));
  A2O1A1Ixp33_ASAP7_75t_L   g14929(.A1(new_n14830), .A2(new_n14823), .B(new_n15021), .C(new_n15185), .Y(new_n15186));
  OR2x4_ASAP7_75t_L         g14930(.A(new_n15186), .B(new_n15183), .Y(new_n15187));
  NAND2xp33_ASAP7_75t_L     g14931(.A(new_n15184), .B(new_n15187), .Y(new_n15188));
  AOI22xp33_ASAP7_75t_L     g14932(.A1(new_n7111), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n7391), .Y(new_n15189));
  OAI221xp5_ASAP7_75t_L     g14933(.A1(new_n8558), .A2(new_n3207), .B1(new_n8237), .B2(new_n3572), .C(new_n15189), .Y(new_n15190));
  XNOR2x2_ASAP7_75t_L       g14934(.A(\a[50] ), .B(new_n15190), .Y(new_n15191));
  AOI21xp33_ASAP7_75t_L     g14935(.A1(new_n15031), .A2(new_n14988), .B(new_n15032), .Y(new_n15192));
  XNOR2x2_ASAP7_75t_L       g14936(.A(new_n15191), .B(new_n15192), .Y(new_n15193));
  XOR2x2_ASAP7_75t_L        g14937(.A(new_n15193), .B(new_n15188), .Y(new_n15194));
  AOI22xp33_ASAP7_75t_L     g14938(.A1(new_n6376), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n6648), .Y(new_n15195));
  OAI221xp5_ASAP7_75t_L     g14939(.A1(new_n6646), .A2(new_n3804), .B1(new_n6636), .B2(new_n4223), .C(new_n15195), .Y(new_n15196));
  XNOR2x2_ASAP7_75t_L       g14940(.A(\a[47] ), .B(new_n15196), .Y(new_n15197));
  NOR2xp33_ASAP7_75t_L      g14941(.A(new_n15197), .B(new_n15194), .Y(new_n15198));
  INVx1_ASAP7_75t_L         g14942(.A(new_n15198), .Y(new_n15199));
  NAND2xp33_ASAP7_75t_L     g14943(.A(new_n15197), .B(new_n15194), .Y(new_n15200));
  NAND2xp33_ASAP7_75t_L     g14944(.A(new_n15200), .B(new_n15199), .Y(new_n15201));
  A2O1A1Ixp33_ASAP7_75t_L   g14945(.A1(new_n15041), .A2(new_n15044), .B(new_n15037), .C(new_n15201), .Y(new_n15202));
  OR3x1_ASAP7_75t_L         g14946(.A(new_n15201), .B(new_n15037), .C(new_n15045), .Y(new_n15203));
  NAND2xp33_ASAP7_75t_L     g14947(.A(new_n15202), .B(new_n15203), .Y(new_n15204));
  AOI22xp33_ASAP7_75t_L     g14948(.A1(new_n5624), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n5901), .Y(new_n15205));
  OAI221xp5_ASAP7_75t_L     g14949(.A1(new_n5900), .A2(new_n4632), .B1(new_n5892), .B2(new_n4858), .C(new_n15205), .Y(new_n15206));
  XNOR2x2_ASAP7_75t_L       g14950(.A(\a[44] ), .B(new_n15206), .Y(new_n15207));
  XNOR2x2_ASAP7_75t_L       g14951(.A(new_n15207), .B(new_n15204), .Y(new_n15208));
  O2A1O1Ixp33_ASAP7_75t_L   g14952(.A1(new_n14981), .A2(new_n15050), .B(new_n15139), .C(new_n15208), .Y(new_n15209));
  AOI21xp33_ASAP7_75t_L     g14953(.A1(new_n15051), .A2(new_n14982), .B(new_n15048), .Y(new_n15210));
  AND2x2_ASAP7_75t_L        g14954(.A(new_n15210), .B(new_n15208), .Y(new_n15211));
  OR3x1_ASAP7_75t_L         g14955(.A(new_n15211), .B(new_n15138), .C(new_n15209), .Y(new_n15212));
  OAI21xp33_ASAP7_75t_L     g14956(.A1(new_n15209), .A2(new_n15211), .B(new_n15138), .Y(new_n15213));
  AO21x2_ASAP7_75t_L        g14957(.A1(new_n15213), .A2(new_n15212), .B(new_n15135), .Y(new_n15214));
  NAND3xp33_ASAP7_75t_L     g14958(.A(new_n15212), .B(new_n15135), .C(new_n15213), .Y(new_n15215));
  NAND2xp33_ASAP7_75t_L     g14959(.A(new_n15215), .B(new_n15214), .Y(new_n15216));
  AOI22xp33_ASAP7_75t_L     g14960(.A1(new_n4283), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n4512), .Y(new_n15217));
  OAI221xp5_ASAP7_75t_L     g14961(.A1(new_n4277), .A2(new_n5829), .B1(new_n4499), .B2(new_n6329), .C(new_n15217), .Y(new_n15218));
  XNOR2x2_ASAP7_75t_L       g14962(.A(\a[38] ), .B(new_n15218), .Y(new_n15219));
  XNOR2x2_ASAP7_75t_L       g14963(.A(new_n15219), .B(new_n15216), .Y(new_n15220));
  A2O1A1Ixp33_ASAP7_75t_L   g14964(.A1(new_n14674), .A2(new_n14616), .B(new_n14778), .C(new_n14871), .Y(new_n15221));
  INVx1_ASAP7_75t_L         g14965(.A(new_n14873), .Y(new_n15222));
  A2O1A1Ixp33_ASAP7_75t_L   g14966(.A1(new_n15222), .A2(new_n15221), .B(new_n15054), .C(new_n15056), .Y(new_n15223));
  INVx1_ASAP7_75t_L         g14967(.A(new_n15223), .Y(new_n15224));
  NAND2xp33_ASAP7_75t_L     g14968(.A(new_n15220), .B(new_n15224), .Y(new_n15225));
  OR2x4_ASAP7_75t_L         g14969(.A(new_n15220), .B(new_n15224), .Y(new_n15226));
  NAND2xp33_ASAP7_75t_L     g14970(.A(new_n15225), .B(new_n15226), .Y(new_n15227));
  AOI22xp33_ASAP7_75t_L     g14971(.A1(new_n3633), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n3858), .Y(new_n15228));
  OAI221xp5_ASAP7_75t_L     g14972(.A1(new_n3853), .A2(new_n6812), .B1(new_n3856), .B2(new_n6837), .C(new_n15228), .Y(new_n15229));
  XNOR2x2_ASAP7_75t_L       g14973(.A(\a[35] ), .B(new_n15229), .Y(new_n15230));
  XOR2x2_ASAP7_75t_L        g14974(.A(new_n15230), .B(new_n15227), .Y(new_n15231));
  INVx1_ASAP7_75t_L         g14975(.A(new_n15231), .Y(new_n15232));
  A2O1A1Ixp33_ASAP7_75t_L   g14976(.A1(new_n15062), .A2(new_n15065), .B(new_n15132), .C(new_n15232), .Y(new_n15233));
  AOI21xp33_ASAP7_75t_L     g14977(.A1(new_n15062), .A2(new_n15065), .B(new_n15132), .Y(new_n15234));
  NAND2xp33_ASAP7_75t_L     g14978(.A(new_n15234), .B(new_n15231), .Y(new_n15235));
  NAND2xp33_ASAP7_75t_L     g14979(.A(new_n15235), .B(new_n15233), .Y(new_n15236));
  AOI22xp33_ASAP7_75t_L     g14980(.A1(new_n3029), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n3258), .Y(new_n15237));
  OAI221xp5_ASAP7_75t_L     g14981(.A1(new_n3024), .A2(new_n7593), .B1(new_n3256), .B2(new_n7623), .C(new_n15237), .Y(new_n15238));
  XNOR2x2_ASAP7_75t_L       g14982(.A(\a[32] ), .B(new_n15238), .Y(new_n15239));
  INVx1_ASAP7_75t_L         g14983(.A(new_n15239), .Y(new_n15240));
  A2O1A1Ixp33_ASAP7_75t_L   g14984(.A1(new_n15066), .A2(new_n14966), .B(new_n14965), .C(new_n15240), .Y(new_n15241));
  AOI21xp33_ASAP7_75t_L     g14985(.A1(new_n15066), .A2(new_n14966), .B(new_n14965), .Y(new_n15242));
  NAND2xp33_ASAP7_75t_L     g14986(.A(new_n15239), .B(new_n15242), .Y(new_n15243));
  NAND2xp33_ASAP7_75t_L     g14987(.A(new_n15241), .B(new_n15243), .Y(new_n15244));
  XNOR2x2_ASAP7_75t_L       g14988(.A(new_n15236), .B(new_n15244), .Y(new_n15245));
  NAND3xp33_ASAP7_75t_L     g14989(.A(new_n15245), .B(new_n15130), .C(new_n15129), .Y(new_n15246));
  AO21x2_ASAP7_75t_L        g14990(.A1(new_n15129), .A2(new_n15130), .B(new_n15245), .Y(new_n15247));
  NAND2xp33_ASAP7_75t_L     g14991(.A(new_n15246), .B(new_n15247), .Y(new_n15248));
  INVx1_ASAP7_75t_L         g14992(.A(new_n15248), .Y(new_n15249));
  AOI22xp33_ASAP7_75t_L     g14993(.A1(new_n2114), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n2259), .Y(new_n15250));
  OAI221xp5_ASAP7_75t_L     g14994(.A1(new_n2109), .A2(new_n9323), .B1(new_n2257), .B2(new_n9627), .C(new_n15250), .Y(new_n15251));
  XNOR2x2_ASAP7_75t_L       g14995(.A(\a[26] ), .B(new_n15251), .Y(new_n15252));
  O2A1O1Ixp33_ASAP7_75t_L   g14996(.A1(new_n14942), .A2(new_n14943), .B(new_n15071), .C(new_n15252), .Y(new_n15253));
  OA211x2_ASAP7_75t_L       g14997(.A1(new_n14942), .A2(new_n14943), .B(new_n15071), .C(new_n15252), .Y(new_n15254));
  NOR2xp33_ASAP7_75t_L      g14998(.A(new_n15253), .B(new_n15254), .Y(new_n15255));
  XNOR2x2_ASAP7_75t_L       g14999(.A(new_n15249), .B(new_n15255), .Y(new_n15256));
  OR2x4_ASAP7_75t_L         g15000(.A(new_n15123), .B(new_n15256), .Y(new_n15257));
  NAND2xp33_ASAP7_75t_L     g15001(.A(new_n15123), .B(new_n15256), .Y(new_n15258));
  NAND2xp33_ASAP7_75t_L     g15002(.A(new_n15258), .B(new_n15257), .Y(new_n15259));
  OAI21xp33_ASAP7_75t_L     g15003(.A1(new_n15112), .A2(new_n15114), .B(new_n15259), .Y(new_n15260));
  INVx1_ASAP7_75t_L         g15004(.A(new_n15260), .Y(new_n15261));
  NOR3xp33_ASAP7_75t_L      g15005(.A(new_n15114), .B(new_n15259), .C(new_n15112), .Y(new_n15262));
  OR3x1_ASAP7_75t_L         g15006(.A(new_n15261), .B(new_n15104), .C(new_n15262), .Y(new_n15263));
  OAI21xp33_ASAP7_75t_L     g15007(.A1(new_n15262), .A2(new_n15261), .B(new_n15104), .Y(new_n15264));
  AND2x2_ASAP7_75t_L        g15008(.A(new_n15264), .B(new_n15263), .Y(new_n15265));
  A2O1A1Ixp33_ASAP7_75t_L   g15009(.A1(new_n15100), .A2(new_n15096), .B(new_n15094), .C(new_n15265), .Y(new_n15266));
  INVx1_ASAP7_75t_L         g15010(.A(new_n15266), .Y(new_n15267));
  INVx1_ASAP7_75t_L         g15011(.A(new_n15094), .Y(new_n15268));
  A2O1A1Ixp33_ASAP7_75t_L   g15012(.A1(new_n14921), .A2(new_n15099), .B(new_n15095), .C(new_n15268), .Y(new_n15269));
  NOR2xp33_ASAP7_75t_L      g15013(.A(new_n15265), .B(new_n15269), .Y(new_n15270));
  NOR2xp33_ASAP7_75t_L      g15014(.A(new_n15270), .B(new_n15267), .Y(\f[81] ));
  INVx1_ASAP7_75t_L         g15015(.A(new_n15263), .Y(new_n15272));
  O2A1O1Ixp33_ASAP7_75t_L   g15016(.A1(new_n15074), .A2(new_n14932), .B(new_n14933), .C(new_n15110), .Y(new_n15273));
  O2A1O1Ixp33_ASAP7_75t_L   g15017(.A1(new_n15112), .A2(new_n15114), .B(new_n15259), .C(new_n15273), .Y(new_n15274));
  INVx1_ASAP7_75t_L         g15018(.A(new_n15253), .Y(new_n15275));
  AOI22xp33_ASAP7_75t_L     g15019(.A1(new_n1704), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1837), .Y(new_n15276));
  OAI221xp5_ASAP7_75t_L     g15020(.A1(new_n1699), .A2(new_n10250), .B1(new_n1827), .B2(new_n10855), .C(new_n15276), .Y(new_n15277));
  XNOR2x2_ASAP7_75t_L       g15021(.A(\a[23] ), .B(new_n15277), .Y(new_n15278));
  A2O1A1Ixp33_ASAP7_75t_L   g15022(.A1(new_n15275), .A2(new_n15249), .B(new_n15254), .C(new_n15278), .Y(new_n15279));
  NOR3xp33_ASAP7_75t_L      g15023(.A(new_n15254), .B(new_n15253), .C(new_n15248), .Y(new_n15280));
  OR3x1_ASAP7_75t_L         g15024(.A(new_n15280), .B(new_n15254), .C(new_n15278), .Y(new_n15281));
  AND2x2_ASAP7_75t_L        g15025(.A(new_n15279), .B(new_n15281), .Y(new_n15282));
  AOI22xp33_ASAP7_75t_L     g15026(.A1(new_n2114), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n2259), .Y(new_n15283));
  OAI221xp5_ASAP7_75t_L     g15027(.A1(new_n2109), .A2(new_n9620), .B1(new_n2257), .B2(new_n9925), .C(new_n15283), .Y(new_n15284));
  XNOR2x2_ASAP7_75t_L       g15028(.A(\a[26] ), .B(new_n15284), .Y(new_n15285));
  NAND2xp33_ASAP7_75t_L     g15029(.A(new_n15129), .B(new_n15246), .Y(new_n15286));
  XNOR2x2_ASAP7_75t_L       g15030(.A(new_n15285), .B(new_n15286), .Y(new_n15287));
  AOI22xp33_ASAP7_75t_L     g15031(.A1(new_n2552), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n2736), .Y(new_n15288));
  OAI221xp5_ASAP7_75t_L     g15032(.A1(new_n2547), .A2(new_n8458), .B1(new_n2734), .B2(new_n8768), .C(new_n15288), .Y(new_n15289));
  XNOR2x2_ASAP7_75t_L       g15033(.A(\a[29] ), .B(new_n15289), .Y(new_n15290));
  A2O1A1Ixp33_ASAP7_75t_L   g15034(.A1(new_n15233), .A2(new_n15235), .B(new_n15244), .C(new_n15243), .Y(new_n15291));
  XNOR2x2_ASAP7_75t_L       g15035(.A(new_n15290), .B(new_n15291), .Y(new_n15292));
  AOI22xp33_ASAP7_75t_L     g15036(.A1(new_n3029), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n3258), .Y(new_n15293));
  OAI221xp5_ASAP7_75t_L     g15037(.A1(new_n3024), .A2(new_n7616), .B1(new_n3256), .B2(new_n7906), .C(new_n15293), .Y(new_n15294));
  XNOR2x2_ASAP7_75t_L       g15038(.A(\a[32] ), .B(new_n15294), .Y(new_n15295));
  OAI211xp5_ASAP7_75t_L     g15039(.A1(new_n15230), .A2(new_n15227), .B(new_n15235), .C(new_n15295), .Y(new_n15296));
  O2A1O1Ixp33_ASAP7_75t_L   g15040(.A1(new_n15227), .A2(new_n15230), .B(new_n15235), .C(new_n15295), .Y(new_n15297));
  INVx1_ASAP7_75t_L         g15041(.A(new_n15297), .Y(new_n15298));
  NAND2xp33_ASAP7_75t_L     g15042(.A(new_n15296), .B(new_n15298), .Y(new_n15299));
  MAJIxp5_ASAP7_75t_L       g15043(.A(new_n15204), .B(new_n15207), .C(new_n15210), .Y(new_n15300));
  AOI22xp33_ASAP7_75t_L     g15044(.A1(new_n5624), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n5901), .Y(new_n15301));
  OAI221xp5_ASAP7_75t_L     g15045(.A1(new_n5900), .A2(new_n4848), .B1(new_n5892), .B2(new_n11686), .C(new_n15301), .Y(new_n15302));
  XNOR2x2_ASAP7_75t_L       g15046(.A(\a[44] ), .B(new_n15302), .Y(new_n15303));
  INVx1_ASAP7_75t_L         g15047(.A(new_n15303), .Y(new_n15304));
  NAND2xp33_ASAP7_75t_L     g15048(.A(new_n15199), .B(new_n15203), .Y(new_n15305));
  INVx1_ASAP7_75t_L         g15049(.A(new_n15170), .Y(new_n15306));
  INVx1_ASAP7_75t_L         g15050(.A(new_n15173), .Y(new_n15307));
  AOI22xp33_ASAP7_75t_L     g15051(.A1(new_n8831), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n9115), .Y(new_n15308));
  OAI221xp5_ASAP7_75t_L     g15052(.A1(new_n10343), .A2(new_n2497), .B1(new_n10016), .B2(new_n2672), .C(new_n15308), .Y(new_n15309));
  XNOR2x2_ASAP7_75t_L       g15053(.A(\a[56] ), .B(new_n15309), .Y(new_n15310));
  INVx1_ASAP7_75t_L         g15054(.A(new_n15310), .Y(new_n15311));
  INVx1_ASAP7_75t_L         g15055(.A(new_n15159), .Y(new_n15312));
  NOR2xp33_ASAP7_75t_L      g15056(.A(new_n1313), .B(new_n11535), .Y(new_n15313));
  INVx1_ASAP7_75t_L         g15057(.A(new_n15149), .Y(new_n15314));
  A2O1A1O1Ixp25_ASAP7_75t_L g15058(.A1(new_n11533), .A2(\b[17] ), .B(new_n14996), .C(new_n15151), .D(new_n15314), .Y(new_n15315));
  A2O1A1Ixp33_ASAP7_75t_L   g15059(.A1(new_n11533), .A2(\b[19] ), .B(new_n15313), .C(new_n15315), .Y(new_n15316));
  O2A1O1Ixp33_ASAP7_75t_L   g15060(.A1(new_n11247), .A2(new_n11249), .B(\b[19] ), .C(new_n15313), .Y(new_n15317));
  INVx1_ASAP7_75t_L         g15061(.A(new_n15317), .Y(new_n15318));
  O2A1O1Ixp33_ASAP7_75t_L   g15062(.A1(new_n14998), .A2(new_n15152), .B(new_n15149), .C(new_n15318), .Y(new_n15319));
  INVx1_ASAP7_75t_L         g15063(.A(new_n15319), .Y(new_n15320));
  NAND2xp33_ASAP7_75t_L     g15064(.A(new_n15316), .B(new_n15320), .Y(new_n15321));
  AOI22xp33_ASAP7_75t_L     g15065(.A1(\b[20] ), .A2(new_n10939), .B1(\b[22] ), .B2(new_n10938), .Y(new_n15322));
  OAI221xp5_ASAP7_75t_L     g15066(.A1(new_n10937), .A2(new_n1655), .B1(new_n10629), .B2(new_n1780), .C(new_n15322), .Y(new_n15323));
  XNOR2x2_ASAP7_75t_L       g15067(.A(\a[62] ), .B(new_n15323), .Y(new_n15324));
  NAND2xp33_ASAP7_75t_L     g15068(.A(new_n15321), .B(new_n15324), .Y(new_n15325));
  NOR2xp33_ASAP7_75t_L      g15069(.A(new_n15321), .B(new_n15324), .Y(new_n15326));
  INVx1_ASAP7_75t_L         g15070(.A(new_n15326), .Y(new_n15327));
  AND2x2_ASAP7_75t_L        g15071(.A(new_n15325), .B(new_n15327), .Y(new_n15328));
  NOR2xp33_ASAP7_75t_L      g15072(.A(new_n15154), .B(new_n15146), .Y(new_n15329));
  A2O1A1Ixp33_ASAP7_75t_L   g15073(.A1(new_n15156), .A2(new_n15312), .B(new_n15329), .C(new_n15328), .Y(new_n15330));
  A2O1A1O1Ixp25_ASAP7_75t_L g15074(.A1(new_n14998), .A2(new_n14798), .B(new_n15157), .C(new_n15156), .D(new_n15329), .Y(new_n15331));
  INVx1_ASAP7_75t_L         g15075(.A(new_n15331), .Y(new_n15332));
  NOR2xp33_ASAP7_75t_L      g15076(.A(new_n15328), .B(new_n15332), .Y(new_n15333));
  INVx1_ASAP7_75t_L         g15077(.A(new_n15333), .Y(new_n15334));
  AOI22xp33_ASAP7_75t_L     g15078(.A1(new_n9700), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n10027), .Y(new_n15335));
  OAI221xp5_ASAP7_75t_L     g15079(.A1(new_n10024), .A2(new_n1929), .B1(new_n9696), .B2(new_n2075), .C(new_n15335), .Y(new_n15336));
  XNOR2x2_ASAP7_75t_L       g15080(.A(\a[59] ), .B(new_n15336), .Y(new_n15337));
  NAND3xp33_ASAP7_75t_L     g15081(.A(new_n15334), .B(new_n15330), .C(new_n15337), .Y(new_n15338));
  AO21x2_ASAP7_75t_L        g15082(.A1(new_n15330), .A2(new_n15334), .B(new_n15337), .Y(new_n15339));
  AND2x2_ASAP7_75t_L        g15083(.A(new_n15338), .B(new_n15339), .Y(new_n15340));
  O2A1O1Ixp33_ASAP7_75t_L   g15084(.A1(new_n15143), .A2(new_n15162), .B(new_n15167), .C(new_n15340), .Y(new_n15341));
  INVx1_ASAP7_75t_L         g15085(.A(new_n15341), .Y(new_n15342));
  O2A1O1Ixp33_ASAP7_75t_L   g15086(.A1(new_n14798), .A2(new_n14795), .B(new_n14808), .C(new_n15001), .Y(new_n15343));
  INVx1_ASAP7_75t_L         g15087(.A(new_n15165), .Y(new_n15344));
  O2A1O1Ixp33_ASAP7_75t_L   g15088(.A1(new_n15343), .A2(new_n15007), .B(new_n15163), .C(new_n15344), .Y(new_n15345));
  NAND2xp33_ASAP7_75t_L     g15089(.A(new_n15345), .B(new_n15340), .Y(new_n15346));
  AOI21xp33_ASAP7_75t_L     g15090(.A1(new_n15342), .A2(new_n15346), .B(new_n15311), .Y(new_n15347));
  AND3x1_ASAP7_75t_L        g15091(.A(new_n15342), .B(new_n15346), .C(new_n15311), .Y(new_n15348));
  NOR2xp33_ASAP7_75t_L      g15092(.A(new_n15347), .B(new_n15348), .Y(new_n15349));
  A2O1A1Ixp33_ASAP7_75t_L   g15093(.A1(new_n15307), .A2(new_n15306), .B(new_n15177), .C(new_n15349), .Y(new_n15350));
  NOR2xp33_ASAP7_75t_L      g15094(.A(new_n15173), .B(new_n15170), .Y(new_n15351));
  O2A1O1Ixp33_ASAP7_75t_L   g15095(.A1(new_n15013), .A2(new_n15015), .B(new_n15175), .C(new_n15351), .Y(new_n15352));
  OAI21xp33_ASAP7_75t_L     g15096(.A1(new_n15347), .A2(new_n15348), .B(new_n15352), .Y(new_n15353));
  NAND2xp33_ASAP7_75t_L     g15097(.A(new_n15350), .B(new_n15353), .Y(new_n15354));
  NAND2xp33_ASAP7_75t_L     g15098(.A(\b[29] ), .B(new_n8537), .Y(new_n15355));
  OAI221xp5_ASAP7_75t_L     g15099(.A1(new_n8243), .A2(new_n3180), .B1(new_n7957), .B2(new_n3187), .C(new_n15355), .Y(new_n15356));
  AOI21xp33_ASAP7_75t_L     g15100(.A1(new_n7963), .A2(\b[30] ), .B(new_n15356), .Y(new_n15357));
  NAND2xp33_ASAP7_75t_L     g15101(.A(\a[53] ), .B(new_n15357), .Y(new_n15358));
  A2O1A1Ixp33_ASAP7_75t_L   g15102(.A1(\b[30] ), .A2(new_n7963), .B(new_n15356), .C(new_n7954), .Y(new_n15359));
  NAND2xp33_ASAP7_75t_L     g15103(.A(new_n15359), .B(new_n15358), .Y(new_n15360));
  XNOR2x2_ASAP7_75t_L       g15104(.A(new_n15360), .B(new_n15354), .Y(new_n15361));
  OAI31xp33_ASAP7_75t_L     g15105(.A1(new_n15176), .A2(new_n15181), .A3(new_n15177), .B(new_n15187), .Y(new_n15362));
  XNOR2x2_ASAP7_75t_L       g15106(.A(new_n15361), .B(new_n15362), .Y(new_n15363));
  AOI22xp33_ASAP7_75t_L     g15107(.A1(new_n7111), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n7391), .Y(new_n15364));
  OAI221xp5_ASAP7_75t_L     g15108(.A1(new_n8558), .A2(new_n3565), .B1(new_n8237), .B2(new_n3591), .C(new_n15364), .Y(new_n15365));
  XNOR2x2_ASAP7_75t_L       g15109(.A(\a[50] ), .B(new_n15365), .Y(new_n15366));
  XNOR2x2_ASAP7_75t_L       g15110(.A(new_n15366), .B(new_n15363), .Y(new_n15367));
  AOI211xp5_ASAP7_75t_L     g15111(.A1(new_n15031), .A2(new_n14988), .B(new_n15032), .C(new_n15191), .Y(new_n15368));
  A2O1A1Ixp33_ASAP7_75t_L   g15112(.A1(new_n15031), .A2(new_n14988), .B(new_n15032), .C(new_n15191), .Y(new_n15369));
  A2O1A1Ixp33_ASAP7_75t_L   g15113(.A1(new_n15187), .A2(new_n15184), .B(new_n15368), .C(new_n15369), .Y(new_n15370));
  NAND2xp33_ASAP7_75t_L     g15114(.A(new_n15370), .B(new_n15367), .Y(new_n15371));
  NOR2xp33_ASAP7_75t_L      g15115(.A(new_n15370), .B(new_n15367), .Y(new_n15372));
  INVx1_ASAP7_75t_L         g15116(.A(new_n15372), .Y(new_n15373));
  AND2x2_ASAP7_75t_L        g15117(.A(new_n15371), .B(new_n15373), .Y(new_n15374));
  AOI22xp33_ASAP7_75t_L     g15118(.A1(new_n6376), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n6648), .Y(new_n15375));
  OAI221xp5_ASAP7_75t_L     g15119(.A1(new_n6646), .A2(new_n4216), .B1(new_n6636), .B2(new_n4431), .C(new_n15375), .Y(new_n15376));
  XNOR2x2_ASAP7_75t_L       g15120(.A(\a[47] ), .B(new_n15376), .Y(new_n15377));
  XNOR2x2_ASAP7_75t_L       g15121(.A(new_n15377), .B(new_n15374), .Y(new_n15378));
  XOR2x2_ASAP7_75t_L        g15122(.A(new_n15305), .B(new_n15378), .Y(new_n15379));
  NAND2xp33_ASAP7_75t_L     g15123(.A(new_n15304), .B(new_n15379), .Y(new_n15380));
  INVx1_ASAP7_75t_L         g15124(.A(new_n15379), .Y(new_n15381));
  NAND2xp33_ASAP7_75t_L     g15125(.A(new_n15303), .B(new_n15381), .Y(new_n15382));
  NAND3xp33_ASAP7_75t_L     g15126(.A(new_n15382), .B(new_n15380), .C(new_n15300), .Y(new_n15383));
  INVx1_ASAP7_75t_L         g15127(.A(new_n15300), .Y(new_n15384));
  INVx1_ASAP7_75t_L         g15128(.A(new_n15380), .Y(new_n15385));
  NOR2xp33_ASAP7_75t_L      g15129(.A(new_n15304), .B(new_n15379), .Y(new_n15386));
  OAI21xp33_ASAP7_75t_L     g15130(.A1(new_n15386), .A2(new_n15385), .B(new_n15384), .Y(new_n15387));
  NAND2xp33_ASAP7_75t_L     g15131(.A(new_n15383), .B(new_n15387), .Y(new_n15388));
  AOI22xp33_ASAP7_75t_L     g15132(.A1(new_n4920), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n5167), .Y(new_n15389));
  OAI221xp5_ASAP7_75t_L     g15133(.A1(new_n5154), .A2(new_n5338), .B1(new_n5158), .B2(new_n6338), .C(new_n15389), .Y(new_n15390));
  XNOR2x2_ASAP7_75t_L       g15134(.A(new_n4915), .B(new_n15390), .Y(new_n15391));
  XNOR2x2_ASAP7_75t_L       g15135(.A(new_n15391), .B(new_n15388), .Y(new_n15392));
  NAND2xp33_ASAP7_75t_L     g15136(.A(new_n15212), .B(new_n15215), .Y(new_n15393));
  XNOR2x2_ASAP7_75t_L       g15137(.A(new_n15393), .B(new_n15392), .Y(new_n15394));
  AOI22xp33_ASAP7_75t_L     g15138(.A1(new_n4283), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n4512), .Y(new_n15395));
  OAI221xp5_ASAP7_75t_L     g15139(.A1(new_n4277), .A2(new_n6321), .B1(new_n4499), .B2(new_n6573), .C(new_n15395), .Y(new_n15396));
  XNOR2x2_ASAP7_75t_L       g15140(.A(\a[38] ), .B(new_n15396), .Y(new_n15397));
  INVx1_ASAP7_75t_L         g15141(.A(new_n15397), .Y(new_n15398));
  XNOR2x2_ASAP7_75t_L       g15142(.A(new_n15398), .B(new_n15394), .Y(new_n15399));
  OAI21xp33_ASAP7_75t_L     g15143(.A1(new_n15216), .A2(new_n15219), .B(new_n15226), .Y(new_n15400));
  NOR2xp33_ASAP7_75t_L      g15144(.A(new_n15400), .B(new_n15399), .Y(new_n15401));
  INVx1_ASAP7_75t_L         g15145(.A(new_n15401), .Y(new_n15402));
  NAND2xp33_ASAP7_75t_L     g15146(.A(new_n15400), .B(new_n15399), .Y(new_n15403));
  AOI22xp33_ASAP7_75t_L     g15147(.A1(new_n3633), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n3858), .Y(new_n15404));
  OAI221xp5_ASAP7_75t_L     g15148(.A1(new_n3853), .A2(new_n6830), .B1(new_n3856), .B2(new_n7323), .C(new_n15404), .Y(new_n15405));
  XNOR2x2_ASAP7_75t_L       g15149(.A(\a[35] ), .B(new_n15405), .Y(new_n15406));
  NAND3xp33_ASAP7_75t_L     g15150(.A(new_n15402), .B(new_n15403), .C(new_n15406), .Y(new_n15407));
  AO21x2_ASAP7_75t_L        g15151(.A1(new_n15403), .A2(new_n15402), .B(new_n15406), .Y(new_n15408));
  AO21x2_ASAP7_75t_L        g15152(.A1(new_n15408), .A2(new_n15407), .B(new_n15299), .Y(new_n15409));
  NAND3xp33_ASAP7_75t_L     g15153(.A(new_n15299), .B(new_n15407), .C(new_n15408), .Y(new_n15410));
  NAND2xp33_ASAP7_75t_L     g15154(.A(new_n15410), .B(new_n15409), .Y(new_n15411));
  XNOR2x2_ASAP7_75t_L       g15155(.A(new_n15292), .B(new_n15411), .Y(new_n15412));
  NOR2xp33_ASAP7_75t_L      g15156(.A(new_n15412), .B(new_n15287), .Y(new_n15413));
  AND2x2_ASAP7_75t_L        g15157(.A(new_n15412), .B(new_n15287), .Y(new_n15414));
  OR2x4_ASAP7_75t_L         g15158(.A(new_n15413), .B(new_n15414), .Y(new_n15415));
  NAND2xp33_ASAP7_75t_L     g15159(.A(new_n15415), .B(new_n15282), .Y(new_n15416));
  OR3x1_ASAP7_75t_L         g15160(.A(new_n15282), .B(new_n15413), .C(new_n15414), .Y(new_n15417));
  NAND2xp33_ASAP7_75t_L     g15161(.A(new_n15416), .B(new_n15417), .Y(new_n15418));
  NOR2xp33_ASAP7_75t_L      g15162(.A(new_n1359), .B(new_n11500), .Y(new_n15419));
  AOI21xp33_ASAP7_75t_L     g15163(.A1(new_n1581), .A2(\b[62] ), .B(new_n15419), .Y(new_n15420));
  OAI211xp5_ASAP7_75t_L     g15164(.A1(new_n11468), .A2(new_n1373), .B(new_n15420), .C(\a[20] ), .Y(new_n15421));
  O2A1O1Ixp33_ASAP7_75t_L   g15165(.A1(new_n11468), .A2(new_n1373), .B(new_n15420), .C(\a[20] ), .Y(new_n15422));
  INVx1_ASAP7_75t_L         g15166(.A(new_n15422), .Y(new_n15423));
  NAND2xp33_ASAP7_75t_L     g15167(.A(new_n15421), .B(new_n15423), .Y(new_n15424));
  NAND3xp33_ASAP7_75t_L     g15168(.A(new_n15257), .B(new_n15121), .C(new_n15424), .Y(new_n15425));
  O2A1O1Ixp33_ASAP7_75t_L   g15169(.A1(new_n15123), .A2(new_n15256), .B(new_n15121), .C(new_n15424), .Y(new_n15426));
  INVx1_ASAP7_75t_L         g15170(.A(new_n15426), .Y(new_n15427));
  NAND3xp33_ASAP7_75t_L     g15171(.A(new_n15418), .B(new_n15425), .C(new_n15427), .Y(new_n15428));
  INVx1_ASAP7_75t_L         g15172(.A(new_n15428), .Y(new_n15429));
  AOI21xp33_ASAP7_75t_L     g15173(.A1(new_n15425), .A2(new_n15427), .B(new_n15418), .Y(new_n15430));
  NOR3xp33_ASAP7_75t_L      g15174(.A(new_n15429), .B(new_n15430), .C(new_n15274), .Y(new_n15431));
  OA21x2_ASAP7_75t_L        g15175(.A1(new_n15430), .A2(new_n15429), .B(new_n15274), .Y(new_n15432));
  NOR2xp33_ASAP7_75t_L      g15176(.A(new_n15431), .B(new_n15432), .Y(new_n15433));
  A2O1A1Ixp33_ASAP7_75t_L   g15177(.A1(new_n15269), .A2(new_n15265), .B(new_n15272), .C(new_n15433), .Y(new_n15434));
  INVx1_ASAP7_75t_L         g15178(.A(new_n15434), .Y(new_n15435));
  NAND2xp33_ASAP7_75t_L     g15179(.A(new_n15264), .B(new_n15263), .Y(new_n15436));
  A2O1A1Ixp33_ASAP7_75t_L   g15180(.A1(new_n15097), .A2(new_n15268), .B(new_n15436), .C(new_n15263), .Y(new_n15437));
  NOR2xp33_ASAP7_75t_L      g15181(.A(new_n15433), .B(new_n15437), .Y(new_n15438));
  NOR2xp33_ASAP7_75t_L      g15182(.A(new_n15438), .B(new_n15435), .Y(\f[82] ));
  INVx1_ASAP7_75t_L         g15183(.A(new_n15418), .Y(new_n15440));
  NAND2xp33_ASAP7_75t_L     g15184(.A(new_n15427), .B(new_n15425), .Y(new_n15441));
  A2O1A1Ixp33_ASAP7_75t_L   g15185(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n1365), .Y(new_n15442));
  A2O1A1Ixp33_ASAP7_75t_L   g15186(.A1(new_n15442), .A2(new_n1483), .B(new_n11468), .C(\a[20] ), .Y(new_n15443));
  O2A1O1Ixp33_ASAP7_75t_L   g15187(.A1(new_n1359), .A2(new_n12060), .B(new_n1483), .C(new_n11468), .Y(new_n15444));
  NAND2xp33_ASAP7_75t_L     g15188(.A(new_n1356), .B(new_n15444), .Y(new_n15445));
  AND2x2_ASAP7_75t_L        g15189(.A(new_n15445), .B(new_n15443), .Y(new_n15446));
  INVx1_ASAP7_75t_L         g15190(.A(new_n15446), .Y(new_n15447));
  INVx1_ASAP7_75t_L         g15191(.A(new_n15279), .Y(new_n15448));
  O2A1O1Ixp33_ASAP7_75t_L   g15192(.A1(new_n15413), .A2(new_n15414), .B(new_n15281), .C(new_n15448), .Y(new_n15449));
  NAND2xp33_ASAP7_75t_L     g15193(.A(new_n15447), .B(new_n15449), .Y(new_n15450));
  A2O1A1Ixp33_ASAP7_75t_L   g15194(.A1(new_n15281), .A2(new_n15415), .B(new_n15448), .C(new_n15446), .Y(new_n15451));
  AOI22xp33_ASAP7_75t_L     g15195(.A1(new_n1704), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n1837), .Y(new_n15452));
  OAI221xp5_ASAP7_75t_L     g15196(.A1(new_n1699), .A2(new_n10847), .B1(new_n1827), .B2(new_n12047), .C(new_n15452), .Y(new_n15453));
  XNOR2x2_ASAP7_75t_L       g15197(.A(\a[23] ), .B(new_n15453), .Y(new_n15454));
  INVx1_ASAP7_75t_L         g15198(.A(new_n15454), .Y(new_n15455));
  NOR2xp33_ASAP7_75t_L      g15199(.A(new_n15285), .B(new_n15286), .Y(new_n15456));
  NOR2xp33_ASAP7_75t_L      g15200(.A(new_n15456), .B(new_n15413), .Y(new_n15457));
  XNOR2x2_ASAP7_75t_L       g15201(.A(new_n15455), .B(new_n15457), .Y(new_n15458));
  AOI22xp33_ASAP7_75t_L     g15202(.A1(new_n2114), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n2259), .Y(new_n15459));
  OAI221xp5_ASAP7_75t_L     g15203(.A1(new_n2109), .A2(new_n9920), .B1(new_n2257), .B2(new_n11152), .C(new_n15459), .Y(new_n15460));
  XNOR2x2_ASAP7_75t_L       g15204(.A(new_n2100), .B(new_n15460), .Y(new_n15461));
  MAJIxp5_ASAP7_75t_L       g15205(.A(new_n15411), .B(new_n15290), .C(new_n15291), .Y(new_n15462));
  OR2x4_ASAP7_75t_L         g15206(.A(new_n15461), .B(new_n15462), .Y(new_n15463));
  NAND2xp33_ASAP7_75t_L     g15207(.A(new_n15461), .B(new_n15462), .Y(new_n15464));
  NAND2xp33_ASAP7_75t_L     g15208(.A(new_n15464), .B(new_n15463), .Y(new_n15465));
  AOI22xp33_ASAP7_75t_L     g15209(.A1(new_n2552), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n2736), .Y(new_n15466));
  OAI221xp5_ASAP7_75t_L     g15210(.A1(new_n2547), .A2(new_n8762), .B1(new_n2734), .B2(new_n9331), .C(new_n15466), .Y(new_n15467));
  XNOR2x2_ASAP7_75t_L       g15211(.A(\a[29] ), .B(new_n15467), .Y(new_n15468));
  A2O1A1Ixp33_ASAP7_75t_L   g15212(.A1(new_n15407), .A2(new_n15408), .B(new_n15299), .C(new_n15298), .Y(new_n15469));
  XNOR2x2_ASAP7_75t_L       g15213(.A(new_n15468), .B(new_n15469), .Y(new_n15470));
  AOI22xp33_ASAP7_75t_L     g15214(.A1(new_n3029), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n3258), .Y(new_n15471));
  OAI221xp5_ASAP7_75t_L     g15215(.A1(new_n3024), .A2(new_n7900), .B1(new_n3256), .B2(new_n8174), .C(new_n15471), .Y(new_n15472));
  XNOR2x2_ASAP7_75t_L       g15216(.A(\a[32] ), .B(new_n15472), .Y(new_n15473));
  AOI21xp33_ASAP7_75t_L     g15217(.A1(new_n15403), .A2(new_n15406), .B(new_n15401), .Y(new_n15474));
  XNOR2x2_ASAP7_75t_L       g15218(.A(new_n15473), .B(new_n15474), .Y(new_n15475));
  AOI22xp33_ASAP7_75t_L     g15219(.A1(new_n4920), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n5167), .Y(new_n15476));
  OAI221xp5_ASAP7_75t_L     g15220(.A1(new_n5154), .A2(new_n5805), .B1(new_n5158), .B2(new_n5835), .C(new_n15476), .Y(new_n15477));
  XNOR2x2_ASAP7_75t_L       g15221(.A(\a[41] ), .B(new_n15477), .Y(new_n15478));
  INVx1_ASAP7_75t_L         g15222(.A(new_n15478), .Y(new_n15479));
  INVx1_ASAP7_75t_L         g15223(.A(new_n15378), .Y(new_n15480));
  A2O1A1Ixp33_ASAP7_75t_L   g15224(.A1(new_n15203), .A2(new_n15199), .B(new_n15480), .C(new_n15380), .Y(new_n15481));
  AOI22xp33_ASAP7_75t_L     g15225(.A1(new_n5624), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n5901), .Y(new_n15482));
  OAI221xp5_ASAP7_75t_L     g15226(.A1(new_n5900), .A2(new_n4869), .B1(new_n5892), .B2(new_n5327), .C(new_n15482), .Y(new_n15483));
  XNOR2x2_ASAP7_75t_L       g15227(.A(\a[44] ), .B(new_n15483), .Y(new_n15484));
  INVx1_ASAP7_75t_L         g15228(.A(new_n15484), .Y(new_n15485));
  INVx1_ASAP7_75t_L         g15229(.A(new_n15374), .Y(new_n15486));
  AOI22xp33_ASAP7_75t_L     g15230(.A1(new_n6376), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n6648), .Y(new_n15487));
  OAI221xp5_ASAP7_75t_L     g15231(.A1(new_n6646), .A2(new_n4424), .B1(new_n6636), .B2(new_n4641), .C(new_n15487), .Y(new_n15488));
  XNOR2x2_ASAP7_75t_L       g15232(.A(\a[47] ), .B(new_n15488), .Y(new_n15489));
  INVx1_ASAP7_75t_L         g15233(.A(new_n15489), .Y(new_n15490));
  AOI22xp33_ASAP7_75t_L     g15234(.A1(new_n7111), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n7391), .Y(new_n15491));
  OAI221xp5_ASAP7_75t_L     g15235(.A1(new_n8558), .A2(new_n3584), .B1(new_n8237), .B2(new_n10137), .C(new_n15491), .Y(new_n15492));
  XNOR2x2_ASAP7_75t_L       g15236(.A(\a[50] ), .B(new_n15492), .Y(new_n15493));
  INVx1_ASAP7_75t_L         g15237(.A(new_n15493), .Y(new_n15494));
  AOI22xp33_ASAP7_75t_L     g15238(.A1(new_n7960), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n8537), .Y(new_n15495));
  OAI221xp5_ASAP7_75t_L     g15239(.A1(new_n8817), .A2(new_n3180), .B1(new_n7957), .B2(new_n11047), .C(new_n15495), .Y(new_n15496));
  XNOR2x2_ASAP7_75t_L       g15240(.A(\a[53] ), .B(new_n15496), .Y(new_n15497));
  AOI22xp33_ASAP7_75t_L     g15241(.A1(new_n9700), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n10027), .Y(new_n15498));
  OAI221xp5_ASAP7_75t_L     g15242(.A1(new_n10024), .A2(new_n2067), .B1(new_n9696), .B2(new_n2355), .C(new_n15498), .Y(new_n15499));
  XNOR2x2_ASAP7_75t_L       g15243(.A(\a[59] ), .B(new_n15499), .Y(new_n15500));
  INVx1_ASAP7_75t_L         g15244(.A(new_n15500), .Y(new_n15501));
  NOR2xp33_ASAP7_75t_L      g15245(.A(new_n1432), .B(new_n11535), .Y(new_n15502));
  O2A1O1Ixp33_ASAP7_75t_L   g15246(.A1(new_n11247), .A2(new_n11249), .B(\b[20] ), .C(new_n15502), .Y(new_n15503));
  A2O1A1Ixp33_ASAP7_75t_L   g15247(.A1(new_n11533), .A2(\b[19] ), .B(new_n15313), .C(new_n15503), .Y(new_n15504));
  A2O1A1Ixp33_ASAP7_75t_L   g15248(.A1(\b[20] ), .A2(new_n11533), .B(new_n15502), .C(new_n15317), .Y(new_n15505));
  NAND2xp33_ASAP7_75t_L     g15249(.A(new_n15505), .B(new_n15504), .Y(new_n15506));
  NOR2xp33_ASAP7_75t_L      g15250(.A(new_n1909), .B(new_n10630), .Y(new_n15507));
  AOI221xp5_ASAP7_75t_L     g15251(.A1(\b[21] ), .A2(new_n10939), .B1(\b[22] ), .B2(new_n10632), .C(new_n15507), .Y(new_n15508));
  OAI211xp5_ASAP7_75t_L     g15252(.A1(new_n10629), .A2(new_n1915), .B(\a[62] ), .C(new_n15508), .Y(new_n15509));
  O2A1O1Ixp33_ASAP7_75t_L   g15253(.A1(new_n10629), .A2(new_n1915), .B(new_n15508), .C(\a[62] ), .Y(new_n15510));
  INVx1_ASAP7_75t_L         g15254(.A(new_n15510), .Y(new_n15511));
  AND2x2_ASAP7_75t_L        g15255(.A(new_n15509), .B(new_n15511), .Y(new_n15512));
  NOR2xp33_ASAP7_75t_L      g15256(.A(new_n15506), .B(new_n15512), .Y(new_n15513));
  AND3x1_ASAP7_75t_L        g15257(.A(new_n15511), .B(new_n15509), .C(new_n15506), .Y(new_n15514));
  NOR2xp33_ASAP7_75t_L      g15258(.A(new_n15514), .B(new_n15513), .Y(new_n15515));
  INVx1_ASAP7_75t_L         g15259(.A(new_n15515), .Y(new_n15516));
  O2A1O1Ixp33_ASAP7_75t_L   g15260(.A1(new_n15321), .A2(new_n15324), .B(new_n15320), .C(new_n15516), .Y(new_n15517));
  INVx1_ASAP7_75t_L         g15261(.A(new_n15517), .Y(new_n15518));
  A2O1A1O1Ixp25_ASAP7_75t_L g15262(.A1(new_n15147), .A2(new_n15151), .B(new_n15314), .C(new_n15317), .D(new_n15326), .Y(new_n15519));
  NAND2xp33_ASAP7_75t_L     g15263(.A(new_n15519), .B(new_n15516), .Y(new_n15520));
  NAND3xp33_ASAP7_75t_L     g15264(.A(new_n15518), .B(new_n15501), .C(new_n15520), .Y(new_n15521));
  AO21x2_ASAP7_75t_L        g15265(.A1(new_n15518), .A2(new_n15520), .B(new_n15501), .Y(new_n15522));
  AND2x2_ASAP7_75t_L        g15266(.A(new_n15521), .B(new_n15522), .Y(new_n15523));
  NAND3xp33_ASAP7_75t_L     g15267(.A(new_n15523), .B(new_n15338), .C(new_n15334), .Y(new_n15524));
  O2A1O1Ixp33_ASAP7_75t_L   g15268(.A1(new_n15328), .A2(new_n15332), .B(new_n15338), .C(new_n15523), .Y(new_n15525));
  INVx1_ASAP7_75t_L         g15269(.A(new_n15525), .Y(new_n15526));
  AOI22xp33_ASAP7_75t_L     g15270(.A1(new_n8831), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n9115), .Y(new_n15527));
  OAI221xp5_ASAP7_75t_L     g15271(.A1(new_n10343), .A2(new_n2666), .B1(new_n10016), .B2(new_n2695), .C(new_n15527), .Y(new_n15528));
  XNOR2x2_ASAP7_75t_L       g15272(.A(\a[56] ), .B(new_n15528), .Y(new_n15529));
  NAND3xp33_ASAP7_75t_L     g15273(.A(new_n15526), .B(new_n15524), .C(new_n15529), .Y(new_n15530));
  AO21x2_ASAP7_75t_L        g15274(.A1(new_n15524), .A2(new_n15526), .B(new_n15529), .Y(new_n15531));
  NAND2xp33_ASAP7_75t_L     g15275(.A(new_n15530), .B(new_n15531), .Y(new_n15532));
  A2O1A1Ixp33_ASAP7_75t_L   g15276(.A1(new_n15346), .A2(new_n15311), .B(new_n15341), .C(new_n15532), .Y(new_n15533));
  OR3x1_ASAP7_75t_L         g15277(.A(new_n15532), .B(new_n15341), .C(new_n15348), .Y(new_n15534));
  NAND3xp33_ASAP7_75t_L     g15278(.A(new_n15534), .B(new_n15533), .C(new_n15497), .Y(new_n15535));
  AO21x2_ASAP7_75t_L        g15279(.A1(new_n15533), .A2(new_n15534), .B(new_n15497), .Y(new_n15536));
  AND2x2_ASAP7_75t_L        g15280(.A(new_n15535), .B(new_n15536), .Y(new_n15537));
  OAI21xp33_ASAP7_75t_L     g15281(.A1(new_n15360), .A2(new_n15354), .B(new_n15353), .Y(new_n15538));
  NOR2xp33_ASAP7_75t_L      g15282(.A(new_n15538), .B(new_n15537), .Y(new_n15539));
  INVx1_ASAP7_75t_L         g15283(.A(new_n15539), .Y(new_n15540));
  NAND2xp33_ASAP7_75t_L     g15284(.A(new_n15538), .B(new_n15537), .Y(new_n15541));
  AND2x2_ASAP7_75t_L        g15285(.A(new_n15541), .B(new_n15540), .Y(new_n15542));
  NAND2xp33_ASAP7_75t_L     g15286(.A(new_n15494), .B(new_n15542), .Y(new_n15543));
  AO21x2_ASAP7_75t_L        g15287(.A1(new_n15541), .A2(new_n15540), .B(new_n15494), .Y(new_n15544));
  NAND2xp33_ASAP7_75t_L     g15288(.A(new_n15544), .B(new_n15543), .Y(new_n15545));
  INVx1_ASAP7_75t_L         g15289(.A(new_n15366), .Y(new_n15546));
  MAJIxp5_ASAP7_75t_L       g15290(.A(new_n15362), .B(new_n15361), .C(new_n15546), .Y(new_n15547));
  NOR2xp33_ASAP7_75t_L      g15291(.A(new_n15547), .B(new_n15545), .Y(new_n15548));
  INVx1_ASAP7_75t_L         g15292(.A(new_n15548), .Y(new_n15549));
  NAND2xp33_ASAP7_75t_L     g15293(.A(new_n15547), .B(new_n15545), .Y(new_n15550));
  AND2x2_ASAP7_75t_L        g15294(.A(new_n15550), .B(new_n15549), .Y(new_n15551));
  NAND2xp33_ASAP7_75t_L     g15295(.A(new_n15490), .B(new_n15551), .Y(new_n15552));
  AO21x2_ASAP7_75t_L        g15296(.A1(new_n15550), .A2(new_n15549), .B(new_n15490), .Y(new_n15553));
  NAND2xp33_ASAP7_75t_L     g15297(.A(new_n15553), .B(new_n15552), .Y(new_n15554));
  O2A1O1Ixp33_ASAP7_75t_L   g15298(.A1(new_n15377), .A2(new_n15486), .B(new_n15373), .C(new_n15554), .Y(new_n15555));
  OA21x2_ASAP7_75t_L        g15299(.A1(new_n15377), .A2(new_n15486), .B(new_n15373), .Y(new_n15556));
  AND2x2_ASAP7_75t_L        g15300(.A(new_n15554), .B(new_n15556), .Y(new_n15557));
  NOR2xp33_ASAP7_75t_L      g15301(.A(new_n15557), .B(new_n15555), .Y(new_n15558));
  XNOR2x2_ASAP7_75t_L       g15302(.A(new_n15485), .B(new_n15558), .Y(new_n15559));
  XNOR2x2_ASAP7_75t_L       g15303(.A(new_n15481), .B(new_n15559), .Y(new_n15560));
  XNOR2x2_ASAP7_75t_L       g15304(.A(new_n15479), .B(new_n15560), .Y(new_n15561));
  NOR2xp33_ASAP7_75t_L      g15305(.A(new_n15391), .B(new_n15388), .Y(new_n15562));
  O2A1O1Ixp33_ASAP7_75t_L   g15306(.A1(new_n15385), .A2(new_n15386), .B(new_n15384), .C(new_n15562), .Y(new_n15563));
  XNOR2x2_ASAP7_75t_L       g15307(.A(new_n15563), .B(new_n15561), .Y(new_n15564));
  AOI22xp33_ASAP7_75t_L     g15308(.A1(new_n4283), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n4512), .Y(new_n15565));
  OAI221xp5_ASAP7_75t_L     g15309(.A1(new_n4277), .A2(new_n6568), .B1(new_n4499), .B2(new_n6820), .C(new_n15565), .Y(new_n15566));
  XNOR2x2_ASAP7_75t_L       g15310(.A(\a[38] ), .B(new_n15566), .Y(new_n15567));
  XNOR2x2_ASAP7_75t_L       g15311(.A(new_n15567), .B(new_n15564), .Y(new_n15568));
  MAJIxp5_ASAP7_75t_L       g15312(.A(new_n15392), .B(new_n15393), .C(new_n15398), .Y(new_n15569));
  XNOR2x2_ASAP7_75t_L       g15313(.A(new_n15569), .B(new_n15568), .Y(new_n15570));
  AOI22xp33_ASAP7_75t_L     g15314(.A1(new_n3633), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n3858), .Y(new_n15571));
  OAI221xp5_ASAP7_75t_L     g15315(.A1(new_n3853), .A2(new_n7317), .B1(new_n3856), .B2(new_n7602), .C(new_n15571), .Y(new_n15572));
  XNOR2x2_ASAP7_75t_L       g15316(.A(\a[35] ), .B(new_n15572), .Y(new_n15573));
  INVx1_ASAP7_75t_L         g15317(.A(new_n15573), .Y(new_n15574));
  NAND2xp33_ASAP7_75t_L     g15318(.A(new_n15574), .B(new_n15570), .Y(new_n15575));
  INVx1_ASAP7_75t_L         g15319(.A(new_n15575), .Y(new_n15576));
  NOR2xp33_ASAP7_75t_L      g15320(.A(new_n15574), .B(new_n15570), .Y(new_n15577));
  NOR2xp33_ASAP7_75t_L      g15321(.A(new_n15576), .B(new_n15577), .Y(new_n15578));
  XNOR2x2_ASAP7_75t_L       g15322(.A(new_n15475), .B(new_n15578), .Y(new_n15579));
  XNOR2x2_ASAP7_75t_L       g15323(.A(new_n15470), .B(new_n15579), .Y(new_n15580));
  XNOR2x2_ASAP7_75t_L       g15324(.A(new_n15580), .B(new_n15465), .Y(new_n15581));
  NAND2xp33_ASAP7_75t_L     g15325(.A(new_n15581), .B(new_n15458), .Y(new_n15582));
  INVx1_ASAP7_75t_L         g15326(.A(new_n15582), .Y(new_n15583));
  NOR2xp33_ASAP7_75t_L      g15327(.A(new_n15581), .B(new_n15458), .Y(new_n15584));
  NOR2xp33_ASAP7_75t_L      g15328(.A(new_n15584), .B(new_n15583), .Y(new_n15585));
  NAND3xp33_ASAP7_75t_L     g15329(.A(new_n15585), .B(new_n15451), .C(new_n15450), .Y(new_n15586));
  NAND2xp33_ASAP7_75t_L     g15330(.A(new_n15451), .B(new_n15450), .Y(new_n15587));
  OAI21xp33_ASAP7_75t_L     g15331(.A1(new_n15584), .A2(new_n15583), .B(new_n15587), .Y(new_n15588));
  NAND2xp33_ASAP7_75t_L     g15332(.A(new_n15588), .B(new_n15586), .Y(new_n15589));
  O2A1O1Ixp33_ASAP7_75t_L   g15333(.A1(new_n15440), .A2(new_n15441), .B(new_n15425), .C(new_n15589), .Y(new_n15590));
  INVx1_ASAP7_75t_L         g15334(.A(new_n15590), .Y(new_n15591));
  NAND3xp33_ASAP7_75t_L     g15335(.A(new_n15589), .B(new_n15428), .C(new_n15425), .Y(new_n15592));
  NAND2xp33_ASAP7_75t_L     g15336(.A(new_n15592), .B(new_n15591), .Y(new_n15593));
  INVx1_ASAP7_75t_L         g15337(.A(new_n15593), .Y(new_n15594));
  A2O1A1Ixp33_ASAP7_75t_L   g15338(.A1(new_n15437), .A2(new_n15433), .B(new_n15431), .C(new_n15594), .Y(new_n15595));
  INVx1_ASAP7_75t_L         g15339(.A(new_n15595), .Y(new_n15596));
  INVx1_ASAP7_75t_L         g15340(.A(new_n15431), .Y(new_n15597));
  A2O1A1Ixp33_ASAP7_75t_L   g15341(.A1(new_n15266), .A2(new_n15263), .B(new_n15432), .C(new_n15597), .Y(new_n15598));
  NOR2xp33_ASAP7_75t_L      g15342(.A(new_n15594), .B(new_n15598), .Y(new_n15599));
  NOR2xp33_ASAP7_75t_L      g15343(.A(new_n15596), .B(new_n15599), .Y(\f[83] ));
  AOI22xp33_ASAP7_75t_L     g15344(.A1(new_n1704), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1837), .Y(new_n15601));
  A2O1A1Ixp33_ASAP7_75t_L   g15345(.A1(new_n11470), .A2(new_n11473), .B(new_n1827), .C(new_n15601), .Y(new_n15602));
  AOI21xp33_ASAP7_75t_L     g15346(.A1(new_n1706), .A2(\b[62] ), .B(new_n15602), .Y(new_n15603));
  NAND2xp33_ASAP7_75t_L     g15347(.A(\a[23] ), .B(new_n15603), .Y(new_n15604));
  A2O1A1Ixp33_ASAP7_75t_L   g15348(.A1(\b[62] ), .A2(new_n1706), .B(new_n15602), .C(new_n1689), .Y(new_n15605));
  AND2x2_ASAP7_75t_L        g15349(.A(new_n15605), .B(new_n15604), .Y(new_n15606));
  INVx1_ASAP7_75t_L         g15350(.A(new_n15606), .Y(new_n15607));
  O2A1O1Ixp33_ASAP7_75t_L   g15351(.A1(new_n15454), .A2(new_n15457), .B(new_n15582), .C(new_n15607), .Y(new_n15608));
  OAI21xp33_ASAP7_75t_L     g15352(.A1(new_n15454), .A2(new_n15457), .B(new_n15582), .Y(new_n15609));
  NOR2xp33_ASAP7_75t_L      g15353(.A(new_n15606), .B(new_n15609), .Y(new_n15610));
  NOR2xp33_ASAP7_75t_L      g15354(.A(new_n15608), .B(new_n15610), .Y(new_n15611));
  INVx1_ASAP7_75t_L         g15355(.A(new_n15611), .Y(new_n15612));
  AOI22xp33_ASAP7_75t_L     g15356(.A1(new_n2114), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n2259), .Y(new_n15613));
  OAI221xp5_ASAP7_75t_L     g15357(.A1(new_n2109), .A2(new_n9947), .B1(new_n2257), .B2(new_n11446), .C(new_n15613), .Y(new_n15614));
  XNOR2x2_ASAP7_75t_L       g15358(.A(\a[26] ), .B(new_n15614), .Y(new_n15615));
  INVx1_ASAP7_75t_L         g15359(.A(new_n15615), .Y(new_n15616));
  O2A1O1Ixp33_ASAP7_75t_L   g15360(.A1(new_n15580), .A2(new_n15465), .B(new_n15463), .C(new_n15616), .Y(new_n15617));
  OA211x2_ASAP7_75t_L       g15361(.A1(new_n15580), .A2(new_n15465), .B(new_n15463), .C(new_n15616), .Y(new_n15618));
  OR2x4_ASAP7_75t_L         g15362(.A(new_n15617), .B(new_n15618), .Y(new_n15619));
  INVx1_ASAP7_75t_L         g15363(.A(new_n15469), .Y(new_n15620));
  MAJIxp5_ASAP7_75t_L       g15364(.A(new_n15579), .B(new_n15468), .C(new_n15620), .Y(new_n15621));
  AOI22xp33_ASAP7_75t_L     g15365(.A1(new_n2552), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n2736), .Y(new_n15622));
  OAI221xp5_ASAP7_75t_L     g15366(.A1(new_n2547), .A2(new_n9323), .B1(new_n2734), .B2(new_n9627), .C(new_n15622), .Y(new_n15623));
  XNOR2x2_ASAP7_75t_L       g15367(.A(\a[29] ), .B(new_n15623), .Y(new_n15624));
  XNOR2x2_ASAP7_75t_L       g15368(.A(new_n15624), .B(new_n15621), .Y(new_n15625));
  AOI22xp33_ASAP7_75t_L     g15369(.A1(new_n3029), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n3258), .Y(new_n15626));
  OAI221xp5_ASAP7_75t_L     g15370(.A1(new_n3024), .A2(new_n8165), .B1(new_n3256), .B2(new_n8465), .C(new_n15626), .Y(new_n15627));
  XNOR2x2_ASAP7_75t_L       g15371(.A(\a[32] ), .B(new_n15627), .Y(new_n15628));
  A2O1A1Ixp33_ASAP7_75t_L   g15372(.A1(new_n15403), .A2(new_n15406), .B(new_n15401), .C(new_n15473), .Y(new_n15629));
  AOI211xp5_ASAP7_75t_L     g15373(.A1(new_n15403), .A2(new_n15406), .B(new_n15473), .C(new_n15401), .Y(new_n15630));
  AOI21xp33_ASAP7_75t_L     g15374(.A1(new_n15578), .A2(new_n15629), .B(new_n15630), .Y(new_n15631));
  XNOR2x2_ASAP7_75t_L       g15375(.A(new_n15628), .B(new_n15631), .Y(new_n15632));
  INVx1_ASAP7_75t_L         g15376(.A(new_n15568), .Y(new_n15633));
  OAI21xp33_ASAP7_75t_L     g15377(.A1(new_n15633), .A2(new_n15569), .B(new_n15575), .Y(new_n15634));
  INVx1_ASAP7_75t_L         g15378(.A(new_n15634), .Y(new_n15635));
  INVx1_ASAP7_75t_L         g15379(.A(new_n15563), .Y(new_n15636));
  AND2x2_ASAP7_75t_L        g15380(.A(new_n15567), .B(new_n15564), .Y(new_n15637));
  A2O1A1Ixp33_ASAP7_75t_L   g15381(.A1(new_n15536), .A2(new_n15535), .B(new_n15538), .C(new_n15543), .Y(new_n15638));
  AOI22xp33_ASAP7_75t_L     g15382(.A1(new_n9700), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n10027), .Y(new_n15639));
  OAI221xp5_ASAP7_75t_L     g15383(.A1(new_n10024), .A2(new_n2348), .B1(new_n9696), .B2(new_n2505), .C(new_n15639), .Y(new_n15640));
  XNOR2x2_ASAP7_75t_L       g15384(.A(\a[59] ), .B(new_n15640), .Y(new_n15641));
  INVx1_ASAP7_75t_L         g15385(.A(new_n15641), .Y(new_n15642));
  NOR2xp33_ASAP7_75t_L      g15386(.A(new_n1539), .B(new_n11535), .Y(new_n15643));
  A2O1A1Ixp33_ASAP7_75t_L   g15387(.A1(new_n11533), .A2(\b[21] ), .B(new_n15643), .C(new_n1356), .Y(new_n15644));
  INVx1_ASAP7_75t_L         g15388(.A(new_n15644), .Y(new_n15645));
  O2A1O1Ixp33_ASAP7_75t_L   g15389(.A1(new_n11247), .A2(new_n11249), .B(\b[21] ), .C(new_n15643), .Y(new_n15646));
  NAND2xp33_ASAP7_75t_L     g15390(.A(\a[20] ), .B(new_n15646), .Y(new_n15647));
  INVx1_ASAP7_75t_L         g15391(.A(new_n15647), .Y(new_n15648));
  NOR2xp33_ASAP7_75t_L      g15392(.A(new_n15645), .B(new_n15648), .Y(new_n15649));
  XNOR2x2_ASAP7_75t_L       g15393(.A(new_n15503), .B(new_n15649), .Y(new_n15650));
  INVx1_ASAP7_75t_L         g15394(.A(new_n15650), .Y(new_n15651));
  AOI22xp33_ASAP7_75t_L     g15395(.A1(\b[22] ), .A2(new_n10939), .B1(\b[24] ), .B2(new_n10938), .Y(new_n15652));
  OAI221xp5_ASAP7_75t_L     g15396(.A1(new_n10937), .A2(new_n1909), .B1(new_n10629), .B2(new_n2477), .C(new_n15652), .Y(new_n15653));
  XNOR2x2_ASAP7_75t_L       g15397(.A(\a[62] ), .B(new_n15653), .Y(new_n15654));
  XNOR2x2_ASAP7_75t_L       g15398(.A(new_n15651), .B(new_n15654), .Y(new_n15655));
  O2A1O1Ixp33_ASAP7_75t_L   g15399(.A1(new_n15506), .A2(new_n15512), .B(new_n15504), .C(new_n15655), .Y(new_n15656));
  INVx1_ASAP7_75t_L         g15400(.A(new_n15655), .Y(new_n15657));
  A2O1A1O1Ixp25_ASAP7_75t_L g15401(.A1(new_n11533), .A2(\b[19] ), .B(new_n15313), .C(new_n15503), .D(new_n15513), .Y(new_n15658));
  INVx1_ASAP7_75t_L         g15402(.A(new_n15658), .Y(new_n15659));
  NOR2xp33_ASAP7_75t_L      g15403(.A(new_n15659), .B(new_n15657), .Y(new_n15660));
  NOR2xp33_ASAP7_75t_L      g15404(.A(new_n15656), .B(new_n15660), .Y(new_n15661));
  XNOR2x2_ASAP7_75t_L       g15405(.A(new_n15642), .B(new_n15661), .Y(new_n15662));
  INVx1_ASAP7_75t_L         g15406(.A(new_n15662), .Y(new_n15663));
  A2O1A1Ixp33_ASAP7_75t_L   g15407(.A1(new_n15327), .A2(new_n15320), .B(new_n15516), .C(new_n15521), .Y(new_n15664));
  NOR2xp33_ASAP7_75t_L      g15408(.A(new_n15664), .B(new_n15663), .Y(new_n15665));
  O2A1O1Ixp33_ASAP7_75t_L   g15409(.A1(new_n15519), .A2(new_n15516), .B(new_n15521), .C(new_n15662), .Y(new_n15666));
  NOR2xp33_ASAP7_75t_L      g15410(.A(new_n15666), .B(new_n15665), .Y(new_n15667));
  AOI22xp33_ASAP7_75t_L     g15411(.A1(new_n8831), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n9115), .Y(new_n15668));
  OAI221xp5_ASAP7_75t_L     g15412(.A1(new_n10343), .A2(new_n2688), .B1(new_n10016), .B2(new_n2990), .C(new_n15668), .Y(new_n15669));
  XNOR2x2_ASAP7_75t_L       g15413(.A(\a[56] ), .B(new_n15669), .Y(new_n15670));
  INVx1_ASAP7_75t_L         g15414(.A(new_n15670), .Y(new_n15671));
  XNOR2x2_ASAP7_75t_L       g15415(.A(new_n15671), .B(new_n15667), .Y(new_n15672));
  A2O1A1Ixp33_ASAP7_75t_L   g15416(.A1(new_n15529), .A2(new_n15524), .B(new_n15525), .C(new_n15672), .Y(new_n15673));
  A2O1A1Ixp33_ASAP7_75t_L   g15417(.A1(new_n15338), .A2(new_n15334), .B(new_n15523), .C(new_n15530), .Y(new_n15674));
  OR2x4_ASAP7_75t_L         g15418(.A(new_n15674), .B(new_n15672), .Y(new_n15675));
  AND2x2_ASAP7_75t_L        g15419(.A(new_n15673), .B(new_n15675), .Y(new_n15676));
  AOI22xp33_ASAP7_75t_L     g15420(.A1(new_n7960), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n8537), .Y(new_n15677));
  OAI221xp5_ASAP7_75t_L     g15421(.A1(new_n8817), .A2(new_n3207), .B1(new_n7957), .B2(new_n3572), .C(new_n15677), .Y(new_n15678));
  XNOR2x2_ASAP7_75t_L       g15422(.A(\a[53] ), .B(new_n15678), .Y(new_n15679));
  INVx1_ASAP7_75t_L         g15423(.A(new_n15679), .Y(new_n15680));
  NAND2xp33_ASAP7_75t_L     g15424(.A(new_n15534), .B(new_n15535), .Y(new_n15681));
  XNOR2x2_ASAP7_75t_L       g15425(.A(new_n15680), .B(new_n15681), .Y(new_n15682));
  XNOR2x2_ASAP7_75t_L       g15426(.A(new_n15676), .B(new_n15682), .Y(new_n15683));
  AOI22xp33_ASAP7_75t_L     g15427(.A1(new_n7111), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n7391), .Y(new_n15684));
  OAI221xp5_ASAP7_75t_L     g15428(.A1(new_n8558), .A2(new_n3804), .B1(new_n8237), .B2(new_n4223), .C(new_n15684), .Y(new_n15685));
  XNOR2x2_ASAP7_75t_L       g15429(.A(\a[50] ), .B(new_n15685), .Y(new_n15686));
  NOR2xp33_ASAP7_75t_L      g15430(.A(new_n15686), .B(new_n15683), .Y(new_n15687));
  INVx1_ASAP7_75t_L         g15431(.A(new_n15687), .Y(new_n15688));
  NAND2xp33_ASAP7_75t_L     g15432(.A(new_n15686), .B(new_n15683), .Y(new_n15689));
  NAND2xp33_ASAP7_75t_L     g15433(.A(new_n15689), .B(new_n15688), .Y(new_n15690));
  XOR2x2_ASAP7_75t_L        g15434(.A(new_n15638), .B(new_n15690), .Y(new_n15691));
  AOI22xp33_ASAP7_75t_L     g15435(.A1(new_n6376), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n6648), .Y(new_n15692));
  OAI221xp5_ASAP7_75t_L     g15436(.A1(new_n6646), .A2(new_n4632), .B1(new_n6636), .B2(new_n4858), .C(new_n15692), .Y(new_n15693));
  XNOR2x2_ASAP7_75t_L       g15437(.A(\a[47] ), .B(new_n15693), .Y(new_n15694));
  XNOR2x2_ASAP7_75t_L       g15438(.A(new_n15694), .B(new_n15691), .Y(new_n15695));
  NAND3xp33_ASAP7_75t_L     g15439(.A(new_n15695), .B(new_n15552), .C(new_n15549), .Y(new_n15696));
  INVx1_ASAP7_75t_L         g15440(.A(new_n15695), .Y(new_n15697));
  A2O1A1Ixp33_ASAP7_75t_L   g15441(.A1(new_n15550), .A2(new_n15490), .B(new_n15548), .C(new_n15697), .Y(new_n15698));
  NAND2xp33_ASAP7_75t_L     g15442(.A(new_n15696), .B(new_n15698), .Y(new_n15699));
  AOI22xp33_ASAP7_75t_L     g15443(.A1(new_n5624), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n5901), .Y(new_n15700));
  OAI221xp5_ASAP7_75t_L     g15444(.A1(new_n5900), .A2(new_n5321), .B1(new_n5892), .B2(new_n5346), .C(new_n15700), .Y(new_n15701));
  XNOR2x2_ASAP7_75t_L       g15445(.A(\a[44] ), .B(new_n15701), .Y(new_n15702));
  XNOR2x2_ASAP7_75t_L       g15446(.A(new_n15702), .B(new_n15699), .Y(new_n15703));
  AOI21xp33_ASAP7_75t_L     g15447(.A1(new_n15558), .A2(new_n15485), .B(new_n15555), .Y(new_n15704));
  NAND2xp33_ASAP7_75t_L     g15448(.A(new_n15703), .B(new_n15704), .Y(new_n15705));
  INVx1_ASAP7_75t_L         g15449(.A(new_n15555), .Y(new_n15706));
  O2A1O1Ixp33_ASAP7_75t_L   g15450(.A1(new_n15484), .A2(new_n15557), .B(new_n15706), .C(new_n15703), .Y(new_n15707));
  INVx1_ASAP7_75t_L         g15451(.A(new_n15707), .Y(new_n15708));
  NAND2xp33_ASAP7_75t_L     g15452(.A(new_n15705), .B(new_n15708), .Y(new_n15709));
  AOI22xp33_ASAP7_75t_L     g15453(.A1(new_n4920), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n5167), .Y(new_n15710));
  OAI221xp5_ASAP7_75t_L     g15454(.A1(new_n5154), .A2(new_n5829), .B1(new_n5158), .B2(new_n6329), .C(new_n15710), .Y(new_n15711));
  XNOR2x2_ASAP7_75t_L       g15455(.A(\a[41] ), .B(new_n15711), .Y(new_n15712));
  XOR2x2_ASAP7_75t_L        g15456(.A(new_n15712), .B(new_n15709), .Y(new_n15713));
  A2O1A1O1Ixp25_ASAP7_75t_L g15457(.A1(new_n15203), .A2(new_n15199), .B(new_n15480), .C(new_n15380), .D(new_n15559), .Y(new_n15714));
  AOI21xp33_ASAP7_75t_L     g15458(.A1(new_n15560), .A2(new_n15479), .B(new_n15714), .Y(new_n15715));
  XOR2x2_ASAP7_75t_L        g15459(.A(new_n15715), .B(new_n15713), .Y(new_n15716));
  AOI22xp33_ASAP7_75t_L     g15460(.A1(new_n4283), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n4512), .Y(new_n15717));
  OAI221xp5_ASAP7_75t_L     g15461(.A1(new_n4277), .A2(new_n6812), .B1(new_n4499), .B2(new_n6837), .C(new_n15717), .Y(new_n15718));
  XNOR2x2_ASAP7_75t_L       g15462(.A(\a[38] ), .B(new_n15718), .Y(new_n15719));
  XNOR2x2_ASAP7_75t_L       g15463(.A(new_n15719), .B(new_n15716), .Y(new_n15720));
  A2O1A1Ixp33_ASAP7_75t_L   g15464(.A1(new_n15636), .A2(new_n15561), .B(new_n15637), .C(new_n15720), .Y(new_n15721));
  INVx1_ASAP7_75t_L         g15465(.A(new_n15720), .Y(new_n15722));
  INVx1_ASAP7_75t_L         g15466(.A(new_n15387), .Y(new_n15723));
  O2A1O1Ixp33_ASAP7_75t_L   g15467(.A1(new_n15723), .A2(new_n15562), .B(new_n15561), .C(new_n15637), .Y(new_n15724));
  NAND2xp33_ASAP7_75t_L     g15468(.A(new_n15724), .B(new_n15722), .Y(new_n15725));
  AND2x2_ASAP7_75t_L        g15469(.A(new_n15721), .B(new_n15725), .Y(new_n15726));
  AOI22xp33_ASAP7_75t_L     g15470(.A1(new_n3633), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n3858), .Y(new_n15727));
  OAI221xp5_ASAP7_75t_L     g15471(.A1(new_n3853), .A2(new_n7593), .B1(new_n3856), .B2(new_n7623), .C(new_n15727), .Y(new_n15728));
  XNOR2x2_ASAP7_75t_L       g15472(.A(\a[35] ), .B(new_n15728), .Y(new_n15729));
  INVx1_ASAP7_75t_L         g15473(.A(new_n15729), .Y(new_n15730));
  NAND2xp33_ASAP7_75t_L     g15474(.A(new_n15730), .B(new_n15726), .Y(new_n15731));
  AO21x2_ASAP7_75t_L        g15475(.A1(new_n15721), .A2(new_n15725), .B(new_n15730), .Y(new_n15732));
  AND2x2_ASAP7_75t_L        g15476(.A(new_n15732), .B(new_n15731), .Y(new_n15733));
  INVx1_ASAP7_75t_L         g15477(.A(new_n15733), .Y(new_n15734));
  NAND2xp33_ASAP7_75t_L     g15478(.A(new_n15635), .B(new_n15734), .Y(new_n15735));
  INVx1_ASAP7_75t_L         g15479(.A(new_n15569), .Y(new_n15736));
  A2O1A1Ixp33_ASAP7_75t_L   g15480(.A1(new_n15736), .A2(new_n15568), .B(new_n15576), .C(new_n15733), .Y(new_n15737));
  NAND2xp33_ASAP7_75t_L     g15481(.A(new_n15737), .B(new_n15735), .Y(new_n15738));
  NOR2xp33_ASAP7_75t_L      g15482(.A(new_n15738), .B(new_n15632), .Y(new_n15739));
  AND2x2_ASAP7_75t_L        g15483(.A(new_n15738), .B(new_n15632), .Y(new_n15740));
  NOR2xp33_ASAP7_75t_L      g15484(.A(new_n15739), .B(new_n15740), .Y(new_n15741));
  XNOR2x2_ASAP7_75t_L       g15485(.A(new_n15625), .B(new_n15741), .Y(new_n15742));
  NOR2xp33_ASAP7_75t_L      g15486(.A(new_n15742), .B(new_n15619), .Y(new_n15743));
  AND2x2_ASAP7_75t_L        g15487(.A(new_n15742), .B(new_n15619), .Y(new_n15744));
  NOR2xp33_ASAP7_75t_L      g15488(.A(new_n15743), .B(new_n15744), .Y(new_n15745));
  NAND2xp33_ASAP7_75t_L     g15489(.A(new_n15745), .B(new_n15612), .Y(new_n15746));
  OAI21xp33_ASAP7_75t_L     g15490(.A1(new_n15743), .A2(new_n15744), .B(new_n15611), .Y(new_n15747));
  NAND2xp33_ASAP7_75t_L     g15491(.A(new_n15747), .B(new_n15746), .Y(new_n15748));
  NAND3xp33_ASAP7_75t_L     g15492(.A(new_n15748), .B(new_n15586), .C(new_n15450), .Y(new_n15749));
  INVx1_ASAP7_75t_L         g15493(.A(new_n15449), .Y(new_n15750));
  O2A1O1Ixp33_ASAP7_75t_L   g15494(.A1(new_n15446), .A2(new_n15750), .B(new_n15586), .C(new_n15748), .Y(new_n15751));
  INVx1_ASAP7_75t_L         g15495(.A(new_n15751), .Y(new_n15752));
  NAND2xp33_ASAP7_75t_L     g15496(.A(new_n15749), .B(new_n15752), .Y(new_n15753));
  INVx1_ASAP7_75t_L         g15497(.A(new_n15753), .Y(new_n15754));
  A2O1A1Ixp33_ASAP7_75t_L   g15498(.A1(new_n15598), .A2(new_n15594), .B(new_n15590), .C(new_n15754), .Y(new_n15755));
  INVx1_ASAP7_75t_L         g15499(.A(new_n15755), .Y(new_n15756));
  A2O1A1Ixp33_ASAP7_75t_L   g15500(.A1(new_n15434), .A2(new_n15597), .B(new_n15593), .C(new_n15591), .Y(new_n15757));
  NOR2xp33_ASAP7_75t_L      g15501(.A(new_n15754), .B(new_n15757), .Y(new_n15758));
  NOR2xp33_ASAP7_75t_L      g15502(.A(new_n15758), .B(new_n15756), .Y(\f[84] ));
  AOI22xp33_ASAP7_75t_L     g15503(.A1(new_n1837), .A2(\b[62] ), .B1(new_n1695), .B2(new_n12322), .Y(new_n15760));
  OA211x2_ASAP7_75t_L       g15504(.A1(new_n1699), .A2(new_n11468), .B(new_n15760), .C(\a[23] ), .Y(new_n15761));
  O2A1O1Ixp33_ASAP7_75t_L   g15505(.A1(new_n11468), .A2(new_n1699), .B(new_n15760), .C(\a[23] ), .Y(new_n15762));
  OAI22xp33_ASAP7_75t_L     g15506(.A1(new_n15743), .A2(new_n15618), .B1(new_n15762), .B2(new_n15761), .Y(new_n15763));
  OR4x2_ASAP7_75t_L         g15507(.A(new_n15762), .B(new_n15743), .C(new_n15761), .D(new_n15618), .Y(new_n15764));
  NAND2xp33_ASAP7_75t_L     g15508(.A(new_n15763), .B(new_n15764), .Y(new_n15765));
  AOI22xp33_ASAP7_75t_L     g15509(.A1(new_n2114), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n2259), .Y(new_n15766));
  OAI221xp5_ASAP7_75t_L     g15510(.A1(new_n2109), .A2(new_n10250), .B1(new_n2257), .B2(new_n10855), .C(new_n15766), .Y(new_n15767));
  XNOR2x2_ASAP7_75t_L       g15511(.A(\a[26] ), .B(new_n15767), .Y(new_n15768));
  INVx1_ASAP7_75t_L         g15512(.A(new_n15624), .Y(new_n15769));
  MAJIxp5_ASAP7_75t_L       g15513(.A(new_n15741), .B(new_n15621), .C(new_n15769), .Y(new_n15770));
  NAND2xp33_ASAP7_75t_L     g15514(.A(new_n15768), .B(new_n15770), .Y(new_n15771));
  NOR2xp33_ASAP7_75t_L      g15515(.A(new_n15768), .B(new_n15770), .Y(new_n15772));
  INVx1_ASAP7_75t_L         g15516(.A(new_n15772), .Y(new_n15773));
  NOR2xp33_ASAP7_75t_L      g15517(.A(new_n15628), .B(new_n15631), .Y(new_n15774));
  NOR2xp33_ASAP7_75t_L      g15518(.A(new_n15774), .B(new_n15739), .Y(new_n15775));
  AOI22xp33_ASAP7_75t_L     g15519(.A1(new_n2552), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n2736), .Y(new_n15776));
  OAI221xp5_ASAP7_75t_L     g15520(.A1(new_n2547), .A2(new_n9620), .B1(new_n2734), .B2(new_n9925), .C(new_n15776), .Y(new_n15777));
  XNOR2x2_ASAP7_75t_L       g15521(.A(\a[29] ), .B(new_n15777), .Y(new_n15778));
  XNOR2x2_ASAP7_75t_L       g15522(.A(new_n15778), .B(new_n15775), .Y(new_n15779));
  AOI22xp33_ASAP7_75t_L     g15523(.A1(new_n3029), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n3258), .Y(new_n15780));
  OAI221xp5_ASAP7_75t_L     g15524(.A1(new_n3024), .A2(new_n8458), .B1(new_n3256), .B2(new_n8768), .C(new_n15780), .Y(new_n15781));
  XNOR2x2_ASAP7_75t_L       g15525(.A(\a[32] ), .B(new_n15781), .Y(new_n15782));
  INVx1_ASAP7_75t_L         g15526(.A(new_n15782), .Y(new_n15783));
  O2A1O1Ixp33_ASAP7_75t_L   g15527(.A1(new_n15635), .A2(new_n15734), .B(new_n15731), .C(new_n15783), .Y(new_n15784));
  INVx1_ASAP7_75t_L         g15528(.A(new_n15784), .Y(new_n15785));
  NAND3xp33_ASAP7_75t_L     g15529(.A(new_n15737), .B(new_n15731), .C(new_n15783), .Y(new_n15786));
  NOR2xp33_ASAP7_75t_L      g15530(.A(new_n15694), .B(new_n15691), .Y(new_n15787));
  A2O1A1O1Ixp25_ASAP7_75t_L g15531(.A1(new_n15490), .A2(new_n15551), .B(new_n15548), .C(new_n15697), .D(new_n15787), .Y(new_n15788));
  AOI22xp33_ASAP7_75t_L     g15532(.A1(new_n6376), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n6648), .Y(new_n15789));
  OAI221xp5_ASAP7_75t_L     g15533(.A1(new_n6646), .A2(new_n4848), .B1(new_n6636), .B2(new_n11686), .C(new_n15789), .Y(new_n15790));
  XNOR2x2_ASAP7_75t_L       g15534(.A(\a[47] ), .B(new_n15790), .Y(new_n15791));
  INVx1_ASAP7_75t_L         g15535(.A(new_n15791), .Y(new_n15792));
  INVx1_ASAP7_75t_L         g15536(.A(new_n15676), .Y(new_n15793));
  NAND2xp33_ASAP7_75t_L     g15537(.A(new_n15793), .B(new_n15682), .Y(new_n15794));
  AOI22xp33_ASAP7_75t_L     g15538(.A1(new_n9700), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n10027), .Y(new_n15795));
  OAI221xp5_ASAP7_75t_L     g15539(.A1(new_n10024), .A2(new_n2497), .B1(new_n9696), .B2(new_n2672), .C(new_n15795), .Y(new_n15796));
  XNOR2x2_ASAP7_75t_L       g15540(.A(\a[59] ), .B(new_n15796), .Y(new_n15797));
  A2O1A1Ixp33_ASAP7_75t_L   g15541(.A1(new_n15503), .A2(new_n15318), .B(new_n15513), .C(new_n15657), .Y(new_n15798));
  NOR2xp33_ASAP7_75t_L      g15542(.A(new_n1655), .B(new_n11535), .Y(new_n15799));
  A2O1A1O1Ixp25_ASAP7_75t_L g15543(.A1(new_n11533), .A2(\b[20] ), .B(new_n15502), .C(new_n15647), .D(new_n15645), .Y(new_n15800));
  A2O1A1Ixp33_ASAP7_75t_L   g15544(.A1(new_n11533), .A2(\b[22] ), .B(new_n15799), .C(new_n15800), .Y(new_n15801));
  O2A1O1Ixp33_ASAP7_75t_L   g15545(.A1(new_n11247), .A2(new_n11249), .B(\b[22] ), .C(new_n15799), .Y(new_n15802));
  INVx1_ASAP7_75t_L         g15546(.A(new_n15802), .Y(new_n15803));
  O2A1O1Ixp33_ASAP7_75t_L   g15547(.A1(new_n15503), .A2(new_n15648), .B(new_n15644), .C(new_n15803), .Y(new_n15804));
  INVx1_ASAP7_75t_L         g15548(.A(new_n15804), .Y(new_n15805));
  NAND2xp33_ASAP7_75t_L     g15549(.A(new_n15801), .B(new_n15805), .Y(new_n15806));
  NOR2xp33_ASAP7_75t_L      g15550(.A(new_n2067), .B(new_n10630), .Y(new_n15807));
  AOI221xp5_ASAP7_75t_L     g15551(.A1(\b[23] ), .A2(new_n10939), .B1(\b[24] ), .B2(new_n10632), .C(new_n15807), .Y(new_n15808));
  OAI211xp5_ASAP7_75t_L     g15552(.A1(new_n10629), .A2(new_n2075), .B(\a[62] ), .C(new_n15808), .Y(new_n15809));
  O2A1O1Ixp33_ASAP7_75t_L   g15553(.A1(new_n10629), .A2(new_n2075), .B(new_n15808), .C(\a[62] ), .Y(new_n15810));
  INVx1_ASAP7_75t_L         g15554(.A(new_n15810), .Y(new_n15811));
  AND2x2_ASAP7_75t_L        g15555(.A(new_n15809), .B(new_n15811), .Y(new_n15812));
  NOR2xp33_ASAP7_75t_L      g15556(.A(new_n15806), .B(new_n15812), .Y(new_n15813));
  INVx1_ASAP7_75t_L         g15557(.A(new_n15813), .Y(new_n15814));
  NAND2xp33_ASAP7_75t_L     g15558(.A(new_n15806), .B(new_n15812), .Y(new_n15815));
  AND2x2_ASAP7_75t_L        g15559(.A(new_n15815), .B(new_n15814), .Y(new_n15816));
  INVx1_ASAP7_75t_L         g15560(.A(new_n15816), .Y(new_n15817));
  O2A1O1Ixp33_ASAP7_75t_L   g15561(.A1(new_n15651), .A2(new_n15654), .B(new_n15798), .C(new_n15817), .Y(new_n15818));
  NOR2xp33_ASAP7_75t_L      g15562(.A(new_n15651), .B(new_n15654), .Y(new_n15819));
  NOR3xp33_ASAP7_75t_L      g15563(.A(new_n15816), .B(new_n15819), .C(new_n15656), .Y(new_n15820));
  OR3x1_ASAP7_75t_L         g15564(.A(new_n15818), .B(new_n15797), .C(new_n15820), .Y(new_n15821));
  OAI21xp33_ASAP7_75t_L     g15565(.A1(new_n15820), .A2(new_n15818), .B(new_n15797), .Y(new_n15822));
  AND2x2_ASAP7_75t_L        g15566(.A(new_n15822), .B(new_n15821), .Y(new_n15823));
  A2O1A1Ixp33_ASAP7_75t_L   g15567(.A1(new_n15661), .A2(new_n15642), .B(new_n15666), .C(new_n15823), .Y(new_n15824));
  NAND2xp33_ASAP7_75t_L     g15568(.A(new_n15642), .B(new_n15661), .Y(new_n15825));
  A2O1A1Ixp33_ASAP7_75t_L   g15569(.A1(new_n15521), .A2(new_n15518), .B(new_n15662), .C(new_n15825), .Y(new_n15826));
  NOR2xp33_ASAP7_75t_L      g15570(.A(new_n15826), .B(new_n15823), .Y(new_n15827));
  INVx1_ASAP7_75t_L         g15571(.A(new_n15827), .Y(new_n15828));
  AOI22xp33_ASAP7_75t_L     g15572(.A1(new_n8831), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n9115), .Y(new_n15829));
  OAI221xp5_ASAP7_75t_L     g15573(.A1(new_n10343), .A2(new_n2982), .B1(new_n10016), .B2(new_n3187), .C(new_n15829), .Y(new_n15830));
  XNOR2x2_ASAP7_75t_L       g15574(.A(\a[56] ), .B(new_n15830), .Y(new_n15831));
  NAND3xp33_ASAP7_75t_L     g15575(.A(new_n15828), .B(new_n15824), .C(new_n15831), .Y(new_n15832));
  INVx1_ASAP7_75t_L         g15576(.A(new_n15832), .Y(new_n15833));
  AOI21xp33_ASAP7_75t_L     g15577(.A1(new_n15828), .A2(new_n15824), .B(new_n15831), .Y(new_n15834));
  NOR2xp33_ASAP7_75t_L      g15578(.A(new_n15834), .B(new_n15833), .Y(new_n15835));
  NAND2xp33_ASAP7_75t_L     g15579(.A(new_n15671), .B(new_n15667), .Y(new_n15836));
  AND2x2_ASAP7_75t_L        g15580(.A(new_n15836), .B(new_n15675), .Y(new_n15837));
  NAND2xp33_ASAP7_75t_L     g15581(.A(new_n15835), .B(new_n15837), .Y(new_n15838));
  INVx1_ASAP7_75t_L         g15582(.A(new_n15838), .Y(new_n15839));
  O2A1O1Ixp33_ASAP7_75t_L   g15583(.A1(new_n15674), .A2(new_n15672), .B(new_n15836), .C(new_n15835), .Y(new_n15840));
  NOR2xp33_ASAP7_75t_L      g15584(.A(new_n15840), .B(new_n15839), .Y(new_n15841));
  AOI22xp33_ASAP7_75t_L     g15585(.A1(new_n7960), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n8537), .Y(new_n15842));
  OAI221xp5_ASAP7_75t_L     g15586(.A1(new_n8817), .A2(new_n3565), .B1(new_n7957), .B2(new_n3591), .C(new_n15842), .Y(new_n15843));
  XNOR2x2_ASAP7_75t_L       g15587(.A(\a[53] ), .B(new_n15843), .Y(new_n15844));
  NAND2xp33_ASAP7_75t_L     g15588(.A(new_n15844), .B(new_n15841), .Y(new_n15845));
  INVx1_ASAP7_75t_L         g15589(.A(new_n15845), .Y(new_n15846));
  NOR2xp33_ASAP7_75t_L      g15590(.A(new_n15844), .B(new_n15841), .Y(new_n15847));
  NOR2xp33_ASAP7_75t_L      g15591(.A(new_n15847), .B(new_n15846), .Y(new_n15848));
  INVx1_ASAP7_75t_L         g15592(.A(new_n15848), .Y(new_n15849));
  A2O1A1O1Ixp25_ASAP7_75t_L g15593(.A1(new_n15535), .A2(new_n15534), .B(new_n15680), .C(new_n15794), .D(new_n15849), .Y(new_n15850));
  A2O1A1Ixp33_ASAP7_75t_L   g15594(.A1(new_n15535), .A2(new_n15534), .B(new_n15680), .C(new_n15794), .Y(new_n15851));
  NOR2xp33_ASAP7_75t_L      g15595(.A(new_n15851), .B(new_n15848), .Y(new_n15852));
  NOR2xp33_ASAP7_75t_L      g15596(.A(new_n15852), .B(new_n15850), .Y(new_n15853));
  INVx1_ASAP7_75t_L         g15597(.A(new_n15853), .Y(new_n15854));
  AOI22xp33_ASAP7_75t_L     g15598(.A1(new_n7111), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n7391), .Y(new_n15855));
  OAI221xp5_ASAP7_75t_L     g15599(.A1(new_n8558), .A2(new_n4216), .B1(new_n8237), .B2(new_n4431), .C(new_n15855), .Y(new_n15856));
  XNOR2x2_ASAP7_75t_L       g15600(.A(\a[50] ), .B(new_n15856), .Y(new_n15857));
  NAND2xp33_ASAP7_75t_L     g15601(.A(new_n15857), .B(new_n15854), .Y(new_n15858));
  NOR2xp33_ASAP7_75t_L      g15602(.A(new_n15857), .B(new_n15854), .Y(new_n15859));
  INVx1_ASAP7_75t_L         g15603(.A(new_n15859), .Y(new_n15860));
  AND2x2_ASAP7_75t_L        g15604(.A(new_n15858), .B(new_n15860), .Y(new_n15861));
  A2O1A1Ixp33_ASAP7_75t_L   g15605(.A1(new_n15689), .A2(new_n15638), .B(new_n15687), .C(new_n15861), .Y(new_n15862));
  A2O1A1O1Ixp25_ASAP7_75t_L g15606(.A1(new_n15494), .A2(new_n15542), .B(new_n15539), .C(new_n15689), .D(new_n15687), .Y(new_n15863));
  INVx1_ASAP7_75t_L         g15607(.A(new_n15861), .Y(new_n15864));
  NAND2xp33_ASAP7_75t_L     g15608(.A(new_n15863), .B(new_n15864), .Y(new_n15865));
  AND2x2_ASAP7_75t_L        g15609(.A(new_n15862), .B(new_n15865), .Y(new_n15866));
  NAND2xp33_ASAP7_75t_L     g15610(.A(new_n15792), .B(new_n15866), .Y(new_n15867));
  INVx1_ASAP7_75t_L         g15611(.A(new_n15867), .Y(new_n15868));
  NOR2xp33_ASAP7_75t_L      g15612(.A(new_n15792), .B(new_n15866), .Y(new_n15869));
  OR3x1_ASAP7_75t_L         g15613(.A(new_n15868), .B(new_n15788), .C(new_n15869), .Y(new_n15870));
  OAI21xp33_ASAP7_75t_L     g15614(.A1(new_n15869), .A2(new_n15868), .B(new_n15788), .Y(new_n15871));
  NAND2xp33_ASAP7_75t_L     g15615(.A(new_n15871), .B(new_n15870), .Y(new_n15872));
  AOI22xp33_ASAP7_75t_L     g15616(.A1(new_n5624), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n5901), .Y(new_n15873));
  OAI221xp5_ASAP7_75t_L     g15617(.A1(new_n5900), .A2(new_n5338), .B1(new_n5892), .B2(new_n6338), .C(new_n15873), .Y(new_n15874));
  XNOR2x2_ASAP7_75t_L       g15618(.A(new_n5619), .B(new_n15874), .Y(new_n15875));
  NOR2xp33_ASAP7_75t_L      g15619(.A(new_n15875), .B(new_n15872), .Y(new_n15876));
  AND2x2_ASAP7_75t_L        g15620(.A(new_n15875), .B(new_n15872), .Y(new_n15877));
  NOR2xp33_ASAP7_75t_L      g15621(.A(new_n15876), .B(new_n15877), .Y(new_n15878));
  OA21x2_ASAP7_75t_L        g15622(.A1(new_n15699), .A2(new_n15702), .B(new_n15708), .Y(new_n15879));
  NAND2xp33_ASAP7_75t_L     g15623(.A(new_n15879), .B(new_n15878), .Y(new_n15880));
  XNOR2x2_ASAP7_75t_L       g15624(.A(new_n15875), .B(new_n15872), .Y(new_n15881));
  INVx1_ASAP7_75t_L         g15625(.A(new_n15879), .Y(new_n15882));
  NAND2xp33_ASAP7_75t_L     g15626(.A(new_n15882), .B(new_n15881), .Y(new_n15883));
  AOI22xp33_ASAP7_75t_L     g15627(.A1(new_n4920), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n5167), .Y(new_n15884));
  OAI221xp5_ASAP7_75t_L     g15628(.A1(new_n5154), .A2(new_n6321), .B1(new_n5158), .B2(new_n6573), .C(new_n15884), .Y(new_n15885));
  XNOR2x2_ASAP7_75t_L       g15629(.A(\a[41] ), .B(new_n15885), .Y(new_n15886));
  NAND3xp33_ASAP7_75t_L     g15630(.A(new_n15880), .B(new_n15883), .C(new_n15886), .Y(new_n15887));
  INVx1_ASAP7_75t_L         g15631(.A(new_n15887), .Y(new_n15888));
  AOI21xp33_ASAP7_75t_L     g15632(.A1(new_n15880), .A2(new_n15883), .B(new_n15886), .Y(new_n15889));
  A2O1A1Ixp33_ASAP7_75t_L   g15633(.A1(new_n15560), .A2(new_n15479), .B(new_n15714), .C(new_n15713), .Y(new_n15890));
  OAI21xp33_ASAP7_75t_L     g15634(.A1(new_n15709), .A2(new_n15712), .B(new_n15890), .Y(new_n15891));
  OR3x1_ASAP7_75t_L         g15635(.A(new_n15888), .B(new_n15889), .C(new_n15891), .Y(new_n15892));
  OAI21xp33_ASAP7_75t_L     g15636(.A1(new_n15889), .A2(new_n15888), .B(new_n15891), .Y(new_n15893));
  AOI22xp33_ASAP7_75t_L     g15637(.A1(new_n4283), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n4512), .Y(new_n15894));
  OAI221xp5_ASAP7_75t_L     g15638(.A1(new_n4277), .A2(new_n6830), .B1(new_n4499), .B2(new_n7323), .C(new_n15894), .Y(new_n15895));
  XNOR2x2_ASAP7_75t_L       g15639(.A(\a[38] ), .B(new_n15895), .Y(new_n15896));
  NAND3xp33_ASAP7_75t_L     g15640(.A(new_n15892), .B(new_n15893), .C(new_n15896), .Y(new_n15897));
  AO21x2_ASAP7_75t_L        g15641(.A1(new_n15893), .A2(new_n15892), .B(new_n15896), .Y(new_n15898));
  NAND2xp33_ASAP7_75t_L     g15642(.A(new_n15897), .B(new_n15898), .Y(new_n15899));
  OAI21xp33_ASAP7_75t_L     g15643(.A1(new_n15716), .A2(new_n15719), .B(new_n15725), .Y(new_n15900));
  XNOR2x2_ASAP7_75t_L       g15644(.A(new_n15900), .B(new_n15899), .Y(new_n15901));
  AOI22xp33_ASAP7_75t_L     g15645(.A1(new_n3633), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n3858), .Y(new_n15902));
  OAI221xp5_ASAP7_75t_L     g15646(.A1(new_n3853), .A2(new_n7616), .B1(new_n3856), .B2(new_n7906), .C(new_n15902), .Y(new_n15903));
  XNOR2x2_ASAP7_75t_L       g15647(.A(\a[35] ), .B(new_n15903), .Y(new_n15904));
  XNOR2x2_ASAP7_75t_L       g15648(.A(new_n15904), .B(new_n15901), .Y(new_n15905));
  AO21x2_ASAP7_75t_L        g15649(.A1(new_n15785), .A2(new_n15786), .B(new_n15905), .Y(new_n15906));
  NAND3xp33_ASAP7_75t_L     g15650(.A(new_n15905), .B(new_n15786), .C(new_n15785), .Y(new_n15907));
  NAND2xp33_ASAP7_75t_L     g15651(.A(new_n15907), .B(new_n15906), .Y(new_n15908));
  XOR2x2_ASAP7_75t_L        g15652(.A(new_n15908), .B(new_n15779), .Y(new_n15909));
  NAND3xp33_ASAP7_75t_L     g15653(.A(new_n15909), .B(new_n15773), .C(new_n15771), .Y(new_n15910));
  NAND2xp33_ASAP7_75t_L     g15654(.A(new_n15771), .B(new_n15773), .Y(new_n15911));
  INVx1_ASAP7_75t_L         g15655(.A(new_n15909), .Y(new_n15912));
  NAND2xp33_ASAP7_75t_L     g15656(.A(new_n15911), .B(new_n15912), .Y(new_n15913));
  NAND2xp33_ASAP7_75t_L     g15657(.A(new_n15910), .B(new_n15913), .Y(new_n15914));
  INVx1_ASAP7_75t_L         g15658(.A(new_n15914), .Y(new_n15915));
  NOR2xp33_ASAP7_75t_L      g15659(.A(new_n15765), .B(new_n15915), .Y(new_n15916));
  INVx1_ASAP7_75t_L         g15660(.A(new_n15916), .Y(new_n15917));
  NAND2xp33_ASAP7_75t_L     g15661(.A(new_n15765), .B(new_n15915), .Y(new_n15918));
  NAND2xp33_ASAP7_75t_L     g15662(.A(new_n15918), .B(new_n15917), .Y(new_n15919));
  O2A1O1Ixp33_ASAP7_75t_L   g15663(.A1(new_n15454), .A2(new_n15457), .B(new_n15582), .C(new_n15606), .Y(new_n15920));
  AOI211xp5_ASAP7_75t_L     g15664(.A1(new_n15745), .A2(new_n15612), .B(new_n15920), .C(new_n15919), .Y(new_n15921));
  A2O1A1Ixp33_ASAP7_75t_L   g15665(.A1(new_n15612), .A2(new_n15745), .B(new_n15920), .C(new_n15919), .Y(new_n15922));
  INVx1_ASAP7_75t_L         g15666(.A(new_n15922), .Y(new_n15923));
  NOR2xp33_ASAP7_75t_L      g15667(.A(new_n15921), .B(new_n15923), .Y(new_n15924));
  A2O1A1Ixp33_ASAP7_75t_L   g15668(.A1(new_n15757), .A2(new_n15754), .B(new_n15751), .C(new_n15924), .Y(new_n15925));
  INVx1_ASAP7_75t_L         g15669(.A(new_n15925), .Y(new_n15926));
  A2O1A1Ixp33_ASAP7_75t_L   g15670(.A1(new_n15595), .A2(new_n15591), .B(new_n15753), .C(new_n15752), .Y(new_n15927));
  NOR2xp33_ASAP7_75t_L      g15671(.A(new_n15924), .B(new_n15927), .Y(new_n15928));
  NOR2xp33_ASAP7_75t_L      g15672(.A(new_n15928), .B(new_n15926), .Y(\f[85] ));
  A2O1A1Ixp33_ASAP7_75t_L   g15673(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n1695), .Y(new_n15930));
  A2O1A1Ixp33_ASAP7_75t_L   g15674(.A1(new_n15930), .A2(new_n1829), .B(new_n11468), .C(\a[23] ), .Y(new_n15931));
  O2A1O1Ixp33_ASAP7_75t_L   g15675(.A1(new_n1827), .A2(new_n12060), .B(new_n1829), .C(new_n11468), .Y(new_n15932));
  NAND2xp33_ASAP7_75t_L     g15676(.A(new_n1689), .B(new_n15932), .Y(new_n15933));
  AND2x2_ASAP7_75t_L        g15677(.A(new_n15933), .B(new_n15931), .Y(new_n15934));
  O2A1O1Ixp33_ASAP7_75t_L   g15678(.A1(new_n15911), .A2(new_n15912), .B(new_n15773), .C(new_n15934), .Y(new_n15935));
  INVx1_ASAP7_75t_L         g15679(.A(new_n15935), .Y(new_n15936));
  NAND3xp33_ASAP7_75t_L     g15680(.A(new_n15910), .B(new_n15773), .C(new_n15934), .Y(new_n15937));
  AOI22xp33_ASAP7_75t_L     g15681(.A1(new_n2114), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n2259), .Y(new_n15938));
  OAI221xp5_ASAP7_75t_L     g15682(.A1(new_n2109), .A2(new_n10847), .B1(new_n2257), .B2(new_n12047), .C(new_n15938), .Y(new_n15939));
  XNOR2x2_ASAP7_75t_L       g15683(.A(\a[26] ), .B(new_n15939), .Y(new_n15940));
  INVx1_ASAP7_75t_L         g15684(.A(new_n15778), .Y(new_n15941));
  NOR2xp33_ASAP7_75t_L      g15685(.A(new_n15908), .B(new_n15779), .Y(new_n15942));
  O2A1O1Ixp33_ASAP7_75t_L   g15686(.A1(new_n15774), .A2(new_n15739), .B(new_n15941), .C(new_n15942), .Y(new_n15943));
  NAND2xp33_ASAP7_75t_L     g15687(.A(new_n15940), .B(new_n15943), .Y(new_n15944));
  OR2x4_ASAP7_75t_L         g15688(.A(new_n15940), .B(new_n15943), .Y(new_n15945));
  NAND2xp33_ASAP7_75t_L     g15689(.A(new_n15944), .B(new_n15945), .Y(new_n15946));
  AOI22xp33_ASAP7_75t_L     g15690(.A1(new_n2552), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n2736), .Y(new_n15947));
  OAI221xp5_ASAP7_75t_L     g15691(.A1(new_n2547), .A2(new_n9920), .B1(new_n2734), .B2(new_n11152), .C(new_n15947), .Y(new_n15948));
  XNOR2x2_ASAP7_75t_L       g15692(.A(\a[29] ), .B(new_n15948), .Y(new_n15949));
  INVx1_ASAP7_75t_L         g15693(.A(new_n15731), .Y(new_n15950));
  A2O1A1Ixp33_ASAP7_75t_L   g15694(.A1(new_n15732), .A2(new_n15634), .B(new_n15950), .C(new_n15783), .Y(new_n15951));
  A2O1A1Ixp33_ASAP7_75t_L   g15695(.A1(new_n15786), .A2(new_n15785), .B(new_n15905), .C(new_n15951), .Y(new_n15952));
  XOR2x2_ASAP7_75t_L        g15696(.A(new_n15949), .B(new_n15952), .Y(new_n15953));
  AOI22xp33_ASAP7_75t_L     g15697(.A1(new_n3029), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n3258), .Y(new_n15954));
  OAI221xp5_ASAP7_75t_L     g15698(.A1(new_n3024), .A2(new_n8762), .B1(new_n3256), .B2(new_n9331), .C(new_n15954), .Y(new_n15955));
  XNOR2x2_ASAP7_75t_L       g15699(.A(new_n3015), .B(new_n15955), .Y(new_n15956));
  INVx1_ASAP7_75t_L         g15700(.A(new_n15904), .Y(new_n15957));
  MAJx2_ASAP7_75t_L         g15701(.A(new_n15899), .B(new_n15900), .C(new_n15957), .Y(new_n15958));
  NOR2xp33_ASAP7_75t_L      g15702(.A(new_n15956), .B(new_n15958), .Y(new_n15959));
  AND2x2_ASAP7_75t_L        g15703(.A(new_n15956), .B(new_n15958), .Y(new_n15960));
  NOR2xp33_ASAP7_75t_L      g15704(.A(new_n15959), .B(new_n15960), .Y(new_n15961));
  AOI22xp33_ASAP7_75t_L     g15705(.A1(new_n3633), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n3858), .Y(new_n15962));
  OAI221xp5_ASAP7_75t_L     g15706(.A1(new_n3853), .A2(new_n7900), .B1(new_n3856), .B2(new_n8174), .C(new_n15962), .Y(new_n15963));
  XNOR2x2_ASAP7_75t_L       g15707(.A(\a[35] ), .B(new_n15963), .Y(new_n15964));
  AOI22xp33_ASAP7_75t_L     g15708(.A1(new_n5624), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n5901), .Y(new_n15965));
  OAI221xp5_ASAP7_75t_L     g15709(.A1(new_n5900), .A2(new_n5805), .B1(new_n5892), .B2(new_n5835), .C(new_n15965), .Y(new_n15966));
  XNOR2x2_ASAP7_75t_L       g15710(.A(\a[44] ), .B(new_n15966), .Y(new_n15967));
  INVx1_ASAP7_75t_L         g15711(.A(new_n15967), .Y(new_n15968));
  AOI22xp33_ASAP7_75t_L     g15712(.A1(new_n6376), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n6648), .Y(new_n15969));
  OAI221xp5_ASAP7_75t_L     g15713(.A1(new_n6646), .A2(new_n4869), .B1(new_n6636), .B2(new_n5327), .C(new_n15969), .Y(new_n15970));
  XNOR2x2_ASAP7_75t_L       g15714(.A(\a[47] ), .B(new_n15970), .Y(new_n15971));
  AOI22xp33_ASAP7_75t_L     g15715(.A1(new_n7960), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n8537), .Y(new_n15972));
  OAI221xp5_ASAP7_75t_L     g15716(.A1(new_n8817), .A2(new_n3584), .B1(new_n7957), .B2(new_n10137), .C(new_n15972), .Y(new_n15973));
  XNOR2x2_ASAP7_75t_L       g15717(.A(\a[53] ), .B(new_n15973), .Y(new_n15974));
  INVx1_ASAP7_75t_L         g15718(.A(new_n15974), .Y(new_n15975));
  INVx1_ASAP7_75t_L         g15719(.A(new_n15812), .Y(new_n15976));
  NOR2xp33_ASAP7_75t_L      g15720(.A(new_n1774), .B(new_n11535), .Y(new_n15977));
  O2A1O1Ixp33_ASAP7_75t_L   g15721(.A1(new_n11247), .A2(new_n11249), .B(\b[23] ), .C(new_n15977), .Y(new_n15978));
  A2O1A1Ixp33_ASAP7_75t_L   g15722(.A1(new_n11533), .A2(\b[22] ), .B(new_n15799), .C(new_n15978), .Y(new_n15979));
  A2O1A1Ixp33_ASAP7_75t_L   g15723(.A1(\b[23] ), .A2(new_n11533), .B(new_n15977), .C(new_n15802), .Y(new_n15980));
  NAND2xp33_ASAP7_75t_L     g15724(.A(new_n15980), .B(new_n15979), .Y(new_n15981));
  NOR2xp33_ASAP7_75t_L      g15725(.A(new_n2348), .B(new_n10630), .Y(new_n15982));
  AOI221xp5_ASAP7_75t_L     g15726(.A1(\b[24] ), .A2(new_n10939), .B1(\b[25] ), .B2(new_n10632), .C(new_n15982), .Y(new_n15983));
  OAI211xp5_ASAP7_75t_L     g15727(.A1(new_n10629), .A2(new_n2355), .B(\a[62] ), .C(new_n15983), .Y(new_n15984));
  INVx1_ASAP7_75t_L         g15728(.A(new_n15984), .Y(new_n15985));
  O2A1O1Ixp33_ASAP7_75t_L   g15729(.A1(new_n10629), .A2(new_n2355), .B(new_n15983), .C(\a[62] ), .Y(new_n15986));
  NOR2xp33_ASAP7_75t_L      g15730(.A(new_n15986), .B(new_n15985), .Y(new_n15987));
  NOR2xp33_ASAP7_75t_L      g15731(.A(new_n15981), .B(new_n15987), .Y(new_n15988));
  INVx1_ASAP7_75t_L         g15732(.A(new_n15988), .Y(new_n15989));
  NAND2xp33_ASAP7_75t_L     g15733(.A(new_n15981), .B(new_n15987), .Y(new_n15990));
  AND2x2_ASAP7_75t_L        g15734(.A(new_n15990), .B(new_n15989), .Y(new_n15991));
  A2O1A1Ixp33_ASAP7_75t_L   g15735(.A1(new_n15976), .A2(new_n15801), .B(new_n15804), .C(new_n15991), .Y(new_n15992));
  A2O1A1Ixp33_ASAP7_75t_L   g15736(.A1(new_n15811), .A2(new_n15809), .B(new_n15806), .C(new_n15805), .Y(new_n15993));
  NOR2xp33_ASAP7_75t_L      g15737(.A(new_n15993), .B(new_n15991), .Y(new_n15994));
  INVx1_ASAP7_75t_L         g15738(.A(new_n15994), .Y(new_n15995));
  AOI22xp33_ASAP7_75t_L     g15739(.A1(new_n9700), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n10027), .Y(new_n15996));
  OAI221xp5_ASAP7_75t_L     g15740(.A1(new_n10024), .A2(new_n2666), .B1(new_n9696), .B2(new_n2695), .C(new_n15996), .Y(new_n15997));
  XNOR2x2_ASAP7_75t_L       g15741(.A(\a[59] ), .B(new_n15997), .Y(new_n15998));
  NAND3xp33_ASAP7_75t_L     g15742(.A(new_n15995), .B(new_n15992), .C(new_n15998), .Y(new_n15999));
  INVx1_ASAP7_75t_L         g15743(.A(new_n15999), .Y(new_n16000));
  AOI21xp33_ASAP7_75t_L     g15744(.A1(new_n15995), .A2(new_n15992), .B(new_n15998), .Y(new_n16001));
  A2O1A1Ixp33_ASAP7_75t_L   g15745(.A1(new_n15659), .A2(new_n15657), .B(new_n15819), .C(new_n15816), .Y(new_n16002));
  NAND2xp33_ASAP7_75t_L     g15746(.A(new_n16002), .B(new_n15821), .Y(new_n16003));
  NOR3xp33_ASAP7_75t_L      g15747(.A(new_n16003), .B(new_n16001), .C(new_n16000), .Y(new_n16004));
  A2O1A1O1Ixp25_ASAP7_75t_L g15748(.A1(new_n15503), .A2(new_n15318), .B(new_n15513), .C(new_n15657), .D(new_n15819), .Y(new_n16005));
  NOR2xp33_ASAP7_75t_L      g15749(.A(new_n16001), .B(new_n16000), .Y(new_n16006));
  O2A1O1Ixp33_ASAP7_75t_L   g15750(.A1(new_n16005), .A2(new_n15817), .B(new_n15821), .C(new_n16006), .Y(new_n16007));
  AOI22xp33_ASAP7_75t_L     g15751(.A1(new_n8831), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n9115), .Y(new_n16008));
  OAI221xp5_ASAP7_75t_L     g15752(.A1(new_n10343), .A2(new_n3180), .B1(new_n10016), .B2(new_n11047), .C(new_n16008), .Y(new_n16009));
  XNOR2x2_ASAP7_75t_L       g15753(.A(\a[56] ), .B(new_n16009), .Y(new_n16010));
  OAI21xp33_ASAP7_75t_L     g15754(.A1(new_n16007), .A2(new_n16004), .B(new_n16010), .Y(new_n16011));
  NOR2xp33_ASAP7_75t_L      g15755(.A(new_n16007), .B(new_n16004), .Y(new_n16012));
  INVx1_ASAP7_75t_L         g15756(.A(new_n16010), .Y(new_n16013));
  NAND2xp33_ASAP7_75t_L     g15757(.A(new_n16013), .B(new_n16012), .Y(new_n16014));
  AND2x2_ASAP7_75t_L        g15758(.A(new_n16011), .B(new_n16014), .Y(new_n16015));
  INVx1_ASAP7_75t_L         g15759(.A(new_n16015), .Y(new_n16016));
  A2O1A1Ixp33_ASAP7_75t_L   g15760(.A1(new_n15821), .A2(new_n15822), .B(new_n15826), .C(new_n15832), .Y(new_n16017));
  NOR2xp33_ASAP7_75t_L      g15761(.A(new_n16017), .B(new_n16016), .Y(new_n16018));
  O2A1O1Ixp33_ASAP7_75t_L   g15762(.A1(new_n15826), .A2(new_n15823), .B(new_n15832), .C(new_n16015), .Y(new_n16019));
  NOR2xp33_ASAP7_75t_L      g15763(.A(new_n16019), .B(new_n16018), .Y(new_n16020));
  NAND2xp33_ASAP7_75t_L     g15764(.A(new_n15975), .B(new_n16020), .Y(new_n16021));
  INVx1_ASAP7_75t_L         g15765(.A(new_n16021), .Y(new_n16022));
  NOR2xp33_ASAP7_75t_L      g15766(.A(new_n15975), .B(new_n16020), .Y(new_n16023));
  NOR2xp33_ASAP7_75t_L      g15767(.A(new_n16023), .B(new_n16022), .Y(new_n16024));
  NAND3xp33_ASAP7_75t_L     g15768(.A(new_n16024), .B(new_n15845), .C(new_n15838), .Y(new_n16025));
  INVx1_ASAP7_75t_L         g15769(.A(new_n15844), .Y(new_n16026));
  O2A1O1Ixp33_ASAP7_75t_L   g15770(.A1(new_n15840), .A2(new_n16026), .B(new_n15838), .C(new_n16024), .Y(new_n16027));
  INVx1_ASAP7_75t_L         g15771(.A(new_n16027), .Y(new_n16028));
  AOI22xp33_ASAP7_75t_L     g15772(.A1(new_n7111), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n7391), .Y(new_n16029));
  OAI221xp5_ASAP7_75t_L     g15773(.A1(new_n8558), .A2(new_n4424), .B1(new_n8237), .B2(new_n4641), .C(new_n16029), .Y(new_n16030));
  XNOR2x2_ASAP7_75t_L       g15774(.A(\a[50] ), .B(new_n16030), .Y(new_n16031));
  NAND3xp33_ASAP7_75t_L     g15775(.A(new_n16028), .B(new_n16025), .C(new_n16031), .Y(new_n16032));
  INVx1_ASAP7_75t_L         g15776(.A(new_n16032), .Y(new_n16033));
  AOI21xp33_ASAP7_75t_L     g15777(.A1(new_n16028), .A2(new_n16025), .B(new_n16031), .Y(new_n16034));
  NOR2xp33_ASAP7_75t_L      g15778(.A(new_n16034), .B(new_n16033), .Y(new_n16035));
  O2A1O1Ixp33_ASAP7_75t_L   g15779(.A1(new_n15848), .A2(new_n15851), .B(new_n15860), .C(new_n16035), .Y(new_n16036));
  INVx1_ASAP7_75t_L         g15780(.A(new_n15851), .Y(new_n16037));
  O2A1O1Ixp33_ASAP7_75t_L   g15781(.A1(new_n15846), .A2(new_n15847), .B(new_n16037), .C(new_n15859), .Y(new_n16038));
  NAND2xp33_ASAP7_75t_L     g15782(.A(new_n16035), .B(new_n16038), .Y(new_n16039));
  INVx1_ASAP7_75t_L         g15783(.A(new_n16039), .Y(new_n16040));
  NOR2xp33_ASAP7_75t_L      g15784(.A(new_n16036), .B(new_n16040), .Y(new_n16041));
  NAND2xp33_ASAP7_75t_L     g15785(.A(new_n15971), .B(new_n16041), .Y(new_n16042));
  INVx1_ASAP7_75t_L         g15786(.A(new_n16042), .Y(new_n16043));
  NOR2xp33_ASAP7_75t_L      g15787(.A(new_n15971), .B(new_n16041), .Y(new_n16044));
  NOR2xp33_ASAP7_75t_L      g15788(.A(new_n16044), .B(new_n16043), .Y(new_n16045));
  O2A1O1Ixp33_ASAP7_75t_L   g15789(.A1(new_n15863), .A2(new_n15864), .B(new_n15867), .C(new_n16045), .Y(new_n16046));
  INVx1_ASAP7_75t_L         g15790(.A(new_n16046), .Y(new_n16047));
  NAND3xp33_ASAP7_75t_L     g15791(.A(new_n16045), .B(new_n15867), .C(new_n15862), .Y(new_n16048));
  NAND3xp33_ASAP7_75t_L     g15792(.A(new_n16047), .B(new_n15968), .C(new_n16048), .Y(new_n16049));
  AO21x2_ASAP7_75t_L        g15793(.A1(new_n16048), .A2(new_n16047), .B(new_n15968), .Y(new_n16050));
  NAND2xp33_ASAP7_75t_L     g15794(.A(new_n16049), .B(new_n16050), .Y(new_n16051));
  O2A1O1Ixp33_ASAP7_75t_L   g15795(.A1(new_n15868), .A2(new_n15869), .B(new_n15788), .C(new_n15876), .Y(new_n16052));
  XNOR2x2_ASAP7_75t_L       g15796(.A(new_n16051), .B(new_n16052), .Y(new_n16053));
  AOI22xp33_ASAP7_75t_L     g15797(.A1(new_n4920), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n5167), .Y(new_n16054));
  OAI221xp5_ASAP7_75t_L     g15798(.A1(new_n5154), .A2(new_n6568), .B1(new_n5158), .B2(new_n6820), .C(new_n16054), .Y(new_n16055));
  XNOR2x2_ASAP7_75t_L       g15799(.A(\a[41] ), .B(new_n16055), .Y(new_n16056));
  XNOR2x2_ASAP7_75t_L       g15800(.A(new_n16056), .B(new_n16053), .Y(new_n16057));
  AO21x2_ASAP7_75t_L        g15801(.A1(new_n15880), .A2(new_n15887), .B(new_n16057), .Y(new_n16058));
  NAND3xp33_ASAP7_75t_L     g15802(.A(new_n16057), .B(new_n15887), .C(new_n15880), .Y(new_n16059));
  NAND2xp33_ASAP7_75t_L     g15803(.A(new_n16058), .B(new_n16059), .Y(new_n16060));
  AOI22xp33_ASAP7_75t_L     g15804(.A1(new_n4283), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n4512), .Y(new_n16061));
  OAI221xp5_ASAP7_75t_L     g15805(.A1(new_n4277), .A2(new_n7317), .B1(new_n4499), .B2(new_n7602), .C(new_n16061), .Y(new_n16062));
  XNOR2x2_ASAP7_75t_L       g15806(.A(\a[38] ), .B(new_n16062), .Y(new_n16063));
  NAND2xp33_ASAP7_75t_L     g15807(.A(new_n16063), .B(new_n16060), .Y(new_n16064));
  INVx1_ASAP7_75t_L         g15808(.A(new_n16063), .Y(new_n16065));
  NAND3xp33_ASAP7_75t_L     g15809(.A(new_n16058), .B(new_n16059), .C(new_n16065), .Y(new_n16066));
  NAND2xp33_ASAP7_75t_L     g15810(.A(new_n16066), .B(new_n16064), .Y(new_n16067));
  NAND2xp33_ASAP7_75t_L     g15811(.A(new_n15892), .B(new_n15897), .Y(new_n16068));
  NOR2xp33_ASAP7_75t_L      g15812(.A(new_n16068), .B(new_n16067), .Y(new_n16069));
  AOI22xp33_ASAP7_75t_L     g15813(.A1(new_n15897), .A2(new_n15892), .B1(new_n16066), .B2(new_n16064), .Y(new_n16070));
  NOR2xp33_ASAP7_75t_L      g15814(.A(new_n16069), .B(new_n16070), .Y(new_n16071));
  XOR2x2_ASAP7_75t_L        g15815(.A(new_n15964), .B(new_n16071), .Y(new_n16072));
  XOR2x2_ASAP7_75t_L        g15816(.A(new_n15961), .B(new_n16072), .Y(new_n16073));
  XNOR2x2_ASAP7_75t_L       g15817(.A(new_n15953), .B(new_n16073), .Y(new_n16074));
  XOR2x2_ASAP7_75t_L        g15818(.A(new_n16074), .B(new_n15946), .Y(new_n16075));
  NAND3xp33_ASAP7_75t_L     g15819(.A(new_n16075), .B(new_n15937), .C(new_n15936), .Y(new_n16076));
  AO21x2_ASAP7_75t_L        g15820(.A1(new_n15936), .A2(new_n15937), .B(new_n16075), .Y(new_n16077));
  AND2x2_ASAP7_75t_L        g15821(.A(new_n16076), .B(new_n16077), .Y(new_n16078));
  NAND3xp33_ASAP7_75t_L     g15822(.A(new_n16078), .B(new_n15917), .C(new_n15764), .Y(new_n16079));
  INVx1_ASAP7_75t_L         g15823(.A(new_n16079), .Y(new_n16080));
  O2A1O1Ixp33_ASAP7_75t_L   g15824(.A1(new_n15765), .A2(new_n15915), .B(new_n15764), .C(new_n16078), .Y(new_n16081));
  NOR2xp33_ASAP7_75t_L      g15825(.A(new_n16081), .B(new_n16080), .Y(new_n16082));
  A2O1A1Ixp33_ASAP7_75t_L   g15826(.A1(new_n15927), .A2(new_n15924), .B(new_n15923), .C(new_n16082), .Y(new_n16083));
  INVx1_ASAP7_75t_L         g15827(.A(new_n16083), .Y(new_n16084));
  A2O1A1Ixp33_ASAP7_75t_L   g15828(.A1(new_n15755), .A2(new_n15752), .B(new_n15921), .C(new_n15922), .Y(new_n16085));
  NOR2xp33_ASAP7_75t_L      g15829(.A(new_n16082), .B(new_n16085), .Y(new_n16086));
  NOR2xp33_ASAP7_75t_L      g15830(.A(new_n16084), .B(new_n16086), .Y(\f[86] ));
  A2O1A1Ixp33_ASAP7_75t_L   g15831(.A1(new_n15910), .A2(new_n15773), .B(new_n15934), .C(new_n16076), .Y(new_n16088));
  OA21x2_ASAP7_75t_L        g15832(.A1(new_n16074), .A2(new_n15946), .B(new_n15945), .Y(new_n16089));
  AOI22xp33_ASAP7_75t_L     g15833(.A1(new_n2114), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n2259), .Y(new_n16090));
  A2O1A1Ixp33_ASAP7_75t_L   g15834(.A1(new_n11470), .A2(new_n11473), .B(new_n2257), .C(new_n16090), .Y(new_n16091));
  AOI21xp33_ASAP7_75t_L     g15835(.A1(new_n2115), .A2(\b[62] ), .B(new_n16091), .Y(new_n16092));
  NAND2xp33_ASAP7_75t_L     g15836(.A(\a[26] ), .B(new_n16092), .Y(new_n16093));
  A2O1A1Ixp33_ASAP7_75t_L   g15837(.A1(\b[62] ), .A2(new_n2115), .B(new_n16091), .C(new_n2100), .Y(new_n16094));
  AND2x2_ASAP7_75t_L        g15838(.A(new_n16094), .B(new_n16093), .Y(new_n16095));
  INVx1_ASAP7_75t_L         g15839(.A(new_n16095), .Y(new_n16096));
  XNOR2x2_ASAP7_75t_L       g15840(.A(new_n16096), .B(new_n16089), .Y(new_n16097));
  INVx1_ASAP7_75t_L         g15841(.A(new_n15952), .Y(new_n16098));
  MAJIxp5_ASAP7_75t_L       g15842(.A(new_n16073), .B(new_n15949), .C(new_n16098), .Y(new_n16099));
  AOI22xp33_ASAP7_75t_L     g15843(.A1(new_n2552), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n2736), .Y(new_n16100));
  OAI221xp5_ASAP7_75t_L     g15844(.A1(new_n2547), .A2(new_n9947), .B1(new_n2734), .B2(new_n11446), .C(new_n16100), .Y(new_n16101));
  XNOR2x2_ASAP7_75t_L       g15845(.A(\a[29] ), .B(new_n16101), .Y(new_n16102));
  INVx1_ASAP7_75t_L         g15846(.A(new_n16102), .Y(new_n16103));
  XNOR2x2_ASAP7_75t_L       g15847(.A(new_n16103), .B(new_n16099), .Y(new_n16104));
  AOI22xp33_ASAP7_75t_L     g15848(.A1(new_n3029), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n3258), .Y(new_n16105));
  OAI221xp5_ASAP7_75t_L     g15849(.A1(new_n3024), .A2(new_n9323), .B1(new_n3256), .B2(new_n9627), .C(new_n16105), .Y(new_n16106));
  XNOR2x2_ASAP7_75t_L       g15850(.A(\a[32] ), .B(new_n16106), .Y(new_n16107));
  NOR2xp33_ASAP7_75t_L      g15851(.A(new_n15959), .B(new_n16072), .Y(new_n16108));
  NOR2xp33_ASAP7_75t_L      g15852(.A(new_n15960), .B(new_n16108), .Y(new_n16109));
  XNOR2x2_ASAP7_75t_L       g15853(.A(new_n16107), .B(new_n16109), .Y(new_n16110));
  AOI22xp33_ASAP7_75t_L     g15854(.A1(new_n3633), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n3858), .Y(new_n16111));
  OAI221xp5_ASAP7_75t_L     g15855(.A1(new_n3853), .A2(new_n8165), .B1(new_n3856), .B2(new_n8465), .C(new_n16111), .Y(new_n16112));
  XNOR2x2_ASAP7_75t_L       g15856(.A(\a[35] ), .B(new_n16112), .Y(new_n16113));
  INVx1_ASAP7_75t_L         g15857(.A(new_n16052), .Y(new_n16114));
  AND2x2_ASAP7_75t_L        g15858(.A(new_n16056), .B(new_n16053), .Y(new_n16115));
  AOI21xp33_ASAP7_75t_L     g15859(.A1(new_n16048), .A2(new_n15968), .B(new_n16046), .Y(new_n16116));
  AOI22xp33_ASAP7_75t_L     g15860(.A1(new_n5624), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n5901), .Y(new_n16117));
  OAI221xp5_ASAP7_75t_L     g15861(.A1(new_n5900), .A2(new_n5829), .B1(new_n5892), .B2(new_n6329), .C(new_n16117), .Y(new_n16118));
  XNOR2x2_ASAP7_75t_L       g15862(.A(\a[44] ), .B(new_n16118), .Y(new_n16119));
  INVx1_ASAP7_75t_L         g15863(.A(new_n16119), .Y(new_n16120));
  AOI22xp33_ASAP7_75t_L     g15864(.A1(new_n9700), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n10027), .Y(new_n16121));
  OAI221xp5_ASAP7_75t_L     g15865(.A1(new_n10024), .A2(new_n2688), .B1(new_n9696), .B2(new_n2990), .C(new_n16121), .Y(new_n16122));
  XNOR2x2_ASAP7_75t_L       g15866(.A(\a[59] ), .B(new_n16122), .Y(new_n16123));
  INVx1_ASAP7_75t_L         g15867(.A(new_n16123), .Y(new_n16124));
  NOR2xp33_ASAP7_75t_L      g15868(.A(new_n1909), .B(new_n11535), .Y(new_n16125));
  A2O1A1Ixp33_ASAP7_75t_L   g15869(.A1(new_n11533), .A2(\b[24] ), .B(new_n16125), .C(new_n1689), .Y(new_n16126));
  INVx1_ASAP7_75t_L         g15870(.A(new_n16126), .Y(new_n16127));
  O2A1O1Ixp33_ASAP7_75t_L   g15871(.A1(new_n11247), .A2(new_n11249), .B(\b[24] ), .C(new_n16125), .Y(new_n16128));
  NAND2xp33_ASAP7_75t_L     g15872(.A(\a[23] ), .B(new_n16128), .Y(new_n16129));
  INVx1_ASAP7_75t_L         g15873(.A(new_n16129), .Y(new_n16130));
  NOR2xp33_ASAP7_75t_L      g15874(.A(new_n16127), .B(new_n16130), .Y(new_n16131));
  A2O1A1Ixp33_ASAP7_75t_L   g15875(.A1(new_n11533), .A2(\b[23] ), .B(new_n15977), .C(new_n16131), .Y(new_n16132));
  OAI21xp33_ASAP7_75t_L     g15876(.A1(new_n16127), .A2(new_n16130), .B(new_n15978), .Y(new_n16133));
  AND2x2_ASAP7_75t_L        g15877(.A(new_n16133), .B(new_n16132), .Y(new_n16134));
  INVx1_ASAP7_75t_L         g15878(.A(new_n16134), .Y(new_n16135));
  AOI22xp33_ASAP7_75t_L     g15879(.A1(\b[25] ), .A2(new_n10939), .B1(\b[27] ), .B2(new_n10938), .Y(new_n16136));
  OAI221xp5_ASAP7_75t_L     g15880(.A1(new_n10937), .A2(new_n2348), .B1(new_n10629), .B2(new_n2505), .C(new_n16136), .Y(new_n16137));
  XNOR2x2_ASAP7_75t_L       g15881(.A(\a[62] ), .B(new_n16137), .Y(new_n16138));
  XNOR2x2_ASAP7_75t_L       g15882(.A(new_n16135), .B(new_n16138), .Y(new_n16139));
  O2A1O1Ixp33_ASAP7_75t_L   g15883(.A1(new_n15981), .A2(new_n15987), .B(new_n15979), .C(new_n16139), .Y(new_n16140));
  INVx1_ASAP7_75t_L         g15884(.A(new_n16140), .Y(new_n16141));
  A2O1A1O1Ixp25_ASAP7_75t_L g15885(.A1(new_n11533), .A2(\b[22] ), .B(new_n15799), .C(new_n15978), .D(new_n15988), .Y(new_n16142));
  NAND2xp33_ASAP7_75t_L     g15886(.A(new_n16142), .B(new_n16139), .Y(new_n16143));
  AND2x2_ASAP7_75t_L        g15887(.A(new_n16143), .B(new_n16141), .Y(new_n16144));
  NAND2xp33_ASAP7_75t_L     g15888(.A(new_n16124), .B(new_n16144), .Y(new_n16145));
  AO21x2_ASAP7_75t_L        g15889(.A1(new_n16143), .A2(new_n16141), .B(new_n16124), .Y(new_n16146));
  AND2x2_ASAP7_75t_L        g15890(.A(new_n16146), .B(new_n16145), .Y(new_n16147));
  O2A1O1Ixp33_ASAP7_75t_L   g15891(.A1(new_n15993), .A2(new_n15991), .B(new_n15999), .C(new_n16147), .Y(new_n16148));
  INVx1_ASAP7_75t_L         g15892(.A(new_n16147), .Y(new_n16149));
  A2O1A1Ixp33_ASAP7_75t_L   g15893(.A1(new_n15989), .A2(new_n15990), .B(new_n15993), .C(new_n15999), .Y(new_n16150));
  NOR2xp33_ASAP7_75t_L      g15894(.A(new_n16150), .B(new_n16149), .Y(new_n16151));
  NOR2xp33_ASAP7_75t_L      g15895(.A(new_n16148), .B(new_n16151), .Y(new_n16152));
  AOI22xp33_ASAP7_75t_L     g15896(.A1(new_n8831), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n9115), .Y(new_n16153));
  OAI221xp5_ASAP7_75t_L     g15897(.A1(new_n10343), .A2(new_n3207), .B1(new_n10016), .B2(new_n3572), .C(new_n16153), .Y(new_n16154));
  XNOR2x2_ASAP7_75t_L       g15898(.A(\a[56] ), .B(new_n16154), .Y(new_n16155));
  A2O1A1O1Ixp25_ASAP7_75t_L g15899(.A1(new_n15821), .A2(new_n16002), .B(new_n16006), .C(new_n16014), .D(new_n16155), .Y(new_n16156));
  INVx1_ASAP7_75t_L         g15900(.A(new_n16155), .Y(new_n16157));
  A2O1A1Ixp33_ASAP7_75t_L   g15901(.A1(new_n15821), .A2(new_n16002), .B(new_n16006), .C(new_n16014), .Y(new_n16158));
  NOR2xp33_ASAP7_75t_L      g15902(.A(new_n16157), .B(new_n16158), .Y(new_n16159));
  NOR2xp33_ASAP7_75t_L      g15903(.A(new_n16156), .B(new_n16159), .Y(new_n16160));
  NAND2xp33_ASAP7_75t_L     g15904(.A(new_n16152), .B(new_n16160), .Y(new_n16161));
  INVx1_ASAP7_75t_L         g15905(.A(new_n16161), .Y(new_n16162));
  NOR2xp33_ASAP7_75t_L      g15906(.A(new_n16152), .B(new_n16160), .Y(new_n16163));
  NOR2xp33_ASAP7_75t_L      g15907(.A(new_n16163), .B(new_n16162), .Y(new_n16164));
  AOI22xp33_ASAP7_75t_L     g15908(.A1(new_n7960), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n8537), .Y(new_n16165));
  OAI221xp5_ASAP7_75t_L     g15909(.A1(new_n8817), .A2(new_n3804), .B1(new_n7957), .B2(new_n4223), .C(new_n16165), .Y(new_n16166));
  XNOR2x2_ASAP7_75t_L       g15910(.A(\a[53] ), .B(new_n16166), .Y(new_n16167));
  INVx1_ASAP7_75t_L         g15911(.A(new_n16167), .Y(new_n16168));
  XNOR2x2_ASAP7_75t_L       g15912(.A(new_n16168), .B(new_n16164), .Y(new_n16169));
  INVx1_ASAP7_75t_L         g15913(.A(new_n16169), .Y(new_n16170));
  NOR3xp33_ASAP7_75t_L      g15914(.A(new_n16170), .B(new_n16022), .C(new_n16018), .Y(new_n16171));
  O2A1O1Ixp33_ASAP7_75t_L   g15915(.A1(new_n16016), .A2(new_n16017), .B(new_n16021), .C(new_n16169), .Y(new_n16172));
  NOR2xp33_ASAP7_75t_L      g15916(.A(new_n16172), .B(new_n16171), .Y(new_n16173));
  AOI22xp33_ASAP7_75t_L     g15917(.A1(new_n7111), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n7391), .Y(new_n16174));
  OAI221xp5_ASAP7_75t_L     g15918(.A1(new_n8558), .A2(new_n4632), .B1(new_n8237), .B2(new_n4858), .C(new_n16174), .Y(new_n16175));
  XNOR2x2_ASAP7_75t_L       g15919(.A(\a[50] ), .B(new_n16175), .Y(new_n16176));
  INVx1_ASAP7_75t_L         g15920(.A(new_n16176), .Y(new_n16177));
  XNOR2x2_ASAP7_75t_L       g15921(.A(new_n16177), .B(new_n16173), .Y(new_n16178));
  A2O1A1Ixp33_ASAP7_75t_L   g15922(.A1(new_n16031), .A2(new_n16025), .B(new_n16027), .C(new_n16178), .Y(new_n16179));
  A2O1A1Ixp33_ASAP7_75t_L   g15923(.A1(new_n15845), .A2(new_n15838), .B(new_n16024), .C(new_n16032), .Y(new_n16180));
  NOR2xp33_ASAP7_75t_L      g15924(.A(new_n16180), .B(new_n16178), .Y(new_n16181));
  INVx1_ASAP7_75t_L         g15925(.A(new_n16181), .Y(new_n16182));
  NAND2xp33_ASAP7_75t_L     g15926(.A(new_n16179), .B(new_n16182), .Y(new_n16183));
  AOI22xp33_ASAP7_75t_L     g15927(.A1(new_n6376), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n6648), .Y(new_n16184));
  OAI221xp5_ASAP7_75t_L     g15928(.A1(new_n6646), .A2(new_n5321), .B1(new_n6636), .B2(new_n5346), .C(new_n16184), .Y(new_n16185));
  XNOR2x2_ASAP7_75t_L       g15929(.A(\a[47] ), .B(new_n16185), .Y(new_n16186));
  XNOR2x2_ASAP7_75t_L       g15930(.A(new_n16186), .B(new_n16183), .Y(new_n16187));
  NOR3xp33_ASAP7_75t_L      g15931(.A(new_n16043), .B(new_n16187), .C(new_n16040), .Y(new_n16188));
  INVx1_ASAP7_75t_L         g15932(.A(new_n16188), .Y(new_n16189));
  A2O1A1Ixp33_ASAP7_75t_L   g15933(.A1(new_n16041), .A2(new_n15971), .B(new_n16040), .C(new_n16187), .Y(new_n16190));
  AND2x2_ASAP7_75t_L        g15934(.A(new_n16190), .B(new_n16189), .Y(new_n16191));
  NAND2xp33_ASAP7_75t_L     g15935(.A(new_n16120), .B(new_n16191), .Y(new_n16192));
  NOR2xp33_ASAP7_75t_L      g15936(.A(new_n16120), .B(new_n16191), .Y(new_n16193));
  INVx1_ASAP7_75t_L         g15937(.A(new_n16193), .Y(new_n16194));
  NAND2xp33_ASAP7_75t_L     g15938(.A(new_n16192), .B(new_n16194), .Y(new_n16195));
  XNOR2x2_ASAP7_75t_L       g15939(.A(new_n16116), .B(new_n16195), .Y(new_n16196));
  AOI22xp33_ASAP7_75t_L     g15940(.A1(new_n4920), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n5167), .Y(new_n16197));
  OAI221xp5_ASAP7_75t_L     g15941(.A1(new_n5154), .A2(new_n6812), .B1(new_n5158), .B2(new_n6837), .C(new_n16197), .Y(new_n16198));
  XNOR2x2_ASAP7_75t_L       g15942(.A(\a[41] ), .B(new_n16198), .Y(new_n16199));
  XNOR2x2_ASAP7_75t_L       g15943(.A(new_n16199), .B(new_n16196), .Y(new_n16200));
  A2O1A1Ixp33_ASAP7_75t_L   g15944(.A1(new_n16114), .A2(new_n16051), .B(new_n16115), .C(new_n16200), .Y(new_n16201));
  INVx1_ASAP7_75t_L         g15945(.A(new_n16200), .Y(new_n16202));
  INVx1_ASAP7_75t_L         g15946(.A(new_n15871), .Y(new_n16203));
  O2A1O1Ixp33_ASAP7_75t_L   g15947(.A1(new_n16203), .A2(new_n15876), .B(new_n16051), .C(new_n16115), .Y(new_n16204));
  NAND2xp33_ASAP7_75t_L     g15948(.A(new_n16204), .B(new_n16202), .Y(new_n16205));
  NAND2xp33_ASAP7_75t_L     g15949(.A(new_n16201), .B(new_n16205), .Y(new_n16206));
  AOI22xp33_ASAP7_75t_L     g15950(.A1(new_n4283), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n4512), .Y(new_n16207));
  OAI221xp5_ASAP7_75t_L     g15951(.A1(new_n4277), .A2(new_n7593), .B1(new_n4499), .B2(new_n7623), .C(new_n16207), .Y(new_n16208));
  XNOR2x2_ASAP7_75t_L       g15952(.A(\a[38] ), .B(new_n16208), .Y(new_n16209));
  XNOR2x2_ASAP7_75t_L       g15953(.A(new_n16209), .B(new_n16206), .Y(new_n16210));
  AND3x1_ASAP7_75t_L        g15954(.A(new_n16210), .B(new_n16066), .C(new_n16059), .Y(new_n16211));
  O2A1O1Ixp33_ASAP7_75t_L   g15955(.A1(new_n15881), .A2(new_n15882), .B(new_n15887), .C(new_n16057), .Y(new_n16212));
  O2A1O1Ixp33_ASAP7_75t_L   g15956(.A1(new_n16212), .A2(new_n16063), .B(new_n16059), .C(new_n16210), .Y(new_n16213));
  NOR2xp33_ASAP7_75t_L      g15957(.A(new_n16213), .B(new_n16211), .Y(new_n16214));
  INVx1_ASAP7_75t_L         g15958(.A(new_n16214), .Y(new_n16215));
  NAND2xp33_ASAP7_75t_L     g15959(.A(new_n16113), .B(new_n16215), .Y(new_n16216));
  OR3x1_ASAP7_75t_L         g15960(.A(new_n16211), .B(new_n16113), .C(new_n16213), .Y(new_n16217));
  AND2x2_ASAP7_75t_L        g15961(.A(new_n16217), .B(new_n16216), .Y(new_n16218));
  AOI21xp33_ASAP7_75t_L     g15962(.A1(new_n16071), .A2(new_n15964), .B(new_n16070), .Y(new_n16219));
  NAND2xp33_ASAP7_75t_L     g15963(.A(new_n16219), .B(new_n16218), .Y(new_n16220));
  INVx1_ASAP7_75t_L         g15964(.A(new_n16218), .Y(new_n16221));
  A2O1A1Ixp33_ASAP7_75t_L   g15965(.A1(new_n16071), .A2(new_n15964), .B(new_n16070), .C(new_n16221), .Y(new_n16222));
  NAND2xp33_ASAP7_75t_L     g15966(.A(new_n16220), .B(new_n16222), .Y(new_n16223));
  XOR2x2_ASAP7_75t_L        g15967(.A(new_n16223), .B(new_n16110), .Y(new_n16224));
  XOR2x2_ASAP7_75t_L        g15968(.A(new_n16104), .B(new_n16224), .Y(new_n16225));
  INVx1_ASAP7_75t_L         g15969(.A(new_n16225), .Y(new_n16226));
  NAND2xp33_ASAP7_75t_L     g15970(.A(new_n16097), .B(new_n16226), .Y(new_n16227));
  NOR2xp33_ASAP7_75t_L      g15971(.A(new_n16097), .B(new_n16226), .Y(new_n16228));
  INVx1_ASAP7_75t_L         g15972(.A(new_n16228), .Y(new_n16229));
  NAND3xp33_ASAP7_75t_L     g15973(.A(new_n16229), .B(new_n16227), .C(new_n16088), .Y(new_n16230));
  AO21x2_ASAP7_75t_L        g15974(.A1(new_n16227), .A2(new_n16229), .B(new_n16088), .Y(new_n16231));
  NAND2xp33_ASAP7_75t_L     g15975(.A(new_n16230), .B(new_n16231), .Y(new_n16232));
  INVx1_ASAP7_75t_L         g15976(.A(new_n16232), .Y(new_n16233));
  A2O1A1Ixp33_ASAP7_75t_L   g15977(.A1(new_n16085), .A2(new_n16082), .B(new_n16080), .C(new_n16233), .Y(new_n16234));
  INVx1_ASAP7_75t_L         g15978(.A(new_n16234), .Y(new_n16235));
  A2O1A1Ixp33_ASAP7_75t_L   g15979(.A1(new_n15925), .A2(new_n15922), .B(new_n16081), .C(new_n16079), .Y(new_n16236));
  NOR2xp33_ASAP7_75t_L      g15980(.A(new_n16233), .B(new_n16236), .Y(new_n16237));
  NOR2xp33_ASAP7_75t_L      g15981(.A(new_n16237), .B(new_n16235), .Y(\f[87] ));
  INVx1_ASAP7_75t_L         g15982(.A(new_n16230), .Y(new_n16239));
  AOI22xp33_ASAP7_75t_L     g15983(.A1(new_n2552), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n2736), .Y(new_n16240));
  OAI221xp5_ASAP7_75t_L     g15984(.A1(new_n2547), .A2(new_n10250), .B1(new_n2734), .B2(new_n10855), .C(new_n16240), .Y(new_n16241));
  XNOR2x2_ASAP7_75t_L       g15985(.A(\a[29] ), .B(new_n16241), .Y(new_n16242));
  MAJIxp5_ASAP7_75t_L       g15986(.A(new_n16223), .B(new_n16107), .C(new_n16109), .Y(new_n16243));
  XNOR2x2_ASAP7_75t_L       g15987(.A(new_n16242), .B(new_n16243), .Y(new_n16244));
  NOR2xp33_ASAP7_75t_L      g15988(.A(new_n9920), .B(new_n3022), .Y(new_n16245));
  AOI221xp5_ASAP7_75t_L     g15989(.A1(\b[56] ), .A2(new_n3258), .B1(\b[57] ), .B2(new_n3030), .C(new_n16245), .Y(new_n16246));
  OAI211xp5_ASAP7_75t_L     g15990(.A1(new_n3256), .A2(new_n9925), .B(\a[32] ), .C(new_n16246), .Y(new_n16247));
  INVx1_ASAP7_75t_L         g15991(.A(new_n16247), .Y(new_n16248));
  O2A1O1Ixp33_ASAP7_75t_L   g15992(.A1(new_n3256), .A2(new_n9925), .B(new_n16246), .C(\a[32] ), .Y(new_n16249));
  NOR2xp33_ASAP7_75t_L      g15993(.A(new_n16249), .B(new_n16248), .Y(new_n16250));
  O2A1O1Ixp33_ASAP7_75t_L   g15994(.A1(new_n16113), .A2(new_n16215), .B(new_n16220), .C(new_n16250), .Y(new_n16251));
  INVx1_ASAP7_75t_L         g15995(.A(new_n16251), .Y(new_n16252));
  NAND3xp33_ASAP7_75t_L     g15996(.A(new_n16220), .B(new_n16217), .C(new_n16250), .Y(new_n16253));
  AOI22xp33_ASAP7_75t_L     g15997(.A1(new_n7111), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n7391), .Y(new_n16254));
  OAI221xp5_ASAP7_75t_L     g15998(.A1(new_n8558), .A2(new_n4848), .B1(new_n8237), .B2(new_n11686), .C(new_n16254), .Y(new_n16255));
  XNOR2x2_ASAP7_75t_L       g15999(.A(\a[50] ), .B(new_n16255), .Y(new_n16256));
  INVx1_ASAP7_75t_L         g16000(.A(new_n16256), .Y(new_n16257));
  INVx1_ASAP7_75t_L         g16001(.A(new_n16138), .Y(new_n16258));
  NOR2xp33_ASAP7_75t_L      g16002(.A(new_n1929), .B(new_n11535), .Y(new_n16259));
  A2O1A1O1Ixp25_ASAP7_75t_L g16003(.A1(new_n11533), .A2(\b[23] ), .B(new_n15977), .C(new_n16129), .D(new_n16127), .Y(new_n16260));
  A2O1A1Ixp33_ASAP7_75t_L   g16004(.A1(new_n11533), .A2(\b[25] ), .B(new_n16259), .C(new_n16260), .Y(new_n16261));
  O2A1O1Ixp33_ASAP7_75t_L   g16005(.A1(new_n11247), .A2(new_n11249), .B(\b[25] ), .C(new_n16259), .Y(new_n16262));
  INVx1_ASAP7_75t_L         g16006(.A(new_n16262), .Y(new_n16263));
  O2A1O1Ixp33_ASAP7_75t_L   g16007(.A1(new_n15978), .A2(new_n16130), .B(new_n16126), .C(new_n16263), .Y(new_n16264));
  INVx1_ASAP7_75t_L         g16008(.A(new_n16264), .Y(new_n16265));
  NAND2xp33_ASAP7_75t_L     g16009(.A(new_n16261), .B(new_n16265), .Y(new_n16266));
  NOR2xp33_ASAP7_75t_L      g16010(.A(new_n2666), .B(new_n10630), .Y(new_n16267));
  AOI221xp5_ASAP7_75t_L     g16011(.A1(\b[26] ), .A2(new_n10939), .B1(\b[27] ), .B2(new_n10632), .C(new_n16267), .Y(new_n16268));
  OAI211xp5_ASAP7_75t_L     g16012(.A1(new_n10629), .A2(new_n2672), .B(\a[62] ), .C(new_n16268), .Y(new_n16269));
  O2A1O1Ixp33_ASAP7_75t_L   g16013(.A1(new_n10629), .A2(new_n2672), .B(new_n16268), .C(\a[62] ), .Y(new_n16270));
  INVx1_ASAP7_75t_L         g16014(.A(new_n16270), .Y(new_n16271));
  AND2x2_ASAP7_75t_L        g16015(.A(new_n16269), .B(new_n16271), .Y(new_n16272));
  NOR2xp33_ASAP7_75t_L      g16016(.A(new_n16266), .B(new_n16272), .Y(new_n16273));
  INVx1_ASAP7_75t_L         g16017(.A(new_n16273), .Y(new_n16274));
  NAND2xp33_ASAP7_75t_L     g16018(.A(new_n16266), .B(new_n16272), .Y(new_n16275));
  AND2x2_ASAP7_75t_L        g16019(.A(new_n16275), .B(new_n16274), .Y(new_n16276));
  A2O1A1Ixp33_ASAP7_75t_L   g16020(.A1(new_n16258), .A2(new_n16134), .B(new_n16140), .C(new_n16276), .Y(new_n16277));
  AOI21xp33_ASAP7_75t_L     g16021(.A1(new_n16258), .A2(new_n16134), .B(new_n16140), .Y(new_n16278));
  INVx1_ASAP7_75t_L         g16022(.A(new_n16278), .Y(new_n16279));
  NOR2xp33_ASAP7_75t_L      g16023(.A(new_n16276), .B(new_n16279), .Y(new_n16280));
  INVx1_ASAP7_75t_L         g16024(.A(new_n16280), .Y(new_n16281));
  AOI22xp33_ASAP7_75t_L     g16025(.A1(new_n9700), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n10027), .Y(new_n16282));
  OAI221xp5_ASAP7_75t_L     g16026(.A1(new_n10024), .A2(new_n2982), .B1(new_n9696), .B2(new_n3187), .C(new_n16282), .Y(new_n16283));
  XNOR2x2_ASAP7_75t_L       g16027(.A(\a[59] ), .B(new_n16283), .Y(new_n16284));
  NAND3xp33_ASAP7_75t_L     g16028(.A(new_n16281), .B(new_n16277), .C(new_n16284), .Y(new_n16285));
  AO21x2_ASAP7_75t_L        g16029(.A1(new_n16277), .A2(new_n16281), .B(new_n16284), .Y(new_n16286));
  AND2x2_ASAP7_75t_L        g16030(.A(new_n16285), .B(new_n16286), .Y(new_n16287));
  OAI211xp5_ASAP7_75t_L     g16031(.A1(new_n16149), .A2(new_n16150), .B(new_n16287), .C(new_n16145), .Y(new_n16288));
  O2A1O1Ixp33_ASAP7_75t_L   g16032(.A1(new_n16149), .A2(new_n16150), .B(new_n16145), .C(new_n16287), .Y(new_n16289));
  INVx1_ASAP7_75t_L         g16033(.A(new_n16289), .Y(new_n16290));
  NAND2xp33_ASAP7_75t_L     g16034(.A(\b[32] ), .B(new_n9115), .Y(new_n16291));
  OAI221xp5_ASAP7_75t_L     g16035(.A1(new_n9113), .A2(new_n3584), .B1(new_n10016), .B2(new_n3591), .C(new_n16291), .Y(new_n16292));
  AOI21xp33_ASAP7_75t_L     g16036(.A1(new_n8835), .A2(\b[33] ), .B(new_n16292), .Y(new_n16293));
  NAND2xp33_ASAP7_75t_L     g16037(.A(\a[56] ), .B(new_n16293), .Y(new_n16294));
  A2O1A1Ixp33_ASAP7_75t_L   g16038(.A1(\b[33] ), .A2(new_n8835), .B(new_n16292), .C(new_n8826), .Y(new_n16295));
  AND2x2_ASAP7_75t_L        g16039(.A(new_n16295), .B(new_n16294), .Y(new_n16296));
  NAND3xp33_ASAP7_75t_L     g16040(.A(new_n16290), .B(new_n16288), .C(new_n16296), .Y(new_n16297));
  AO21x2_ASAP7_75t_L        g16041(.A1(new_n16288), .A2(new_n16290), .B(new_n16296), .Y(new_n16298));
  AND2x2_ASAP7_75t_L        g16042(.A(new_n16297), .B(new_n16298), .Y(new_n16299));
  A2O1A1O1Ixp25_ASAP7_75t_L g16043(.A1(new_n16012), .A2(new_n16013), .B(new_n16007), .C(new_n16157), .D(new_n16162), .Y(new_n16300));
  NAND2xp33_ASAP7_75t_L     g16044(.A(new_n16299), .B(new_n16300), .Y(new_n16301));
  INVx1_ASAP7_75t_L         g16045(.A(new_n16299), .Y(new_n16302));
  A2O1A1Ixp33_ASAP7_75t_L   g16046(.A1(new_n16160), .A2(new_n16152), .B(new_n16156), .C(new_n16302), .Y(new_n16303));
  AND2x2_ASAP7_75t_L        g16047(.A(new_n16303), .B(new_n16301), .Y(new_n16304));
  INVx1_ASAP7_75t_L         g16048(.A(new_n16304), .Y(new_n16305));
  AOI22xp33_ASAP7_75t_L     g16049(.A1(new_n7960), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n8537), .Y(new_n16306));
  OAI221xp5_ASAP7_75t_L     g16050(.A1(new_n8817), .A2(new_n4216), .B1(new_n7957), .B2(new_n4431), .C(new_n16306), .Y(new_n16307));
  XNOR2x2_ASAP7_75t_L       g16051(.A(\a[53] ), .B(new_n16307), .Y(new_n16308));
  NAND2xp33_ASAP7_75t_L     g16052(.A(new_n16308), .B(new_n16305), .Y(new_n16309));
  NOR2xp33_ASAP7_75t_L      g16053(.A(new_n16308), .B(new_n16305), .Y(new_n16310));
  INVx1_ASAP7_75t_L         g16054(.A(new_n16310), .Y(new_n16311));
  AND2x2_ASAP7_75t_L        g16055(.A(new_n16309), .B(new_n16311), .Y(new_n16312));
  A2O1A1Ixp33_ASAP7_75t_L   g16056(.A1(new_n16168), .A2(new_n16164), .B(new_n16172), .C(new_n16312), .Y(new_n16313));
  NOR3xp33_ASAP7_75t_L      g16057(.A(new_n16162), .B(new_n16163), .C(new_n16167), .Y(new_n16314));
  O2A1O1Ixp33_ASAP7_75t_L   g16058(.A1(new_n16018), .A2(new_n16022), .B(new_n16170), .C(new_n16314), .Y(new_n16315));
  INVx1_ASAP7_75t_L         g16059(.A(new_n16312), .Y(new_n16316));
  NAND2xp33_ASAP7_75t_L     g16060(.A(new_n16315), .B(new_n16316), .Y(new_n16317));
  AND2x2_ASAP7_75t_L        g16061(.A(new_n16313), .B(new_n16317), .Y(new_n16318));
  NAND2xp33_ASAP7_75t_L     g16062(.A(new_n16257), .B(new_n16318), .Y(new_n16319));
  AO21x2_ASAP7_75t_L        g16063(.A1(new_n16313), .A2(new_n16317), .B(new_n16257), .Y(new_n16320));
  AND2x2_ASAP7_75t_L        g16064(.A(new_n16320), .B(new_n16319), .Y(new_n16321));
  A2O1A1Ixp33_ASAP7_75t_L   g16065(.A1(new_n16177), .A2(new_n16173), .B(new_n16181), .C(new_n16321), .Y(new_n16322));
  AOI21xp33_ASAP7_75t_L     g16066(.A1(new_n16177), .A2(new_n16173), .B(new_n16181), .Y(new_n16323));
  INVx1_ASAP7_75t_L         g16067(.A(new_n16323), .Y(new_n16324));
  NOR2xp33_ASAP7_75t_L      g16068(.A(new_n16324), .B(new_n16321), .Y(new_n16325));
  INVx1_ASAP7_75t_L         g16069(.A(new_n16325), .Y(new_n16326));
  AOI22xp33_ASAP7_75t_L     g16070(.A1(new_n6376), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n6648), .Y(new_n16327));
  OAI221xp5_ASAP7_75t_L     g16071(.A1(new_n6646), .A2(new_n5338), .B1(new_n6636), .B2(new_n6338), .C(new_n16327), .Y(new_n16328));
  XNOR2x2_ASAP7_75t_L       g16072(.A(\a[47] ), .B(new_n16328), .Y(new_n16329));
  NAND3xp33_ASAP7_75t_L     g16073(.A(new_n16326), .B(new_n16322), .C(new_n16329), .Y(new_n16330));
  AO21x2_ASAP7_75t_L        g16074(.A1(new_n16322), .A2(new_n16326), .B(new_n16329), .Y(new_n16331));
  NAND2xp33_ASAP7_75t_L     g16075(.A(new_n16330), .B(new_n16331), .Y(new_n16332));
  OAI21xp33_ASAP7_75t_L     g16076(.A1(new_n16183), .A2(new_n16186), .B(new_n16189), .Y(new_n16333));
  NOR2xp33_ASAP7_75t_L      g16077(.A(new_n16333), .B(new_n16332), .Y(new_n16334));
  INVx1_ASAP7_75t_L         g16078(.A(new_n16334), .Y(new_n16335));
  NAND2xp33_ASAP7_75t_L     g16079(.A(new_n16333), .B(new_n16332), .Y(new_n16336));
  AOI22xp33_ASAP7_75t_L     g16080(.A1(new_n5624), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n5901), .Y(new_n16337));
  OAI221xp5_ASAP7_75t_L     g16081(.A1(new_n5900), .A2(new_n6321), .B1(new_n5892), .B2(new_n6573), .C(new_n16337), .Y(new_n16338));
  XNOR2x2_ASAP7_75t_L       g16082(.A(\a[44] ), .B(new_n16338), .Y(new_n16339));
  NAND3xp33_ASAP7_75t_L     g16083(.A(new_n16335), .B(new_n16336), .C(new_n16339), .Y(new_n16340));
  AO21x2_ASAP7_75t_L        g16084(.A1(new_n16336), .A2(new_n16335), .B(new_n16339), .Y(new_n16341));
  NAND2xp33_ASAP7_75t_L     g16085(.A(new_n16340), .B(new_n16341), .Y(new_n16342));
  A2O1A1Ixp33_ASAP7_75t_L   g16086(.A1(new_n16049), .A2(new_n16047), .B(new_n16193), .C(new_n16192), .Y(new_n16343));
  NOR2xp33_ASAP7_75t_L      g16087(.A(new_n16343), .B(new_n16342), .Y(new_n16344));
  INVx1_ASAP7_75t_L         g16088(.A(new_n16344), .Y(new_n16345));
  A2O1A1O1Ixp25_ASAP7_75t_L g16089(.A1(new_n15867), .A2(new_n15862), .B(new_n16045), .C(new_n16049), .D(new_n16195), .Y(new_n16346));
  A2O1A1Ixp33_ASAP7_75t_L   g16090(.A1(new_n16191), .A2(new_n16120), .B(new_n16346), .C(new_n16342), .Y(new_n16347));
  AOI22xp33_ASAP7_75t_L     g16091(.A1(new_n4920), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n5167), .Y(new_n16348));
  OAI221xp5_ASAP7_75t_L     g16092(.A1(new_n5154), .A2(new_n6830), .B1(new_n5158), .B2(new_n7323), .C(new_n16348), .Y(new_n16349));
  XNOR2x2_ASAP7_75t_L       g16093(.A(\a[41] ), .B(new_n16349), .Y(new_n16350));
  AND3x1_ASAP7_75t_L        g16094(.A(new_n16345), .B(new_n16350), .C(new_n16347), .Y(new_n16351));
  AOI21xp33_ASAP7_75t_L     g16095(.A1(new_n16345), .A2(new_n16347), .B(new_n16350), .Y(new_n16352));
  OR2x4_ASAP7_75t_L         g16096(.A(new_n16352), .B(new_n16351), .Y(new_n16353));
  OAI21xp33_ASAP7_75t_L     g16097(.A1(new_n16196), .A2(new_n16199), .B(new_n16205), .Y(new_n16354));
  NOR2xp33_ASAP7_75t_L      g16098(.A(new_n16353), .B(new_n16354), .Y(new_n16355));
  INVx1_ASAP7_75t_L         g16099(.A(new_n16355), .Y(new_n16356));
  NOR2xp33_ASAP7_75t_L      g16100(.A(new_n16199), .B(new_n16196), .Y(new_n16357));
  A2O1A1Ixp33_ASAP7_75t_L   g16101(.A1(new_n16202), .A2(new_n16204), .B(new_n16357), .C(new_n16353), .Y(new_n16358));
  NAND2xp33_ASAP7_75t_L     g16102(.A(new_n16358), .B(new_n16356), .Y(new_n16359));
  AOI22xp33_ASAP7_75t_L     g16103(.A1(new_n4283), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n4512), .Y(new_n16360));
  OAI221xp5_ASAP7_75t_L     g16104(.A1(new_n4277), .A2(new_n7616), .B1(new_n4499), .B2(new_n7906), .C(new_n16360), .Y(new_n16361));
  XNOR2x2_ASAP7_75t_L       g16105(.A(\a[38] ), .B(new_n16361), .Y(new_n16362));
  XNOR2x2_ASAP7_75t_L       g16106(.A(new_n16362), .B(new_n16359), .Y(new_n16363));
  NOR2xp33_ASAP7_75t_L      g16107(.A(new_n16209), .B(new_n16206), .Y(new_n16364));
  NOR2xp33_ASAP7_75t_L      g16108(.A(new_n16364), .B(new_n16213), .Y(new_n16365));
  XOR2x2_ASAP7_75t_L        g16109(.A(new_n16365), .B(new_n16363), .Y(new_n16366));
  AOI22xp33_ASAP7_75t_L     g16110(.A1(new_n3633), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n3858), .Y(new_n16367));
  OAI221xp5_ASAP7_75t_L     g16111(.A1(new_n3853), .A2(new_n8458), .B1(new_n3856), .B2(new_n8768), .C(new_n16367), .Y(new_n16368));
  XNOR2x2_ASAP7_75t_L       g16112(.A(\a[35] ), .B(new_n16368), .Y(new_n16369));
  XNOR2x2_ASAP7_75t_L       g16113(.A(new_n16369), .B(new_n16366), .Y(new_n16370));
  NAND3xp33_ASAP7_75t_L     g16114(.A(new_n16252), .B(new_n16253), .C(new_n16370), .Y(new_n16371));
  INVx1_ASAP7_75t_L         g16115(.A(new_n16253), .Y(new_n16372));
  INVx1_ASAP7_75t_L         g16116(.A(new_n16370), .Y(new_n16373));
  OAI21xp33_ASAP7_75t_L     g16117(.A1(new_n16251), .A2(new_n16372), .B(new_n16373), .Y(new_n16374));
  NAND2xp33_ASAP7_75t_L     g16118(.A(new_n16374), .B(new_n16371), .Y(new_n16375));
  XNOR2x2_ASAP7_75t_L       g16119(.A(new_n16375), .B(new_n16244), .Y(new_n16376));
  MAJIxp5_ASAP7_75t_L       g16120(.A(new_n16224), .B(new_n16099), .C(new_n16103), .Y(new_n16377));
  NOR2xp33_ASAP7_75t_L      g16121(.A(new_n2257), .B(new_n11500), .Y(new_n16378));
  AOI21xp33_ASAP7_75t_L     g16122(.A1(new_n2259), .A2(\b[62] ), .B(new_n16378), .Y(new_n16379));
  OAI211xp5_ASAP7_75t_L     g16123(.A1(new_n11468), .A2(new_n2109), .B(new_n16379), .C(\a[26] ), .Y(new_n16380));
  O2A1O1Ixp33_ASAP7_75t_L   g16124(.A1(new_n11468), .A2(new_n2109), .B(new_n16379), .C(\a[26] ), .Y(new_n16381));
  INVx1_ASAP7_75t_L         g16125(.A(new_n16381), .Y(new_n16382));
  AND2x2_ASAP7_75t_L        g16126(.A(new_n16380), .B(new_n16382), .Y(new_n16383));
  XOR2x2_ASAP7_75t_L        g16127(.A(new_n16383), .B(new_n16377), .Y(new_n16384));
  XNOR2x2_ASAP7_75t_L       g16128(.A(new_n16376), .B(new_n16384), .Y(new_n16385));
  O2A1O1Ixp33_ASAP7_75t_L   g16129(.A1(new_n16089), .A2(new_n16095), .B(new_n16227), .C(new_n16385), .Y(new_n16386));
  A2O1A1Ixp33_ASAP7_75t_L   g16130(.A1(new_n16093), .A2(new_n16094), .B(new_n16089), .C(new_n16227), .Y(new_n16387));
  INVx1_ASAP7_75t_L         g16131(.A(new_n16385), .Y(new_n16388));
  NOR2xp33_ASAP7_75t_L      g16132(.A(new_n16387), .B(new_n16388), .Y(new_n16389));
  NOR2xp33_ASAP7_75t_L      g16133(.A(new_n16386), .B(new_n16389), .Y(new_n16390));
  A2O1A1Ixp33_ASAP7_75t_L   g16134(.A1(new_n16236), .A2(new_n16233), .B(new_n16239), .C(new_n16390), .Y(new_n16391));
  INVx1_ASAP7_75t_L         g16135(.A(new_n16391), .Y(new_n16392));
  A2O1A1Ixp33_ASAP7_75t_L   g16136(.A1(new_n16083), .A2(new_n16079), .B(new_n16232), .C(new_n16230), .Y(new_n16393));
  NOR2xp33_ASAP7_75t_L      g16137(.A(new_n16390), .B(new_n16393), .Y(new_n16394));
  NOR2xp33_ASAP7_75t_L      g16138(.A(new_n16394), .B(new_n16392), .Y(\f[88] ));
  NOR2xp33_ASAP7_75t_L      g16139(.A(new_n16383), .B(new_n16377), .Y(new_n16396));
  AOI21xp33_ASAP7_75t_L     g16140(.A1(new_n16384), .A2(new_n16376), .B(new_n16396), .Y(new_n16397));
  AOI22xp33_ASAP7_75t_L     g16141(.A1(new_n2552), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n2736), .Y(new_n16398));
  OAI221xp5_ASAP7_75t_L     g16142(.A1(new_n2547), .A2(new_n10847), .B1(new_n2734), .B2(new_n12047), .C(new_n16398), .Y(new_n16399));
  XNOR2x2_ASAP7_75t_L       g16143(.A(\a[29] ), .B(new_n16399), .Y(new_n16400));
  INVx1_ASAP7_75t_L         g16144(.A(new_n16400), .Y(new_n16401));
  A2O1A1Ixp33_ASAP7_75t_L   g16145(.A1(new_n16220), .A2(new_n16217), .B(new_n16250), .C(new_n16371), .Y(new_n16402));
  NOR2xp33_ASAP7_75t_L      g16146(.A(new_n16401), .B(new_n16402), .Y(new_n16403));
  O2A1O1Ixp33_ASAP7_75t_L   g16147(.A1(new_n16373), .A2(new_n16372), .B(new_n16252), .C(new_n16400), .Y(new_n16404));
  AOI22xp33_ASAP7_75t_L     g16148(.A1(new_n3029), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n3258), .Y(new_n16405));
  OAI221xp5_ASAP7_75t_L     g16149(.A1(new_n3024), .A2(new_n9920), .B1(new_n3256), .B2(new_n11152), .C(new_n16405), .Y(new_n16406));
  XNOR2x2_ASAP7_75t_L       g16150(.A(\a[32] ), .B(new_n16406), .Y(new_n16407));
  MAJx2_ASAP7_75t_L         g16151(.A(new_n16363), .B(new_n16365), .C(new_n16369), .Y(new_n16408));
  AND2x2_ASAP7_75t_L        g16152(.A(new_n16407), .B(new_n16408), .Y(new_n16409));
  NOR2xp33_ASAP7_75t_L      g16153(.A(new_n16407), .B(new_n16408), .Y(new_n16410));
  NOR2xp33_ASAP7_75t_L      g16154(.A(new_n16410), .B(new_n16409), .Y(new_n16411));
  AOI22xp33_ASAP7_75t_L     g16155(.A1(new_n3633), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n3858), .Y(new_n16412));
  OAI221xp5_ASAP7_75t_L     g16156(.A1(new_n3853), .A2(new_n8762), .B1(new_n3856), .B2(new_n9331), .C(new_n16412), .Y(new_n16413));
  XNOR2x2_ASAP7_75t_L       g16157(.A(\a[35] ), .B(new_n16413), .Y(new_n16414));
  AOI22xp33_ASAP7_75t_L     g16158(.A1(new_n4283), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n4512), .Y(new_n16415));
  OAI221xp5_ASAP7_75t_L     g16159(.A1(new_n4277), .A2(new_n7900), .B1(new_n4499), .B2(new_n8174), .C(new_n16415), .Y(new_n16416));
  XNOR2x2_ASAP7_75t_L       g16160(.A(\a[38] ), .B(new_n16416), .Y(new_n16417));
  INVx1_ASAP7_75t_L         g16161(.A(new_n16417), .Y(new_n16418));
  AOI22xp33_ASAP7_75t_L     g16162(.A1(new_n6376), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n6648), .Y(new_n16419));
  OAI221xp5_ASAP7_75t_L     g16163(.A1(new_n6646), .A2(new_n5805), .B1(new_n6636), .B2(new_n5835), .C(new_n16419), .Y(new_n16420));
  XNOR2x2_ASAP7_75t_L       g16164(.A(\a[47] ), .B(new_n16420), .Y(new_n16421));
  INVx1_ASAP7_75t_L         g16165(.A(new_n16421), .Y(new_n16422));
  AOI22xp33_ASAP7_75t_L     g16166(.A1(new_n7111), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n7391), .Y(new_n16423));
  OAI221xp5_ASAP7_75t_L     g16167(.A1(new_n8558), .A2(new_n4869), .B1(new_n8237), .B2(new_n5327), .C(new_n16423), .Y(new_n16424));
  XNOR2x2_ASAP7_75t_L       g16168(.A(\a[50] ), .B(new_n16424), .Y(new_n16425));
  AOI22xp33_ASAP7_75t_L     g16169(.A1(new_n8831), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n9115), .Y(new_n16426));
  OAI221xp5_ASAP7_75t_L     g16170(.A1(new_n10343), .A2(new_n3584), .B1(new_n10016), .B2(new_n10137), .C(new_n16426), .Y(new_n16427));
  XNOR2x2_ASAP7_75t_L       g16171(.A(\a[56] ), .B(new_n16427), .Y(new_n16428));
  INVx1_ASAP7_75t_L         g16172(.A(new_n16428), .Y(new_n16429));
  AOI22xp33_ASAP7_75t_L     g16173(.A1(new_n9700), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n10027), .Y(new_n16430));
  OAI221xp5_ASAP7_75t_L     g16174(.A1(new_n10024), .A2(new_n3180), .B1(new_n9696), .B2(new_n11047), .C(new_n16430), .Y(new_n16431));
  XNOR2x2_ASAP7_75t_L       g16175(.A(\a[59] ), .B(new_n16431), .Y(new_n16432));
  INVx1_ASAP7_75t_L         g16176(.A(new_n16432), .Y(new_n16433));
  NOR2xp33_ASAP7_75t_L      g16177(.A(new_n2067), .B(new_n11535), .Y(new_n16434));
  O2A1O1Ixp33_ASAP7_75t_L   g16178(.A1(new_n11247), .A2(new_n11249), .B(\b[26] ), .C(new_n16434), .Y(new_n16435));
  A2O1A1Ixp33_ASAP7_75t_L   g16179(.A1(new_n11533), .A2(\b[25] ), .B(new_n16259), .C(new_n16435), .Y(new_n16436));
  A2O1A1Ixp33_ASAP7_75t_L   g16180(.A1(\b[26] ), .A2(new_n11533), .B(new_n16434), .C(new_n16262), .Y(new_n16437));
  NAND2xp33_ASAP7_75t_L     g16181(.A(new_n16437), .B(new_n16436), .Y(new_n16438));
  NOR2xp33_ASAP7_75t_L      g16182(.A(new_n2688), .B(new_n10630), .Y(new_n16439));
  AOI221xp5_ASAP7_75t_L     g16183(.A1(\b[27] ), .A2(new_n10939), .B1(\b[28] ), .B2(new_n10632), .C(new_n16439), .Y(new_n16440));
  OAI211xp5_ASAP7_75t_L     g16184(.A1(new_n10629), .A2(new_n2695), .B(\a[62] ), .C(new_n16440), .Y(new_n16441));
  O2A1O1Ixp33_ASAP7_75t_L   g16185(.A1(new_n10629), .A2(new_n2695), .B(new_n16440), .C(\a[62] ), .Y(new_n16442));
  INVx1_ASAP7_75t_L         g16186(.A(new_n16442), .Y(new_n16443));
  AND2x2_ASAP7_75t_L        g16187(.A(new_n16441), .B(new_n16443), .Y(new_n16444));
  NOR2xp33_ASAP7_75t_L      g16188(.A(new_n16438), .B(new_n16444), .Y(new_n16445));
  AND3x1_ASAP7_75t_L        g16189(.A(new_n16443), .B(new_n16441), .C(new_n16438), .Y(new_n16446));
  NOR2xp33_ASAP7_75t_L      g16190(.A(new_n16446), .B(new_n16445), .Y(new_n16447));
  INVx1_ASAP7_75t_L         g16191(.A(new_n16447), .Y(new_n16448));
  O2A1O1Ixp33_ASAP7_75t_L   g16192(.A1(new_n16266), .A2(new_n16272), .B(new_n16265), .C(new_n16448), .Y(new_n16449));
  INVx1_ASAP7_75t_L         g16193(.A(new_n16449), .Y(new_n16450));
  NAND3xp33_ASAP7_75t_L     g16194(.A(new_n16448), .B(new_n16274), .C(new_n16265), .Y(new_n16451));
  NAND3xp33_ASAP7_75t_L     g16195(.A(new_n16450), .B(new_n16433), .C(new_n16451), .Y(new_n16452));
  AO21x2_ASAP7_75t_L        g16196(.A1(new_n16450), .A2(new_n16451), .B(new_n16433), .Y(new_n16453));
  AND2x2_ASAP7_75t_L        g16197(.A(new_n16452), .B(new_n16453), .Y(new_n16454));
  INVx1_ASAP7_75t_L         g16198(.A(new_n16454), .Y(new_n16455));
  A2O1A1Ixp33_ASAP7_75t_L   g16199(.A1(new_n16274), .A2(new_n16275), .B(new_n16279), .C(new_n16285), .Y(new_n16456));
  NOR2xp33_ASAP7_75t_L      g16200(.A(new_n16456), .B(new_n16455), .Y(new_n16457));
  O2A1O1Ixp33_ASAP7_75t_L   g16201(.A1(new_n16279), .A2(new_n16276), .B(new_n16285), .C(new_n16454), .Y(new_n16458));
  NOR2xp33_ASAP7_75t_L      g16202(.A(new_n16458), .B(new_n16457), .Y(new_n16459));
  NAND2xp33_ASAP7_75t_L     g16203(.A(new_n16429), .B(new_n16459), .Y(new_n16460));
  INVx1_ASAP7_75t_L         g16204(.A(new_n16460), .Y(new_n16461));
  NOR2xp33_ASAP7_75t_L      g16205(.A(new_n16429), .B(new_n16459), .Y(new_n16462));
  NOR2xp33_ASAP7_75t_L      g16206(.A(new_n16462), .B(new_n16461), .Y(new_n16463));
  NAND3xp33_ASAP7_75t_L     g16207(.A(new_n16463), .B(new_n16297), .C(new_n16288), .Y(new_n16464));
  INVx1_ASAP7_75t_L         g16208(.A(new_n16296), .Y(new_n16465));
  O2A1O1Ixp33_ASAP7_75t_L   g16209(.A1(new_n16289), .A2(new_n16465), .B(new_n16288), .C(new_n16463), .Y(new_n16466));
  INVx1_ASAP7_75t_L         g16210(.A(new_n16466), .Y(new_n16467));
  AOI22xp33_ASAP7_75t_L     g16211(.A1(new_n7960), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n8537), .Y(new_n16468));
  OAI221xp5_ASAP7_75t_L     g16212(.A1(new_n8817), .A2(new_n4424), .B1(new_n7957), .B2(new_n4641), .C(new_n16468), .Y(new_n16469));
  XNOR2x2_ASAP7_75t_L       g16213(.A(\a[53] ), .B(new_n16469), .Y(new_n16470));
  NAND3xp33_ASAP7_75t_L     g16214(.A(new_n16467), .B(new_n16464), .C(new_n16470), .Y(new_n16471));
  AO21x2_ASAP7_75t_L        g16215(.A1(new_n16464), .A2(new_n16467), .B(new_n16470), .Y(new_n16472));
  AND2x2_ASAP7_75t_L        g16216(.A(new_n16471), .B(new_n16472), .Y(new_n16473));
  O2A1O1Ixp33_ASAP7_75t_L   g16217(.A1(new_n16308), .A2(new_n16305), .B(new_n16303), .C(new_n16473), .Y(new_n16474));
  AND3x1_ASAP7_75t_L        g16218(.A(new_n16311), .B(new_n16473), .C(new_n16303), .Y(new_n16475));
  NOR2xp33_ASAP7_75t_L      g16219(.A(new_n16474), .B(new_n16475), .Y(new_n16476));
  XOR2x2_ASAP7_75t_L        g16220(.A(new_n16425), .B(new_n16476), .Y(new_n16477));
  O2A1O1Ixp33_ASAP7_75t_L   g16221(.A1(new_n16315), .A2(new_n16316), .B(new_n16319), .C(new_n16477), .Y(new_n16478));
  INVx1_ASAP7_75t_L         g16222(.A(new_n16478), .Y(new_n16479));
  NAND3xp33_ASAP7_75t_L     g16223(.A(new_n16319), .B(new_n16313), .C(new_n16477), .Y(new_n16480));
  NAND3xp33_ASAP7_75t_L     g16224(.A(new_n16479), .B(new_n16422), .C(new_n16480), .Y(new_n16481));
  INVx1_ASAP7_75t_L         g16225(.A(new_n16481), .Y(new_n16482));
  AOI21xp33_ASAP7_75t_L     g16226(.A1(new_n16479), .A2(new_n16480), .B(new_n16422), .Y(new_n16483));
  NOR2xp33_ASAP7_75t_L      g16227(.A(new_n16483), .B(new_n16482), .Y(new_n16484));
  NAND3xp33_ASAP7_75t_L     g16228(.A(new_n16484), .B(new_n16330), .C(new_n16326), .Y(new_n16485));
  O2A1O1Ixp33_ASAP7_75t_L   g16229(.A1(new_n16324), .A2(new_n16321), .B(new_n16330), .C(new_n16484), .Y(new_n16486));
  INVx1_ASAP7_75t_L         g16230(.A(new_n16486), .Y(new_n16487));
  AOI22xp33_ASAP7_75t_L     g16231(.A1(new_n5624), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n5901), .Y(new_n16488));
  OAI221xp5_ASAP7_75t_L     g16232(.A1(new_n5900), .A2(new_n6568), .B1(new_n5892), .B2(new_n6820), .C(new_n16488), .Y(new_n16489));
  XNOR2x2_ASAP7_75t_L       g16233(.A(\a[44] ), .B(new_n16489), .Y(new_n16490));
  NAND3xp33_ASAP7_75t_L     g16234(.A(new_n16487), .B(new_n16485), .C(new_n16490), .Y(new_n16491));
  INVx1_ASAP7_75t_L         g16235(.A(new_n16491), .Y(new_n16492));
  AOI21xp33_ASAP7_75t_L     g16236(.A1(new_n16487), .A2(new_n16485), .B(new_n16490), .Y(new_n16493));
  NOR2xp33_ASAP7_75t_L      g16237(.A(new_n16493), .B(new_n16492), .Y(new_n16494));
  A2O1A1Ixp33_ASAP7_75t_L   g16238(.A1(new_n16336), .A2(new_n16339), .B(new_n16334), .C(new_n16494), .Y(new_n16495));
  AOI211xp5_ASAP7_75t_L     g16239(.A1(new_n16336), .A2(new_n16339), .B(new_n16334), .C(new_n16494), .Y(new_n16496));
  INVx1_ASAP7_75t_L         g16240(.A(new_n16496), .Y(new_n16497));
  NAND2xp33_ASAP7_75t_L     g16241(.A(new_n16495), .B(new_n16497), .Y(new_n16498));
  AOI22xp33_ASAP7_75t_L     g16242(.A1(new_n4920), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n5167), .Y(new_n16499));
  OAI221xp5_ASAP7_75t_L     g16243(.A1(new_n5154), .A2(new_n7317), .B1(new_n5158), .B2(new_n7602), .C(new_n16499), .Y(new_n16500));
  XNOR2x2_ASAP7_75t_L       g16244(.A(\a[41] ), .B(new_n16500), .Y(new_n16501));
  XNOR2x2_ASAP7_75t_L       g16245(.A(new_n16501), .B(new_n16498), .Y(new_n16502));
  INVx1_ASAP7_75t_L         g16246(.A(new_n16502), .Y(new_n16503));
  NOR2xp33_ASAP7_75t_L      g16247(.A(new_n16344), .B(new_n16351), .Y(new_n16504));
  NAND2xp33_ASAP7_75t_L     g16248(.A(new_n16504), .B(new_n16503), .Y(new_n16505));
  INVx1_ASAP7_75t_L         g16249(.A(new_n16505), .Y(new_n16506));
  INVx1_ASAP7_75t_L         g16250(.A(new_n16351), .Y(new_n16507));
  O2A1O1Ixp33_ASAP7_75t_L   g16251(.A1(new_n16342), .A2(new_n16343), .B(new_n16507), .C(new_n16503), .Y(new_n16508));
  NOR2xp33_ASAP7_75t_L      g16252(.A(new_n16506), .B(new_n16508), .Y(new_n16509));
  NAND2xp33_ASAP7_75t_L     g16253(.A(new_n16418), .B(new_n16509), .Y(new_n16510));
  INVx1_ASAP7_75t_L         g16254(.A(new_n16510), .Y(new_n16511));
  NOR2xp33_ASAP7_75t_L      g16255(.A(new_n16418), .B(new_n16509), .Y(new_n16512));
  NOR2xp33_ASAP7_75t_L      g16256(.A(new_n16512), .B(new_n16511), .Y(new_n16513));
  AOI21xp33_ASAP7_75t_L     g16257(.A1(new_n16358), .A2(new_n16362), .B(new_n16355), .Y(new_n16514));
  AND2x2_ASAP7_75t_L        g16258(.A(new_n16514), .B(new_n16513), .Y(new_n16515));
  INVx1_ASAP7_75t_L         g16259(.A(new_n16362), .Y(new_n16516));
  O2A1O1Ixp33_ASAP7_75t_L   g16260(.A1(new_n16359), .A2(new_n16516), .B(new_n16356), .C(new_n16513), .Y(new_n16517));
  NOR2xp33_ASAP7_75t_L      g16261(.A(new_n16517), .B(new_n16515), .Y(new_n16518));
  XNOR2x2_ASAP7_75t_L       g16262(.A(new_n16414), .B(new_n16518), .Y(new_n16519));
  XNOR2x2_ASAP7_75t_L       g16263(.A(new_n16411), .B(new_n16519), .Y(new_n16520));
  OAI21xp33_ASAP7_75t_L     g16264(.A1(new_n16404), .A2(new_n16403), .B(new_n16520), .Y(new_n16521));
  OR3x1_ASAP7_75t_L         g16265(.A(new_n16403), .B(new_n16404), .C(new_n16520), .Y(new_n16522));
  NAND2xp33_ASAP7_75t_L     g16266(.A(new_n16521), .B(new_n16522), .Y(new_n16523));
  INVx1_ASAP7_75t_L         g16267(.A(new_n16523), .Y(new_n16524));
  INVx1_ASAP7_75t_L         g16268(.A(new_n16243), .Y(new_n16525));
  MAJIxp5_ASAP7_75t_L       g16269(.A(new_n16375), .B(new_n16242), .C(new_n16525), .Y(new_n16526));
  A2O1A1O1Ixp25_ASAP7_75t_L g16270(.A1(new_n2106), .A2(new_n12061), .B(new_n2259), .C(\b[63] ), .D(new_n2100), .Y(new_n16527));
  A2O1A1O1Ixp25_ASAP7_75t_L g16271(.A1(\b[61] ), .A2(new_n11471), .B(\b[62] ), .C(new_n2106), .D(new_n2259), .Y(new_n16528));
  NOR3xp33_ASAP7_75t_L      g16272(.A(new_n16528), .B(new_n11468), .C(\a[26] ), .Y(new_n16529));
  NOR2xp33_ASAP7_75t_L      g16273(.A(new_n16527), .B(new_n16529), .Y(new_n16530));
  INVx1_ASAP7_75t_L         g16274(.A(new_n16530), .Y(new_n16531));
  NAND2xp33_ASAP7_75t_L     g16275(.A(new_n16531), .B(new_n16526), .Y(new_n16532));
  INVx1_ASAP7_75t_L         g16276(.A(new_n16532), .Y(new_n16533));
  NOR2xp33_ASAP7_75t_L      g16277(.A(new_n16531), .B(new_n16526), .Y(new_n16534));
  NOR2xp33_ASAP7_75t_L      g16278(.A(new_n16534), .B(new_n16533), .Y(new_n16535));
  NAND2xp33_ASAP7_75t_L     g16279(.A(new_n16535), .B(new_n16524), .Y(new_n16536));
  OAI21xp33_ASAP7_75t_L     g16280(.A1(new_n16533), .A2(new_n16534), .B(new_n16523), .Y(new_n16537));
  NAND2xp33_ASAP7_75t_L     g16281(.A(new_n16537), .B(new_n16536), .Y(new_n16538));
  XOR2x2_ASAP7_75t_L        g16282(.A(new_n16397), .B(new_n16538), .Y(new_n16539));
  A2O1A1Ixp33_ASAP7_75t_L   g16283(.A1(new_n16393), .A2(new_n16390), .B(new_n16386), .C(new_n16539), .Y(new_n16540));
  INVx1_ASAP7_75t_L         g16284(.A(new_n16540), .Y(new_n16541));
  INVx1_ASAP7_75t_L         g16285(.A(new_n16386), .Y(new_n16542));
  A2O1A1Ixp33_ASAP7_75t_L   g16286(.A1(new_n16234), .A2(new_n16230), .B(new_n16389), .C(new_n16542), .Y(new_n16543));
  NOR2xp33_ASAP7_75t_L      g16287(.A(new_n16539), .B(new_n16543), .Y(new_n16544));
  NOR2xp33_ASAP7_75t_L      g16288(.A(new_n16541), .B(new_n16544), .Y(\f[89] ));
  INVx1_ASAP7_75t_L         g16289(.A(new_n16538), .Y(new_n16546));
  A2O1A1Ixp33_ASAP7_75t_L   g16290(.A1(new_n16384), .A2(new_n16376), .B(new_n16396), .C(new_n16546), .Y(new_n16547));
  INVx1_ASAP7_75t_L         g16291(.A(new_n16547), .Y(new_n16548));
  INVx1_ASAP7_75t_L         g16292(.A(new_n16404), .Y(new_n16549));
  AOI22xp33_ASAP7_75t_L     g16293(.A1(new_n2552), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n2736), .Y(new_n16550));
  A2O1A1Ixp33_ASAP7_75t_L   g16294(.A1(new_n11470), .A2(new_n11473), .B(new_n2734), .C(new_n16550), .Y(new_n16551));
  AOI21xp33_ASAP7_75t_L     g16295(.A1(new_n2553), .A2(\b[62] ), .B(new_n16551), .Y(new_n16552));
  NAND2xp33_ASAP7_75t_L     g16296(.A(\a[29] ), .B(new_n16552), .Y(new_n16553));
  A2O1A1Ixp33_ASAP7_75t_L   g16297(.A1(\b[62] ), .A2(new_n2553), .B(new_n16551), .C(new_n2538), .Y(new_n16554));
  AND2x2_ASAP7_75t_L        g16298(.A(new_n16554), .B(new_n16553), .Y(new_n16555));
  INVx1_ASAP7_75t_L         g16299(.A(new_n16555), .Y(new_n16556));
  O2A1O1Ixp33_ASAP7_75t_L   g16300(.A1(new_n16520), .A2(new_n16403), .B(new_n16549), .C(new_n16556), .Y(new_n16557));
  A2O1A1Ixp33_ASAP7_75t_L   g16301(.A1(new_n16371), .A2(new_n16252), .B(new_n16400), .C(new_n16522), .Y(new_n16558));
  NOR2xp33_ASAP7_75t_L      g16302(.A(new_n16555), .B(new_n16558), .Y(new_n16559));
  OR2x4_ASAP7_75t_L         g16303(.A(new_n16557), .B(new_n16559), .Y(new_n16560));
  A2O1A1Ixp33_ASAP7_75t_L   g16304(.A1(new_n16347), .A2(new_n16350), .B(new_n16344), .C(new_n16502), .Y(new_n16561));
  AOI22xp33_ASAP7_75t_L     g16305(.A1(new_n4283), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n4512), .Y(new_n16562));
  OAI221xp5_ASAP7_75t_L     g16306(.A1(new_n4277), .A2(new_n8165), .B1(new_n4499), .B2(new_n8465), .C(new_n16562), .Y(new_n16563));
  XNOR2x2_ASAP7_75t_L       g16307(.A(\a[38] ), .B(new_n16563), .Y(new_n16564));
  OAI21xp33_ASAP7_75t_L     g16308(.A1(new_n16501), .A2(new_n16498), .B(new_n16497), .Y(new_n16565));
  A2O1A1Ixp33_ASAP7_75t_L   g16309(.A1(new_n16319), .A2(new_n16313), .B(new_n16477), .C(new_n16481), .Y(new_n16566));
  AOI22xp33_ASAP7_75t_L     g16310(.A1(new_n6376), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n6648), .Y(new_n16567));
  OAI221xp5_ASAP7_75t_L     g16311(.A1(new_n6646), .A2(new_n5829), .B1(new_n6636), .B2(new_n6329), .C(new_n16567), .Y(new_n16568));
  XNOR2x2_ASAP7_75t_L       g16312(.A(\a[47] ), .B(new_n16568), .Y(new_n16569));
  INVx1_ASAP7_75t_L         g16313(.A(new_n16569), .Y(new_n16570));
  AOI22xp33_ASAP7_75t_L     g16314(.A1(new_n9700), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n10027), .Y(new_n16571));
  OAI221xp5_ASAP7_75t_L     g16315(.A1(new_n10024), .A2(new_n3207), .B1(new_n9696), .B2(new_n3572), .C(new_n16571), .Y(new_n16572));
  XNOR2x2_ASAP7_75t_L       g16316(.A(\a[59] ), .B(new_n16572), .Y(new_n16573));
  INVx1_ASAP7_75t_L         g16317(.A(new_n16573), .Y(new_n16574));
  A2O1A1Ixp33_ASAP7_75t_L   g16318(.A1(new_n16274), .A2(new_n16265), .B(new_n16448), .C(new_n16452), .Y(new_n16575));
  NOR2xp33_ASAP7_75t_L      g16319(.A(new_n16574), .B(new_n16575), .Y(new_n16576));
  A2O1A1O1Ixp25_ASAP7_75t_L g16320(.A1(new_n16274), .A2(new_n16265), .B(new_n16448), .C(new_n16452), .D(new_n16573), .Y(new_n16577));
  NOR2xp33_ASAP7_75t_L      g16321(.A(new_n16577), .B(new_n16576), .Y(new_n16578));
  NOR2xp33_ASAP7_75t_L      g16322(.A(new_n2348), .B(new_n11535), .Y(new_n16579));
  A2O1A1Ixp33_ASAP7_75t_L   g16323(.A1(new_n11533), .A2(\b[27] ), .B(new_n16579), .C(new_n2100), .Y(new_n16580));
  INVx1_ASAP7_75t_L         g16324(.A(new_n16580), .Y(new_n16581));
  O2A1O1Ixp33_ASAP7_75t_L   g16325(.A1(new_n11247), .A2(new_n11249), .B(\b[27] ), .C(new_n16579), .Y(new_n16582));
  NAND2xp33_ASAP7_75t_L     g16326(.A(\a[26] ), .B(new_n16582), .Y(new_n16583));
  INVx1_ASAP7_75t_L         g16327(.A(new_n16583), .Y(new_n16584));
  NOR2xp33_ASAP7_75t_L      g16328(.A(new_n16581), .B(new_n16584), .Y(new_n16585));
  A2O1A1Ixp33_ASAP7_75t_L   g16329(.A1(new_n11533), .A2(\b[26] ), .B(new_n16434), .C(new_n16585), .Y(new_n16586));
  OAI21xp33_ASAP7_75t_L     g16330(.A1(new_n16581), .A2(new_n16584), .B(new_n16435), .Y(new_n16587));
  NAND2xp33_ASAP7_75t_L     g16331(.A(new_n16587), .B(new_n16586), .Y(new_n16588));
  A2O1A1O1Ixp25_ASAP7_75t_L g16332(.A1(new_n16441), .A2(new_n16443), .B(new_n16438), .C(new_n16436), .D(new_n16588), .Y(new_n16589));
  INVx1_ASAP7_75t_L         g16333(.A(new_n16589), .Y(new_n16590));
  OAI211xp5_ASAP7_75t_L     g16334(.A1(new_n16438), .A2(new_n16444), .B(new_n16436), .C(new_n16588), .Y(new_n16591));
  AND2x2_ASAP7_75t_L        g16335(.A(new_n16590), .B(new_n16591), .Y(new_n16592));
  AOI22xp33_ASAP7_75t_L     g16336(.A1(\b[28] ), .A2(new_n10939), .B1(\b[30] ), .B2(new_n10938), .Y(new_n16593));
  OAI221xp5_ASAP7_75t_L     g16337(.A1(new_n10937), .A2(new_n2688), .B1(new_n10629), .B2(new_n2990), .C(new_n16593), .Y(new_n16594));
  XNOR2x2_ASAP7_75t_L       g16338(.A(\a[62] ), .B(new_n16594), .Y(new_n16595));
  NAND2xp33_ASAP7_75t_L     g16339(.A(new_n16595), .B(new_n16592), .Y(new_n16596));
  AO21x2_ASAP7_75t_L        g16340(.A1(new_n16590), .A2(new_n16591), .B(new_n16595), .Y(new_n16597));
  AND2x2_ASAP7_75t_L        g16341(.A(new_n16597), .B(new_n16596), .Y(new_n16598));
  XOR2x2_ASAP7_75t_L        g16342(.A(new_n16578), .B(new_n16598), .Y(new_n16599));
  NAND2xp33_ASAP7_75t_L     g16343(.A(\b[34] ), .B(new_n9115), .Y(new_n16600));
  OAI221xp5_ASAP7_75t_L     g16344(.A1(new_n9113), .A2(new_n4216), .B1(new_n10016), .B2(new_n4223), .C(new_n16600), .Y(new_n16601));
  AOI21xp33_ASAP7_75t_L     g16345(.A1(new_n8835), .A2(\b[35] ), .B(new_n16601), .Y(new_n16602));
  NAND2xp33_ASAP7_75t_L     g16346(.A(\a[56] ), .B(new_n16602), .Y(new_n16603));
  A2O1A1Ixp33_ASAP7_75t_L   g16347(.A1(\b[35] ), .A2(new_n8835), .B(new_n16601), .C(new_n8826), .Y(new_n16604));
  AND2x2_ASAP7_75t_L        g16348(.A(new_n16604), .B(new_n16603), .Y(new_n16605));
  XNOR2x2_ASAP7_75t_L       g16349(.A(new_n16605), .B(new_n16599), .Y(new_n16606));
  INVx1_ASAP7_75t_L         g16350(.A(new_n16606), .Y(new_n16607));
  NOR3xp33_ASAP7_75t_L      g16351(.A(new_n16607), .B(new_n16461), .C(new_n16457), .Y(new_n16608));
  O2A1O1Ixp33_ASAP7_75t_L   g16352(.A1(new_n16455), .A2(new_n16456), .B(new_n16460), .C(new_n16606), .Y(new_n16609));
  NOR2xp33_ASAP7_75t_L      g16353(.A(new_n16609), .B(new_n16608), .Y(new_n16610));
  AOI22xp33_ASAP7_75t_L     g16354(.A1(new_n7960), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n8537), .Y(new_n16611));
  OAI221xp5_ASAP7_75t_L     g16355(.A1(new_n8817), .A2(new_n4632), .B1(new_n7957), .B2(new_n4858), .C(new_n16611), .Y(new_n16612));
  XNOR2x2_ASAP7_75t_L       g16356(.A(\a[53] ), .B(new_n16612), .Y(new_n16613));
  INVx1_ASAP7_75t_L         g16357(.A(new_n16613), .Y(new_n16614));
  XNOR2x2_ASAP7_75t_L       g16358(.A(new_n16614), .B(new_n16610), .Y(new_n16615));
  A2O1A1Ixp33_ASAP7_75t_L   g16359(.A1(new_n16470), .A2(new_n16464), .B(new_n16466), .C(new_n16615), .Y(new_n16616));
  A2O1A1Ixp33_ASAP7_75t_L   g16360(.A1(new_n16297), .A2(new_n16288), .B(new_n16463), .C(new_n16471), .Y(new_n16617));
  NOR2xp33_ASAP7_75t_L      g16361(.A(new_n16617), .B(new_n16615), .Y(new_n16618));
  INVx1_ASAP7_75t_L         g16362(.A(new_n16618), .Y(new_n16619));
  NAND2xp33_ASAP7_75t_L     g16363(.A(new_n16616), .B(new_n16619), .Y(new_n16620));
  AOI22xp33_ASAP7_75t_L     g16364(.A1(new_n7111), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n7391), .Y(new_n16621));
  OAI221xp5_ASAP7_75t_L     g16365(.A1(new_n8558), .A2(new_n5321), .B1(new_n8237), .B2(new_n5346), .C(new_n16621), .Y(new_n16622));
  XNOR2x2_ASAP7_75t_L       g16366(.A(\a[50] ), .B(new_n16622), .Y(new_n16623));
  XNOR2x2_ASAP7_75t_L       g16367(.A(new_n16623), .B(new_n16620), .Y(new_n16624));
  AOI211xp5_ASAP7_75t_L     g16368(.A1(new_n16476), .A2(new_n16425), .B(new_n16475), .C(new_n16624), .Y(new_n16625));
  INVx1_ASAP7_75t_L         g16369(.A(new_n16625), .Y(new_n16626));
  A2O1A1Ixp33_ASAP7_75t_L   g16370(.A1(new_n16476), .A2(new_n16425), .B(new_n16475), .C(new_n16624), .Y(new_n16627));
  AND2x2_ASAP7_75t_L        g16371(.A(new_n16627), .B(new_n16626), .Y(new_n16628));
  NAND2xp33_ASAP7_75t_L     g16372(.A(new_n16570), .B(new_n16628), .Y(new_n16629));
  NOR2xp33_ASAP7_75t_L      g16373(.A(new_n16570), .B(new_n16628), .Y(new_n16630));
  INVx1_ASAP7_75t_L         g16374(.A(new_n16630), .Y(new_n16631));
  AO21x2_ASAP7_75t_L        g16375(.A1(new_n16631), .A2(new_n16629), .B(new_n16566), .Y(new_n16632));
  NAND3xp33_ASAP7_75t_L     g16376(.A(new_n16566), .B(new_n16629), .C(new_n16631), .Y(new_n16633));
  NAND2xp33_ASAP7_75t_L     g16377(.A(new_n16633), .B(new_n16632), .Y(new_n16634));
  AOI22xp33_ASAP7_75t_L     g16378(.A1(new_n5624), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n5901), .Y(new_n16635));
  OAI221xp5_ASAP7_75t_L     g16379(.A1(new_n5900), .A2(new_n6812), .B1(new_n5892), .B2(new_n6837), .C(new_n16635), .Y(new_n16636));
  XNOR2x2_ASAP7_75t_L       g16380(.A(\a[44] ), .B(new_n16636), .Y(new_n16637));
  XNOR2x2_ASAP7_75t_L       g16381(.A(new_n16637), .B(new_n16634), .Y(new_n16638));
  A2O1A1Ixp33_ASAP7_75t_L   g16382(.A1(new_n16490), .A2(new_n16485), .B(new_n16486), .C(new_n16638), .Y(new_n16639));
  OR3x1_ASAP7_75t_L         g16383(.A(new_n16492), .B(new_n16638), .C(new_n16486), .Y(new_n16640));
  NAND2xp33_ASAP7_75t_L     g16384(.A(new_n16639), .B(new_n16640), .Y(new_n16641));
  AOI22xp33_ASAP7_75t_L     g16385(.A1(new_n4920), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n5167), .Y(new_n16642));
  OAI221xp5_ASAP7_75t_L     g16386(.A1(new_n5154), .A2(new_n7593), .B1(new_n5158), .B2(new_n7623), .C(new_n16642), .Y(new_n16643));
  XNOR2x2_ASAP7_75t_L       g16387(.A(\a[41] ), .B(new_n16643), .Y(new_n16644));
  XNOR2x2_ASAP7_75t_L       g16388(.A(new_n16644), .B(new_n16641), .Y(new_n16645));
  XNOR2x2_ASAP7_75t_L       g16389(.A(new_n16645), .B(new_n16565), .Y(new_n16646));
  INVx1_ASAP7_75t_L         g16390(.A(new_n16646), .Y(new_n16647));
  NAND2xp33_ASAP7_75t_L     g16391(.A(new_n16564), .B(new_n16647), .Y(new_n16648));
  INVx1_ASAP7_75t_L         g16392(.A(new_n16564), .Y(new_n16649));
  NAND2xp33_ASAP7_75t_L     g16393(.A(new_n16649), .B(new_n16646), .Y(new_n16650));
  NAND2xp33_ASAP7_75t_L     g16394(.A(new_n16650), .B(new_n16648), .Y(new_n16651));
  INVx1_ASAP7_75t_L         g16395(.A(new_n16651), .Y(new_n16652));
  A2O1A1Ixp33_ASAP7_75t_L   g16396(.A1(new_n16561), .A2(new_n16418), .B(new_n16506), .C(new_n16652), .Y(new_n16653));
  NAND3xp33_ASAP7_75t_L     g16397(.A(new_n16510), .B(new_n16505), .C(new_n16651), .Y(new_n16654));
  NAND2xp33_ASAP7_75t_L     g16398(.A(new_n16654), .B(new_n16653), .Y(new_n16655));
  AOI22xp33_ASAP7_75t_L     g16399(.A1(new_n3633), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n3858), .Y(new_n16656));
  OAI221xp5_ASAP7_75t_L     g16400(.A1(new_n3853), .A2(new_n9323), .B1(new_n3856), .B2(new_n9627), .C(new_n16656), .Y(new_n16657));
  XNOR2x2_ASAP7_75t_L       g16401(.A(\a[35] ), .B(new_n16657), .Y(new_n16658));
  INVx1_ASAP7_75t_L         g16402(.A(new_n16658), .Y(new_n16659));
  XNOR2x2_ASAP7_75t_L       g16403(.A(new_n16659), .B(new_n16655), .Y(new_n16660));
  INVx1_ASAP7_75t_L         g16404(.A(new_n16660), .Y(new_n16661));
  A2O1A1Ixp33_ASAP7_75t_L   g16405(.A1(new_n16518), .A2(new_n16414), .B(new_n16517), .C(new_n16661), .Y(new_n16662));
  AOI21xp33_ASAP7_75t_L     g16406(.A1(new_n16518), .A2(new_n16414), .B(new_n16517), .Y(new_n16663));
  NAND2xp33_ASAP7_75t_L     g16407(.A(new_n16660), .B(new_n16663), .Y(new_n16664));
  NAND2xp33_ASAP7_75t_L     g16408(.A(new_n16662), .B(new_n16664), .Y(new_n16665));
  INVx1_ASAP7_75t_L         g16409(.A(new_n16665), .Y(new_n16666));
  NAND2xp33_ASAP7_75t_L     g16410(.A(new_n16407), .B(new_n16408), .Y(new_n16667));
  AOI22xp33_ASAP7_75t_L     g16411(.A1(new_n3029), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n3258), .Y(new_n16668));
  OAI221xp5_ASAP7_75t_L     g16412(.A1(new_n3024), .A2(new_n9947), .B1(new_n3256), .B2(new_n11446), .C(new_n16668), .Y(new_n16669));
  XNOR2x2_ASAP7_75t_L       g16413(.A(\a[32] ), .B(new_n16669), .Y(new_n16670));
  INVx1_ASAP7_75t_L         g16414(.A(new_n16670), .Y(new_n16671));
  O2A1O1Ixp33_ASAP7_75t_L   g16415(.A1(new_n16410), .A2(new_n16519), .B(new_n16667), .C(new_n16671), .Y(new_n16672));
  INVx1_ASAP7_75t_L         g16416(.A(new_n16672), .Y(new_n16673));
  OAI211xp5_ASAP7_75t_L     g16417(.A1(new_n16410), .A2(new_n16519), .B(new_n16667), .C(new_n16671), .Y(new_n16674));
  AND2x2_ASAP7_75t_L        g16418(.A(new_n16674), .B(new_n16673), .Y(new_n16675));
  INVx1_ASAP7_75t_L         g16419(.A(new_n16675), .Y(new_n16676));
  NAND2xp33_ASAP7_75t_L     g16420(.A(new_n16666), .B(new_n16676), .Y(new_n16677));
  NAND2xp33_ASAP7_75t_L     g16421(.A(new_n16665), .B(new_n16675), .Y(new_n16678));
  AND2x2_ASAP7_75t_L        g16422(.A(new_n16678), .B(new_n16677), .Y(new_n16679));
  INVx1_ASAP7_75t_L         g16423(.A(new_n16679), .Y(new_n16680));
  NAND2xp33_ASAP7_75t_L     g16424(.A(new_n16680), .B(new_n16560), .Y(new_n16681));
  OR3x1_ASAP7_75t_L         g16425(.A(new_n16680), .B(new_n16557), .C(new_n16559), .Y(new_n16682));
  NAND2xp33_ASAP7_75t_L     g16426(.A(new_n16682), .B(new_n16681), .Y(new_n16683));
  AND3x1_ASAP7_75t_L        g16427(.A(new_n16683), .B(new_n16536), .C(new_n16532), .Y(new_n16684));
  O2A1O1Ixp33_ASAP7_75t_L   g16428(.A1(new_n16523), .A2(new_n16534), .B(new_n16532), .C(new_n16683), .Y(new_n16685));
  NOR2xp33_ASAP7_75t_L      g16429(.A(new_n16685), .B(new_n16684), .Y(new_n16686));
  A2O1A1Ixp33_ASAP7_75t_L   g16430(.A1(new_n16543), .A2(new_n16539), .B(new_n16548), .C(new_n16686), .Y(new_n16687));
  INVx1_ASAP7_75t_L         g16431(.A(new_n16687), .Y(new_n16688));
  AND2x2_ASAP7_75t_L        g16432(.A(new_n16397), .B(new_n16538), .Y(new_n16689));
  A2O1A1Ixp33_ASAP7_75t_L   g16433(.A1(new_n16391), .A2(new_n16542), .B(new_n16689), .C(new_n16547), .Y(new_n16690));
  NOR2xp33_ASAP7_75t_L      g16434(.A(new_n16686), .B(new_n16690), .Y(new_n16691));
  NOR2xp33_ASAP7_75t_L      g16435(.A(new_n16691), .B(new_n16688), .Y(\f[90] ));
  O2A1O1Ixp33_ASAP7_75t_L   g16436(.A1(new_n16520), .A2(new_n16403), .B(new_n16549), .C(new_n16555), .Y(new_n16693));
  O2A1O1Ixp33_ASAP7_75t_L   g16437(.A1(new_n16557), .A2(new_n16559), .B(new_n16680), .C(new_n16693), .Y(new_n16694));
  NOR2xp33_ASAP7_75t_L      g16438(.A(new_n11172), .B(new_n2747), .Y(new_n16695));
  AOI221xp5_ASAP7_75t_L     g16439(.A1(\b[63] ), .A2(new_n2553), .B1(new_n2544), .B2(new_n12322), .C(new_n16695), .Y(new_n16696));
  XNOR2x2_ASAP7_75t_L       g16440(.A(new_n2538), .B(new_n16696), .Y(new_n16697));
  A2O1A1Ixp33_ASAP7_75t_L   g16441(.A1(new_n16662), .A2(new_n16664), .B(new_n16676), .C(new_n16673), .Y(new_n16698));
  NOR2xp33_ASAP7_75t_L      g16442(.A(new_n16697), .B(new_n16698), .Y(new_n16699));
  INVx1_ASAP7_75t_L         g16443(.A(new_n16699), .Y(new_n16700));
  A2O1A1Ixp33_ASAP7_75t_L   g16444(.A1(new_n16674), .A2(new_n16665), .B(new_n16672), .C(new_n16697), .Y(new_n16701));
  AND2x2_ASAP7_75t_L        g16445(.A(new_n16701), .B(new_n16700), .Y(new_n16702));
  AOI22xp33_ASAP7_75t_L     g16446(.A1(new_n3029), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n3258), .Y(new_n16703));
  OAI221xp5_ASAP7_75t_L     g16447(.A1(new_n3024), .A2(new_n10250), .B1(new_n3256), .B2(new_n10855), .C(new_n16703), .Y(new_n16704));
  XNOR2x2_ASAP7_75t_L       g16448(.A(\a[32] ), .B(new_n16704), .Y(new_n16705));
  NOR2xp33_ASAP7_75t_L      g16449(.A(new_n16658), .B(new_n16655), .Y(new_n16706));
  AOI21xp33_ASAP7_75t_L     g16450(.A1(new_n16663), .A2(new_n16660), .B(new_n16706), .Y(new_n16707));
  NAND2xp33_ASAP7_75t_L     g16451(.A(new_n16705), .B(new_n16707), .Y(new_n16708));
  O2A1O1Ixp33_ASAP7_75t_L   g16452(.A1(new_n16655), .A2(new_n16658), .B(new_n16664), .C(new_n16705), .Y(new_n16709));
  INVx1_ASAP7_75t_L         g16453(.A(new_n16709), .Y(new_n16710));
  AOI22xp33_ASAP7_75t_L     g16454(.A1(new_n7960), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n8537), .Y(new_n16711));
  OAI221xp5_ASAP7_75t_L     g16455(.A1(new_n8817), .A2(new_n4848), .B1(new_n7957), .B2(new_n11686), .C(new_n16711), .Y(new_n16712));
  XNOR2x2_ASAP7_75t_L       g16456(.A(\a[53] ), .B(new_n16712), .Y(new_n16713));
  INVx1_ASAP7_75t_L         g16457(.A(new_n16713), .Y(new_n16714));
  INVx1_ASAP7_75t_L         g16458(.A(new_n16609), .Y(new_n16715));
  AOI22xp33_ASAP7_75t_L     g16459(.A1(new_n8831), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n9115), .Y(new_n16716));
  OAI221xp5_ASAP7_75t_L     g16460(.A1(new_n10343), .A2(new_n4216), .B1(new_n10016), .B2(new_n4431), .C(new_n16716), .Y(new_n16717));
  XNOR2x2_ASAP7_75t_L       g16461(.A(\a[56] ), .B(new_n16717), .Y(new_n16718));
  A2O1A1Ixp33_ASAP7_75t_L   g16462(.A1(new_n16451), .A2(new_n16433), .B(new_n16449), .C(new_n16574), .Y(new_n16719));
  NOR2xp33_ASAP7_75t_L      g16463(.A(new_n2497), .B(new_n11535), .Y(new_n16720));
  A2O1A1O1Ixp25_ASAP7_75t_L g16464(.A1(new_n11533), .A2(\b[26] ), .B(new_n16434), .C(new_n16583), .D(new_n16581), .Y(new_n16721));
  A2O1A1Ixp33_ASAP7_75t_L   g16465(.A1(new_n11533), .A2(\b[28] ), .B(new_n16720), .C(new_n16721), .Y(new_n16722));
  O2A1O1Ixp33_ASAP7_75t_L   g16466(.A1(new_n11247), .A2(new_n11249), .B(\b[28] ), .C(new_n16720), .Y(new_n16723));
  INVx1_ASAP7_75t_L         g16467(.A(new_n16723), .Y(new_n16724));
  O2A1O1Ixp33_ASAP7_75t_L   g16468(.A1(new_n16435), .A2(new_n16584), .B(new_n16580), .C(new_n16724), .Y(new_n16725));
  INVx1_ASAP7_75t_L         g16469(.A(new_n16725), .Y(new_n16726));
  NAND2xp33_ASAP7_75t_L     g16470(.A(new_n16722), .B(new_n16726), .Y(new_n16727));
  NAND2xp33_ASAP7_75t_L     g16471(.A(\b[29] ), .B(new_n10939), .Y(new_n16728));
  OAI221xp5_ASAP7_75t_L     g16472(.A1(new_n10630), .A2(new_n3180), .B1(new_n10629), .B2(new_n3187), .C(new_n16728), .Y(new_n16729));
  AOI21xp33_ASAP7_75t_L     g16473(.A1(new_n10632), .A2(\b[30] ), .B(new_n16729), .Y(new_n16730));
  NAND2xp33_ASAP7_75t_L     g16474(.A(\a[62] ), .B(new_n16730), .Y(new_n16731));
  A2O1A1Ixp33_ASAP7_75t_L   g16475(.A1(\b[30] ), .A2(new_n10632), .B(new_n16729), .C(new_n10622), .Y(new_n16732));
  AND2x2_ASAP7_75t_L        g16476(.A(new_n16732), .B(new_n16731), .Y(new_n16733));
  NAND2xp33_ASAP7_75t_L     g16477(.A(new_n16727), .B(new_n16733), .Y(new_n16734));
  NOR2xp33_ASAP7_75t_L      g16478(.A(new_n16727), .B(new_n16733), .Y(new_n16735));
  INVx1_ASAP7_75t_L         g16479(.A(new_n16735), .Y(new_n16736));
  AND2x2_ASAP7_75t_L        g16480(.A(new_n16734), .B(new_n16736), .Y(new_n16737));
  A2O1A1Ixp33_ASAP7_75t_L   g16481(.A1(new_n16443), .A2(new_n16441), .B(new_n16438), .C(new_n16436), .Y(new_n16738));
  A2O1A1Ixp33_ASAP7_75t_L   g16482(.A1(new_n16586), .A2(new_n16587), .B(new_n16738), .C(new_n16596), .Y(new_n16739));
  INVx1_ASAP7_75t_L         g16483(.A(new_n16739), .Y(new_n16740));
  NAND2xp33_ASAP7_75t_L     g16484(.A(new_n16740), .B(new_n16737), .Y(new_n16741));
  A2O1A1O1Ixp25_ASAP7_75t_L g16485(.A1(new_n16586), .A2(new_n16587), .B(new_n16738), .C(new_n16596), .D(new_n16737), .Y(new_n16742));
  INVx1_ASAP7_75t_L         g16486(.A(new_n16742), .Y(new_n16743));
  AOI22xp33_ASAP7_75t_L     g16487(.A1(new_n9700), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n10027), .Y(new_n16744));
  OAI221xp5_ASAP7_75t_L     g16488(.A1(new_n10024), .A2(new_n3565), .B1(new_n9696), .B2(new_n3591), .C(new_n16744), .Y(new_n16745));
  XNOR2x2_ASAP7_75t_L       g16489(.A(\a[59] ), .B(new_n16745), .Y(new_n16746));
  NAND3xp33_ASAP7_75t_L     g16490(.A(new_n16743), .B(new_n16741), .C(new_n16746), .Y(new_n16747));
  AO21x2_ASAP7_75t_L        g16491(.A1(new_n16741), .A2(new_n16743), .B(new_n16746), .Y(new_n16748));
  AND2x2_ASAP7_75t_L        g16492(.A(new_n16747), .B(new_n16748), .Y(new_n16749));
  O2A1O1Ixp33_ASAP7_75t_L   g16493(.A1(new_n16576), .A2(new_n16598), .B(new_n16719), .C(new_n16749), .Y(new_n16750));
  INVx1_ASAP7_75t_L         g16494(.A(new_n16749), .Y(new_n16751));
  A2O1A1Ixp33_ASAP7_75t_L   g16495(.A1(new_n16596), .A2(new_n16597), .B(new_n16576), .C(new_n16719), .Y(new_n16752));
  NOR2xp33_ASAP7_75t_L      g16496(.A(new_n16752), .B(new_n16751), .Y(new_n16753));
  NOR2xp33_ASAP7_75t_L      g16497(.A(new_n16750), .B(new_n16753), .Y(new_n16754));
  NAND2xp33_ASAP7_75t_L     g16498(.A(new_n16718), .B(new_n16754), .Y(new_n16755));
  INVx1_ASAP7_75t_L         g16499(.A(new_n16718), .Y(new_n16756));
  OAI21xp33_ASAP7_75t_L     g16500(.A1(new_n16750), .A2(new_n16753), .B(new_n16756), .Y(new_n16757));
  AND2x2_ASAP7_75t_L        g16501(.A(new_n16757), .B(new_n16755), .Y(new_n16758));
  INVx1_ASAP7_75t_L         g16502(.A(new_n16758), .Y(new_n16759));
  O2A1O1Ixp33_ASAP7_75t_L   g16503(.A1(new_n16599), .A2(new_n16605), .B(new_n16715), .C(new_n16759), .Y(new_n16760));
  A2O1A1Ixp33_ASAP7_75t_L   g16504(.A1(new_n16603), .A2(new_n16604), .B(new_n16599), .C(new_n16715), .Y(new_n16761));
  NOR2xp33_ASAP7_75t_L      g16505(.A(new_n16761), .B(new_n16758), .Y(new_n16762));
  NOR2xp33_ASAP7_75t_L      g16506(.A(new_n16762), .B(new_n16760), .Y(new_n16763));
  XNOR2x2_ASAP7_75t_L       g16507(.A(new_n16714), .B(new_n16763), .Y(new_n16764));
  A2O1A1Ixp33_ASAP7_75t_L   g16508(.A1(new_n16614), .A2(new_n16610), .B(new_n16618), .C(new_n16764), .Y(new_n16765));
  AOI211xp5_ASAP7_75t_L     g16509(.A1(new_n16610), .A2(new_n16614), .B(new_n16618), .C(new_n16764), .Y(new_n16766));
  INVx1_ASAP7_75t_L         g16510(.A(new_n16766), .Y(new_n16767));
  NAND2xp33_ASAP7_75t_L     g16511(.A(new_n16765), .B(new_n16767), .Y(new_n16768));
  AOI22xp33_ASAP7_75t_L     g16512(.A1(new_n7111), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n7391), .Y(new_n16769));
  OAI221xp5_ASAP7_75t_L     g16513(.A1(new_n8558), .A2(new_n5338), .B1(new_n8237), .B2(new_n6338), .C(new_n16769), .Y(new_n16770));
  XNOR2x2_ASAP7_75t_L       g16514(.A(new_n7106), .B(new_n16770), .Y(new_n16771));
  NOR2xp33_ASAP7_75t_L      g16515(.A(new_n16771), .B(new_n16768), .Y(new_n16772));
  AND2x2_ASAP7_75t_L        g16516(.A(new_n16771), .B(new_n16768), .Y(new_n16773));
  NOR2xp33_ASAP7_75t_L      g16517(.A(new_n16772), .B(new_n16773), .Y(new_n16774));
  INVx1_ASAP7_75t_L         g16518(.A(new_n16774), .Y(new_n16775));
  OAI21xp33_ASAP7_75t_L     g16519(.A1(new_n16620), .A2(new_n16623), .B(new_n16626), .Y(new_n16776));
  NOR2xp33_ASAP7_75t_L      g16520(.A(new_n16776), .B(new_n16775), .Y(new_n16777));
  O2A1O1Ixp33_ASAP7_75t_L   g16521(.A1(new_n16620), .A2(new_n16623), .B(new_n16626), .C(new_n16774), .Y(new_n16778));
  NOR2xp33_ASAP7_75t_L      g16522(.A(new_n16778), .B(new_n16777), .Y(new_n16779));
  INVx1_ASAP7_75t_L         g16523(.A(new_n16779), .Y(new_n16780));
  AOI22xp33_ASAP7_75t_L     g16524(.A1(new_n6376), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n6648), .Y(new_n16781));
  OAI221xp5_ASAP7_75t_L     g16525(.A1(new_n6646), .A2(new_n6321), .B1(new_n6636), .B2(new_n6573), .C(new_n16781), .Y(new_n16782));
  XNOR2x2_ASAP7_75t_L       g16526(.A(\a[47] ), .B(new_n16782), .Y(new_n16783));
  INVx1_ASAP7_75t_L         g16527(.A(new_n16783), .Y(new_n16784));
  NOR2xp33_ASAP7_75t_L      g16528(.A(new_n16784), .B(new_n16780), .Y(new_n16785));
  INVx1_ASAP7_75t_L         g16529(.A(new_n16785), .Y(new_n16786));
  NAND2xp33_ASAP7_75t_L     g16530(.A(new_n16784), .B(new_n16780), .Y(new_n16787));
  AND2x2_ASAP7_75t_L        g16531(.A(new_n16787), .B(new_n16786), .Y(new_n16788));
  INVx1_ASAP7_75t_L         g16532(.A(new_n16788), .Y(new_n16789));
  A2O1A1Ixp33_ASAP7_75t_L   g16533(.A1(new_n16481), .A2(new_n16479), .B(new_n16630), .C(new_n16629), .Y(new_n16790));
  NOR2xp33_ASAP7_75t_L      g16534(.A(new_n16790), .B(new_n16789), .Y(new_n16791));
  A2O1A1O1Ixp25_ASAP7_75t_L g16535(.A1(new_n16481), .A2(new_n16479), .B(new_n16630), .C(new_n16629), .D(new_n16788), .Y(new_n16792));
  NOR2xp33_ASAP7_75t_L      g16536(.A(new_n16792), .B(new_n16791), .Y(new_n16793));
  AOI22xp33_ASAP7_75t_L     g16537(.A1(new_n5624), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n5901), .Y(new_n16794));
  OAI221xp5_ASAP7_75t_L     g16538(.A1(new_n5900), .A2(new_n6830), .B1(new_n5892), .B2(new_n7323), .C(new_n16794), .Y(new_n16795));
  XNOR2x2_ASAP7_75t_L       g16539(.A(\a[44] ), .B(new_n16795), .Y(new_n16796));
  NAND2xp33_ASAP7_75t_L     g16540(.A(new_n16796), .B(new_n16793), .Y(new_n16797));
  INVx1_ASAP7_75t_L         g16541(.A(new_n16796), .Y(new_n16798));
  OAI21xp33_ASAP7_75t_L     g16542(.A1(new_n16792), .A2(new_n16791), .B(new_n16798), .Y(new_n16799));
  AND2x2_ASAP7_75t_L        g16543(.A(new_n16799), .B(new_n16797), .Y(new_n16800));
  OA211x2_ASAP7_75t_L       g16544(.A1(new_n16637), .A2(new_n16634), .B(new_n16800), .C(new_n16640), .Y(new_n16801));
  O2A1O1Ixp33_ASAP7_75t_L   g16545(.A1(new_n16634), .A2(new_n16637), .B(new_n16640), .C(new_n16800), .Y(new_n16802));
  NOR2xp33_ASAP7_75t_L      g16546(.A(new_n16802), .B(new_n16801), .Y(new_n16803));
  AOI22xp33_ASAP7_75t_L     g16547(.A1(new_n4920), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n5167), .Y(new_n16804));
  OAI221xp5_ASAP7_75t_L     g16548(.A1(new_n5154), .A2(new_n7616), .B1(new_n5158), .B2(new_n7906), .C(new_n16804), .Y(new_n16805));
  XNOR2x2_ASAP7_75t_L       g16549(.A(\a[41] ), .B(new_n16805), .Y(new_n16806));
  XNOR2x2_ASAP7_75t_L       g16550(.A(new_n16806), .B(new_n16803), .Y(new_n16807));
  NOR2xp33_ASAP7_75t_L      g16551(.A(new_n16644), .B(new_n16641), .Y(new_n16808));
  O2A1O1Ixp33_ASAP7_75t_L   g16552(.A1(new_n16501), .A2(new_n16498), .B(new_n16497), .C(new_n16645), .Y(new_n16809));
  NOR2xp33_ASAP7_75t_L      g16553(.A(new_n16808), .B(new_n16809), .Y(new_n16810));
  INVx1_ASAP7_75t_L         g16554(.A(new_n16810), .Y(new_n16811));
  XNOR2x2_ASAP7_75t_L       g16555(.A(new_n16811), .B(new_n16807), .Y(new_n16812));
  AOI22xp33_ASAP7_75t_L     g16556(.A1(new_n4283), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n4512), .Y(new_n16813));
  OAI221xp5_ASAP7_75t_L     g16557(.A1(new_n4277), .A2(new_n8458), .B1(new_n4499), .B2(new_n8768), .C(new_n16813), .Y(new_n16814));
  XNOR2x2_ASAP7_75t_L       g16558(.A(\a[38] ), .B(new_n16814), .Y(new_n16815));
  XNOR2x2_ASAP7_75t_L       g16559(.A(new_n16815), .B(new_n16812), .Y(new_n16816));
  O2A1O1Ixp33_ASAP7_75t_L   g16560(.A1(new_n16564), .A2(new_n16647), .B(new_n16653), .C(new_n16816), .Y(new_n16817));
  A2O1A1Ixp33_ASAP7_75t_L   g16561(.A1(new_n16510), .A2(new_n16505), .B(new_n16651), .C(new_n16650), .Y(new_n16818));
  INVx1_ASAP7_75t_L         g16562(.A(new_n16816), .Y(new_n16819));
  NOR2xp33_ASAP7_75t_L      g16563(.A(new_n16818), .B(new_n16819), .Y(new_n16820));
  NOR2xp33_ASAP7_75t_L      g16564(.A(new_n16817), .B(new_n16820), .Y(new_n16821));
  AOI22xp33_ASAP7_75t_L     g16565(.A1(new_n3633), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n3858), .Y(new_n16822));
  OAI221xp5_ASAP7_75t_L     g16566(.A1(new_n3853), .A2(new_n9620), .B1(new_n3856), .B2(new_n9925), .C(new_n16822), .Y(new_n16823));
  XNOR2x2_ASAP7_75t_L       g16567(.A(\a[35] ), .B(new_n16823), .Y(new_n16824));
  XNOR2x2_ASAP7_75t_L       g16568(.A(new_n16824), .B(new_n16821), .Y(new_n16825));
  NAND3xp33_ASAP7_75t_L     g16569(.A(new_n16710), .B(new_n16825), .C(new_n16708), .Y(new_n16826));
  AO21x2_ASAP7_75t_L        g16570(.A1(new_n16708), .A2(new_n16710), .B(new_n16825), .Y(new_n16827));
  NAND2xp33_ASAP7_75t_L     g16571(.A(new_n16826), .B(new_n16827), .Y(new_n16828));
  XNOR2x2_ASAP7_75t_L       g16572(.A(new_n16828), .B(new_n16702), .Y(new_n16829));
  XNOR2x2_ASAP7_75t_L       g16573(.A(new_n16694), .B(new_n16829), .Y(new_n16830));
  A2O1A1Ixp33_ASAP7_75t_L   g16574(.A1(new_n16690), .A2(new_n16686), .B(new_n16685), .C(new_n16830), .Y(new_n16831));
  INVx1_ASAP7_75t_L         g16575(.A(new_n16831), .Y(new_n16832));
  INVx1_ASAP7_75t_L         g16576(.A(new_n16685), .Y(new_n16833));
  A2O1A1Ixp33_ASAP7_75t_L   g16577(.A1(new_n16540), .A2(new_n16547), .B(new_n16684), .C(new_n16833), .Y(new_n16834));
  NOR2xp33_ASAP7_75t_L      g16578(.A(new_n16830), .B(new_n16834), .Y(new_n16835));
  NOR2xp33_ASAP7_75t_L      g16579(.A(new_n16835), .B(new_n16832), .Y(\f[91] ));
  INVx1_ASAP7_75t_L         g16580(.A(new_n16829), .Y(new_n16837));
  A2O1A1O1Ixp25_ASAP7_75t_L g16581(.A1(new_n16522), .A2(new_n16549), .B(new_n16555), .C(new_n16681), .D(new_n16837), .Y(new_n16838));
  INVx1_ASAP7_75t_L         g16582(.A(new_n16828), .Y(new_n16839));
  AOI21xp33_ASAP7_75t_L     g16583(.A1(new_n16839), .A2(new_n16701), .B(new_n16699), .Y(new_n16840));
  AOI22xp33_ASAP7_75t_L     g16584(.A1(new_n3029), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n3258), .Y(new_n16841));
  OAI221xp5_ASAP7_75t_L     g16585(.A1(new_n3024), .A2(new_n10847), .B1(new_n3256), .B2(new_n12047), .C(new_n16841), .Y(new_n16842));
  XNOR2x2_ASAP7_75t_L       g16586(.A(\a[32] ), .B(new_n16842), .Y(new_n16843));
  A2O1A1Ixp33_ASAP7_75t_L   g16587(.A1(new_n16821), .A2(new_n16824), .B(new_n16820), .C(new_n16843), .Y(new_n16844));
  AOI211xp5_ASAP7_75t_L     g16588(.A1(new_n16821), .A2(new_n16824), .B(new_n16843), .C(new_n16820), .Y(new_n16845));
  INVx1_ASAP7_75t_L         g16589(.A(new_n16845), .Y(new_n16846));
  NAND2xp33_ASAP7_75t_L     g16590(.A(new_n16844), .B(new_n16846), .Y(new_n16847));
  NOR2xp33_ASAP7_75t_L      g16591(.A(new_n16815), .B(new_n16812), .Y(new_n16848));
  AOI22xp33_ASAP7_75t_L     g16592(.A1(new_n4283), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n4512), .Y(new_n16849));
  OAI221xp5_ASAP7_75t_L     g16593(.A1(new_n4277), .A2(new_n8762), .B1(new_n4499), .B2(new_n9331), .C(new_n16849), .Y(new_n16850));
  XNOR2x2_ASAP7_75t_L       g16594(.A(\a[38] ), .B(new_n16850), .Y(new_n16851));
  INVx1_ASAP7_75t_L         g16595(.A(new_n16851), .Y(new_n16852));
  AOI22xp33_ASAP7_75t_L     g16596(.A1(new_n4920), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n5167), .Y(new_n16853));
  OAI221xp5_ASAP7_75t_L     g16597(.A1(new_n5154), .A2(new_n7900), .B1(new_n5158), .B2(new_n8174), .C(new_n16853), .Y(new_n16854));
  XNOR2x2_ASAP7_75t_L       g16598(.A(\a[41] ), .B(new_n16854), .Y(new_n16855));
  INVx1_ASAP7_75t_L         g16599(.A(new_n16855), .Y(new_n16856));
  AOI22xp33_ASAP7_75t_L     g16600(.A1(new_n7111), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n7391), .Y(new_n16857));
  OAI221xp5_ASAP7_75t_L     g16601(.A1(new_n8558), .A2(new_n5805), .B1(new_n8237), .B2(new_n5835), .C(new_n16857), .Y(new_n16858));
  XNOR2x2_ASAP7_75t_L       g16602(.A(\a[50] ), .B(new_n16858), .Y(new_n16859));
  INVx1_ASAP7_75t_L         g16603(.A(new_n16859), .Y(new_n16860));
  O2A1O1Ixp33_ASAP7_75t_L   g16604(.A1(new_n16599), .A2(new_n16605), .B(new_n16715), .C(new_n16758), .Y(new_n16861));
  O2A1O1Ixp33_ASAP7_75t_L   g16605(.A1(new_n16762), .A2(new_n16760), .B(new_n16714), .C(new_n16861), .Y(new_n16862));
  AOI22xp33_ASAP7_75t_L     g16606(.A1(new_n7960), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n8537), .Y(new_n16863));
  OAI221xp5_ASAP7_75t_L     g16607(.A1(new_n8817), .A2(new_n4869), .B1(new_n7957), .B2(new_n5327), .C(new_n16863), .Y(new_n16864));
  XNOR2x2_ASAP7_75t_L       g16608(.A(\a[53] ), .B(new_n16864), .Y(new_n16865));
  AOI22xp33_ASAP7_75t_L     g16609(.A1(new_n9700), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n10027), .Y(new_n16866));
  OAI221xp5_ASAP7_75t_L     g16610(.A1(new_n10024), .A2(new_n3584), .B1(new_n9696), .B2(new_n10137), .C(new_n16866), .Y(new_n16867));
  XNOR2x2_ASAP7_75t_L       g16611(.A(\a[59] ), .B(new_n16867), .Y(new_n16868));
  AOI22xp33_ASAP7_75t_L     g16612(.A1(\b[30] ), .A2(new_n10939), .B1(\b[32] ), .B2(new_n10938), .Y(new_n16869));
  OAI221xp5_ASAP7_75t_L     g16613(.A1(new_n10937), .A2(new_n3180), .B1(new_n10629), .B2(new_n11047), .C(new_n16869), .Y(new_n16870));
  XNOR2x2_ASAP7_75t_L       g16614(.A(\a[62] ), .B(new_n16870), .Y(new_n16871));
  A2O1A1Ixp33_ASAP7_75t_L   g16615(.A1(new_n16731), .A2(new_n16732), .B(new_n16727), .C(new_n16726), .Y(new_n16872));
  NOR2xp33_ASAP7_75t_L      g16616(.A(new_n2666), .B(new_n11535), .Y(new_n16873));
  A2O1A1Ixp33_ASAP7_75t_L   g16617(.A1(\b[29] ), .A2(new_n11533), .B(new_n16873), .C(new_n16723), .Y(new_n16874));
  INVx1_ASAP7_75t_L         g16618(.A(new_n16874), .Y(new_n16875));
  O2A1O1Ixp33_ASAP7_75t_L   g16619(.A1(new_n11247), .A2(new_n11249), .B(\b[29] ), .C(new_n16873), .Y(new_n16876));
  A2O1A1Ixp33_ASAP7_75t_L   g16620(.A1(new_n11533), .A2(\b[28] ), .B(new_n16720), .C(new_n16876), .Y(new_n16877));
  INVx1_ASAP7_75t_L         g16621(.A(new_n16877), .Y(new_n16878));
  NOR3xp33_ASAP7_75t_L      g16622(.A(new_n16872), .B(new_n16875), .C(new_n16878), .Y(new_n16879));
  NOR2xp33_ASAP7_75t_L      g16623(.A(new_n16875), .B(new_n16878), .Y(new_n16880));
  A2O1A1O1Ixp25_ASAP7_75t_L g16624(.A1(new_n16732), .A2(new_n16731), .B(new_n16727), .C(new_n16726), .D(new_n16880), .Y(new_n16881));
  NOR2xp33_ASAP7_75t_L      g16625(.A(new_n16881), .B(new_n16879), .Y(new_n16882));
  NOR2xp33_ASAP7_75t_L      g16626(.A(new_n16871), .B(new_n16882), .Y(new_n16883));
  INVx1_ASAP7_75t_L         g16627(.A(new_n16883), .Y(new_n16884));
  NAND2xp33_ASAP7_75t_L     g16628(.A(new_n16871), .B(new_n16882), .Y(new_n16885));
  NAND2xp33_ASAP7_75t_L     g16629(.A(new_n16885), .B(new_n16884), .Y(new_n16886));
  NOR2xp33_ASAP7_75t_L      g16630(.A(new_n16868), .B(new_n16886), .Y(new_n16887));
  AND2x2_ASAP7_75t_L        g16631(.A(new_n16868), .B(new_n16886), .Y(new_n16888));
  NOR2xp33_ASAP7_75t_L      g16632(.A(new_n16887), .B(new_n16888), .Y(new_n16889));
  NAND3xp33_ASAP7_75t_L     g16633(.A(new_n16889), .B(new_n16747), .C(new_n16743), .Y(new_n16890));
  O2A1O1Ixp33_ASAP7_75t_L   g16634(.A1(new_n16737), .A2(new_n16740), .B(new_n16747), .C(new_n16889), .Y(new_n16891));
  INVx1_ASAP7_75t_L         g16635(.A(new_n16891), .Y(new_n16892));
  AOI22xp33_ASAP7_75t_L     g16636(.A1(new_n8831), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n9115), .Y(new_n16893));
  OAI221xp5_ASAP7_75t_L     g16637(.A1(new_n10343), .A2(new_n4424), .B1(new_n10016), .B2(new_n4641), .C(new_n16893), .Y(new_n16894));
  XNOR2x2_ASAP7_75t_L       g16638(.A(\a[56] ), .B(new_n16894), .Y(new_n16895));
  NAND3xp33_ASAP7_75t_L     g16639(.A(new_n16892), .B(new_n16890), .C(new_n16895), .Y(new_n16896));
  INVx1_ASAP7_75t_L         g16640(.A(new_n16896), .Y(new_n16897));
  AOI21xp33_ASAP7_75t_L     g16641(.A1(new_n16892), .A2(new_n16890), .B(new_n16895), .Y(new_n16898));
  NOR2xp33_ASAP7_75t_L      g16642(.A(new_n16898), .B(new_n16897), .Y(new_n16899));
  INVx1_ASAP7_75t_L         g16643(.A(new_n16899), .Y(new_n16900));
  OAI211xp5_ASAP7_75t_L     g16644(.A1(new_n16751), .A2(new_n16752), .B(new_n16900), .C(new_n16755), .Y(new_n16901));
  O2A1O1Ixp33_ASAP7_75t_L   g16645(.A1(new_n16751), .A2(new_n16752), .B(new_n16755), .C(new_n16900), .Y(new_n16902));
  INVx1_ASAP7_75t_L         g16646(.A(new_n16902), .Y(new_n16903));
  AND2x2_ASAP7_75t_L        g16647(.A(new_n16901), .B(new_n16903), .Y(new_n16904));
  NAND2xp33_ASAP7_75t_L     g16648(.A(new_n16865), .B(new_n16904), .Y(new_n16905));
  AO21x2_ASAP7_75t_L        g16649(.A1(new_n16901), .A2(new_n16903), .B(new_n16865), .Y(new_n16906));
  AND2x2_ASAP7_75t_L        g16650(.A(new_n16906), .B(new_n16905), .Y(new_n16907));
  NOR2xp33_ASAP7_75t_L      g16651(.A(new_n16862), .B(new_n16907), .Y(new_n16908));
  INVx1_ASAP7_75t_L         g16652(.A(new_n16908), .Y(new_n16909));
  NAND2xp33_ASAP7_75t_L     g16653(.A(new_n16862), .B(new_n16907), .Y(new_n16910));
  NAND3xp33_ASAP7_75t_L     g16654(.A(new_n16909), .B(new_n16860), .C(new_n16910), .Y(new_n16911));
  INVx1_ASAP7_75t_L         g16655(.A(new_n16911), .Y(new_n16912));
  AOI21xp33_ASAP7_75t_L     g16656(.A1(new_n16909), .A2(new_n16910), .B(new_n16860), .Y(new_n16913));
  NOR4xp25_ASAP7_75t_L      g16657(.A(new_n16912), .B(new_n16772), .C(new_n16766), .D(new_n16913), .Y(new_n16914));
  NOR2xp33_ASAP7_75t_L      g16658(.A(new_n16913), .B(new_n16912), .Y(new_n16915));
  O2A1O1Ixp33_ASAP7_75t_L   g16659(.A1(new_n16768), .A2(new_n16771), .B(new_n16767), .C(new_n16915), .Y(new_n16916));
  NOR2xp33_ASAP7_75t_L      g16660(.A(new_n16914), .B(new_n16916), .Y(new_n16917));
  AOI22xp33_ASAP7_75t_L     g16661(.A1(new_n6376), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n6648), .Y(new_n16918));
  OAI221xp5_ASAP7_75t_L     g16662(.A1(new_n6646), .A2(new_n6568), .B1(new_n6636), .B2(new_n6820), .C(new_n16918), .Y(new_n16919));
  XNOR2x2_ASAP7_75t_L       g16663(.A(\a[47] ), .B(new_n16919), .Y(new_n16920));
  AND2x2_ASAP7_75t_L        g16664(.A(new_n16920), .B(new_n16917), .Y(new_n16921));
  NOR2xp33_ASAP7_75t_L      g16665(.A(new_n16920), .B(new_n16917), .Y(new_n16922));
  NOR2xp33_ASAP7_75t_L      g16666(.A(new_n16922), .B(new_n16921), .Y(new_n16923));
  A2O1A1Ixp33_ASAP7_75t_L   g16667(.A1(new_n16779), .A2(new_n16783), .B(new_n16777), .C(new_n16923), .Y(new_n16924));
  INVx1_ASAP7_75t_L         g16668(.A(new_n16923), .Y(new_n16925));
  NOR2xp33_ASAP7_75t_L      g16669(.A(new_n16777), .B(new_n16785), .Y(new_n16926));
  NAND2xp33_ASAP7_75t_L     g16670(.A(new_n16925), .B(new_n16926), .Y(new_n16927));
  AND2x2_ASAP7_75t_L        g16671(.A(new_n16924), .B(new_n16927), .Y(new_n16928));
  INVx1_ASAP7_75t_L         g16672(.A(new_n16928), .Y(new_n16929));
  AOI22xp33_ASAP7_75t_L     g16673(.A1(new_n5624), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n5901), .Y(new_n16930));
  OAI221xp5_ASAP7_75t_L     g16674(.A1(new_n5900), .A2(new_n7317), .B1(new_n5892), .B2(new_n7602), .C(new_n16930), .Y(new_n16931));
  XNOR2x2_ASAP7_75t_L       g16675(.A(\a[44] ), .B(new_n16931), .Y(new_n16932));
  AND2x2_ASAP7_75t_L        g16676(.A(new_n16932), .B(new_n16929), .Y(new_n16933));
  NOR2xp33_ASAP7_75t_L      g16677(.A(new_n16932), .B(new_n16929), .Y(new_n16934));
  NOR2xp33_ASAP7_75t_L      g16678(.A(new_n16934), .B(new_n16933), .Y(new_n16935));
  AOI21xp33_ASAP7_75t_L     g16679(.A1(new_n16793), .A2(new_n16796), .B(new_n16791), .Y(new_n16936));
  NAND2xp33_ASAP7_75t_L     g16680(.A(new_n16936), .B(new_n16935), .Y(new_n16937));
  INVx1_ASAP7_75t_L         g16681(.A(new_n16937), .Y(new_n16938));
  O2A1O1Ixp33_ASAP7_75t_L   g16682(.A1(new_n16789), .A2(new_n16790), .B(new_n16797), .C(new_n16935), .Y(new_n16939));
  NOR2xp33_ASAP7_75t_L      g16683(.A(new_n16939), .B(new_n16938), .Y(new_n16940));
  NAND2xp33_ASAP7_75t_L     g16684(.A(new_n16856), .B(new_n16940), .Y(new_n16941));
  OAI21xp33_ASAP7_75t_L     g16685(.A1(new_n16939), .A2(new_n16938), .B(new_n16855), .Y(new_n16942));
  AND2x2_ASAP7_75t_L        g16686(.A(new_n16942), .B(new_n16941), .Y(new_n16943));
  AOI21xp33_ASAP7_75t_L     g16687(.A1(new_n16803), .A2(new_n16806), .B(new_n16801), .Y(new_n16944));
  NAND2xp33_ASAP7_75t_L     g16688(.A(new_n16944), .B(new_n16943), .Y(new_n16945));
  INVx1_ASAP7_75t_L         g16689(.A(new_n16943), .Y(new_n16946));
  A2O1A1Ixp33_ASAP7_75t_L   g16690(.A1(new_n16803), .A2(new_n16806), .B(new_n16801), .C(new_n16946), .Y(new_n16947));
  NAND3xp33_ASAP7_75t_L     g16691(.A(new_n16947), .B(new_n16945), .C(new_n16852), .Y(new_n16948));
  AO21x2_ASAP7_75t_L        g16692(.A1(new_n16945), .A2(new_n16947), .B(new_n16852), .Y(new_n16949));
  AND2x2_ASAP7_75t_L        g16693(.A(new_n16948), .B(new_n16949), .Y(new_n16950));
  A2O1A1Ixp33_ASAP7_75t_L   g16694(.A1(new_n16811), .A2(new_n16807), .B(new_n16848), .C(new_n16950), .Y(new_n16951));
  O2A1O1Ixp33_ASAP7_75t_L   g16695(.A1(new_n16808), .A2(new_n16809), .B(new_n16807), .C(new_n16848), .Y(new_n16952));
  INVx1_ASAP7_75t_L         g16696(.A(new_n16952), .Y(new_n16953));
  NOR2xp33_ASAP7_75t_L      g16697(.A(new_n16950), .B(new_n16953), .Y(new_n16954));
  INVx1_ASAP7_75t_L         g16698(.A(new_n16954), .Y(new_n16955));
  AOI22xp33_ASAP7_75t_L     g16699(.A1(new_n3633), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n3858), .Y(new_n16956));
  OAI221xp5_ASAP7_75t_L     g16700(.A1(new_n3853), .A2(new_n9920), .B1(new_n3856), .B2(new_n11152), .C(new_n16956), .Y(new_n16957));
  XNOR2x2_ASAP7_75t_L       g16701(.A(\a[35] ), .B(new_n16957), .Y(new_n16958));
  AND3x1_ASAP7_75t_L        g16702(.A(new_n16955), .B(new_n16958), .C(new_n16951), .Y(new_n16959));
  INVx1_ASAP7_75t_L         g16703(.A(new_n16959), .Y(new_n16960));
  AO21x2_ASAP7_75t_L        g16704(.A1(new_n16951), .A2(new_n16955), .B(new_n16958), .Y(new_n16961));
  NAND3xp33_ASAP7_75t_L     g16705(.A(new_n16847), .B(new_n16960), .C(new_n16961), .Y(new_n16962));
  AO21x2_ASAP7_75t_L        g16706(.A1(new_n16961), .A2(new_n16960), .B(new_n16847), .Y(new_n16963));
  AND2x2_ASAP7_75t_L        g16707(.A(new_n16962), .B(new_n16963), .Y(new_n16964));
  A2O1A1Ixp33_ASAP7_75t_L   g16708(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n2544), .Y(new_n16965));
  A2O1A1Ixp33_ASAP7_75t_L   g16709(.A1(new_n16965), .A2(new_n2747), .B(new_n11468), .C(\a[29] ), .Y(new_n16966));
  O2A1O1Ixp33_ASAP7_75t_L   g16710(.A1(new_n2734), .A2(new_n12060), .B(new_n2747), .C(new_n11468), .Y(new_n16967));
  NAND2xp33_ASAP7_75t_L     g16711(.A(new_n2538), .B(new_n16967), .Y(new_n16968));
  AND2x2_ASAP7_75t_L        g16712(.A(new_n16968), .B(new_n16966), .Y(new_n16969));
  O2A1O1Ixp33_ASAP7_75t_L   g16713(.A1(new_n16705), .A2(new_n16707), .B(new_n16826), .C(new_n16969), .Y(new_n16970));
  INVx1_ASAP7_75t_L         g16714(.A(new_n16970), .Y(new_n16971));
  NAND3xp33_ASAP7_75t_L     g16715(.A(new_n16826), .B(new_n16710), .C(new_n16969), .Y(new_n16972));
  NAND3xp33_ASAP7_75t_L     g16716(.A(new_n16964), .B(new_n16971), .C(new_n16972), .Y(new_n16973));
  AO21x2_ASAP7_75t_L        g16717(.A1(new_n16972), .A2(new_n16971), .B(new_n16964), .Y(new_n16974));
  AND2x2_ASAP7_75t_L        g16718(.A(new_n16973), .B(new_n16974), .Y(new_n16975));
  XNOR2x2_ASAP7_75t_L       g16719(.A(new_n16840), .B(new_n16975), .Y(new_n16976));
  A2O1A1Ixp33_ASAP7_75t_L   g16720(.A1(new_n16834), .A2(new_n16830), .B(new_n16838), .C(new_n16976), .Y(new_n16977));
  INVx1_ASAP7_75t_L         g16721(.A(new_n16838), .Y(new_n16978));
  INVx1_ASAP7_75t_L         g16722(.A(new_n16976), .Y(new_n16979));
  NAND3xp33_ASAP7_75t_L     g16723(.A(new_n16831), .B(new_n16978), .C(new_n16979), .Y(new_n16980));
  AND2x2_ASAP7_75t_L        g16724(.A(new_n16977), .B(new_n16980), .Y(\f[92] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16725(.A1(new_n16701), .A2(new_n16839), .B(new_n16699), .C(new_n16975), .Y(new_n16982));
  AOI22xp33_ASAP7_75t_L     g16726(.A1(new_n4920), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n5167), .Y(new_n16983));
  OAI221xp5_ASAP7_75t_L     g16727(.A1(new_n5154), .A2(new_n8165), .B1(new_n5158), .B2(new_n8465), .C(new_n16983), .Y(new_n16984));
  XNOR2x2_ASAP7_75t_L       g16728(.A(\a[41] ), .B(new_n16984), .Y(new_n16985));
  O2A1O1Ixp33_ASAP7_75t_L   g16729(.A1(new_n16921), .A2(new_n16922), .B(new_n16926), .C(new_n16934), .Y(new_n16986));
  A2O1A1Ixp33_ASAP7_75t_L   g16730(.A1(new_n16905), .A2(new_n16906), .B(new_n16862), .C(new_n16911), .Y(new_n16987));
  AOI22xp33_ASAP7_75t_L     g16731(.A1(new_n7111), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n7391), .Y(new_n16988));
  OAI221xp5_ASAP7_75t_L     g16732(.A1(new_n8558), .A2(new_n5829), .B1(new_n8237), .B2(new_n6329), .C(new_n16988), .Y(new_n16989));
  XNOR2x2_ASAP7_75t_L       g16733(.A(\a[50] ), .B(new_n16989), .Y(new_n16990));
  INVx1_ASAP7_75t_L         g16734(.A(new_n16990), .Y(new_n16991));
  AOI22xp33_ASAP7_75t_L     g16735(.A1(new_n9700), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n10027), .Y(new_n16992));
  OAI221xp5_ASAP7_75t_L     g16736(.A1(new_n10024), .A2(new_n3804), .B1(new_n9696), .B2(new_n4223), .C(new_n16992), .Y(new_n16993));
  XNOR2x2_ASAP7_75t_L       g16737(.A(\a[59] ), .B(new_n16993), .Y(new_n16994));
  INVx1_ASAP7_75t_L         g16738(.A(new_n16994), .Y(new_n16995));
  AOI22xp33_ASAP7_75t_L     g16739(.A1(\b[31] ), .A2(new_n10939), .B1(\b[33] ), .B2(new_n10938), .Y(new_n16996));
  OAI221xp5_ASAP7_75t_L     g16740(.A1(new_n10937), .A2(new_n3207), .B1(new_n10629), .B2(new_n3572), .C(new_n16996), .Y(new_n16997));
  XNOR2x2_ASAP7_75t_L       g16741(.A(\a[62] ), .B(new_n16997), .Y(new_n16998));
  NOR2xp33_ASAP7_75t_L      g16742(.A(new_n2688), .B(new_n11535), .Y(new_n16999));
  A2O1A1Ixp33_ASAP7_75t_L   g16743(.A1(new_n11533), .A2(\b[30] ), .B(new_n16999), .C(new_n2538), .Y(new_n17000));
  INVx1_ASAP7_75t_L         g16744(.A(new_n17000), .Y(new_n17001));
  O2A1O1Ixp33_ASAP7_75t_L   g16745(.A1(new_n11247), .A2(new_n11249), .B(\b[30] ), .C(new_n16999), .Y(new_n17002));
  NAND2xp33_ASAP7_75t_L     g16746(.A(\a[29] ), .B(new_n17002), .Y(new_n17003));
  INVx1_ASAP7_75t_L         g16747(.A(new_n17003), .Y(new_n17004));
  OAI21xp33_ASAP7_75t_L     g16748(.A1(new_n17001), .A2(new_n17004), .B(new_n16876), .Y(new_n17005));
  NOR2xp33_ASAP7_75t_L      g16749(.A(new_n17001), .B(new_n17004), .Y(new_n17006));
  A2O1A1Ixp33_ASAP7_75t_L   g16750(.A1(new_n11533), .A2(\b[29] ), .B(new_n16873), .C(new_n17006), .Y(new_n17007));
  AND2x2_ASAP7_75t_L        g16751(.A(new_n17005), .B(new_n17007), .Y(new_n17008));
  INVx1_ASAP7_75t_L         g16752(.A(new_n17008), .Y(new_n17009));
  A2O1A1O1Ixp25_ASAP7_75t_L g16753(.A1(new_n16726), .A2(new_n16736), .B(new_n16875), .C(new_n16877), .D(new_n17009), .Y(new_n17010));
  INVx1_ASAP7_75t_L         g16754(.A(new_n17010), .Y(new_n17011));
  A2O1A1O1Ixp25_ASAP7_75t_L g16755(.A1(new_n16732), .A2(new_n16731), .B(new_n16727), .C(new_n16726), .D(new_n16875), .Y(new_n17012));
  A2O1A1O1Ixp25_ASAP7_75t_L g16756(.A1(new_n11533), .A2(\b[28] ), .B(new_n16720), .C(new_n16876), .D(new_n17012), .Y(new_n17013));
  NAND2xp33_ASAP7_75t_L     g16757(.A(new_n17009), .B(new_n17013), .Y(new_n17014));
  NAND2xp33_ASAP7_75t_L     g16758(.A(new_n17014), .B(new_n17011), .Y(new_n17015));
  NOR2xp33_ASAP7_75t_L      g16759(.A(new_n16998), .B(new_n17015), .Y(new_n17016));
  INVx1_ASAP7_75t_L         g16760(.A(new_n17016), .Y(new_n17017));
  NAND2xp33_ASAP7_75t_L     g16761(.A(new_n16998), .B(new_n17015), .Y(new_n17018));
  NAND3xp33_ASAP7_75t_L     g16762(.A(new_n17017), .B(new_n16995), .C(new_n17018), .Y(new_n17019));
  INVx1_ASAP7_75t_L         g16763(.A(new_n17019), .Y(new_n17020));
  AOI21xp33_ASAP7_75t_L     g16764(.A1(new_n17017), .A2(new_n17018), .B(new_n16995), .Y(new_n17021));
  NOR2xp33_ASAP7_75t_L      g16765(.A(new_n17021), .B(new_n17020), .Y(new_n17022));
  INVx1_ASAP7_75t_L         g16766(.A(new_n17022), .Y(new_n17023));
  O2A1O1Ixp33_ASAP7_75t_L   g16767(.A1(new_n16868), .A2(new_n16886), .B(new_n16884), .C(new_n17023), .Y(new_n17024));
  NOR3xp33_ASAP7_75t_L      g16768(.A(new_n17022), .B(new_n16887), .C(new_n16883), .Y(new_n17025));
  NOR2xp33_ASAP7_75t_L      g16769(.A(new_n17025), .B(new_n17024), .Y(new_n17026));
  AOI22xp33_ASAP7_75t_L     g16770(.A1(new_n8831), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n9115), .Y(new_n17027));
  OAI221xp5_ASAP7_75t_L     g16771(.A1(new_n10343), .A2(new_n4632), .B1(new_n10016), .B2(new_n4858), .C(new_n17027), .Y(new_n17028));
  XNOR2x2_ASAP7_75t_L       g16772(.A(\a[56] ), .B(new_n17028), .Y(new_n17029));
  INVx1_ASAP7_75t_L         g16773(.A(new_n17029), .Y(new_n17030));
  XNOR2x2_ASAP7_75t_L       g16774(.A(new_n17030), .B(new_n17026), .Y(new_n17031));
  A2O1A1Ixp33_ASAP7_75t_L   g16775(.A1(new_n16895), .A2(new_n16890), .B(new_n16891), .C(new_n17031), .Y(new_n17032));
  A2O1A1Ixp33_ASAP7_75t_L   g16776(.A1(new_n16747), .A2(new_n16743), .B(new_n16889), .C(new_n16896), .Y(new_n17033));
  NOR2xp33_ASAP7_75t_L      g16777(.A(new_n17033), .B(new_n17031), .Y(new_n17034));
  INVx1_ASAP7_75t_L         g16778(.A(new_n17034), .Y(new_n17035));
  NAND2xp33_ASAP7_75t_L     g16779(.A(new_n17032), .B(new_n17035), .Y(new_n17036));
  AOI22xp33_ASAP7_75t_L     g16780(.A1(new_n7960), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n8537), .Y(new_n17037));
  OAI221xp5_ASAP7_75t_L     g16781(.A1(new_n8817), .A2(new_n5321), .B1(new_n7957), .B2(new_n5346), .C(new_n17037), .Y(new_n17038));
  XNOR2x2_ASAP7_75t_L       g16782(.A(\a[53] ), .B(new_n17038), .Y(new_n17039));
  XNOR2x2_ASAP7_75t_L       g16783(.A(new_n17039), .B(new_n17036), .Y(new_n17040));
  AOI211xp5_ASAP7_75t_L     g16784(.A1(new_n16865), .A2(new_n16901), .B(new_n16902), .C(new_n17040), .Y(new_n17041));
  INVx1_ASAP7_75t_L         g16785(.A(new_n17041), .Y(new_n17042));
  A2O1A1Ixp33_ASAP7_75t_L   g16786(.A1(new_n16901), .A2(new_n16865), .B(new_n16902), .C(new_n17040), .Y(new_n17043));
  AND2x2_ASAP7_75t_L        g16787(.A(new_n17043), .B(new_n17042), .Y(new_n17044));
  NAND2xp33_ASAP7_75t_L     g16788(.A(new_n16991), .B(new_n17044), .Y(new_n17045));
  NOR2xp33_ASAP7_75t_L      g16789(.A(new_n16991), .B(new_n17044), .Y(new_n17046));
  INVx1_ASAP7_75t_L         g16790(.A(new_n17046), .Y(new_n17047));
  AO21x2_ASAP7_75t_L        g16791(.A1(new_n17045), .A2(new_n17047), .B(new_n16987), .Y(new_n17048));
  NAND3xp33_ASAP7_75t_L     g16792(.A(new_n17047), .B(new_n17045), .C(new_n16987), .Y(new_n17049));
  NAND2xp33_ASAP7_75t_L     g16793(.A(new_n17049), .B(new_n17048), .Y(new_n17050));
  AOI22xp33_ASAP7_75t_L     g16794(.A1(new_n6376), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n6648), .Y(new_n17051));
  OAI221xp5_ASAP7_75t_L     g16795(.A1(new_n6646), .A2(new_n6812), .B1(new_n6636), .B2(new_n6837), .C(new_n17051), .Y(new_n17052));
  XNOR2x2_ASAP7_75t_L       g16796(.A(\a[47] ), .B(new_n17052), .Y(new_n17053));
  XNOR2x2_ASAP7_75t_L       g16797(.A(new_n17053), .B(new_n17050), .Y(new_n17054));
  A2O1A1Ixp33_ASAP7_75t_L   g16798(.A1(new_n16917), .A2(new_n16920), .B(new_n16916), .C(new_n17054), .Y(new_n17055));
  OR3x1_ASAP7_75t_L         g16799(.A(new_n17054), .B(new_n16916), .C(new_n16921), .Y(new_n17056));
  NAND2xp33_ASAP7_75t_L     g16800(.A(new_n17055), .B(new_n17056), .Y(new_n17057));
  AOI22xp33_ASAP7_75t_L     g16801(.A1(new_n5624), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n5901), .Y(new_n17058));
  OAI221xp5_ASAP7_75t_L     g16802(.A1(new_n5900), .A2(new_n7593), .B1(new_n5892), .B2(new_n7623), .C(new_n17058), .Y(new_n17059));
  XNOR2x2_ASAP7_75t_L       g16803(.A(\a[44] ), .B(new_n17059), .Y(new_n17060));
  XNOR2x2_ASAP7_75t_L       g16804(.A(new_n17060), .B(new_n17057), .Y(new_n17061));
  AND2x2_ASAP7_75t_L        g16805(.A(new_n17061), .B(new_n16986), .Y(new_n17062));
  O2A1O1Ixp33_ASAP7_75t_L   g16806(.A1(new_n16775), .A2(new_n16776), .B(new_n16786), .C(new_n16925), .Y(new_n17063));
  O2A1O1Ixp33_ASAP7_75t_L   g16807(.A1(new_n17063), .A2(new_n16932), .B(new_n16927), .C(new_n17061), .Y(new_n17064));
  OAI21xp33_ASAP7_75t_L     g16808(.A1(new_n17064), .A2(new_n17062), .B(new_n16985), .Y(new_n17065));
  INVx1_ASAP7_75t_L         g16809(.A(new_n16985), .Y(new_n17066));
  NOR2xp33_ASAP7_75t_L      g16810(.A(new_n17064), .B(new_n17062), .Y(new_n17067));
  NAND2xp33_ASAP7_75t_L     g16811(.A(new_n17066), .B(new_n17067), .Y(new_n17068));
  AND2x2_ASAP7_75t_L        g16812(.A(new_n17065), .B(new_n17068), .Y(new_n17069));
  INVx1_ASAP7_75t_L         g16813(.A(new_n17069), .Y(new_n17070));
  O2A1O1Ixp33_ASAP7_75t_L   g16814(.A1(new_n16855), .A2(new_n16939), .B(new_n16937), .C(new_n17070), .Y(new_n17071));
  INVx1_ASAP7_75t_L         g16815(.A(new_n17071), .Y(new_n17072));
  NAND3xp33_ASAP7_75t_L     g16816(.A(new_n17070), .B(new_n16941), .C(new_n16937), .Y(new_n17073));
  NAND2xp33_ASAP7_75t_L     g16817(.A(new_n17073), .B(new_n17072), .Y(new_n17074));
  AOI22xp33_ASAP7_75t_L     g16818(.A1(new_n4283), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n4512), .Y(new_n17075));
  OAI221xp5_ASAP7_75t_L     g16819(.A1(new_n4277), .A2(new_n9323), .B1(new_n4499), .B2(new_n9627), .C(new_n17075), .Y(new_n17076));
  XNOR2x2_ASAP7_75t_L       g16820(.A(\a[38] ), .B(new_n17076), .Y(new_n17077));
  XNOR2x2_ASAP7_75t_L       g16821(.A(new_n17077), .B(new_n17074), .Y(new_n17078));
  NAND3xp33_ASAP7_75t_L     g16822(.A(new_n17078), .B(new_n16948), .C(new_n16945), .Y(new_n17079));
  AO21x2_ASAP7_75t_L        g16823(.A1(new_n16945), .A2(new_n16948), .B(new_n17078), .Y(new_n17080));
  AND2x2_ASAP7_75t_L        g16824(.A(new_n17079), .B(new_n17080), .Y(new_n17081));
  AOI22xp33_ASAP7_75t_L     g16825(.A1(new_n3633), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n3858), .Y(new_n17082));
  OAI221xp5_ASAP7_75t_L     g16826(.A1(new_n3853), .A2(new_n9947), .B1(new_n3856), .B2(new_n11446), .C(new_n17082), .Y(new_n17083));
  XNOR2x2_ASAP7_75t_L       g16827(.A(\a[35] ), .B(new_n17083), .Y(new_n17084));
  INVx1_ASAP7_75t_L         g16828(.A(new_n17084), .Y(new_n17085));
  XNOR2x2_ASAP7_75t_L       g16829(.A(new_n17085), .B(new_n17081), .Y(new_n17086));
  A2O1A1Ixp33_ASAP7_75t_L   g16830(.A1(new_n16958), .A2(new_n16951), .B(new_n16954), .C(new_n17086), .Y(new_n17087));
  INVx1_ASAP7_75t_L         g16831(.A(new_n17086), .Y(new_n17088));
  NAND3xp33_ASAP7_75t_L     g16832(.A(new_n17088), .B(new_n16960), .C(new_n16955), .Y(new_n17089));
  AND2x2_ASAP7_75t_L        g16833(.A(new_n17087), .B(new_n17089), .Y(new_n17090));
  INVx1_ASAP7_75t_L         g16834(.A(new_n17090), .Y(new_n17091));
  AOI22xp33_ASAP7_75t_L     g16835(.A1(new_n3029), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n3258), .Y(new_n17092));
  A2O1A1Ixp33_ASAP7_75t_L   g16836(.A1(new_n11470), .A2(new_n11473), .B(new_n3256), .C(new_n17092), .Y(new_n17093));
  AOI21xp33_ASAP7_75t_L     g16837(.A1(new_n3030), .A2(\b[62] ), .B(new_n17093), .Y(new_n17094));
  NAND2xp33_ASAP7_75t_L     g16838(.A(\a[32] ), .B(new_n17094), .Y(new_n17095));
  A2O1A1Ixp33_ASAP7_75t_L   g16839(.A1(\b[62] ), .A2(new_n3030), .B(new_n17093), .C(new_n3015), .Y(new_n17096));
  AND2x2_ASAP7_75t_L        g16840(.A(new_n17096), .B(new_n17095), .Y(new_n17097));
  INVx1_ASAP7_75t_L         g16841(.A(new_n17097), .Y(new_n17098));
  A2O1A1O1Ixp25_ASAP7_75t_L g16842(.A1(new_n16961), .A2(new_n16960), .B(new_n16847), .C(new_n16846), .D(new_n17098), .Y(new_n17099));
  A2O1A1Ixp33_ASAP7_75t_L   g16843(.A1(new_n16960), .A2(new_n16961), .B(new_n16847), .C(new_n16846), .Y(new_n17100));
  NOR2xp33_ASAP7_75t_L      g16844(.A(new_n17097), .B(new_n17100), .Y(new_n17101));
  NOR2xp33_ASAP7_75t_L      g16845(.A(new_n17099), .B(new_n17101), .Y(new_n17102));
  NAND2xp33_ASAP7_75t_L     g16846(.A(new_n17091), .B(new_n17102), .Y(new_n17103));
  NOR2xp33_ASAP7_75t_L      g16847(.A(new_n17091), .B(new_n17102), .Y(new_n17104));
  INVx1_ASAP7_75t_L         g16848(.A(new_n17104), .Y(new_n17105));
  NAND2xp33_ASAP7_75t_L     g16849(.A(new_n17103), .B(new_n17105), .Y(new_n17106));
  A2O1A1O1Ixp25_ASAP7_75t_L g16850(.A1(new_n16826), .A2(new_n16710), .B(new_n16969), .C(new_n16973), .D(new_n17106), .Y(new_n17107));
  INVx1_ASAP7_75t_L         g16851(.A(new_n17107), .Y(new_n17108));
  NAND3xp33_ASAP7_75t_L     g16852(.A(new_n17106), .B(new_n16973), .C(new_n16971), .Y(new_n17109));
  NAND2xp33_ASAP7_75t_L     g16853(.A(new_n17109), .B(new_n17108), .Y(new_n17110));
  A2O1A1O1Ixp25_ASAP7_75t_L g16854(.A1(new_n16978), .A2(new_n16831), .B(new_n16979), .C(new_n16982), .D(new_n17110), .Y(new_n17111));
  A2O1A1Ixp33_ASAP7_75t_L   g16855(.A1(new_n16831), .A2(new_n16978), .B(new_n16979), .C(new_n16982), .Y(new_n17112));
  INVx1_ASAP7_75t_L         g16856(.A(new_n17110), .Y(new_n17113));
  NOR2xp33_ASAP7_75t_L      g16857(.A(new_n17113), .B(new_n17112), .Y(new_n17114));
  NOR2xp33_ASAP7_75t_L      g16858(.A(new_n17111), .B(new_n17114), .Y(\f[93] ));
  INVx1_ASAP7_75t_L         g16859(.A(new_n17081), .Y(new_n17116));
  NOR2xp33_ASAP7_75t_L      g16860(.A(new_n11172), .B(new_n3402), .Y(new_n17117));
  AOI221xp5_ASAP7_75t_L     g16861(.A1(\b[63] ), .A2(new_n3030), .B1(new_n3021), .B2(new_n12322), .C(new_n17117), .Y(new_n17118));
  XNOR2x2_ASAP7_75t_L       g16862(.A(new_n3015), .B(new_n17118), .Y(new_n17119));
  O2A1O1Ixp33_ASAP7_75t_L   g16863(.A1(new_n17116), .A2(new_n17084), .B(new_n17089), .C(new_n17119), .Y(new_n17120));
  INVx1_ASAP7_75t_L         g16864(.A(new_n17120), .Y(new_n17121));
  OAI211xp5_ASAP7_75t_L     g16865(.A1(new_n17084), .A2(new_n17116), .B(new_n17089), .C(new_n17119), .Y(new_n17122));
  NAND2xp33_ASAP7_75t_L     g16866(.A(new_n17122), .B(new_n17121), .Y(new_n17123));
  AOI22xp33_ASAP7_75t_L     g16867(.A1(new_n8831), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n9115), .Y(new_n17124));
  OAI221xp5_ASAP7_75t_L     g16868(.A1(new_n10343), .A2(new_n4848), .B1(new_n10016), .B2(new_n11686), .C(new_n17124), .Y(new_n17125));
  XNOR2x2_ASAP7_75t_L       g16869(.A(\a[56] ), .B(new_n17125), .Y(new_n17126));
  INVx1_ASAP7_75t_L         g16870(.A(new_n17126), .Y(new_n17127));
  INVx1_ASAP7_75t_L         g16871(.A(new_n16871), .Y(new_n17128));
  O2A1O1Ixp33_ASAP7_75t_L   g16872(.A1(new_n16879), .A2(new_n16881), .B(new_n17128), .C(new_n16887), .Y(new_n17129));
  AOI22xp33_ASAP7_75t_L     g16873(.A1(new_n9700), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n10027), .Y(new_n17130));
  OAI221xp5_ASAP7_75t_L     g16874(.A1(new_n10024), .A2(new_n4216), .B1(new_n9696), .B2(new_n4431), .C(new_n17130), .Y(new_n17131));
  XNOR2x2_ASAP7_75t_L       g16875(.A(\a[59] ), .B(new_n17131), .Y(new_n17132));
  INVx1_ASAP7_75t_L         g16876(.A(new_n17132), .Y(new_n17133));
  NOR2xp33_ASAP7_75t_L      g16877(.A(new_n2982), .B(new_n11535), .Y(new_n17134));
  A2O1A1O1Ixp25_ASAP7_75t_L g16878(.A1(new_n11533), .A2(\b[29] ), .B(new_n16873), .C(new_n17003), .D(new_n17001), .Y(new_n17135));
  A2O1A1Ixp33_ASAP7_75t_L   g16879(.A1(new_n11533), .A2(\b[31] ), .B(new_n17134), .C(new_n17135), .Y(new_n17136));
  O2A1O1Ixp33_ASAP7_75t_L   g16880(.A1(new_n11247), .A2(new_n11249), .B(\b[31] ), .C(new_n17134), .Y(new_n17137));
  INVx1_ASAP7_75t_L         g16881(.A(new_n17137), .Y(new_n17138));
  O2A1O1Ixp33_ASAP7_75t_L   g16882(.A1(new_n16876), .A2(new_n17004), .B(new_n17000), .C(new_n17138), .Y(new_n17139));
  INVx1_ASAP7_75t_L         g16883(.A(new_n17139), .Y(new_n17140));
  NAND2xp33_ASAP7_75t_L     g16884(.A(new_n17136), .B(new_n17140), .Y(new_n17141));
  NAND2xp33_ASAP7_75t_L     g16885(.A(\b[32] ), .B(new_n10939), .Y(new_n17142));
  OAI221xp5_ASAP7_75t_L     g16886(.A1(new_n10630), .A2(new_n3584), .B1(new_n10629), .B2(new_n3591), .C(new_n17142), .Y(new_n17143));
  AOI21xp33_ASAP7_75t_L     g16887(.A1(new_n10632), .A2(\b[33] ), .B(new_n17143), .Y(new_n17144));
  NAND2xp33_ASAP7_75t_L     g16888(.A(\a[62] ), .B(new_n17144), .Y(new_n17145));
  A2O1A1Ixp33_ASAP7_75t_L   g16889(.A1(\b[33] ), .A2(new_n10632), .B(new_n17143), .C(new_n10622), .Y(new_n17146));
  AND2x2_ASAP7_75t_L        g16890(.A(new_n17146), .B(new_n17145), .Y(new_n17147));
  XOR2x2_ASAP7_75t_L        g16891(.A(new_n17141), .B(new_n17147), .Y(new_n17148));
  INVx1_ASAP7_75t_L         g16892(.A(new_n17148), .Y(new_n17149));
  O2A1O1Ixp33_ASAP7_75t_L   g16893(.A1(new_n16998), .A2(new_n17015), .B(new_n17011), .C(new_n17149), .Y(new_n17150));
  INVx1_ASAP7_75t_L         g16894(.A(new_n17150), .Y(new_n17151));
  O2A1O1Ixp33_ASAP7_75t_L   g16895(.A1(new_n16878), .A2(new_n17012), .B(new_n17008), .C(new_n17016), .Y(new_n17152));
  NAND2xp33_ASAP7_75t_L     g16896(.A(new_n17149), .B(new_n17152), .Y(new_n17153));
  NAND3xp33_ASAP7_75t_L     g16897(.A(new_n17153), .B(new_n17151), .C(new_n17133), .Y(new_n17154));
  INVx1_ASAP7_75t_L         g16898(.A(new_n17154), .Y(new_n17155));
  AOI21xp33_ASAP7_75t_L     g16899(.A1(new_n17153), .A2(new_n17151), .B(new_n17133), .Y(new_n17156));
  NOR2xp33_ASAP7_75t_L      g16900(.A(new_n17156), .B(new_n17155), .Y(new_n17157));
  INVx1_ASAP7_75t_L         g16901(.A(new_n17157), .Y(new_n17158));
  O2A1O1Ixp33_ASAP7_75t_L   g16902(.A1(new_n17129), .A2(new_n17023), .B(new_n17019), .C(new_n17158), .Y(new_n17159));
  INVx1_ASAP7_75t_L         g16903(.A(new_n17159), .Y(new_n17160));
  INVx1_ASAP7_75t_L         g16904(.A(new_n17024), .Y(new_n17161));
  NAND3xp33_ASAP7_75t_L     g16905(.A(new_n17161), .B(new_n17019), .C(new_n17158), .Y(new_n17162));
  AND2x2_ASAP7_75t_L        g16906(.A(new_n17162), .B(new_n17160), .Y(new_n17163));
  NAND2xp33_ASAP7_75t_L     g16907(.A(new_n17127), .B(new_n17163), .Y(new_n17164));
  INVx1_ASAP7_75t_L         g16908(.A(new_n17164), .Y(new_n17165));
  NOR2xp33_ASAP7_75t_L      g16909(.A(new_n17127), .B(new_n17163), .Y(new_n17166));
  NOR2xp33_ASAP7_75t_L      g16910(.A(new_n17166), .B(new_n17165), .Y(new_n17167));
  A2O1A1Ixp33_ASAP7_75t_L   g16911(.A1(new_n17030), .A2(new_n17026), .B(new_n17034), .C(new_n17167), .Y(new_n17168));
  AOI211xp5_ASAP7_75t_L     g16912(.A1(new_n17026), .A2(new_n17030), .B(new_n17034), .C(new_n17167), .Y(new_n17169));
  INVx1_ASAP7_75t_L         g16913(.A(new_n17169), .Y(new_n17170));
  NAND2xp33_ASAP7_75t_L     g16914(.A(new_n17168), .B(new_n17170), .Y(new_n17171));
  NAND2xp33_ASAP7_75t_L     g16915(.A(\b[41] ), .B(new_n8537), .Y(new_n17172));
  OAI221xp5_ASAP7_75t_L     g16916(.A1(new_n8243), .A2(new_n5805), .B1(new_n7957), .B2(new_n6338), .C(new_n17172), .Y(new_n17173));
  AOI21xp33_ASAP7_75t_L     g16917(.A1(new_n7963), .A2(\b[42] ), .B(new_n17173), .Y(new_n17174));
  NAND2xp33_ASAP7_75t_L     g16918(.A(\a[53] ), .B(new_n17174), .Y(new_n17175));
  A2O1A1Ixp33_ASAP7_75t_L   g16919(.A1(\b[42] ), .A2(new_n7963), .B(new_n17173), .C(new_n7954), .Y(new_n17176));
  NAND2xp33_ASAP7_75t_L     g16920(.A(new_n17176), .B(new_n17175), .Y(new_n17177));
  NOR2xp33_ASAP7_75t_L      g16921(.A(new_n17177), .B(new_n17171), .Y(new_n17178));
  INVx1_ASAP7_75t_L         g16922(.A(new_n17178), .Y(new_n17179));
  NAND2xp33_ASAP7_75t_L     g16923(.A(new_n17177), .B(new_n17171), .Y(new_n17180));
  AND2x2_ASAP7_75t_L        g16924(.A(new_n17180), .B(new_n17179), .Y(new_n17181));
  INVx1_ASAP7_75t_L         g16925(.A(new_n17181), .Y(new_n17182));
  OAI21xp33_ASAP7_75t_L     g16926(.A1(new_n17036), .A2(new_n17039), .B(new_n17042), .Y(new_n17183));
  NOR2xp33_ASAP7_75t_L      g16927(.A(new_n17183), .B(new_n17182), .Y(new_n17184));
  O2A1O1Ixp33_ASAP7_75t_L   g16928(.A1(new_n17036), .A2(new_n17039), .B(new_n17042), .C(new_n17181), .Y(new_n17185));
  NOR2xp33_ASAP7_75t_L      g16929(.A(new_n17185), .B(new_n17184), .Y(new_n17186));
  INVx1_ASAP7_75t_L         g16930(.A(new_n17186), .Y(new_n17187));
  AOI22xp33_ASAP7_75t_L     g16931(.A1(new_n7111), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n7391), .Y(new_n17188));
  OAI221xp5_ASAP7_75t_L     g16932(.A1(new_n8558), .A2(new_n6321), .B1(new_n8237), .B2(new_n6573), .C(new_n17188), .Y(new_n17189));
  XNOR2x2_ASAP7_75t_L       g16933(.A(\a[50] ), .B(new_n17189), .Y(new_n17190));
  INVx1_ASAP7_75t_L         g16934(.A(new_n17190), .Y(new_n17191));
  NOR2xp33_ASAP7_75t_L      g16935(.A(new_n17191), .B(new_n17187), .Y(new_n17192));
  INVx1_ASAP7_75t_L         g16936(.A(new_n17192), .Y(new_n17193));
  NAND2xp33_ASAP7_75t_L     g16937(.A(new_n17191), .B(new_n17187), .Y(new_n17194));
  AND2x2_ASAP7_75t_L        g16938(.A(new_n17194), .B(new_n17193), .Y(new_n17195));
  INVx1_ASAP7_75t_L         g16939(.A(new_n17195), .Y(new_n17196));
  A2O1A1Ixp33_ASAP7_75t_L   g16940(.A1(new_n16911), .A2(new_n16909), .B(new_n17046), .C(new_n17045), .Y(new_n17197));
  NOR2xp33_ASAP7_75t_L      g16941(.A(new_n17197), .B(new_n17196), .Y(new_n17198));
  A2O1A1O1Ixp25_ASAP7_75t_L g16942(.A1(new_n16911), .A2(new_n16909), .B(new_n17046), .C(new_n17045), .D(new_n17195), .Y(new_n17199));
  NOR2xp33_ASAP7_75t_L      g16943(.A(new_n17199), .B(new_n17198), .Y(new_n17200));
  AOI22xp33_ASAP7_75t_L     g16944(.A1(new_n6376), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n6648), .Y(new_n17201));
  OAI221xp5_ASAP7_75t_L     g16945(.A1(new_n6646), .A2(new_n6830), .B1(new_n6636), .B2(new_n7323), .C(new_n17201), .Y(new_n17202));
  XNOR2x2_ASAP7_75t_L       g16946(.A(\a[47] ), .B(new_n17202), .Y(new_n17203));
  NAND2xp33_ASAP7_75t_L     g16947(.A(new_n17203), .B(new_n17200), .Y(new_n17204));
  INVx1_ASAP7_75t_L         g16948(.A(new_n17203), .Y(new_n17205));
  OAI21xp33_ASAP7_75t_L     g16949(.A1(new_n17199), .A2(new_n17198), .B(new_n17205), .Y(new_n17206));
  AND2x2_ASAP7_75t_L        g16950(.A(new_n17206), .B(new_n17204), .Y(new_n17207));
  OA211x2_ASAP7_75t_L       g16951(.A1(new_n17053), .A2(new_n17050), .B(new_n17207), .C(new_n17056), .Y(new_n17208));
  O2A1O1Ixp33_ASAP7_75t_L   g16952(.A1(new_n17050), .A2(new_n17053), .B(new_n17056), .C(new_n17207), .Y(new_n17209));
  NOR2xp33_ASAP7_75t_L      g16953(.A(new_n17209), .B(new_n17208), .Y(new_n17210));
  AOI22xp33_ASAP7_75t_L     g16954(.A1(new_n5624), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n5901), .Y(new_n17211));
  OAI221xp5_ASAP7_75t_L     g16955(.A1(new_n5900), .A2(new_n7616), .B1(new_n5892), .B2(new_n7906), .C(new_n17211), .Y(new_n17212));
  XNOR2x2_ASAP7_75t_L       g16956(.A(\a[44] ), .B(new_n17212), .Y(new_n17213));
  XNOR2x2_ASAP7_75t_L       g16957(.A(new_n17213), .B(new_n17210), .Y(new_n17214));
  MAJIxp5_ASAP7_75t_L       g16958(.A(new_n16986), .B(new_n17057), .C(new_n17060), .Y(new_n17215));
  XNOR2x2_ASAP7_75t_L       g16959(.A(new_n17215), .B(new_n17214), .Y(new_n17216));
  AOI22xp33_ASAP7_75t_L     g16960(.A1(new_n4920), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n5167), .Y(new_n17217));
  OAI221xp5_ASAP7_75t_L     g16961(.A1(new_n5154), .A2(new_n8458), .B1(new_n5158), .B2(new_n8768), .C(new_n17217), .Y(new_n17218));
  XNOR2x2_ASAP7_75t_L       g16962(.A(\a[41] ), .B(new_n17218), .Y(new_n17219));
  INVx1_ASAP7_75t_L         g16963(.A(new_n17219), .Y(new_n17220));
  XNOR2x2_ASAP7_75t_L       g16964(.A(new_n17220), .B(new_n17216), .Y(new_n17221));
  A2O1A1Ixp33_ASAP7_75t_L   g16965(.A1(new_n17067), .A2(new_n17066), .B(new_n17071), .C(new_n17221), .Y(new_n17222));
  A2O1A1Ixp33_ASAP7_75t_L   g16966(.A1(new_n16937), .A2(new_n16941), .B(new_n17070), .C(new_n17068), .Y(new_n17223));
  NOR2xp33_ASAP7_75t_L      g16967(.A(new_n17223), .B(new_n17221), .Y(new_n17224));
  INVx1_ASAP7_75t_L         g16968(.A(new_n17224), .Y(new_n17225));
  AND2x2_ASAP7_75t_L        g16969(.A(new_n17222), .B(new_n17225), .Y(new_n17226));
  AOI22xp33_ASAP7_75t_L     g16970(.A1(new_n4283), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n4512), .Y(new_n17227));
  OAI221xp5_ASAP7_75t_L     g16971(.A1(new_n4277), .A2(new_n9620), .B1(new_n4499), .B2(new_n9925), .C(new_n17227), .Y(new_n17228));
  XNOR2x2_ASAP7_75t_L       g16972(.A(\a[38] ), .B(new_n17228), .Y(new_n17229));
  NAND2xp33_ASAP7_75t_L     g16973(.A(new_n17229), .B(new_n17226), .Y(new_n17230));
  AO21x2_ASAP7_75t_L        g16974(.A1(new_n17222), .A2(new_n17225), .B(new_n17229), .Y(new_n17231));
  NAND2xp33_ASAP7_75t_L     g16975(.A(new_n17231), .B(new_n17230), .Y(new_n17232));
  OAI21xp33_ASAP7_75t_L     g16976(.A1(new_n17074), .A2(new_n17077), .B(new_n17080), .Y(new_n17233));
  NOR2xp33_ASAP7_75t_L      g16977(.A(new_n17233), .B(new_n17232), .Y(new_n17234));
  AND2x2_ASAP7_75t_L        g16978(.A(new_n17233), .B(new_n17232), .Y(new_n17235));
  NAND2xp33_ASAP7_75t_L     g16979(.A(\b[59] ), .B(new_n3858), .Y(new_n17236));
  OAI221xp5_ASAP7_75t_L     g16980(.A1(new_n4061), .A2(new_n10847), .B1(new_n3856), .B2(new_n10855), .C(new_n17236), .Y(new_n17237));
  AOI21xp33_ASAP7_75t_L     g16981(.A1(new_n3639), .A2(\b[60] ), .B(new_n17237), .Y(new_n17238));
  NAND2xp33_ASAP7_75t_L     g16982(.A(\a[35] ), .B(new_n17238), .Y(new_n17239));
  A2O1A1Ixp33_ASAP7_75t_L   g16983(.A1(\b[60] ), .A2(new_n3639), .B(new_n17237), .C(new_n3628), .Y(new_n17240));
  AOI211xp5_ASAP7_75t_L     g16984(.A1(new_n17240), .A2(new_n17239), .B(new_n17234), .C(new_n17235), .Y(new_n17241));
  INVx1_ASAP7_75t_L         g16985(.A(new_n17241), .Y(new_n17242));
  OAI211xp5_ASAP7_75t_L     g16986(.A1(new_n17234), .A2(new_n17235), .B(new_n17239), .C(new_n17240), .Y(new_n17243));
  NAND2xp33_ASAP7_75t_L     g16987(.A(new_n17243), .B(new_n17242), .Y(new_n17244));
  NOR2xp33_ASAP7_75t_L      g16988(.A(new_n17123), .B(new_n17244), .Y(new_n17245));
  INVx1_ASAP7_75t_L         g16989(.A(new_n17245), .Y(new_n17246));
  NAND2xp33_ASAP7_75t_L     g16990(.A(new_n17123), .B(new_n17244), .Y(new_n17247));
  NAND2xp33_ASAP7_75t_L     g16991(.A(new_n17247), .B(new_n17246), .Y(new_n17248));
  A2O1A1O1Ixp25_ASAP7_75t_L g16992(.A1(new_n16963), .A2(new_n16846), .B(new_n17097), .C(new_n17105), .D(new_n17248), .Y(new_n17249));
  A2O1A1O1Ixp25_ASAP7_75t_L g16993(.A1(new_n16961), .A2(new_n16960), .B(new_n16847), .C(new_n16846), .D(new_n17097), .Y(new_n17250));
  AOI211xp5_ASAP7_75t_L     g16994(.A1(new_n17246), .A2(new_n17247), .B(new_n17250), .C(new_n17104), .Y(new_n17251));
  NOR2xp33_ASAP7_75t_L      g16995(.A(new_n17251), .B(new_n17249), .Y(new_n17252));
  A2O1A1Ixp33_ASAP7_75t_L   g16996(.A1(new_n17112), .A2(new_n17113), .B(new_n17107), .C(new_n17252), .Y(new_n17253));
  INVx1_ASAP7_75t_L         g16997(.A(new_n17253), .Y(new_n17254));
  A2O1A1Ixp33_ASAP7_75t_L   g16998(.A1(new_n16977), .A2(new_n16982), .B(new_n17110), .C(new_n17108), .Y(new_n17255));
  NOR2xp33_ASAP7_75t_L      g16999(.A(new_n17252), .B(new_n17255), .Y(new_n17256));
  NOR2xp33_ASAP7_75t_L      g17000(.A(new_n17256), .B(new_n17254), .Y(\f[94] ));
  MAJIxp5_ASAP7_75t_L       g17001(.A(new_n17214), .B(new_n17215), .C(new_n17220), .Y(new_n17258));
  INVx1_ASAP7_75t_L         g17002(.A(new_n17258), .Y(new_n17259));
  AOI22xp33_ASAP7_75t_L     g17003(.A1(new_n4920), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n5167), .Y(new_n17260));
  OAI221xp5_ASAP7_75t_L     g17004(.A1(new_n5154), .A2(new_n8762), .B1(new_n5158), .B2(new_n9331), .C(new_n17260), .Y(new_n17261));
  XNOR2x2_ASAP7_75t_L       g17005(.A(\a[41] ), .B(new_n17261), .Y(new_n17262));
  INVx1_ASAP7_75t_L         g17006(.A(new_n17262), .Y(new_n17263));
  AOI22xp33_ASAP7_75t_L     g17007(.A1(new_n5624), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n5901), .Y(new_n17264));
  OAI221xp5_ASAP7_75t_L     g17008(.A1(new_n5900), .A2(new_n7900), .B1(new_n5892), .B2(new_n8174), .C(new_n17264), .Y(new_n17265));
  XNOR2x2_ASAP7_75t_L       g17009(.A(\a[44] ), .B(new_n17265), .Y(new_n17266));
  INVx1_ASAP7_75t_L         g17010(.A(new_n17266), .Y(new_n17267));
  AOI22xp33_ASAP7_75t_L     g17011(.A1(new_n7960), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n8537), .Y(new_n17268));
  OAI221xp5_ASAP7_75t_L     g17012(.A1(new_n8817), .A2(new_n5805), .B1(new_n7957), .B2(new_n5835), .C(new_n17268), .Y(new_n17269));
  XNOR2x2_ASAP7_75t_L       g17013(.A(\a[53] ), .B(new_n17269), .Y(new_n17270));
  INVx1_ASAP7_75t_L         g17014(.A(new_n17270), .Y(new_n17271));
  AOI22xp33_ASAP7_75t_L     g17015(.A1(new_n8831), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n9115), .Y(new_n17272));
  OAI221xp5_ASAP7_75t_L     g17016(.A1(new_n10343), .A2(new_n4869), .B1(new_n10016), .B2(new_n5327), .C(new_n17272), .Y(new_n17273));
  XNOR2x2_ASAP7_75t_L       g17017(.A(\a[56] ), .B(new_n17273), .Y(new_n17274));
  INVx1_ASAP7_75t_L         g17018(.A(new_n17274), .Y(new_n17275));
  AOI22xp33_ASAP7_75t_L     g17019(.A1(new_n9700), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n10027), .Y(new_n17276));
  OAI221xp5_ASAP7_75t_L     g17020(.A1(new_n10024), .A2(new_n4424), .B1(new_n9696), .B2(new_n4641), .C(new_n17276), .Y(new_n17277));
  XNOR2x2_ASAP7_75t_L       g17021(.A(\a[59] ), .B(new_n17277), .Y(new_n17278));
  AOI22xp33_ASAP7_75t_L     g17022(.A1(\b[33] ), .A2(new_n10939), .B1(\b[35] ), .B2(new_n10938), .Y(new_n17279));
  OAI221xp5_ASAP7_75t_L     g17023(.A1(new_n10937), .A2(new_n3584), .B1(new_n10629), .B2(new_n10137), .C(new_n17279), .Y(new_n17280));
  XNOR2x2_ASAP7_75t_L       g17024(.A(\a[62] ), .B(new_n17280), .Y(new_n17281));
  A2O1A1Ixp33_ASAP7_75t_L   g17025(.A1(new_n17145), .A2(new_n17146), .B(new_n17141), .C(new_n17140), .Y(new_n17282));
  NOR2xp33_ASAP7_75t_L      g17026(.A(new_n3180), .B(new_n11535), .Y(new_n17283));
  A2O1A1Ixp33_ASAP7_75t_L   g17027(.A1(\b[32] ), .A2(new_n11533), .B(new_n17283), .C(new_n17137), .Y(new_n17284));
  O2A1O1Ixp33_ASAP7_75t_L   g17028(.A1(new_n11247), .A2(new_n11249), .B(\b[32] ), .C(new_n17283), .Y(new_n17285));
  A2O1A1Ixp33_ASAP7_75t_L   g17029(.A1(new_n11533), .A2(\b[31] ), .B(new_n17134), .C(new_n17285), .Y(new_n17286));
  NAND2xp33_ASAP7_75t_L     g17030(.A(new_n17286), .B(new_n17284), .Y(new_n17287));
  XNOR2x2_ASAP7_75t_L       g17031(.A(new_n17287), .B(new_n17282), .Y(new_n17288));
  INVx1_ASAP7_75t_L         g17032(.A(new_n17288), .Y(new_n17289));
  NOR2xp33_ASAP7_75t_L      g17033(.A(new_n17281), .B(new_n17289), .Y(new_n17290));
  INVx1_ASAP7_75t_L         g17034(.A(new_n17290), .Y(new_n17291));
  NAND2xp33_ASAP7_75t_L     g17035(.A(new_n17281), .B(new_n17289), .Y(new_n17292));
  NAND2xp33_ASAP7_75t_L     g17036(.A(new_n17292), .B(new_n17291), .Y(new_n17293));
  NOR2xp33_ASAP7_75t_L      g17037(.A(new_n17278), .B(new_n17293), .Y(new_n17294));
  AND2x2_ASAP7_75t_L        g17038(.A(new_n17278), .B(new_n17293), .Y(new_n17295));
  NOR2xp33_ASAP7_75t_L      g17039(.A(new_n17294), .B(new_n17295), .Y(new_n17296));
  INVx1_ASAP7_75t_L         g17040(.A(new_n17296), .Y(new_n17297));
  O2A1O1Ixp33_ASAP7_75t_L   g17041(.A1(new_n17152), .A2(new_n17149), .B(new_n17154), .C(new_n17297), .Y(new_n17298));
  INVx1_ASAP7_75t_L         g17042(.A(new_n17298), .Y(new_n17299));
  NAND3xp33_ASAP7_75t_L     g17043(.A(new_n17297), .B(new_n17154), .C(new_n17151), .Y(new_n17300));
  NAND3xp33_ASAP7_75t_L     g17044(.A(new_n17299), .B(new_n17275), .C(new_n17300), .Y(new_n17301));
  AO21x2_ASAP7_75t_L        g17045(.A1(new_n17300), .A2(new_n17299), .B(new_n17275), .Y(new_n17302));
  AND2x2_ASAP7_75t_L        g17046(.A(new_n17301), .B(new_n17302), .Y(new_n17303));
  A2O1A1Ixp33_ASAP7_75t_L   g17047(.A1(new_n17162), .A2(new_n17127), .B(new_n17159), .C(new_n17303), .Y(new_n17304));
  OR3x1_ASAP7_75t_L         g17048(.A(new_n17165), .B(new_n17159), .C(new_n17303), .Y(new_n17305));
  AND2x2_ASAP7_75t_L        g17049(.A(new_n17304), .B(new_n17305), .Y(new_n17306));
  NAND2xp33_ASAP7_75t_L     g17050(.A(new_n17271), .B(new_n17306), .Y(new_n17307));
  INVx1_ASAP7_75t_L         g17051(.A(new_n17307), .Y(new_n17308));
  NOR2xp33_ASAP7_75t_L      g17052(.A(new_n17271), .B(new_n17306), .Y(new_n17309));
  NOR2xp33_ASAP7_75t_L      g17053(.A(new_n17309), .B(new_n17308), .Y(new_n17310));
  NAND3xp33_ASAP7_75t_L     g17054(.A(new_n17179), .B(new_n17310), .C(new_n17170), .Y(new_n17311));
  O2A1O1Ixp33_ASAP7_75t_L   g17055(.A1(new_n17171), .A2(new_n17177), .B(new_n17170), .C(new_n17310), .Y(new_n17312));
  INVx1_ASAP7_75t_L         g17056(.A(new_n17312), .Y(new_n17313));
  AOI22xp33_ASAP7_75t_L     g17057(.A1(new_n7111), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n7391), .Y(new_n17314));
  OAI221xp5_ASAP7_75t_L     g17058(.A1(new_n8558), .A2(new_n6568), .B1(new_n8237), .B2(new_n6820), .C(new_n17314), .Y(new_n17315));
  XNOR2x2_ASAP7_75t_L       g17059(.A(\a[50] ), .B(new_n17315), .Y(new_n17316));
  NAND3xp33_ASAP7_75t_L     g17060(.A(new_n17313), .B(new_n17311), .C(new_n17316), .Y(new_n17317));
  AO21x2_ASAP7_75t_L        g17061(.A1(new_n17311), .A2(new_n17313), .B(new_n17316), .Y(new_n17318));
  AND2x2_ASAP7_75t_L        g17062(.A(new_n17317), .B(new_n17318), .Y(new_n17319));
  INVx1_ASAP7_75t_L         g17063(.A(new_n17319), .Y(new_n17320));
  O2A1O1Ixp33_ASAP7_75t_L   g17064(.A1(new_n17182), .A2(new_n17183), .B(new_n17193), .C(new_n17320), .Y(new_n17321));
  NOR2xp33_ASAP7_75t_L      g17065(.A(new_n17184), .B(new_n17192), .Y(new_n17322));
  NAND2xp33_ASAP7_75t_L     g17066(.A(new_n17320), .B(new_n17322), .Y(new_n17323));
  INVx1_ASAP7_75t_L         g17067(.A(new_n17323), .Y(new_n17324));
  NOR2xp33_ASAP7_75t_L      g17068(.A(new_n17321), .B(new_n17324), .Y(new_n17325));
  INVx1_ASAP7_75t_L         g17069(.A(new_n17325), .Y(new_n17326));
  AOI22xp33_ASAP7_75t_L     g17070(.A1(new_n6376), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n6648), .Y(new_n17327));
  OAI221xp5_ASAP7_75t_L     g17071(.A1(new_n6646), .A2(new_n7317), .B1(new_n6636), .B2(new_n7602), .C(new_n17327), .Y(new_n17328));
  XNOR2x2_ASAP7_75t_L       g17072(.A(\a[47] ), .B(new_n17328), .Y(new_n17329));
  AND2x2_ASAP7_75t_L        g17073(.A(new_n17329), .B(new_n17326), .Y(new_n17330));
  NOR2xp33_ASAP7_75t_L      g17074(.A(new_n17329), .B(new_n17326), .Y(new_n17331));
  NOR2xp33_ASAP7_75t_L      g17075(.A(new_n17331), .B(new_n17330), .Y(new_n17332));
  AOI21xp33_ASAP7_75t_L     g17076(.A1(new_n17200), .A2(new_n17203), .B(new_n17198), .Y(new_n17333));
  NAND2xp33_ASAP7_75t_L     g17077(.A(new_n17333), .B(new_n17332), .Y(new_n17334));
  INVx1_ASAP7_75t_L         g17078(.A(new_n17334), .Y(new_n17335));
  O2A1O1Ixp33_ASAP7_75t_L   g17079(.A1(new_n17196), .A2(new_n17197), .B(new_n17204), .C(new_n17332), .Y(new_n17336));
  NOR2xp33_ASAP7_75t_L      g17080(.A(new_n17336), .B(new_n17335), .Y(new_n17337));
  NAND2xp33_ASAP7_75t_L     g17081(.A(new_n17267), .B(new_n17337), .Y(new_n17338));
  OAI21xp33_ASAP7_75t_L     g17082(.A1(new_n17336), .A2(new_n17335), .B(new_n17266), .Y(new_n17339));
  AND2x2_ASAP7_75t_L        g17083(.A(new_n17339), .B(new_n17338), .Y(new_n17340));
  AOI21xp33_ASAP7_75t_L     g17084(.A1(new_n17210), .A2(new_n17213), .B(new_n17208), .Y(new_n17341));
  NAND2xp33_ASAP7_75t_L     g17085(.A(new_n17341), .B(new_n17340), .Y(new_n17342));
  INVx1_ASAP7_75t_L         g17086(.A(new_n17340), .Y(new_n17343));
  A2O1A1Ixp33_ASAP7_75t_L   g17087(.A1(new_n17210), .A2(new_n17213), .B(new_n17208), .C(new_n17343), .Y(new_n17344));
  NAND3xp33_ASAP7_75t_L     g17088(.A(new_n17344), .B(new_n17342), .C(new_n17263), .Y(new_n17345));
  AO21x2_ASAP7_75t_L        g17089(.A1(new_n17342), .A2(new_n17344), .B(new_n17263), .Y(new_n17346));
  AND2x2_ASAP7_75t_L        g17090(.A(new_n17345), .B(new_n17346), .Y(new_n17347));
  NAND2xp33_ASAP7_75t_L     g17091(.A(new_n17259), .B(new_n17347), .Y(new_n17348));
  NOR2xp33_ASAP7_75t_L      g17092(.A(new_n17259), .B(new_n17347), .Y(new_n17349));
  INVx1_ASAP7_75t_L         g17093(.A(new_n17349), .Y(new_n17350));
  AOI22xp33_ASAP7_75t_L     g17094(.A1(new_n4283), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n4512), .Y(new_n17351));
  OAI221xp5_ASAP7_75t_L     g17095(.A1(new_n4277), .A2(new_n9920), .B1(new_n4499), .B2(new_n11152), .C(new_n17351), .Y(new_n17352));
  XNOR2x2_ASAP7_75t_L       g17096(.A(\a[38] ), .B(new_n17352), .Y(new_n17353));
  NAND3xp33_ASAP7_75t_L     g17097(.A(new_n17350), .B(new_n17348), .C(new_n17353), .Y(new_n17354));
  AO21x2_ASAP7_75t_L        g17098(.A1(new_n17348), .A2(new_n17350), .B(new_n17353), .Y(new_n17355));
  NAND2xp33_ASAP7_75t_L     g17099(.A(new_n17354), .B(new_n17355), .Y(new_n17356));
  O2A1O1Ixp33_ASAP7_75t_L   g17100(.A1(new_n17223), .A2(new_n17221), .B(new_n17230), .C(new_n17356), .Y(new_n17357));
  INVx1_ASAP7_75t_L         g17101(.A(new_n17357), .Y(new_n17358));
  NAND3xp33_ASAP7_75t_L     g17102(.A(new_n17356), .B(new_n17230), .C(new_n17225), .Y(new_n17359));
  AOI22xp33_ASAP7_75t_L     g17103(.A1(new_n3633), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n3858), .Y(new_n17360));
  OAI221xp5_ASAP7_75t_L     g17104(.A1(new_n3853), .A2(new_n10847), .B1(new_n3856), .B2(new_n12047), .C(new_n17360), .Y(new_n17361));
  XNOR2x2_ASAP7_75t_L       g17105(.A(\a[35] ), .B(new_n17361), .Y(new_n17362));
  AND3x1_ASAP7_75t_L        g17106(.A(new_n17358), .B(new_n17362), .C(new_n17359), .Y(new_n17363));
  INVx1_ASAP7_75t_L         g17107(.A(new_n17363), .Y(new_n17364));
  AO21x2_ASAP7_75t_L        g17108(.A1(new_n17359), .A2(new_n17358), .B(new_n17362), .Y(new_n17365));
  NAND2xp33_ASAP7_75t_L     g17109(.A(new_n17365), .B(new_n17364), .Y(new_n17366));
  A2O1A1Ixp33_ASAP7_75t_L   g17110(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n3021), .Y(new_n17367));
  A2O1A1Ixp33_ASAP7_75t_L   g17111(.A1(new_n17367), .A2(new_n3402), .B(new_n11468), .C(\a[32] ), .Y(new_n17368));
  O2A1O1Ixp33_ASAP7_75t_L   g17112(.A1(new_n3256), .A2(new_n12060), .B(new_n3402), .C(new_n11468), .Y(new_n17369));
  NAND2xp33_ASAP7_75t_L     g17113(.A(new_n3015), .B(new_n17369), .Y(new_n17370));
  AND2x2_ASAP7_75t_L        g17114(.A(new_n17370), .B(new_n17368), .Y(new_n17371));
  INVx1_ASAP7_75t_L         g17115(.A(new_n17371), .Y(new_n17372));
  A2O1A1Ixp33_ASAP7_75t_L   g17116(.A1(new_n17233), .A2(new_n17232), .B(new_n17241), .C(new_n17372), .Y(new_n17373));
  NOR2xp33_ASAP7_75t_L      g17117(.A(new_n17235), .B(new_n17241), .Y(new_n17374));
  NAND2xp33_ASAP7_75t_L     g17118(.A(new_n17371), .B(new_n17374), .Y(new_n17375));
  NAND2xp33_ASAP7_75t_L     g17119(.A(new_n17373), .B(new_n17375), .Y(new_n17376));
  XOR2x2_ASAP7_75t_L        g17120(.A(new_n17366), .B(new_n17376), .Y(new_n17377));
  O2A1O1Ixp33_ASAP7_75t_L   g17121(.A1(new_n17123), .A2(new_n17244), .B(new_n17121), .C(new_n17377), .Y(new_n17378));
  INVx1_ASAP7_75t_L         g17122(.A(new_n17378), .Y(new_n17379));
  NAND3xp33_ASAP7_75t_L     g17123(.A(new_n17377), .B(new_n17246), .C(new_n17121), .Y(new_n17380));
  NAND2xp33_ASAP7_75t_L     g17124(.A(new_n17380), .B(new_n17379), .Y(new_n17381));
  INVx1_ASAP7_75t_L         g17125(.A(new_n17381), .Y(new_n17382));
  A2O1A1Ixp33_ASAP7_75t_L   g17126(.A1(new_n17255), .A2(new_n17252), .B(new_n17249), .C(new_n17382), .Y(new_n17383));
  A2O1A1O1Ixp25_ASAP7_75t_L g17127(.A1(new_n17113), .A2(new_n17112), .B(new_n17107), .C(new_n17252), .D(new_n17249), .Y(new_n17384));
  NAND2xp33_ASAP7_75t_L     g17128(.A(new_n17381), .B(new_n17384), .Y(new_n17385));
  AND2x2_ASAP7_75t_L        g17129(.A(new_n17383), .B(new_n17385), .Y(\f[95] ));
  INVx1_ASAP7_75t_L         g17130(.A(new_n17249), .Y(new_n17387));
  INVx1_ASAP7_75t_L         g17131(.A(new_n17375), .Y(new_n17388));
  AOI22xp33_ASAP7_75t_L     g17132(.A1(new_n5624), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n5901), .Y(new_n17389));
  OAI221xp5_ASAP7_75t_L     g17133(.A1(new_n5900), .A2(new_n8165), .B1(new_n5892), .B2(new_n8465), .C(new_n17389), .Y(new_n17390));
  XNOR2x2_ASAP7_75t_L       g17134(.A(\a[44] ), .B(new_n17390), .Y(new_n17391));
  OAI21xp33_ASAP7_75t_L     g17135(.A1(new_n17329), .A2(new_n17321), .B(new_n17323), .Y(new_n17392));
  AOI22xp33_ASAP7_75t_L     g17136(.A1(new_n9700), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n10027), .Y(new_n17393));
  OAI221xp5_ASAP7_75t_L     g17137(.A1(new_n10024), .A2(new_n4632), .B1(new_n9696), .B2(new_n4858), .C(new_n17393), .Y(new_n17394));
  XNOR2x2_ASAP7_75t_L       g17138(.A(\a[59] ), .B(new_n17394), .Y(new_n17395));
  INVx1_ASAP7_75t_L         g17139(.A(new_n17395), .Y(new_n17396));
  AOI22xp33_ASAP7_75t_L     g17140(.A1(\b[34] ), .A2(new_n10939), .B1(\b[36] ), .B2(new_n10938), .Y(new_n17397));
  OAI221xp5_ASAP7_75t_L     g17141(.A1(new_n10937), .A2(new_n3804), .B1(new_n10629), .B2(new_n4223), .C(new_n17397), .Y(new_n17398));
  XNOR2x2_ASAP7_75t_L       g17142(.A(\a[62] ), .B(new_n17398), .Y(new_n17399));
  A2O1A1O1Ixp25_ASAP7_75t_L g17143(.A1(new_n11533), .A2(\b[31] ), .B(new_n17134), .C(new_n17285), .D(new_n17282), .Y(new_n17400));
  A2O1A1O1Ixp25_ASAP7_75t_L g17144(.A1(new_n11533), .A2(\b[32] ), .B(new_n17283), .C(new_n17137), .D(new_n17400), .Y(new_n17401));
  NOR2xp33_ASAP7_75t_L      g17145(.A(new_n3207), .B(new_n11535), .Y(new_n17402));
  A2O1A1Ixp33_ASAP7_75t_L   g17146(.A1(new_n11533), .A2(\b[33] ), .B(new_n17402), .C(new_n3015), .Y(new_n17403));
  INVx1_ASAP7_75t_L         g17147(.A(new_n17403), .Y(new_n17404));
  O2A1O1Ixp33_ASAP7_75t_L   g17148(.A1(new_n11247), .A2(new_n11249), .B(\b[33] ), .C(new_n17402), .Y(new_n17405));
  NAND2xp33_ASAP7_75t_L     g17149(.A(\a[32] ), .B(new_n17405), .Y(new_n17406));
  INVx1_ASAP7_75t_L         g17150(.A(new_n17406), .Y(new_n17407));
  NOR2xp33_ASAP7_75t_L      g17151(.A(new_n17404), .B(new_n17407), .Y(new_n17408));
  XNOR2x2_ASAP7_75t_L       g17152(.A(new_n17285), .B(new_n17408), .Y(new_n17409));
  NAND2xp33_ASAP7_75t_L     g17153(.A(new_n17409), .B(new_n17401), .Y(new_n17410));
  INVx1_ASAP7_75t_L         g17154(.A(new_n17410), .Y(new_n17411));
  INVx1_ASAP7_75t_L         g17155(.A(new_n17286), .Y(new_n17412));
  O2A1O1Ixp33_ASAP7_75t_L   g17156(.A1(new_n17412), .A2(new_n17282), .B(new_n17284), .C(new_n17409), .Y(new_n17413));
  NOR2xp33_ASAP7_75t_L      g17157(.A(new_n17413), .B(new_n17411), .Y(new_n17414));
  INVx1_ASAP7_75t_L         g17158(.A(new_n17414), .Y(new_n17415));
  NOR2xp33_ASAP7_75t_L      g17159(.A(new_n17399), .B(new_n17415), .Y(new_n17416));
  INVx1_ASAP7_75t_L         g17160(.A(new_n17416), .Y(new_n17417));
  NAND2xp33_ASAP7_75t_L     g17161(.A(new_n17399), .B(new_n17415), .Y(new_n17418));
  AND2x2_ASAP7_75t_L        g17162(.A(new_n17418), .B(new_n17417), .Y(new_n17419));
  NAND2xp33_ASAP7_75t_L     g17163(.A(new_n17396), .B(new_n17419), .Y(new_n17420));
  INVx1_ASAP7_75t_L         g17164(.A(new_n17420), .Y(new_n17421));
  NOR2xp33_ASAP7_75t_L      g17165(.A(new_n17396), .B(new_n17419), .Y(new_n17422));
  NOR2xp33_ASAP7_75t_L      g17166(.A(new_n17422), .B(new_n17421), .Y(new_n17423));
  INVx1_ASAP7_75t_L         g17167(.A(new_n17423), .Y(new_n17424));
  O2A1O1Ixp33_ASAP7_75t_L   g17168(.A1(new_n17278), .A2(new_n17293), .B(new_n17291), .C(new_n17424), .Y(new_n17425));
  NOR3xp33_ASAP7_75t_L      g17169(.A(new_n17423), .B(new_n17294), .C(new_n17290), .Y(new_n17426));
  NOR2xp33_ASAP7_75t_L      g17170(.A(new_n17426), .B(new_n17425), .Y(new_n17427));
  AOI22xp33_ASAP7_75t_L     g17171(.A1(new_n8831), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n9115), .Y(new_n17428));
  OAI221xp5_ASAP7_75t_L     g17172(.A1(new_n10343), .A2(new_n5321), .B1(new_n10016), .B2(new_n5346), .C(new_n17428), .Y(new_n17429));
  XNOR2x2_ASAP7_75t_L       g17173(.A(\a[56] ), .B(new_n17429), .Y(new_n17430));
  INVx1_ASAP7_75t_L         g17174(.A(new_n17430), .Y(new_n17431));
  XNOR2x2_ASAP7_75t_L       g17175(.A(new_n17431), .B(new_n17427), .Y(new_n17432));
  A2O1A1Ixp33_ASAP7_75t_L   g17176(.A1(new_n17154), .A2(new_n17151), .B(new_n17297), .C(new_n17301), .Y(new_n17433));
  INVx1_ASAP7_75t_L         g17177(.A(new_n17433), .Y(new_n17434));
  AND2x2_ASAP7_75t_L        g17178(.A(new_n17434), .B(new_n17432), .Y(new_n17435));
  A2O1A1O1Ixp25_ASAP7_75t_L g17179(.A1(new_n17154), .A2(new_n17151), .B(new_n17297), .C(new_n17301), .D(new_n17432), .Y(new_n17436));
  NOR2xp33_ASAP7_75t_L      g17180(.A(new_n17436), .B(new_n17435), .Y(new_n17437));
  AOI22xp33_ASAP7_75t_L     g17181(.A1(new_n7960), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n8537), .Y(new_n17438));
  OAI221xp5_ASAP7_75t_L     g17182(.A1(new_n8817), .A2(new_n5829), .B1(new_n7957), .B2(new_n6329), .C(new_n17438), .Y(new_n17439));
  XNOR2x2_ASAP7_75t_L       g17183(.A(\a[53] ), .B(new_n17439), .Y(new_n17440));
  INVx1_ASAP7_75t_L         g17184(.A(new_n17440), .Y(new_n17441));
  XNOR2x2_ASAP7_75t_L       g17185(.A(new_n17441), .B(new_n17437), .Y(new_n17442));
  O2A1O1Ixp33_ASAP7_75t_L   g17186(.A1(new_n17159), .A2(new_n17165), .B(new_n17303), .C(new_n17308), .Y(new_n17443));
  XOR2x2_ASAP7_75t_L        g17187(.A(new_n17443), .B(new_n17442), .Y(new_n17444));
  AOI22xp33_ASAP7_75t_L     g17188(.A1(new_n7111), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n7391), .Y(new_n17445));
  OAI221xp5_ASAP7_75t_L     g17189(.A1(new_n8558), .A2(new_n6812), .B1(new_n8237), .B2(new_n6837), .C(new_n17445), .Y(new_n17446));
  XNOR2x2_ASAP7_75t_L       g17190(.A(\a[50] ), .B(new_n17446), .Y(new_n17447));
  INVx1_ASAP7_75t_L         g17191(.A(new_n17447), .Y(new_n17448));
  XNOR2x2_ASAP7_75t_L       g17192(.A(new_n17448), .B(new_n17444), .Y(new_n17449));
  A2O1A1Ixp33_ASAP7_75t_L   g17193(.A1(new_n17316), .A2(new_n17311), .B(new_n17312), .C(new_n17449), .Y(new_n17450));
  A2O1A1Ixp33_ASAP7_75t_L   g17194(.A1(new_n17179), .A2(new_n17170), .B(new_n17310), .C(new_n17317), .Y(new_n17451));
  NOR2xp33_ASAP7_75t_L      g17195(.A(new_n17451), .B(new_n17449), .Y(new_n17452));
  INVx1_ASAP7_75t_L         g17196(.A(new_n17452), .Y(new_n17453));
  NAND2xp33_ASAP7_75t_L     g17197(.A(new_n17450), .B(new_n17453), .Y(new_n17454));
  AOI22xp33_ASAP7_75t_L     g17198(.A1(new_n6376), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n6648), .Y(new_n17455));
  OAI221xp5_ASAP7_75t_L     g17199(.A1(new_n6646), .A2(new_n7593), .B1(new_n6636), .B2(new_n7623), .C(new_n17455), .Y(new_n17456));
  XNOR2x2_ASAP7_75t_L       g17200(.A(\a[47] ), .B(new_n17456), .Y(new_n17457));
  NOR2xp33_ASAP7_75t_L      g17201(.A(new_n17457), .B(new_n17454), .Y(new_n17458));
  INVx1_ASAP7_75t_L         g17202(.A(new_n17458), .Y(new_n17459));
  NAND2xp33_ASAP7_75t_L     g17203(.A(new_n17457), .B(new_n17454), .Y(new_n17460));
  AND2x2_ASAP7_75t_L        g17204(.A(new_n17460), .B(new_n17459), .Y(new_n17461));
  NOR2xp33_ASAP7_75t_L      g17205(.A(new_n17392), .B(new_n17461), .Y(new_n17462));
  A2O1A1Ixp33_ASAP7_75t_L   g17206(.A1(new_n17322), .A2(new_n17320), .B(new_n17331), .C(new_n17461), .Y(new_n17463));
  INVx1_ASAP7_75t_L         g17207(.A(new_n17463), .Y(new_n17464));
  OAI21xp33_ASAP7_75t_L     g17208(.A1(new_n17462), .A2(new_n17464), .B(new_n17391), .Y(new_n17465));
  INVx1_ASAP7_75t_L         g17209(.A(new_n17391), .Y(new_n17466));
  NOR2xp33_ASAP7_75t_L      g17210(.A(new_n17462), .B(new_n17464), .Y(new_n17467));
  NAND2xp33_ASAP7_75t_L     g17211(.A(new_n17466), .B(new_n17467), .Y(new_n17468));
  AND2x2_ASAP7_75t_L        g17212(.A(new_n17465), .B(new_n17468), .Y(new_n17469));
  INVx1_ASAP7_75t_L         g17213(.A(new_n17469), .Y(new_n17470));
  O2A1O1Ixp33_ASAP7_75t_L   g17214(.A1(new_n17266), .A2(new_n17336), .B(new_n17334), .C(new_n17470), .Y(new_n17471));
  INVx1_ASAP7_75t_L         g17215(.A(new_n17471), .Y(new_n17472));
  NAND3xp33_ASAP7_75t_L     g17216(.A(new_n17470), .B(new_n17338), .C(new_n17334), .Y(new_n17473));
  NAND2xp33_ASAP7_75t_L     g17217(.A(new_n17473), .B(new_n17472), .Y(new_n17474));
  AOI22xp33_ASAP7_75t_L     g17218(.A1(new_n4920), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n5167), .Y(new_n17475));
  OAI221xp5_ASAP7_75t_L     g17219(.A1(new_n5154), .A2(new_n9323), .B1(new_n5158), .B2(new_n9627), .C(new_n17475), .Y(new_n17476));
  XNOR2x2_ASAP7_75t_L       g17220(.A(\a[41] ), .B(new_n17476), .Y(new_n17477));
  XNOR2x2_ASAP7_75t_L       g17221(.A(new_n17477), .B(new_n17474), .Y(new_n17478));
  NAND3xp33_ASAP7_75t_L     g17222(.A(new_n17478), .B(new_n17345), .C(new_n17342), .Y(new_n17479));
  AO21x2_ASAP7_75t_L        g17223(.A1(new_n17342), .A2(new_n17345), .B(new_n17478), .Y(new_n17480));
  AND2x2_ASAP7_75t_L        g17224(.A(new_n17479), .B(new_n17480), .Y(new_n17481));
  AOI22xp33_ASAP7_75t_L     g17225(.A1(new_n4283), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n4512), .Y(new_n17482));
  OAI221xp5_ASAP7_75t_L     g17226(.A1(new_n4277), .A2(new_n9947), .B1(new_n4499), .B2(new_n11446), .C(new_n17482), .Y(new_n17483));
  XNOR2x2_ASAP7_75t_L       g17227(.A(\a[38] ), .B(new_n17483), .Y(new_n17484));
  INVx1_ASAP7_75t_L         g17228(.A(new_n17484), .Y(new_n17485));
  XNOR2x2_ASAP7_75t_L       g17229(.A(new_n17485), .B(new_n17481), .Y(new_n17486));
  A2O1A1Ixp33_ASAP7_75t_L   g17230(.A1(new_n17353), .A2(new_n17348), .B(new_n17349), .C(new_n17486), .Y(new_n17487));
  A2O1A1Ixp33_ASAP7_75t_L   g17231(.A1(new_n17345), .A2(new_n17346), .B(new_n17259), .C(new_n17354), .Y(new_n17488));
  OR2x4_ASAP7_75t_L         g17232(.A(new_n17488), .B(new_n17486), .Y(new_n17489));
  AOI22xp33_ASAP7_75t_L     g17233(.A1(new_n3633), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n3858), .Y(new_n17490));
  A2O1A1Ixp33_ASAP7_75t_L   g17234(.A1(new_n11470), .A2(new_n11473), .B(new_n3856), .C(new_n17490), .Y(new_n17491));
  AOI21xp33_ASAP7_75t_L     g17235(.A1(new_n3639), .A2(\b[62] ), .B(new_n17491), .Y(new_n17492));
  NAND2xp33_ASAP7_75t_L     g17236(.A(\a[35] ), .B(new_n17492), .Y(new_n17493));
  A2O1A1Ixp33_ASAP7_75t_L   g17237(.A1(\b[62] ), .A2(new_n3639), .B(new_n17491), .C(new_n3628), .Y(new_n17494));
  NAND2xp33_ASAP7_75t_L     g17238(.A(new_n17494), .B(new_n17493), .Y(new_n17495));
  INVx1_ASAP7_75t_L         g17239(.A(new_n17356), .Y(new_n17496));
  A2O1A1O1Ixp25_ASAP7_75t_L g17240(.A1(new_n17226), .A2(new_n17229), .B(new_n17224), .C(new_n17496), .D(new_n17363), .Y(new_n17497));
  NAND2xp33_ASAP7_75t_L     g17241(.A(new_n17495), .B(new_n17497), .Y(new_n17498));
  INVx1_ASAP7_75t_L         g17242(.A(new_n17495), .Y(new_n17499));
  A2O1A1Ixp33_ASAP7_75t_L   g17243(.A1(new_n17359), .A2(new_n17362), .B(new_n17357), .C(new_n17499), .Y(new_n17500));
  AO22x1_ASAP7_75t_L        g17244(.A1(new_n17487), .A2(new_n17489), .B1(new_n17500), .B2(new_n17498), .Y(new_n17501));
  NAND4xp25_ASAP7_75t_L     g17245(.A(new_n17498), .B(new_n17487), .C(new_n17489), .D(new_n17500), .Y(new_n17502));
  NAND2xp33_ASAP7_75t_L     g17246(.A(new_n17502), .B(new_n17501), .Y(new_n17503));
  A2O1A1O1Ixp25_ASAP7_75t_L g17247(.A1(new_n17365), .A2(new_n17364), .B(new_n17388), .C(new_n17373), .D(new_n17503), .Y(new_n17504));
  INVx1_ASAP7_75t_L         g17248(.A(new_n17504), .Y(new_n17505));
  A2O1A1Ixp33_ASAP7_75t_L   g17249(.A1(new_n17364), .A2(new_n17365), .B(new_n17388), .C(new_n17373), .Y(new_n17506));
  AO21x2_ASAP7_75t_L        g17250(.A1(new_n17502), .A2(new_n17501), .B(new_n17506), .Y(new_n17507));
  NAND2xp33_ASAP7_75t_L     g17251(.A(new_n17507), .B(new_n17505), .Y(new_n17508));
  A2O1A1O1Ixp25_ASAP7_75t_L g17252(.A1(new_n17387), .A2(new_n17253), .B(new_n17381), .C(new_n17379), .D(new_n17508), .Y(new_n17509));
  A2O1A1Ixp33_ASAP7_75t_L   g17253(.A1(new_n17253), .A2(new_n17387), .B(new_n17381), .C(new_n17379), .Y(new_n17510));
  INVx1_ASAP7_75t_L         g17254(.A(new_n17508), .Y(new_n17511));
  NOR2xp33_ASAP7_75t_L      g17255(.A(new_n17511), .B(new_n17510), .Y(new_n17512));
  NOR2xp33_ASAP7_75t_L      g17256(.A(new_n17509), .B(new_n17512), .Y(\f[96] ));
  INVx1_ASAP7_75t_L         g17257(.A(new_n17497), .Y(new_n17514));
  NAND2xp33_ASAP7_75t_L     g17258(.A(new_n17485), .B(new_n17481), .Y(new_n17515));
  NOR2xp33_ASAP7_75t_L      g17259(.A(new_n11172), .B(new_n4052), .Y(new_n17516));
  AOI221xp5_ASAP7_75t_L     g17260(.A1(\b[63] ), .A2(new_n3639), .B1(new_n3630), .B2(new_n12322), .C(new_n17516), .Y(new_n17517));
  XNOR2x2_ASAP7_75t_L       g17261(.A(new_n3628), .B(new_n17517), .Y(new_n17518));
  O2A1O1Ixp33_ASAP7_75t_L   g17262(.A1(new_n17488), .A2(new_n17486), .B(new_n17515), .C(new_n17518), .Y(new_n17519));
  AND3x1_ASAP7_75t_L        g17263(.A(new_n17489), .B(new_n17518), .C(new_n17515), .Y(new_n17520));
  NOR2xp33_ASAP7_75t_L      g17264(.A(new_n17519), .B(new_n17520), .Y(new_n17521));
  INVx1_ASAP7_75t_L         g17265(.A(new_n17521), .Y(new_n17522));
  AOI22xp33_ASAP7_75t_L     g17266(.A1(new_n9700), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n10027), .Y(new_n17523));
  OAI221xp5_ASAP7_75t_L     g17267(.A1(new_n10024), .A2(new_n4848), .B1(new_n9696), .B2(new_n11686), .C(new_n17523), .Y(new_n17524));
  XNOR2x2_ASAP7_75t_L       g17268(.A(\a[59] ), .B(new_n17524), .Y(new_n17525));
  INVx1_ASAP7_75t_L         g17269(.A(new_n17525), .Y(new_n17526));
  NOR2xp33_ASAP7_75t_L      g17270(.A(new_n3565), .B(new_n11535), .Y(new_n17527));
  A2O1A1O1Ixp25_ASAP7_75t_L g17271(.A1(new_n11533), .A2(\b[32] ), .B(new_n17283), .C(new_n17406), .D(new_n17404), .Y(new_n17528));
  A2O1A1Ixp33_ASAP7_75t_L   g17272(.A1(new_n11533), .A2(\b[34] ), .B(new_n17527), .C(new_n17528), .Y(new_n17529));
  O2A1O1Ixp33_ASAP7_75t_L   g17273(.A1(new_n11247), .A2(new_n11249), .B(\b[34] ), .C(new_n17527), .Y(new_n17530));
  INVx1_ASAP7_75t_L         g17274(.A(new_n17530), .Y(new_n17531));
  O2A1O1Ixp33_ASAP7_75t_L   g17275(.A1(new_n17285), .A2(new_n17407), .B(new_n17403), .C(new_n17531), .Y(new_n17532));
  INVx1_ASAP7_75t_L         g17276(.A(new_n17532), .Y(new_n17533));
  NAND2xp33_ASAP7_75t_L     g17277(.A(new_n17529), .B(new_n17533), .Y(new_n17534));
  NAND2xp33_ASAP7_75t_L     g17278(.A(\b[35] ), .B(new_n10939), .Y(new_n17535));
  OAI221xp5_ASAP7_75t_L     g17279(.A1(new_n10630), .A2(new_n4424), .B1(new_n10629), .B2(new_n4431), .C(new_n17535), .Y(new_n17536));
  AOI21xp33_ASAP7_75t_L     g17280(.A1(new_n10632), .A2(\b[36] ), .B(new_n17536), .Y(new_n17537));
  NAND2xp33_ASAP7_75t_L     g17281(.A(\a[62] ), .B(new_n17537), .Y(new_n17538));
  A2O1A1Ixp33_ASAP7_75t_L   g17282(.A1(\b[36] ), .A2(new_n10632), .B(new_n17536), .C(new_n10622), .Y(new_n17539));
  AND2x2_ASAP7_75t_L        g17283(.A(new_n17539), .B(new_n17538), .Y(new_n17540));
  XOR2x2_ASAP7_75t_L        g17284(.A(new_n17534), .B(new_n17540), .Y(new_n17541));
  INVx1_ASAP7_75t_L         g17285(.A(new_n17541), .Y(new_n17542));
  O2A1O1Ixp33_ASAP7_75t_L   g17286(.A1(new_n17399), .A2(new_n17413), .B(new_n17410), .C(new_n17542), .Y(new_n17543));
  INVx1_ASAP7_75t_L         g17287(.A(new_n17543), .Y(new_n17544));
  NOR2xp33_ASAP7_75t_L      g17288(.A(new_n17411), .B(new_n17416), .Y(new_n17545));
  NAND2xp33_ASAP7_75t_L     g17289(.A(new_n17542), .B(new_n17545), .Y(new_n17546));
  NAND3xp33_ASAP7_75t_L     g17290(.A(new_n17546), .B(new_n17544), .C(new_n17526), .Y(new_n17547));
  AO21x2_ASAP7_75t_L        g17291(.A1(new_n17544), .A2(new_n17546), .B(new_n17526), .Y(new_n17548));
  AND2x2_ASAP7_75t_L        g17292(.A(new_n17547), .B(new_n17548), .Y(new_n17549));
  A2O1A1Ixp33_ASAP7_75t_L   g17293(.A1(new_n17419), .A2(new_n17396), .B(new_n17425), .C(new_n17549), .Y(new_n17550));
  INVx1_ASAP7_75t_L         g17294(.A(new_n17294), .Y(new_n17551));
  A2O1A1Ixp33_ASAP7_75t_L   g17295(.A1(new_n17291), .A2(new_n17551), .B(new_n17422), .C(new_n17420), .Y(new_n17552));
  NOR2xp33_ASAP7_75t_L      g17296(.A(new_n17552), .B(new_n17549), .Y(new_n17553));
  INVx1_ASAP7_75t_L         g17297(.A(new_n17553), .Y(new_n17554));
  AOI22xp33_ASAP7_75t_L     g17298(.A1(new_n8831), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n9115), .Y(new_n17555));
  OAI221xp5_ASAP7_75t_L     g17299(.A1(new_n10343), .A2(new_n5338), .B1(new_n10016), .B2(new_n6338), .C(new_n17555), .Y(new_n17556));
  XNOR2x2_ASAP7_75t_L       g17300(.A(\a[56] ), .B(new_n17556), .Y(new_n17557));
  NAND3xp33_ASAP7_75t_L     g17301(.A(new_n17554), .B(new_n17550), .C(new_n17557), .Y(new_n17558));
  AO21x2_ASAP7_75t_L        g17302(.A1(new_n17554), .A2(new_n17550), .B(new_n17557), .Y(new_n17559));
  AND2x2_ASAP7_75t_L        g17303(.A(new_n17558), .B(new_n17559), .Y(new_n17560));
  INVx1_ASAP7_75t_L         g17304(.A(new_n17560), .Y(new_n17561));
  NAND2xp33_ASAP7_75t_L     g17305(.A(new_n17431), .B(new_n17427), .Y(new_n17562));
  A2O1A1Ixp33_ASAP7_75t_L   g17306(.A1(new_n17301), .A2(new_n17299), .B(new_n17432), .C(new_n17562), .Y(new_n17563));
  NOR2xp33_ASAP7_75t_L      g17307(.A(new_n17563), .B(new_n17561), .Y(new_n17564));
  INVx1_ASAP7_75t_L         g17308(.A(new_n17564), .Y(new_n17565));
  O2A1O1Ixp33_ASAP7_75t_L   g17309(.A1(new_n17434), .A2(new_n17432), .B(new_n17562), .C(new_n17560), .Y(new_n17566));
  INVx1_ASAP7_75t_L         g17310(.A(new_n17566), .Y(new_n17567));
  AOI22xp33_ASAP7_75t_L     g17311(.A1(new_n7960), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n8537), .Y(new_n17568));
  OAI221xp5_ASAP7_75t_L     g17312(.A1(new_n8817), .A2(new_n6321), .B1(new_n7957), .B2(new_n6573), .C(new_n17568), .Y(new_n17569));
  XNOR2x2_ASAP7_75t_L       g17313(.A(\a[53] ), .B(new_n17569), .Y(new_n17570));
  NAND3xp33_ASAP7_75t_L     g17314(.A(new_n17565), .B(new_n17567), .C(new_n17570), .Y(new_n17571));
  AO21x2_ASAP7_75t_L        g17315(.A1(new_n17567), .A2(new_n17565), .B(new_n17570), .Y(new_n17572));
  AND2x2_ASAP7_75t_L        g17316(.A(new_n17571), .B(new_n17572), .Y(new_n17573));
  INVx1_ASAP7_75t_L         g17317(.A(new_n17573), .Y(new_n17574));
  NAND2xp33_ASAP7_75t_L     g17318(.A(new_n17441), .B(new_n17437), .Y(new_n17575));
  A2O1A1Ixp33_ASAP7_75t_L   g17319(.A1(new_n17307), .A2(new_n17304), .B(new_n17442), .C(new_n17575), .Y(new_n17576));
  NOR2xp33_ASAP7_75t_L      g17320(.A(new_n17576), .B(new_n17574), .Y(new_n17577));
  O2A1O1Ixp33_ASAP7_75t_L   g17321(.A1(new_n17443), .A2(new_n17442), .B(new_n17575), .C(new_n17573), .Y(new_n17578));
  NOR2xp33_ASAP7_75t_L      g17322(.A(new_n17578), .B(new_n17577), .Y(new_n17579));
  AOI22xp33_ASAP7_75t_L     g17323(.A1(new_n7111), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n7391), .Y(new_n17580));
  OAI221xp5_ASAP7_75t_L     g17324(.A1(new_n8558), .A2(new_n6830), .B1(new_n8237), .B2(new_n7323), .C(new_n17580), .Y(new_n17581));
  XNOR2x2_ASAP7_75t_L       g17325(.A(\a[50] ), .B(new_n17581), .Y(new_n17582));
  NAND2xp33_ASAP7_75t_L     g17326(.A(new_n17582), .B(new_n17579), .Y(new_n17583));
  INVx1_ASAP7_75t_L         g17327(.A(new_n17583), .Y(new_n17584));
  NOR2xp33_ASAP7_75t_L      g17328(.A(new_n17582), .B(new_n17579), .Y(new_n17585));
  NOR2xp33_ASAP7_75t_L      g17329(.A(new_n17585), .B(new_n17584), .Y(new_n17586));
  INVx1_ASAP7_75t_L         g17330(.A(new_n17586), .Y(new_n17587));
  AOI21xp33_ASAP7_75t_L     g17331(.A1(new_n17448), .A2(new_n17444), .B(new_n17452), .Y(new_n17588));
  INVx1_ASAP7_75t_L         g17332(.A(new_n17588), .Y(new_n17589));
  NOR2xp33_ASAP7_75t_L      g17333(.A(new_n17589), .B(new_n17587), .Y(new_n17590));
  INVx1_ASAP7_75t_L         g17334(.A(new_n17590), .Y(new_n17591));
  A2O1A1Ixp33_ASAP7_75t_L   g17335(.A1(new_n17448), .A2(new_n17444), .B(new_n17452), .C(new_n17587), .Y(new_n17592));
  AOI22xp33_ASAP7_75t_L     g17336(.A1(new_n6376), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n6648), .Y(new_n17593));
  OAI221xp5_ASAP7_75t_L     g17337(.A1(new_n6646), .A2(new_n7616), .B1(new_n6636), .B2(new_n7906), .C(new_n17593), .Y(new_n17594));
  XNOR2x2_ASAP7_75t_L       g17338(.A(\a[47] ), .B(new_n17594), .Y(new_n17595));
  NAND3xp33_ASAP7_75t_L     g17339(.A(new_n17591), .B(new_n17592), .C(new_n17595), .Y(new_n17596));
  AO21x2_ASAP7_75t_L        g17340(.A1(new_n17592), .A2(new_n17591), .B(new_n17595), .Y(new_n17597));
  AND2x2_ASAP7_75t_L        g17341(.A(new_n17596), .B(new_n17597), .Y(new_n17598));
  A2O1A1Ixp33_ASAP7_75t_L   g17342(.A1(new_n17460), .A2(new_n17392), .B(new_n17458), .C(new_n17598), .Y(new_n17599));
  INVx1_ASAP7_75t_L         g17343(.A(new_n17598), .Y(new_n17600));
  O2A1O1Ixp33_ASAP7_75t_L   g17344(.A1(new_n17324), .A2(new_n17331), .B(new_n17460), .C(new_n17458), .Y(new_n17601));
  NAND2xp33_ASAP7_75t_L     g17345(.A(new_n17601), .B(new_n17600), .Y(new_n17602));
  AND2x2_ASAP7_75t_L        g17346(.A(new_n17599), .B(new_n17602), .Y(new_n17603));
  NAND2xp33_ASAP7_75t_L     g17347(.A(\b[53] ), .B(new_n5901), .Y(new_n17604));
  OAI221xp5_ASAP7_75t_L     g17348(.A1(new_n5894), .A2(new_n8762), .B1(new_n5892), .B2(new_n8768), .C(new_n17604), .Y(new_n17605));
  AOI21xp33_ASAP7_75t_L     g17349(.A1(new_n5628), .A2(\b[54] ), .B(new_n17605), .Y(new_n17606));
  NAND2xp33_ASAP7_75t_L     g17350(.A(\a[44] ), .B(new_n17606), .Y(new_n17607));
  A2O1A1Ixp33_ASAP7_75t_L   g17351(.A1(\b[54] ), .A2(new_n5628), .B(new_n17605), .C(new_n5619), .Y(new_n17608));
  AND2x2_ASAP7_75t_L        g17352(.A(new_n17608), .B(new_n17607), .Y(new_n17609));
  INVx1_ASAP7_75t_L         g17353(.A(new_n17609), .Y(new_n17610));
  XNOR2x2_ASAP7_75t_L       g17354(.A(new_n17610), .B(new_n17603), .Y(new_n17611));
  A2O1A1Ixp33_ASAP7_75t_L   g17355(.A1(new_n17467), .A2(new_n17466), .B(new_n17471), .C(new_n17611), .Y(new_n17612));
  A2O1A1Ixp33_ASAP7_75t_L   g17356(.A1(new_n17334), .A2(new_n17338), .B(new_n17470), .C(new_n17468), .Y(new_n17613));
  NOR2xp33_ASAP7_75t_L      g17357(.A(new_n17613), .B(new_n17611), .Y(new_n17614));
  INVx1_ASAP7_75t_L         g17358(.A(new_n17614), .Y(new_n17615));
  AOI22xp33_ASAP7_75t_L     g17359(.A1(new_n4920), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n5167), .Y(new_n17616));
  OAI221xp5_ASAP7_75t_L     g17360(.A1(new_n5154), .A2(new_n9620), .B1(new_n5158), .B2(new_n9925), .C(new_n17616), .Y(new_n17617));
  XNOR2x2_ASAP7_75t_L       g17361(.A(\a[41] ), .B(new_n17617), .Y(new_n17618));
  NAND3xp33_ASAP7_75t_L     g17362(.A(new_n17615), .B(new_n17612), .C(new_n17618), .Y(new_n17619));
  AO21x2_ASAP7_75t_L        g17363(.A1(new_n17612), .A2(new_n17615), .B(new_n17618), .Y(new_n17620));
  NAND2xp33_ASAP7_75t_L     g17364(.A(new_n17619), .B(new_n17620), .Y(new_n17621));
  OAI21xp33_ASAP7_75t_L     g17365(.A1(new_n17474), .A2(new_n17477), .B(new_n17480), .Y(new_n17622));
  NOR2xp33_ASAP7_75t_L      g17366(.A(new_n17621), .B(new_n17622), .Y(new_n17623));
  NAND2xp33_ASAP7_75t_L     g17367(.A(new_n17621), .B(new_n17622), .Y(new_n17624));
  INVx1_ASAP7_75t_L         g17368(.A(new_n17624), .Y(new_n17625));
  NOR2xp33_ASAP7_75t_L      g17369(.A(new_n17623), .B(new_n17625), .Y(new_n17626));
  NAND2xp33_ASAP7_75t_L     g17370(.A(\b[59] ), .B(new_n4512), .Y(new_n17627));
  OAI221xp5_ASAP7_75t_L     g17371(.A1(new_n4275), .A2(new_n10847), .B1(new_n4499), .B2(new_n10855), .C(new_n17627), .Y(new_n17628));
  AOI21xp33_ASAP7_75t_L     g17372(.A1(new_n4285), .A2(\b[60] ), .B(new_n17628), .Y(new_n17629));
  NAND2xp33_ASAP7_75t_L     g17373(.A(\a[38] ), .B(new_n17629), .Y(new_n17630));
  A2O1A1Ixp33_ASAP7_75t_L   g17374(.A1(\b[60] ), .A2(new_n4285), .B(new_n17628), .C(new_n4268), .Y(new_n17631));
  NAND2xp33_ASAP7_75t_L     g17375(.A(new_n17631), .B(new_n17630), .Y(new_n17632));
  NAND2xp33_ASAP7_75t_L     g17376(.A(new_n17632), .B(new_n17626), .Y(new_n17633));
  INVx1_ASAP7_75t_L         g17377(.A(new_n17633), .Y(new_n17634));
  NOR2xp33_ASAP7_75t_L      g17378(.A(new_n17632), .B(new_n17626), .Y(new_n17635));
  NOR2xp33_ASAP7_75t_L      g17379(.A(new_n17635), .B(new_n17634), .Y(new_n17636));
  INVx1_ASAP7_75t_L         g17380(.A(new_n17636), .Y(new_n17637));
  NOR2xp33_ASAP7_75t_L      g17381(.A(new_n17637), .B(new_n17522), .Y(new_n17638));
  INVx1_ASAP7_75t_L         g17382(.A(new_n17638), .Y(new_n17639));
  NAND2xp33_ASAP7_75t_L     g17383(.A(new_n17637), .B(new_n17522), .Y(new_n17640));
  NAND2xp33_ASAP7_75t_L     g17384(.A(new_n17640), .B(new_n17639), .Y(new_n17641));
  O2A1O1Ixp33_ASAP7_75t_L   g17385(.A1(new_n17499), .A2(new_n17514), .B(new_n17502), .C(new_n17641), .Y(new_n17642));
  A2O1A1Ixp33_ASAP7_75t_L   g17386(.A1(new_n17494), .A2(new_n17493), .B(new_n17514), .C(new_n17502), .Y(new_n17643));
  AOI21xp33_ASAP7_75t_L     g17387(.A1(new_n17640), .A2(new_n17639), .B(new_n17643), .Y(new_n17644));
  NOR2xp33_ASAP7_75t_L      g17388(.A(new_n17644), .B(new_n17642), .Y(new_n17645));
  A2O1A1Ixp33_ASAP7_75t_L   g17389(.A1(new_n17510), .A2(new_n17511), .B(new_n17504), .C(new_n17645), .Y(new_n17646));
  INVx1_ASAP7_75t_L         g17390(.A(new_n17646), .Y(new_n17647));
  A2O1A1Ixp33_ASAP7_75t_L   g17391(.A1(new_n17383), .A2(new_n17379), .B(new_n17508), .C(new_n17505), .Y(new_n17648));
  NOR2xp33_ASAP7_75t_L      g17392(.A(new_n17645), .B(new_n17648), .Y(new_n17649));
  NOR2xp33_ASAP7_75t_L      g17393(.A(new_n17649), .B(new_n17647), .Y(\f[97] ));
  INVx1_ASAP7_75t_L         g17394(.A(new_n17603), .Y(new_n17651));
  O2A1O1Ixp33_ASAP7_75t_L   g17395(.A1(new_n17454), .A2(new_n17457), .B(new_n17463), .C(new_n17598), .Y(new_n17652));
  AOI22xp33_ASAP7_75t_L     g17396(.A1(new_n5624), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n5901), .Y(new_n17653));
  OAI221xp5_ASAP7_75t_L     g17397(.A1(new_n5900), .A2(new_n8762), .B1(new_n5892), .B2(new_n9331), .C(new_n17653), .Y(new_n17654));
  XNOR2x2_ASAP7_75t_L       g17398(.A(\a[44] ), .B(new_n17654), .Y(new_n17655));
  INVx1_ASAP7_75t_L         g17399(.A(new_n17655), .Y(new_n17656));
  AOI22xp33_ASAP7_75t_L     g17400(.A1(new_n6376), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n6648), .Y(new_n17657));
  OAI221xp5_ASAP7_75t_L     g17401(.A1(new_n6646), .A2(new_n7900), .B1(new_n6636), .B2(new_n8174), .C(new_n17657), .Y(new_n17658));
  XNOR2x2_ASAP7_75t_L       g17402(.A(\a[47] ), .B(new_n17658), .Y(new_n17659));
  INVx1_ASAP7_75t_L         g17403(.A(new_n17659), .Y(new_n17660));
  AOI22xp33_ASAP7_75t_L     g17404(.A1(new_n8831), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n9115), .Y(new_n17661));
  OAI221xp5_ASAP7_75t_L     g17405(.A1(new_n10343), .A2(new_n5805), .B1(new_n10016), .B2(new_n5835), .C(new_n17661), .Y(new_n17662));
  XNOR2x2_ASAP7_75t_L       g17406(.A(\a[56] ), .B(new_n17662), .Y(new_n17663));
  INVx1_ASAP7_75t_L         g17407(.A(new_n17663), .Y(new_n17664));
  AOI22xp33_ASAP7_75t_L     g17408(.A1(new_n9700), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n10027), .Y(new_n17665));
  OAI221xp5_ASAP7_75t_L     g17409(.A1(new_n10024), .A2(new_n4869), .B1(new_n9696), .B2(new_n5327), .C(new_n17665), .Y(new_n17666));
  XNOR2x2_ASAP7_75t_L       g17410(.A(\a[59] ), .B(new_n17666), .Y(new_n17667));
  AOI22xp33_ASAP7_75t_L     g17411(.A1(\b[36] ), .A2(new_n10939), .B1(\b[38] ), .B2(new_n10938), .Y(new_n17668));
  OAI221xp5_ASAP7_75t_L     g17412(.A1(new_n10937), .A2(new_n4424), .B1(new_n10629), .B2(new_n4641), .C(new_n17668), .Y(new_n17669));
  XNOR2x2_ASAP7_75t_L       g17413(.A(\a[62] ), .B(new_n17669), .Y(new_n17670));
  A2O1A1Ixp33_ASAP7_75t_L   g17414(.A1(new_n17538), .A2(new_n17539), .B(new_n17534), .C(new_n17533), .Y(new_n17671));
  NOR2xp33_ASAP7_75t_L      g17415(.A(new_n3584), .B(new_n11535), .Y(new_n17672));
  INVx1_ASAP7_75t_L         g17416(.A(new_n17672), .Y(new_n17673));
  O2A1O1Ixp33_ASAP7_75t_L   g17417(.A1(new_n11253), .A2(new_n3804), .B(new_n17673), .C(new_n17531), .Y(new_n17674));
  INVx1_ASAP7_75t_L         g17418(.A(new_n17674), .Y(new_n17675));
  O2A1O1Ixp33_ASAP7_75t_L   g17419(.A1(new_n11247), .A2(new_n11249), .B(\b[35] ), .C(new_n17672), .Y(new_n17676));
  A2O1A1Ixp33_ASAP7_75t_L   g17420(.A1(new_n11533), .A2(\b[34] ), .B(new_n17527), .C(new_n17676), .Y(new_n17677));
  NAND2xp33_ASAP7_75t_L     g17421(.A(new_n17677), .B(new_n17675), .Y(new_n17678));
  XNOR2x2_ASAP7_75t_L       g17422(.A(new_n17678), .B(new_n17671), .Y(new_n17679));
  INVx1_ASAP7_75t_L         g17423(.A(new_n17679), .Y(new_n17680));
  NOR2xp33_ASAP7_75t_L      g17424(.A(new_n17670), .B(new_n17680), .Y(new_n17681));
  INVx1_ASAP7_75t_L         g17425(.A(new_n17681), .Y(new_n17682));
  NAND2xp33_ASAP7_75t_L     g17426(.A(new_n17670), .B(new_n17680), .Y(new_n17683));
  NAND2xp33_ASAP7_75t_L     g17427(.A(new_n17683), .B(new_n17682), .Y(new_n17684));
  NOR2xp33_ASAP7_75t_L      g17428(.A(new_n17667), .B(new_n17684), .Y(new_n17685));
  INVx1_ASAP7_75t_L         g17429(.A(new_n17667), .Y(new_n17686));
  AOI21xp33_ASAP7_75t_L     g17430(.A1(new_n17682), .A2(new_n17683), .B(new_n17686), .Y(new_n17687));
  NOR2xp33_ASAP7_75t_L      g17431(.A(new_n17687), .B(new_n17685), .Y(new_n17688));
  INVx1_ASAP7_75t_L         g17432(.A(new_n17688), .Y(new_n17689));
  O2A1O1Ixp33_ASAP7_75t_L   g17433(.A1(new_n17545), .A2(new_n17542), .B(new_n17547), .C(new_n17689), .Y(new_n17690));
  INVx1_ASAP7_75t_L         g17434(.A(new_n17690), .Y(new_n17691));
  A2O1A1Ixp33_ASAP7_75t_L   g17435(.A1(new_n17417), .A2(new_n17410), .B(new_n17542), .C(new_n17547), .Y(new_n17692));
  INVx1_ASAP7_75t_L         g17436(.A(new_n17692), .Y(new_n17693));
  NAND2xp33_ASAP7_75t_L     g17437(.A(new_n17689), .B(new_n17693), .Y(new_n17694));
  NAND3xp33_ASAP7_75t_L     g17438(.A(new_n17694), .B(new_n17691), .C(new_n17664), .Y(new_n17695));
  INVx1_ASAP7_75t_L         g17439(.A(new_n17695), .Y(new_n17696));
  AOI21xp33_ASAP7_75t_L     g17440(.A1(new_n17694), .A2(new_n17691), .B(new_n17664), .Y(new_n17697));
  NOR2xp33_ASAP7_75t_L      g17441(.A(new_n17697), .B(new_n17696), .Y(new_n17698));
  NAND3xp33_ASAP7_75t_L     g17442(.A(new_n17558), .B(new_n17554), .C(new_n17698), .Y(new_n17699));
  O2A1O1Ixp33_ASAP7_75t_L   g17443(.A1(new_n17552), .A2(new_n17549), .B(new_n17558), .C(new_n17698), .Y(new_n17700));
  INVx1_ASAP7_75t_L         g17444(.A(new_n17700), .Y(new_n17701));
  AOI22xp33_ASAP7_75t_L     g17445(.A1(new_n7960), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n8537), .Y(new_n17702));
  OAI221xp5_ASAP7_75t_L     g17446(.A1(new_n8817), .A2(new_n6568), .B1(new_n7957), .B2(new_n6820), .C(new_n17702), .Y(new_n17703));
  XNOR2x2_ASAP7_75t_L       g17447(.A(\a[53] ), .B(new_n17703), .Y(new_n17704));
  NAND3xp33_ASAP7_75t_L     g17448(.A(new_n17701), .B(new_n17699), .C(new_n17704), .Y(new_n17705));
  AO21x2_ASAP7_75t_L        g17449(.A1(new_n17699), .A2(new_n17701), .B(new_n17704), .Y(new_n17706));
  AND2x2_ASAP7_75t_L        g17450(.A(new_n17705), .B(new_n17706), .Y(new_n17707));
  A2O1A1Ixp33_ASAP7_75t_L   g17451(.A1(new_n17567), .A2(new_n17570), .B(new_n17564), .C(new_n17707), .Y(new_n17708));
  NAND2xp33_ASAP7_75t_L     g17452(.A(new_n17565), .B(new_n17571), .Y(new_n17709));
  NOR2xp33_ASAP7_75t_L      g17453(.A(new_n17707), .B(new_n17709), .Y(new_n17710));
  INVx1_ASAP7_75t_L         g17454(.A(new_n17710), .Y(new_n17711));
  NAND2xp33_ASAP7_75t_L     g17455(.A(new_n17708), .B(new_n17711), .Y(new_n17712));
  AOI22xp33_ASAP7_75t_L     g17456(.A1(new_n7111), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n7391), .Y(new_n17713));
  OAI221xp5_ASAP7_75t_L     g17457(.A1(new_n8558), .A2(new_n7317), .B1(new_n8237), .B2(new_n7602), .C(new_n17713), .Y(new_n17714));
  XNOR2x2_ASAP7_75t_L       g17458(.A(\a[50] ), .B(new_n17714), .Y(new_n17715));
  NAND2xp33_ASAP7_75t_L     g17459(.A(new_n17715), .B(new_n17712), .Y(new_n17716));
  NOR2xp33_ASAP7_75t_L      g17460(.A(new_n17715), .B(new_n17712), .Y(new_n17717));
  INVx1_ASAP7_75t_L         g17461(.A(new_n17717), .Y(new_n17718));
  AND2x2_ASAP7_75t_L        g17462(.A(new_n17716), .B(new_n17718), .Y(new_n17719));
  INVx1_ASAP7_75t_L         g17463(.A(new_n17719), .Y(new_n17720));
  NOR2xp33_ASAP7_75t_L      g17464(.A(new_n17577), .B(new_n17584), .Y(new_n17721));
  INVx1_ASAP7_75t_L         g17465(.A(new_n17721), .Y(new_n17722));
  NOR2xp33_ASAP7_75t_L      g17466(.A(new_n17720), .B(new_n17722), .Y(new_n17723));
  O2A1O1Ixp33_ASAP7_75t_L   g17467(.A1(new_n17574), .A2(new_n17576), .B(new_n17583), .C(new_n17719), .Y(new_n17724));
  NOR2xp33_ASAP7_75t_L      g17468(.A(new_n17724), .B(new_n17723), .Y(new_n17725));
  NAND2xp33_ASAP7_75t_L     g17469(.A(new_n17660), .B(new_n17725), .Y(new_n17726));
  OAI21xp33_ASAP7_75t_L     g17470(.A1(new_n17724), .A2(new_n17723), .B(new_n17659), .Y(new_n17727));
  AND2x2_ASAP7_75t_L        g17471(.A(new_n17727), .B(new_n17726), .Y(new_n17728));
  AND3x1_ASAP7_75t_L        g17472(.A(new_n17728), .B(new_n17596), .C(new_n17591), .Y(new_n17729));
  O2A1O1Ixp33_ASAP7_75t_L   g17473(.A1(new_n17587), .A2(new_n17589), .B(new_n17596), .C(new_n17728), .Y(new_n17730));
  NOR2xp33_ASAP7_75t_L      g17474(.A(new_n17730), .B(new_n17729), .Y(new_n17731));
  NAND2xp33_ASAP7_75t_L     g17475(.A(new_n17656), .B(new_n17731), .Y(new_n17732));
  OAI21xp33_ASAP7_75t_L     g17476(.A1(new_n17730), .A2(new_n17729), .B(new_n17655), .Y(new_n17733));
  AND2x2_ASAP7_75t_L        g17477(.A(new_n17733), .B(new_n17732), .Y(new_n17734));
  A2O1A1Ixp33_ASAP7_75t_L   g17478(.A1(new_n17651), .A2(new_n17610), .B(new_n17652), .C(new_n17734), .Y(new_n17735));
  INVx1_ASAP7_75t_L         g17479(.A(new_n17652), .Y(new_n17736));
  A2O1A1Ixp33_ASAP7_75t_L   g17480(.A1(new_n17602), .A2(new_n17599), .B(new_n17609), .C(new_n17736), .Y(new_n17737));
  NOR2xp33_ASAP7_75t_L      g17481(.A(new_n17737), .B(new_n17734), .Y(new_n17738));
  INVx1_ASAP7_75t_L         g17482(.A(new_n17738), .Y(new_n17739));
  AOI22xp33_ASAP7_75t_L     g17483(.A1(new_n4920), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n5167), .Y(new_n17740));
  OAI221xp5_ASAP7_75t_L     g17484(.A1(new_n5154), .A2(new_n9920), .B1(new_n5158), .B2(new_n11152), .C(new_n17740), .Y(new_n17741));
  XNOR2x2_ASAP7_75t_L       g17485(.A(\a[41] ), .B(new_n17741), .Y(new_n17742));
  NAND3xp33_ASAP7_75t_L     g17486(.A(new_n17739), .B(new_n17735), .C(new_n17742), .Y(new_n17743));
  INVx1_ASAP7_75t_L         g17487(.A(new_n17743), .Y(new_n17744));
  AOI21xp33_ASAP7_75t_L     g17488(.A1(new_n17739), .A2(new_n17735), .B(new_n17742), .Y(new_n17745));
  NOR2xp33_ASAP7_75t_L      g17489(.A(new_n17745), .B(new_n17744), .Y(new_n17746));
  INVx1_ASAP7_75t_L         g17490(.A(new_n17746), .Y(new_n17747));
  O2A1O1Ixp33_ASAP7_75t_L   g17491(.A1(new_n17613), .A2(new_n17611), .B(new_n17619), .C(new_n17747), .Y(new_n17748));
  INVx1_ASAP7_75t_L         g17492(.A(new_n17748), .Y(new_n17749));
  NAND3xp33_ASAP7_75t_L     g17493(.A(new_n17747), .B(new_n17619), .C(new_n17615), .Y(new_n17750));
  AOI22xp33_ASAP7_75t_L     g17494(.A1(new_n4283), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n4512), .Y(new_n17751));
  OAI221xp5_ASAP7_75t_L     g17495(.A1(new_n4277), .A2(new_n10847), .B1(new_n4499), .B2(new_n12047), .C(new_n17751), .Y(new_n17752));
  XNOR2x2_ASAP7_75t_L       g17496(.A(\a[38] ), .B(new_n17752), .Y(new_n17753));
  NAND3xp33_ASAP7_75t_L     g17497(.A(new_n17749), .B(new_n17750), .C(new_n17753), .Y(new_n17754));
  INVx1_ASAP7_75t_L         g17498(.A(new_n17754), .Y(new_n17755));
  AOI21xp33_ASAP7_75t_L     g17499(.A1(new_n17749), .A2(new_n17750), .B(new_n17753), .Y(new_n17756));
  NOR2xp33_ASAP7_75t_L      g17500(.A(new_n17756), .B(new_n17755), .Y(new_n17757));
  A2O1A1O1Ixp25_ASAP7_75t_L g17501(.A1(new_n3630), .A2(new_n12061), .B(new_n3858), .C(\b[63] ), .D(new_n3628), .Y(new_n17758));
  A2O1A1O1Ixp25_ASAP7_75t_L g17502(.A1(\b[61] ), .A2(new_n11471), .B(\b[62] ), .C(new_n3630), .D(new_n3858), .Y(new_n17759));
  NOR3xp33_ASAP7_75t_L      g17503(.A(new_n17759), .B(new_n11468), .C(\a[35] ), .Y(new_n17760));
  NOR2xp33_ASAP7_75t_L      g17504(.A(new_n17758), .B(new_n17760), .Y(new_n17761));
  A2O1A1O1Ixp25_ASAP7_75t_L g17505(.A1(new_n17630), .A2(new_n17631), .B(new_n17623), .C(new_n17624), .D(new_n17761), .Y(new_n17762));
  INVx1_ASAP7_75t_L         g17506(.A(new_n17762), .Y(new_n17763));
  NAND3xp33_ASAP7_75t_L     g17507(.A(new_n17633), .B(new_n17624), .C(new_n17761), .Y(new_n17764));
  NAND2xp33_ASAP7_75t_L     g17508(.A(new_n17763), .B(new_n17764), .Y(new_n17765));
  XNOR2x2_ASAP7_75t_L       g17509(.A(new_n17757), .B(new_n17765), .Y(new_n17766));
  A2O1A1O1Ixp25_ASAP7_75t_L g17510(.A1(new_n17515), .A2(new_n17489), .B(new_n17518), .C(new_n17639), .D(new_n17766), .Y(new_n17767));
  INVx1_ASAP7_75t_L         g17511(.A(new_n17767), .Y(new_n17768));
  NOR2xp33_ASAP7_75t_L      g17512(.A(new_n17519), .B(new_n17638), .Y(new_n17769));
  NAND2xp33_ASAP7_75t_L     g17513(.A(new_n17766), .B(new_n17769), .Y(new_n17770));
  AND2x2_ASAP7_75t_L        g17514(.A(new_n17770), .B(new_n17768), .Y(new_n17771));
  A2O1A1Ixp33_ASAP7_75t_L   g17515(.A1(new_n17648), .A2(new_n17645), .B(new_n17642), .C(new_n17771), .Y(new_n17772));
  A2O1A1O1Ixp25_ASAP7_75t_L g17516(.A1(new_n17511), .A2(new_n17510), .B(new_n17504), .C(new_n17645), .D(new_n17642), .Y(new_n17773));
  INVx1_ASAP7_75t_L         g17517(.A(new_n17771), .Y(new_n17774));
  NAND2xp33_ASAP7_75t_L     g17518(.A(new_n17774), .B(new_n17773), .Y(new_n17775));
  AND2x2_ASAP7_75t_L        g17519(.A(new_n17772), .B(new_n17775), .Y(\f[98] ));
  INVx1_ASAP7_75t_L         g17520(.A(new_n17642), .Y(new_n17777));
  INVx1_ASAP7_75t_L         g17521(.A(new_n17764), .Y(new_n17778));
  INVx1_ASAP7_75t_L         g17522(.A(new_n17729), .Y(new_n17779));
  AOI22xp33_ASAP7_75t_L     g17523(.A1(new_n6376), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n6648), .Y(new_n17780));
  OAI221xp5_ASAP7_75t_L     g17524(.A1(new_n6646), .A2(new_n8165), .B1(new_n6636), .B2(new_n8465), .C(new_n17780), .Y(new_n17781));
  XNOR2x2_ASAP7_75t_L       g17525(.A(\a[47] ), .B(new_n17781), .Y(new_n17782));
  INVx1_ASAP7_75t_L         g17526(.A(new_n17782), .Y(new_n17783));
  AOI22xp33_ASAP7_75t_L     g17527(.A1(new_n8831), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n9115), .Y(new_n17784));
  OAI221xp5_ASAP7_75t_L     g17528(.A1(new_n10343), .A2(new_n5829), .B1(new_n10016), .B2(new_n6329), .C(new_n17784), .Y(new_n17785));
  XNOR2x2_ASAP7_75t_L       g17529(.A(\a[56] ), .B(new_n17785), .Y(new_n17786));
  INVx1_ASAP7_75t_L         g17530(.A(new_n17786), .Y(new_n17787));
  NOR2xp33_ASAP7_75t_L      g17531(.A(new_n3804), .B(new_n11535), .Y(new_n17788));
  O2A1O1Ixp33_ASAP7_75t_L   g17532(.A1(new_n3804), .A2(new_n11253), .B(new_n17673), .C(new_n3628), .Y(new_n17789));
  AOI211xp5_ASAP7_75t_L     g17533(.A1(new_n11533), .A2(\b[35] ), .B(new_n17672), .C(\a[35] ), .Y(new_n17790));
  NOR2xp33_ASAP7_75t_L      g17534(.A(new_n17790), .B(new_n17789), .Y(new_n17791));
  INVx1_ASAP7_75t_L         g17535(.A(new_n17791), .Y(new_n17792));
  A2O1A1Ixp33_ASAP7_75t_L   g17536(.A1(new_n11533), .A2(\b[36] ), .B(new_n17788), .C(new_n17792), .Y(new_n17793));
  O2A1O1Ixp33_ASAP7_75t_L   g17537(.A1(new_n11247), .A2(new_n11249), .B(\b[36] ), .C(new_n17788), .Y(new_n17794));
  NAND2xp33_ASAP7_75t_L     g17538(.A(new_n17794), .B(new_n17791), .Y(new_n17795));
  AND2x2_ASAP7_75t_L        g17539(.A(new_n17795), .B(new_n17793), .Y(new_n17796));
  A2O1A1O1Ixp25_ASAP7_75t_L g17540(.A1(new_n11533), .A2(\b[34] ), .B(new_n17527), .C(new_n17676), .D(new_n17671), .Y(new_n17797));
  A2O1A1O1Ixp25_ASAP7_75t_L g17541(.A1(new_n11533), .A2(\b[35] ), .B(new_n17672), .C(new_n17530), .D(new_n17797), .Y(new_n17798));
  NAND2xp33_ASAP7_75t_L     g17542(.A(new_n17796), .B(new_n17798), .Y(new_n17799));
  INVx1_ASAP7_75t_L         g17543(.A(new_n17799), .Y(new_n17800));
  INVx1_ASAP7_75t_L         g17544(.A(new_n17677), .Y(new_n17801));
  O2A1O1Ixp33_ASAP7_75t_L   g17545(.A1(new_n17801), .A2(new_n17671), .B(new_n17675), .C(new_n17796), .Y(new_n17802));
  NOR2xp33_ASAP7_75t_L      g17546(.A(new_n17802), .B(new_n17800), .Y(new_n17803));
  INVx1_ASAP7_75t_L         g17547(.A(new_n17803), .Y(new_n17804));
  AOI22xp33_ASAP7_75t_L     g17548(.A1(\b[37] ), .A2(new_n10939), .B1(\b[39] ), .B2(new_n10938), .Y(new_n17805));
  OAI221xp5_ASAP7_75t_L     g17549(.A1(new_n10937), .A2(new_n4632), .B1(new_n10629), .B2(new_n4858), .C(new_n17805), .Y(new_n17806));
  XNOR2x2_ASAP7_75t_L       g17550(.A(\a[62] ), .B(new_n17806), .Y(new_n17807));
  AND2x2_ASAP7_75t_L        g17551(.A(new_n17807), .B(new_n17804), .Y(new_n17808));
  NOR2xp33_ASAP7_75t_L      g17552(.A(new_n17807), .B(new_n17804), .Y(new_n17809));
  NOR2xp33_ASAP7_75t_L      g17553(.A(new_n17809), .B(new_n17808), .Y(new_n17810));
  AOI22xp33_ASAP7_75t_L     g17554(.A1(new_n9700), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n10027), .Y(new_n17811));
  OAI221xp5_ASAP7_75t_L     g17555(.A1(new_n10024), .A2(new_n5321), .B1(new_n9696), .B2(new_n5346), .C(new_n17811), .Y(new_n17812));
  XNOR2x2_ASAP7_75t_L       g17556(.A(\a[59] ), .B(new_n17812), .Y(new_n17813));
  INVx1_ASAP7_75t_L         g17557(.A(new_n17813), .Y(new_n17814));
  XNOR2x2_ASAP7_75t_L       g17558(.A(new_n17814), .B(new_n17810), .Y(new_n17815));
  O2A1O1Ixp33_ASAP7_75t_L   g17559(.A1(new_n17667), .A2(new_n17684), .B(new_n17682), .C(new_n17815), .Y(new_n17816));
  NOR2xp33_ASAP7_75t_L      g17560(.A(new_n17681), .B(new_n17685), .Y(new_n17817));
  AND2x2_ASAP7_75t_L        g17561(.A(new_n17817), .B(new_n17815), .Y(new_n17818));
  NOR2xp33_ASAP7_75t_L      g17562(.A(new_n17816), .B(new_n17818), .Y(new_n17819));
  XNOR2x2_ASAP7_75t_L       g17563(.A(new_n17787), .B(new_n17819), .Y(new_n17820));
  A2O1A1Ixp33_ASAP7_75t_L   g17564(.A1(new_n17547), .A2(new_n17544), .B(new_n17689), .C(new_n17695), .Y(new_n17821));
  INVx1_ASAP7_75t_L         g17565(.A(new_n17821), .Y(new_n17822));
  AND2x2_ASAP7_75t_L        g17566(.A(new_n17822), .B(new_n17820), .Y(new_n17823));
  O2A1O1Ixp33_ASAP7_75t_L   g17567(.A1(new_n17693), .A2(new_n17689), .B(new_n17695), .C(new_n17820), .Y(new_n17824));
  NOR2xp33_ASAP7_75t_L      g17568(.A(new_n17824), .B(new_n17823), .Y(new_n17825));
  AOI22xp33_ASAP7_75t_L     g17569(.A1(new_n7960), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n8537), .Y(new_n17826));
  OAI221xp5_ASAP7_75t_L     g17570(.A1(new_n8817), .A2(new_n6812), .B1(new_n7957), .B2(new_n6837), .C(new_n17826), .Y(new_n17827));
  XNOR2x2_ASAP7_75t_L       g17571(.A(\a[53] ), .B(new_n17827), .Y(new_n17828));
  INVx1_ASAP7_75t_L         g17572(.A(new_n17828), .Y(new_n17829));
  XNOR2x2_ASAP7_75t_L       g17573(.A(new_n17829), .B(new_n17825), .Y(new_n17830));
  A2O1A1Ixp33_ASAP7_75t_L   g17574(.A1(new_n17704), .A2(new_n17699), .B(new_n17700), .C(new_n17830), .Y(new_n17831));
  A2O1A1Ixp33_ASAP7_75t_L   g17575(.A1(new_n17558), .A2(new_n17554), .B(new_n17698), .C(new_n17705), .Y(new_n17832));
  NOR2xp33_ASAP7_75t_L      g17576(.A(new_n17832), .B(new_n17830), .Y(new_n17833));
  INVx1_ASAP7_75t_L         g17577(.A(new_n17833), .Y(new_n17834));
  NAND2xp33_ASAP7_75t_L     g17578(.A(new_n17831), .B(new_n17834), .Y(new_n17835));
  AOI22xp33_ASAP7_75t_L     g17579(.A1(new_n7111), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n7391), .Y(new_n17836));
  OAI221xp5_ASAP7_75t_L     g17580(.A1(new_n8558), .A2(new_n7593), .B1(new_n8237), .B2(new_n7623), .C(new_n17836), .Y(new_n17837));
  XNOR2x2_ASAP7_75t_L       g17581(.A(\a[50] ), .B(new_n17837), .Y(new_n17838));
  NAND2xp33_ASAP7_75t_L     g17582(.A(new_n17838), .B(new_n17835), .Y(new_n17839));
  NOR2xp33_ASAP7_75t_L      g17583(.A(new_n17838), .B(new_n17835), .Y(new_n17840));
  INVx1_ASAP7_75t_L         g17584(.A(new_n17840), .Y(new_n17841));
  AND2x2_ASAP7_75t_L        g17585(.A(new_n17839), .B(new_n17841), .Y(new_n17842));
  INVx1_ASAP7_75t_L         g17586(.A(new_n17842), .Y(new_n17843));
  O2A1O1Ixp33_ASAP7_75t_L   g17587(.A1(new_n17707), .A2(new_n17709), .B(new_n17718), .C(new_n17843), .Y(new_n17844));
  A2O1A1Ixp33_ASAP7_75t_L   g17588(.A1(new_n17706), .A2(new_n17705), .B(new_n17709), .C(new_n17718), .Y(new_n17845));
  NOR2xp33_ASAP7_75t_L      g17589(.A(new_n17842), .B(new_n17845), .Y(new_n17846));
  NOR2xp33_ASAP7_75t_L      g17590(.A(new_n17846), .B(new_n17844), .Y(new_n17847));
  NAND2xp33_ASAP7_75t_L     g17591(.A(new_n17783), .B(new_n17847), .Y(new_n17848));
  OAI21xp33_ASAP7_75t_L     g17592(.A1(new_n17846), .A2(new_n17844), .B(new_n17782), .Y(new_n17849));
  AND2x2_ASAP7_75t_L        g17593(.A(new_n17849), .B(new_n17848), .Y(new_n17850));
  A2O1A1Ixp33_ASAP7_75t_L   g17594(.A1(new_n17725), .A2(new_n17660), .B(new_n17723), .C(new_n17850), .Y(new_n17851));
  INVx1_ASAP7_75t_L         g17595(.A(new_n17726), .Y(new_n17852));
  OR3x1_ASAP7_75t_L         g17596(.A(new_n17852), .B(new_n17850), .C(new_n17723), .Y(new_n17853));
  NAND2xp33_ASAP7_75t_L     g17597(.A(new_n17851), .B(new_n17853), .Y(new_n17854));
  AOI22xp33_ASAP7_75t_L     g17598(.A1(new_n5624), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n5901), .Y(new_n17855));
  OAI221xp5_ASAP7_75t_L     g17599(.A1(new_n5900), .A2(new_n9323), .B1(new_n5892), .B2(new_n9627), .C(new_n17855), .Y(new_n17856));
  XNOR2x2_ASAP7_75t_L       g17600(.A(\a[44] ), .B(new_n17856), .Y(new_n17857));
  XNOR2x2_ASAP7_75t_L       g17601(.A(new_n17857), .B(new_n17854), .Y(new_n17858));
  AND3x1_ASAP7_75t_L        g17602(.A(new_n17858), .B(new_n17732), .C(new_n17779), .Y(new_n17859));
  O2A1O1Ixp33_ASAP7_75t_L   g17603(.A1(new_n17655), .A2(new_n17730), .B(new_n17779), .C(new_n17858), .Y(new_n17860));
  NOR2xp33_ASAP7_75t_L      g17604(.A(new_n17860), .B(new_n17859), .Y(new_n17861));
  AOI22xp33_ASAP7_75t_L     g17605(.A1(new_n4920), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n5167), .Y(new_n17862));
  OAI221xp5_ASAP7_75t_L     g17606(.A1(new_n5154), .A2(new_n9947), .B1(new_n5158), .B2(new_n11446), .C(new_n17862), .Y(new_n17863));
  XNOR2x2_ASAP7_75t_L       g17607(.A(\a[41] ), .B(new_n17863), .Y(new_n17864));
  INVx1_ASAP7_75t_L         g17608(.A(new_n17864), .Y(new_n17865));
  XNOR2x2_ASAP7_75t_L       g17609(.A(new_n17865), .B(new_n17861), .Y(new_n17866));
  A2O1A1Ixp33_ASAP7_75t_L   g17610(.A1(new_n17742), .A2(new_n17735), .B(new_n17738), .C(new_n17866), .Y(new_n17867));
  A2O1A1Ixp33_ASAP7_75t_L   g17611(.A1(new_n17732), .A2(new_n17733), .B(new_n17737), .C(new_n17743), .Y(new_n17868));
  NOR2xp33_ASAP7_75t_L      g17612(.A(new_n17866), .B(new_n17868), .Y(new_n17869));
  INVx1_ASAP7_75t_L         g17613(.A(new_n17869), .Y(new_n17870));
  NAND2xp33_ASAP7_75t_L     g17614(.A(new_n17867), .B(new_n17870), .Y(new_n17871));
  AOI22xp33_ASAP7_75t_L     g17615(.A1(new_n4283), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n4512), .Y(new_n17872));
  A2O1A1Ixp33_ASAP7_75t_L   g17616(.A1(new_n11470), .A2(new_n11473), .B(new_n4499), .C(new_n17872), .Y(new_n17873));
  AOI21xp33_ASAP7_75t_L     g17617(.A1(new_n4285), .A2(\b[62] ), .B(new_n17873), .Y(new_n17874));
  NAND2xp33_ASAP7_75t_L     g17618(.A(\a[38] ), .B(new_n17874), .Y(new_n17875));
  A2O1A1Ixp33_ASAP7_75t_L   g17619(.A1(\b[62] ), .A2(new_n4285), .B(new_n17873), .C(new_n4268), .Y(new_n17876));
  NAND2xp33_ASAP7_75t_L     g17620(.A(new_n17876), .B(new_n17875), .Y(new_n17877));
  XOR2x2_ASAP7_75t_L        g17621(.A(new_n17877), .B(new_n17871), .Y(new_n17878));
  A2O1A1Ixp33_ASAP7_75t_L   g17622(.A1(new_n17750), .A2(new_n17753), .B(new_n17748), .C(new_n17878), .Y(new_n17879));
  A2O1A1Ixp33_ASAP7_75t_L   g17623(.A1(new_n17619), .A2(new_n17615), .B(new_n17747), .C(new_n17754), .Y(new_n17880));
  NOR2xp33_ASAP7_75t_L      g17624(.A(new_n17878), .B(new_n17880), .Y(new_n17881));
  INVx1_ASAP7_75t_L         g17625(.A(new_n17881), .Y(new_n17882));
  NAND2xp33_ASAP7_75t_L     g17626(.A(new_n17879), .B(new_n17882), .Y(new_n17883));
  O2A1O1Ixp33_ASAP7_75t_L   g17627(.A1(new_n17757), .A2(new_n17778), .B(new_n17763), .C(new_n17883), .Y(new_n17884));
  INVx1_ASAP7_75t_L         g17628(.A(new_n17884), .Y(new_n17885));
  OAI211xp5_ASAP7_75t_L     g17629(.A1(new_n17757), .A2(new_n17778), .B(new_n17883), .C(new_n17763), .Y(new_n17886));
  AND2x2_ASAP7_75t_L        g17630(.A(new_n17886), .B(new_n17885), .Y(new_n17887));
  INVx1_ASAP7_75t_L         g17631(.A(new_n17887), .Y(new_n17888));
  A2O1A1O1Ixp25_ASAP7_75t_L g17632(.A1(new_n17777), .A2(new_n17646), .B(new_n17774), .C(new_n17768), .D(new_n17888), .Y(new_n17889));
  A2O1A1Ixp33_ASAP7_75t_L   g17633(.A1(new_n17646), .A2(new_n17777), .B(new_n17774), .C(new_n17768), .Y(new_n17890));
  NOR2xp33_ASAP7_75t_L      g17634(.A(new_n17887), .B(new_n17890), .Y(new_n17891));
  NOR2xp33_ASAP7_75t_L      g17635(.A(new_n17889), .B(new_n17891), .Y(\f[99] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17636(.A1(new_n17875), .A2(new_n17876), .B(new_n17871), .C(new_n17882), .Y(new_n17893));
  NOR2xp33_ASAP7_75t_L      g17637(.A(new_n11172), .B(new_n4501), .Y(new_n17894));
  AOI221xp5_ASAP7_75t_L     g17638(.A1(\b[63] ), .A2(new_n4285), .B1(new_n4274), .B2(new_n12322), .C(new_n17894), .Y(new_n17895));
  XNOR2x2_ASAP7_75t_L       g17639(.A(new_n4268), .B(new_n17895), .Y(new_n17896));
  INVx1_ASAP7_75t_L         g17640(.A(new_n17896), .Y(new_n17897));
  A2O1A1Ixp33_ASAP7_75t_L   g17641(.A1(new_n17865), .A2(new_n17861), .B(new_n17869), .C(new_n17897), .Y(new_n17898));
  AOI21xp33_ASAP7_75t_L     g17642(.A1(new_n17865), .A2(new_n17861), .B(new_n17869), .Y(new_n17899));
  NAND2xp33_ASAP7_75t_L     g17643(.A(new_n17896), .B(new_n17899), .Y(new_n17900));
  AND2x2_ASAP7_75t_L        g17644(.A(new_n17898), .B(new_n17900), .Y(new_n17901));
  NAND2xp33_ASAP7_75t_L     g17645(.A(new_n17848), .B(new_n17851), .Y(new_n17902));
  NAND2xp33_ASAP7_75t_L     g17646(.A(\b[38] ), .B(new_n10939), .Y(new_n17903));
  OAI221xp5_ASAP7_75t_L     g17647(.A1(new_n10630), .A2(new_n4869), .B1(new_n10629), .B2(new_n11686), .C(new_n17903), .Y(new_n17904));
  AOI21xp33_ASAP7_75t_L     g17648(.A1(new_n10632), .A2(\b[39] ), .B(new_n17904), .Y(new_n17905));
  NAND2xp33_ASAP7_75t_L     g17649(.A(\a[62] ), .B(new_n17905), .Y(new_n17906));
  A2O1A1Ixp33_ASAP7_75t_L   g17650(.A1(\b[39] ), .A2(new_n10632), .B(new_n17904), .C(new_n10622), .Y(new_n17907));
  NAND2xp33_ASAP7_75t_L     g17651(.A(new_n17907), .B(new_n17906), .Y(new_n17908));
  NOR2xp33_ASAP7_75t_L      g17652(.A(new_n4216), .B(new_n11535), .Y(new_n17909));
  O2A1O1Ixp33_ASAP7_75t_L   g17653(.A1(new_n11247), .A2(new_n11249), .B(\b[37] ), .C(new_n17909), .Y(new_n17910));
  INVx1_ASAP7_75t_L         g17654(.A(new_n17794), .Y(new_n17911));
  O2A1O1Ixp33_ASAP7_75t_L   g17655(.A1(new_n3804), .A2(new_n11253), .B(new_n17673), .C(\a[35] ), .Y(new_n17912));
  O2A1O1Ixp33_ASAP7_75t_L   g17656(.A1(new_n17790), .A2(new_n17789), .B(new_n17911), .C(new_n17912), .Y(new_n17913));
  NAND2xp33_ASAP7_75t_L     g17657(.A(new_n17910), .B(new_n17913), .Y(new_n17914));
  INVx1_ASAP7_75t_L         g17658(.A(new_n17910), .Y(new_n17915));
  A2O1A1Ixp33_ASAP7_75t_L   g17659(.A1(new_n17792), .A2(new_n17911), .B(new_n17912), .C(new_n17915), .Y(new_n17916));
  AND2x2_ASAP7_75t_L        g17660(.A(new_n17914), .B(new_n17916), .Y(new_n17917));
  XOR2x2_ASAP7_75t_L        g17661(.A(new_n17917), .B(new_n17908), .Y(new_n17918));
  INVx1_ASAP7_75t_L         g17662(.A(new_n17918), .Y(new_n17919));
  NOR2xp33_ASAP7_75t_L      g17663(.A(new_n17800), .B(new_n17809), .Y(new_n17920));
  INVx1_ASAP7_75t_L         g17664(.A(new_n17920), .Y(new_n17921));
  NOR2xp33_ASAP7_75t_L      g17665(.A(new_n17919), .B(new_n17921), .Y(new_n17922));
  INVx1_ASAP7_75t_L         g17666(.A(new_n17922), .Y(new_n17923));
  O2A1O1Ixp33_ASAP7_75t_L   g17667(.A1(new_n17802), .A2(new_n17807), .B(new_n17799), .C(new_n17918), .Y(new_n17924));
  INVx1_ASAP7_75t_L         g17668(.A(new_n17924), .Y(new_n17925));
  AOI22xp33_ASAP7_75t_L     g17669(.A1(new_n9700), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n10027), .Y(new_n17926));
  OAI221xp5_ASAP7_75t_L     g17670(.A1(new_n10024), .A2(new_n5338), .B1(new_n9696), .B2(new_n6338), .C(new_n17926), .Y(new_n17927));
  XNOR2x2_ASAP7_75t_L       g17671(.A(\a[59] ), .B(new_n17927), .Y(new_n17928));
  NAND3xp33_ASAP7_75t_L     g17672(.A(new_n17923), .B(new_n17925), .C(new_n17928), .Y(new_n17929));
  AO21x2_ASAP7_75t_L        g17673(.A1(new_n17925), .A2(new_n17923), .B(new_n17928), .Y(new_n17930));
  AND2x2_ASAP7_75t_L        g17674(.A(new_n17929), .B(new_n17930), .Y(new_n17931));
  INVx1_ASAP7_75t_L         g17675(.A(new_n17931), .Y(new_n17932));
  INVx1_ASAP7_75t_L         g17676(.A(new_n17685), .Y(new_n17933));
  NAND2xp33_ASAP7_75t_L     g17677(.A(new_n17814), .B(new_n17810), .Y(new_n17934));
  A2O1A1Ixp33_ASAP7_75t_L   g17678(.A1(new_n17933), .A2(new_n17682), .B(new_n17815), .C(new_n17934), .Y(new_n17935));
  NOR2xp33_ASAP7_75t_L      g17679(.A(new_n17935), .B(new_n17932), .Y(new_n17936));
  INVx1_ASAP7_75t_L         g17680(.A(new_n17936), .Y(new_n17937));
  O2A1O1Ixp33_ASAP7_75t_L   g17681(.A1(new_n17817), .A2(new_n17815), .B(new_n17934), .C(new_n17931), .Y(new_n17938));
  INVx1_ASAP7_75t_L         g17682(.A(new_n17938), .Y(new_n17939));
  AOI22xp33_ASAP7_75t_L     g17683(.A1(new_n8831), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n9115), .Y(new_n17940));
  OAI221xp5_ASAP7_75t_L     g17684(.A1(new_n10343), .A2(new_n6321), .B1(new_n10016), .B2(new_n6573), .C(new_n17940), .Y(new_n17941));
  XNOR2x2_ASAP7_75t_L       g17685(.A(\a[56] ), .B(new_n17941), .Y(new_n17942));
  NAND3xp33_ASAP7_75t_L     g17686(.A(new_n17937), .B(new_n17939), .C(new_n17942), .Y(new_n17943));
  AO21x2_ASAP7_75t_L        g17687(.A1(new_n17939), .A2(new_n17937), .B(new_n17942), .Y(new_n17944));
  AND2x2_ASAP7_75t_L        g17688(.A(new_n17943), .B(new_n17944), .Y(new_n17945));
  INVx1_ASAP7_75t_L         g17689(.A(new_n17945), .Y(new_n17946));
  NAND2xp33_ASAP7_75t_L     g17690(.A(new_n17787), .B(new_n17819), .Y(new_n17947));
  A2O1A1Ixp33_ASAP7_75t_L   g17691(.A1(new_n17695), .A2(new_n17691), .B(new_n17820), .C(new_n17947), .Y(new_n17948));
  NOR2xp33_ASAP7_75t_L      g17692(.A(new_n17948), .B(new_n17946), .Y(new_n17949));
  INVx1_ASAP7_75t_L         g17693(.A(new_n17949), .Y(new_n17950));
  O2A1O1Ixp33_ASAP7_75t_L   g17694(.A1(new_n17822), .A2(new_n17820), .B(new_n17947), .C(new_n17945), .Y(new_n17951));
  INVx1_ASAP7_75t_L         g17695(.A(new_n17951), .Y(new_n17952));
  AOI22xp33_ASAP7_75t_L     g17696(.A1(new_n7960), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n8537), .Y(new_n17953));
  OAI221xp5_ASAP7_75t_L     g17697(.A1(new_n8817), .A2(new_n6830), .B1(new_n7957), .B2(new_n7323), .C(new_n17953), .Y(new_n17954));
  XNOR2x2_ASAP7_75t_L       g17698(.A(\a[53] ), .B(new_n17954), .Y(new_n17955));
  NAND3xp33_ASAP7_75t_L     g17699(.A(new_n17950), .B(new_n17952), .C(new_n17955), .Y(new_n17956));
  AO21x2_ASAP7_75t_L        g17700(.A1(new_n17952), .A2(new_n17950), .B(new_n17955), .Y(new_n17957));
  AND2x2_ASAP7_75t_L        g17701(.A(new_n17956), .B(new_n17957), .Y(new_n17958));
  AOI21xp33_ASAP7_75t_L     g17702(.A1(new_n17829), .A2(new_n17825), .B(new_n17833), .Y(new_n17959));
  NAND2xp33_ASAP7_75t_L     g17703(.A(new_n17959), .B(new_n17958), .Y(new_n17960));
  INVx1_ASAP7_75t_L         g17704(.A(new_n17958), .Y(new_n17961));
  A2O1A1Ixp33_ASAP7_75t_L   g17705(.A1(new_n17829), .A2(new_n17825), .B(new_n17833), .C(new_n17961), .Y(new_n17962));
  AOI22xp33_ASAP7_75t_L     g17706(.A1(new_n7111), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n7391), .Y(new_n17963));
  OAI221xp5_ASAP7_75t_L     g17707(.A1(new_n8558), .A2(new_n7616), .B1(new_n8237), .B2(new_n7906), .C(new_n17963), .Y(new_n17964));
  XNOR2x2_ASAP7_75t_L       g17708(.A(\a[50] ), .B(new_n17964), .Y(new_n17965));
  NAND3xp33_ASAP7_75t_L     g17709(.A(new_n17962), .B(new_n17960), .C(new_n17965), .Y(new_n17966));
  AO21x2_ASAP7_75t_L        g17710(.A1(new_n17960), .A2(new_n17962), .B(new_n17965), .Y(new_n17967));
  AND2x2_ASAP7_75t_L        g17711(.A(new_n17966), .B(new_n17967), .Y(new_n17968));
  INVx1_ASAP7_75t_L         g17712(.A(new_n17968), .Y(new_n17969));
  O2A1O1Ixp33_ASAP7_75t_L   g17713(.A1(new_n17710), .A2(new_n17717), .B(new_n17839), .C(new_n17840), .Y(new_n17970));
  NAND2xp33_ASAP7_75t_L     g17714(.A(new_n17970), .B(new_n17969), .Y(new_n17971));
  A2O1A1Ixp33_ASAP7_75t_L   g17715(.A1(new_n17839), .A2(new_n17845), .B(new_n17840), .C(new_n17968), .Y(new_n17972));
  AND2x2_ASAP7_75t_L        g17716(.A(new_n17972), .B(new_n17971), .Y(new_n17973));
  NAND2xp33_ASAP7_75t_L     g17717(.A(\b[53] ), .B(new_n6648), .Y(new_n17974));
  OAI221xp5_ASAP7_75t_L     g17718(.A1(new_n6880), .A2(new_n8762), .B1(new_n6636), .B2(new_n8768), .C(new_n17974), .Y(new_n17975));
  AOI21xp33_ASAP7_75t_L     g17719(.A1(new_n6380), .A2(\b[54] ), .B(new_n17975), .Y(new_n17976));
  NAND2xp33_ASAP7_75t_L     g17720(.A(\a[47] ), .B(new_n17976), .Y(new_n17977));
  A2O1A1Ixp33_ASAP7_75t_L   g17721(.A1(\b[54] ), .A2(new_n6380), .B(new_n17975), .C(new_n6371), .Y(new_n17978));
  AND2x2_ASAP7_75t_L        g17722(.A(new_n17978), .B(new_n17977), .Y(new_n17979));
  INVx1_ASAP7_75t_L         g17723(.A(new_n17979), .Y(new_n17980));
  XNOR2x2_ASAP7_75t_L       g17724(.A(new_n17980), .B(new_n17973), .Y(new_n17981));
  OR2x4_ASAP7_75t_L         g17725(.A(new_n17902), .B(new_n17981), .Y(new_n17982));
  INVx1_ASAP7_75t_L         g17726(.A(new_n17851), .Y(new_n17983));
  A2O1A1Ixp33_ASAP7_75t_L   g17727(.A1(new_n17847), .A2(new_n17783), .B(new_n17983), .C(new_n17981), .Y(new_n17984));
  NAND2xp33_ASAP7_75t_L     g17728(.A(\b[56] ), .B(new_n5901), .Y(new_n17985));
  OAI221xp5_ASAP7_75t_L     g17729(.A1(new_n5894), .A2(new_n9920), .B1(new_n5892), .B2(new_n9925), .C(new_n17985), .Y(new_n17986));
  AOI21xp33_ASAP7_75t_L     g17730(.A1(new_n5628), .A2(\b[57] ), .B(new_n17986), .Y(new_n17987));
  NAND2xp33_ASAP7_75t_L     g17731(.A(\a[44] ), .B(new_n17987), .Y(new_n17988));
  A2O1A1Ixp33_ASAP7_75t_L   g17732(.A1(\b[57] ), .A2(new_n5628), .B(new_n17986), .C(new_n5619), .Y(new_n17989));
  AND2x2_ASAP7_75t_L        g17733(.A(new_n17989), .B(new_n17988), .Y(new_n17990));
  NAND3xp33_ASAP7_75t_L     g17734(.A(new_n17982), .B(new_n17984), .C(new_n17990), .Y(new_n17991));
  AO21x2_ASAP7_75t_L        g17735(.A1(new_n17984), .A2(new_n17982), .B(new_n17990), .Y(new_n17992));
  NAND2xp33_ASAP7_75t_L     g17736(.A(new_n17991), .B(new_n17992), .Y(new_n17993));
  OR2x4_ASAP7_75t_L         g17737(.A(new_n17857), .B(new_n17854), .Y(new_n17994));
  A2O1A1Ixp33_ASAP7_75t_L   g17738(.A1(new_n17732), .A2(new_n17779), .B(new_n17858), .C(new_n17994), .Y(new_n17995));
  NOR2xp33_ASAP7_75t_L      g17739(.A(new_n17995), .B(new_n17993), .Y(new_n17996));
  NAND2xp33_ASAP7_75t_L     g17740(.A(new_n17995), .B(new_n17993), .Y(new_n17997));
  INVx1_ASAP7_75t_L         g17741(.A(new_n17997), .Y(new_n17998));
  NOR2xp33_ASAP7_75t_L      g17742(.A(new_n17996), .B(new_n17998), .Y(new_n17999));
  NAND2xp33_ASAP7_75t_L     g17743(.A(\b[59] ), .B(new_n5167), .Y(new_n18000));
  OAI221xp5_ASAP7_75t_L     g17744(.A1(new_n5153), .A2(new_n10847), .B1(new_n5158), .B2(new_n10855), .C(new_n18000), .Y(new_n18001));
  AOI21xp33_ASAP7_75t_L     g17745(.A1(new_n4924), .A2(\b[60] ), .B(new_n18001), .Y(new_n18002));
  NAND2xp33_ASAP7_75t_L     g17746(.A(\a[41] ), .B(new_n18002), .Y(new_n18003));
  A2O1A1Ixp33_ASAP7_75t_L   g17747(.A1(\b[60] ), .A2(new_n4924), .B(new_n18001), .C(new_n4915), .Y(new_n18004));
  NAND2xp33_ASAP7_75t_L     g17748(.A(new_n18004), .B(new_n18003), .Y(new_n18005));
  NAND2xp33_ASAP7_75t_L     g17749(.A(new_n18005), .B(new_n17999), .Y(new_n18006));
  INVx1_ASAP7_75t_L         g17750(.A(new_n18006), .Y(new_n18007));
  NOR2xp33_ASAP7_75t_L      g17751(.A(new_n18005), .B(new_n17999), .Y(new_n18008));
  NOR2xp33_ASAP7_75t_L      g17752(.A(new_n18008), .B(new_n18007), .Y(new_n18009));
  NAND2xp33_ASAP7_75t_L     g17753(.A(new_n18009), .B(new_n17901), .Y(new_n18010));
  INVx1_ASAP7_75t_L         g17754(.A(new_n18010), .Y(new_n18011));
  NOR2xp33_ASAP7_75t_L      g17755(.A(new_n18009), .B(new_n17901), .Y(new_n18012));
  NOR2xp33_ASAP7_75t_L      g17756(.A(new_n18012), .B(new_n18011), .Y(new_n18013));
  NOR2xp33_ASAP7_75t_L      g17757(.A(new_n18013), .B(new_n17893), .Y(new_n18014));
  INVx1_ASAP7_75t_L         g17758(.A(new_n18013), .Y(new_n18015));
  A2O1A1O1Ixp25_ASAP7_75t_L g17759(.A1(new_n17875), .A2(new_n17876), .B(new_n17871), .C(new_n17882), .D(new_n18015), .Y(new_n18016));
  NOR2xp33_ASAP7_75t_L      g17760(.A(new_n18016), .B(new_n18014), .Y(new_n18017));
  A2O1A1Ixp33_ASAP7_75t_L   g17761(.A1(new_n17890), .A2(new_n17887), .B(new_n17884), .C(new_n18017), .Y(new_n18018));
  INVx1_ASAP7_75t_L         g17762(.A(new_n18018), .Y(new_n18019));
  A2O1A1Ixp33_ASAP7_75t_L   g17763(.A1(new_n17772), .A2(new_n17768), .B(new_n17888), .C(new_n17885), .Y(new_n18020));
  NOR2xp33_ASAP7_75t_L      g17764(.A(new_n18017), .B(new_n18020), .Y(new_n18021));
  NOR2xp33_ASAP7_75t_L      g17765(.A(new_n18021), .B(new_n18019), .Y(\f[100] ));
  INVx1_ASAP7_75t_L         g17766(.A(new_n17973), .Y(new_n18023));
  A2O1A1O1Ixp25_ASAP7_75t_L g17767(.A1(new_n17718), .A2(new_n17711), .B(new_n17843), .C(new_n17841), .D(new_n17968), .Y(new_n18024));
  AOI22xp33_ASAP7_75t_L     g17768(.A1(new_n6376), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n6648), .Y(new_n18025));
  OAI221xp5_ASAP7_75t_L     g17769(.A1(new_n6646), .A2(new_n8762), .B1(new_n6636), .B2(new_n9331), .C(new_n18025), .Y(new_n18026));
  XNOR2x2_ASAP7_75t_L       g17770(.A(\a[47] ), .B(new_n18026), .Y(new_n18027));
  INVx1_ASAP7_75t_L         g17771(.A(new_n18027), .Y(new_n18028));
  AOI22xp33_ASAP7_75t_L     g17772(.A1(new_n7111), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n7391), .Y(new_n18029));
  OAI221xp5_ASAP7_75t_L     g17773(.A1(new_n8558), .A2(new_n7900), .B1(new_n8237), .B2(new_n8174), .C(new_n18029), .Y(new_n18030));
  XNOR2x2_ASAP7_75t_L       g17774(.A(\a[50] ), .B(new_n18030), .Y(new_n18031));
  INVx1_ASAP7_75t_L         g17775(.A(new_n18031), .Y(new_n18032));
  AOI22xp33_ASAP7_75t_L     g17776(.A1(new_n9700), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n10027), .Y(new_n18033));
  OAI221xp5_ASAP7_75t_L     g17777(.A1(new_n10024), .A2(new_n5805), .B1(new_n9696), .B2(new_n5835), .C(new_n18033), .Y(new_n18034));
  XNOR2x2_ASAP7_75t_L       g17778(.A(\a[59] ), .B(new_n18034), .Y(new_n18035));
  A2O1A1Ixp33_ASAP7_75t_L   g17779(.A1(new_n17792), .A2(new_n17911), .B(new_n17912), .C(new_n17910), .Y(new_n18036));
  NAND2xp33_ASAP7_75t_L     g17780(.A(\b[37] ), .B(new_n11534), .Y(new_n18037));
  OAI211xp5_ASAP7_75t_L     g17781(.A1(new_n11253), .A2(new_n4632), .B(new_n17910), .C(new_n18037), .Y(new_n18038));
  A2O1A1Ixp33_ASAP7_75t_L   g17782(.A1(new_n14788), .A2(new_n14789), .B(new_n4632), .C(new_n18037), .Y(new_n18039));
  A2O1A1Ixp33_ASAP7_75t_L   g17783(.A1(new_n11533), .A2(\b[37] ), .B(new_n17909), .C(new_n18039), .Y(new_n18040));
  AND2x2_ASAP7_75t_L        g17784(.A(new_n18040), .B(new_n18038), .Y(new_n18041));
  INVx1_ASAP7_75t_L         g17785(.A(new_n18041), .Y(new_n18042));
  A2O1A1O1Ixp25_ASAP7_75t_L g17786(.A1(new_n17907), .A2(new_n17906), .B(new_n17917), .C(new_n18036), .D(new_n18042), .Y(new_n18043));
  A2O1A1Ixp33_ASAP7_75t_L   g17787(.A1(new_n17906), .A2(new_n17907), .B(new_n17917), .C(new_n18036), .Y(new_n18044));
  NOR2xp33_ASAP7_75t_L      g17788(.A(new_n18041), .B(new_n18044), .Y(new_n18045));
  NOR2xp33_ASAP7_75t_L      g17789(.A(new_n18043), .B(new_n18045), .Y(new_n18046));
  INVx1_ASAP7_75t_L         g17790(.A(new_n18046), .Y(new_n18047));
  AOI22xp33_ASAP7_75t_L     g17791(.A1(\b[39] ), .A2(new_n10939), .B1(\b[41] ), .B2(new_n10938), .Y(new_n18048));
  OAI221xp5_ASAP7_75t_L     g17792(.A1(new_n10937), .A2(new_n4869), .B1(new_n10629), .B2(new_n5327), .C(new_n18048), .Y(new_n18049));
  XNOR2x2_ASAP7_75t_L       g17793(.A(\a[62] ), .B(new_n18049), .Y(new_n18050));
  INVx1_ASAP7_75t_L         g17794(.A(new_n18050), .Y(new_n18051));
  NAND2xp33_ASAP7_75t_L     g17795(.A(new_n18051), .B(new_n18047), .Y(new_n18052));
  NAND2xp33_ASAP7_75t_L     g17796(.A(new_n18050), .B(new_n18046), .Y(new_n18053));
  NAND3xp33_ASAP7_75t_L     g17797(.A(new_n18052), .B(new_n18035), .C(new_n18053), .Y(new_n18054));
  INVx1_ASAP7_75t_L         g17798(.A(new_n18054), .Y(new_n18055));
  AOI21xp33_ASAP7_75t_L     g17799(.A1(new_n18052), .A2(new_n18053), .B(new_n18035), .Y(new_n18056));
  NOR2xp33_ASAP7_75t_L      g17800(.A(new_n18056), .B(new_n18055), .Y(new_n18057));
  INVx1_ASAP7_75t_L         g17801(.A(new_n18057), .Y(new_n18058));
  O2A1O1Ixp33_ASAP7_75t_L   g17802(.A1(new_n17919), .A2(new_n17921), .B(new_n17929), .C(new_n18058), .Y(new_n18059));
  INVx1_ASAP7_75t_L         g17803(.A(new_n18059), .Y(new_n18060));
  NAND3xp33_ASAP7_75t_L     g17804(.A(new_n17929), .B(new_n18058), .C(new_n17923), .Y(new_n18061));
  AOI22xp33_ASAP7_75t_L     g17805(.A1(new_n8831), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n9115), .Y(new_n18062));
  OAI221xp5_ASAP7_75t_L     g17806(.A1(new_n10343), .A2(new_n6568), .B1(new_n10016), .B2(new_n6820), .C(new_n18062), .Y(new_n18063));
  XNOR2x2_ASAP7_75t_L       g17807(.A(\a[56] ), .B(new_n18063), .Y(new_n18064));
  NAND3xp33_ASAP7_75t_L     g17808(.A(new_n18060), .B(new_n18061), .C(new_n18064), .Y(new_n18065));
  AO21x2_ASAP7_75t_L        g17809(.A1(new_n18061), .A2(new_n18060), .B(new_n18064), .Y(new_n18066));
  AND2x2_ASAP7_75t_L        g17810(.A(new_n18065), .B(new_n18066), .Y(new_n18067));
  A2O1A1Ixp33_ASAP7_75t_L   g17811(.A1(new_n17939), .A2(new_n17942), .B(new_n17936), .C(new_n18067), .Y(new_n18068));
  NAND2xp33_ASAP7_75t_L     g17812(.A(new_n17937), .B(new_n17943), .Y(new_n18069));
  NOR2xp33_ASAP7_75t_L      g17813(.A(new_n18067), .B(new_n18069), .Y(new_n18070));
  INVx1_ASAP7_75t_L         g17814(.A(new_n18070), .Y(new_n18071));
  NAND2xp33_ASAP7_75t_L     g17815(.A(new_n18068), .B(new_n18071), .Y(new_n18072));
  AOI22xp33_ASAP7_75t_L     g17816(.A1(new_n7960), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n8537), .Y(new_n18073));
  OAI221xp5_ASAP7_75t_L     g17817(.A1(new_n8817), .A2(new_n7317), .B1(new_n7957), .B2(new_n7602), .C(new_n18073), .Y(new_n18074));
  XNOR2x2_ASAP7_75t_L       g17818(.A(\a[53] ), .B(new_n18074), .Y(new_n18075));
  NAND2xp33_ASAP7_75t_L     g17819(.A(new_n18075), .B(new_n18072), .Y(new_n18076));
  NOR2xp33_ASAP7_75t_L      g17820(.A(new_n18075), .B(new_n18072), .Y(new_n18077));
  INVx1_ASAP7_75t_L         g17821(.A(new_n18077), .Y(new_n18078));
  AND2x2_ASAP7_75t_L        g17822(.A(new_n18076), .B(new_n18078), .Y(new_n18079));
  INVx1_ASAP7_75t_L         g17823(.A(new_n18079), .Y(new_n18080));
  NAND2xp33_ASAP7_75t_L     g17824(.A(new_n17950), .B(new_n17956), .Y(new_n18081));
  NOR2xp33_ASAP7_75t_L      g17825(.A(new_n18081), .B(new_n18080), .Y(new_n18082));
  O2A1O1Ixp33_ASAP7_75t_L   g17826(.A1(new_n17946), .A2(new_n17948), .B(new_n17956), .C(new_n18079), .Y(new_n18083));
  NOR2xp33_ASAP7_75t_L      g17827(.A(new_n18083), .B(new_n18082), .Y(new_n18084));
  NAND2xp33_ASAP7_75t_L     g17828(.A(new_n18032), .B(new_n18084), .Y(new_n18085));
  INVx1_ASAP7_75t_L         g17829(.A(new_n18085), .Y(new_n18086));
  NOR2xp33_ASAP7_75t_L      g17830(.A(new_n18032), .B(new_n18084), .Y(new_n18087));
  NOR2xp33_ASAP7_75t_L      g17831(.A(new_n18087), .B(new_n18086), .Y(new_n18088));
  INVx1_ASAP7_75t_L         g17832(.A(new_n18088), .Y(new_n18089));
  NAND2xp33_ASAP7_75t_L     g17833(.A(new_n17960), .B(new_n17966), .Y(new_n18090));
  NOR2xp33_ASAP7_75t_L      g17834(.A(new_n18090), .B(new_n18089), .Y(new_n18091));
  INVx1_ASAP7_75t_L         g17835(.A(new_n18091), .Y(new_n18092));
  INVx1_ASAP7_75t_L         g17836(.A(new_n17960), .Y(new_n18093));
  A2O1A1Ixp33_ASAP7_75t_L   g17837(.A1(new_n17962), .A2(new_n17965), .B(new_n18093), .C(new_n18089), .Y(new_n18094));
  NAND3xp33_ASAP7_75t_L     g17838(.A(new_n18092), .B(new_n18028), .C(new_n18094), .Y(new_n18095));
  AO21x2_ASAP7_75t_L        g17839(.A1(new_n18094), .A2(new_n18092), .B(new_n18028), .Y(new_n18096));
  AND2x2_ASAP7_75t_L        g17840(.A(new_n18095), .B(new_n18096), .Y(new_n18097));
  A2O1A1Ixp33_ASAP7_75t_L   g17841(.A1(new_n17980), .A2(new_n18023), .B(new_n18024), .C(new_n18097), .Y(new_n18098));
  INVx1_ASAP7_75t_L         g17842(.A(new_n18024), .Y(new_n18099));
  A2O1A1Ixp33_ASAP7_75t_L   g17843(.A1(new_n17971), .A2(new_n17972), .B(new_n17979), .C(new_n18099), .Y(new_n18100));
  NOR2xp33_ASAP7_75t_L      g17844(.A(new_n18100), .B(new_n18097), .Y(new_n18101));
  INVx1_ASAP7_75t_L         g17845(.A(new_n18101), .Y(new_n18102));
  AOI22xp33_ASAP7_75t_L     g17846(.A1(new_n5624), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n5901), .Y(new_n18103));
  OAI221xp5_ASAP7_75t_L     g17847(.A1(new_n5900), .A2(new_n9920), .B1(new_n5892), .B2(new_n11152), .C(new_n18103), .Y(new_n18104));
  XNOR2x2_ASAP7_75t_L       g17848(.A(\a[44] ), .B(new_n18104), .Y(new_n18105));
  NAND3xp33_ASAP7_75t_L     g17849(.A(new_n18102), .B(new_n18098), .C(new_n18105), .Y(new_n18106));
  INVx1_ASAP7_75t_L         g17850(.A(new_n18106), .Y(new_n18107));
  AOI21xp33_ASAP7_75t_L     g17851(.A1(new_n18102), .A2(new_n18098), .B(new_n18105), .Y(new_n18108));
  NOR2xp33_ASAP7_75t_L      g17852(.A(new_n18108), .B(new_n18107), .Y(new_n18109));
  INVx1_ASAP7_75t_L         g17853(.A(new_n18109), .Y(new_n18110));
  O2A1O1Ixp33_ASAP7_75t_L   g17854(.A1(new_n17902), .A2(new_n17981), .B(new_n17991), .C(new_n18110), .Y(new_n18111));
  INVx1_ASAP7_75t_L         g17855(.A(new_n18111), .Y(new_n18112));
  NAND3xp33_ASAP7_75t_L     g17856(.A(new_n18110), .B(new_n17991), .C(new_n17982), .Y(new_n18113));
  AOI22xp33_ASAP7_75t_L     g17857(.A1(new_n4920), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n5167), .Y(new_n18114));
  OAI221xp5_ASAP7_75t_L     g17858(.A1(new_n5154), .A2(new_n10847), .B1(new_n5158), .B2(new_n12047), .C(new_n18114), .Y(new_n18115));
  XNOR2x2_ASAP7_75t_L       g17859(.A(\a[41] ), .B(new_n18115), .Y(new_n18116));
  NAND3xp33_ASAP7_75t_L     g17860(.A(new_n18112), .B(new_n18113), .C(new_n18116), .Y(new_n18117));
  INVx1_ASAP7_75t_L         g17861(.A(new_n18117), .Y(new_n18118));
  AOI21xp33_ASAP7_75t_L     g17862(.A1(new_n18112), .A2(new_n18113), .B(new_n18116), .Y(new_n18119));
  NOR2xp33_ASAP7_75t_L      g17863(.A(new_n18119), .B(new_n18118), .Y(new_n18120));
  A2O1A1O1Ixp25_ASAP7_75t_L g17864(.A1(new_n4274), .A2(new_n12061), .B(new_n4512), .C(\b[63] ), .D(new_n4268), .Y(new_n18121));
  A2O1A1O1Ixp25_ASAP7_75t_L g17865(.A1(\b[61] ), .A2(new_n11471), .B(\b[62] ), .C(new_n4274), .D(new_n4512), .Y(new_n18122));
  NOR3xp33_ASAP7_75t_L      g17866(.A(new_n18122), .B(new_n11468), .C(\a[38] ), .Y(new_n18123));
  NOR2xp33_ASAP7_75t_L      g17867(.A(new_n18121), .B(new_n18123), .Y(new_n18124));
  A2O1A1O1Ixp25_ASAP7_75t_L g17868(.A1(new_n18003), .A2(new_n18004), .B(new_n17996), .C(new_n17997), .D(new_n18124), .Y(new_n18125));
  INVx1_ASAP7_75t_L         g17869(.A(new_n18125), .Y(new_n18126));
  NAND3xp33_ASAP7_75t_L     g17870(.A(new_n18006), .B(new_n17997), .C(new_n18124), .Y(new_n18127));
  NAND2xp33_ASAP7_75t_L     g17871(.A(new_n18126), .B(new_n18127), .Y(new_n18128));
  XNOR2x2_ASAP7_75t_L       g17872(.A(new_n18128), .B(new_n18120), .Y(new_n18129));
  O2A1O1Ixp33_ASAP7_75t_L   g17873(.A1(new_n17899), .A2(new_n17896), .B(new_n18010), .C(new_n18129), .Y(new_n18130));
  INVx1_ASAP7_75t_L         g17874(.A(new_n18130), .Y(new_n18131));
  A2O1A1O1Ixp25_ASAP7_75t_L g17875(.A1(new_n17865), .A2(new_n17861), .B(new_n17869), .C(new_n17897), .D(new_n18011), .Y(new_n18132));
  NAND2xp33_ASAP7_75t_L     g17876(.A(new_n18129), .B(new_n18132), .Y(new_n18133));
  AND2x2_ASAP7_75t_L        g17877(.A(new_n18133), .B(new_n18131), .Y(new_n18134));
  A2O1A1Ixp33_ASAP7_75t_L   g17878(.A1(new_n18020), .A2(new_n18017), .B(new_n18016), .C(new_n18134), .Y(new_n18135));
  A2O1A1O1Ixp25_ASAP7_75t_L g17879(.A1(new_n17887), .A2(new_n17890), .B(new_n17884), .C(new_n18017), .D(new_n18016), .Y(new_n18136));
  INVx1_ASAP7_75t_L         g17880(.A(new_n18134), .Y(new_n18137));
  NAND2xp33_ASAP7_75t_L     g17881(.A(new_n18137), .B(new_n18136), .Y(new_n18138));
  AND2x2_ASAP7_75t_L        g17882(.A(new_n18135), .B(new_n18138), .Y(\f[101] ));
  INVx1_ASAP7_75t_L         g17883(.A(new_n18016), .Y(new_n18140));
  INVx1_ASAP7_75t_L         g17884(.A(new_n18127), .Y(new_n18141));
  AOI22xp33_ASAP7_75t_L     g17885(.A1(new_n7111), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n7391), .Y(new_n18142));
  OAI221xp5_ASAP7_75t_L     g17886(.A1(new_n8558), .A2(new_n8165), .B1(new_n8237), .B2(new_n8465), .C(new_n18142), .Y(new_n18143));
  XNOR2x2_ASAP7_75t_L       g17887(.A(\a[50] ), .B(new_n18143), .Y(new_n18144));
  INVx1_ASAP7_75t_L         g17888(.A(new_n18144), .Y(new_n18145));
  AOI22xp33_ASAP7_75t_L     g17889(.A1(new_n8831), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n9115), .Y(new_n18146));
  OAI221xp5_ASAP7_75t_L     g17890(.A1(new_n10343), .A2(new_n6812), .B1(new_n10016), .B2(new_n6837), .C(new_n18146), .Y(new_n18147));
  XNOR2x2_ASAP7_75t_L       g17891(.A(\a[56] ), .B(new_n18147), .Y(new_n18148));
  INVx1_ASAP7_75t_L         g17892(.A(new_n18148), .Y(new_n18149));
  O2A1O1Ixp33_ASAP7_75t_L   g17893(.A1(new_n11253), .A2(new_n4632), .B(new_n18037), .C(new_n17915), .Y(new_n18150));
  NOR2xp33_ASAP7_75t_L      g17894(.A(new_n4632), .B(new_n11535), .Y(new_n18151));
  A2O1A1Ixp33_ASAP7_75t_L   g17895(.A1(new_n11533), .A2(\b[37] ), .B(new_n17909), .C(\a[38] ), .Y(new_n18152));
  NOR2xp33_ASAP7_75t_L      g17896(.A(\a[38] ), .B(new_n17915), .Y(new_n18153));
  INVx1_ASAP7_75t_L         g17897(.A(new_n18153), .Y(new_n18154));
  NAND2xp33_ASAP7_75t_L     g17898(.A(new_n18152), .B(new_n18154), .Y(new_n18155));
  A2O1A1Ixp33_ASAP7_75t_L   g17899(.A1(new_n11533), .A2(\b[39] ), .B(new_n18151), .C(new_n18155), .Y(new_n18156));
  INVx1_ASAP7_75t_L         g17900(.A(new_n18156), .Y(new_n18157));
  O2A1O1Ixp33_ASAP7_75t_L   g17901(.A1(new_n11247), .A2(new_n11249), .B(\b[39] ), .C(new_n18151), .Y(new_n18158));
  AND3x1_ASAP7_75t_L        g17902(.A(new_n18154), .B(new_n18152), .C(new_n18158), .Y(new_n18159));
  NOR2xp33_ASAP7_75t_L      g17903(.A(new_n18159), .B(new_n18157), .Y(new_n18160));
  A2O1A1Ixp33_ASAP7_75t_L   g17904(.A1(new_n18044), .A2(new_n18042), .B(new_n18150), .C(new_n18160), .Y(new_n18161));
  A2O1A1O1Ixp25_ASAP7_75t_L g17905(.A1(new_n17907), .A2(new_n17906), .B(new_n17917), .C(new_n18036), .D(new_n18041), .Y(new_n18162));
  OR3x1_ASAP7_75t_L         g17906(.A(new_n18162), .B(new_n18150), .C(new_n18160), .Y(new_n18163));
  NAND2xp33_ASAP7_75t_L     g17907(.A(\b[40] ), .B(new_n10939), .Y(new_n18164));
  OAI221xp5_ASAP7_75t_L     g17908(.A1(new_n10630), .A2(new_n5338), .B1(new_n10629), .B2(new_n5346), .C(new_n18164), .Y(new_n18165));
  AOI21xp33_ASAP7_75t_L     g17909(.A1(new_n10632), .A2(\b[41] ), .B(new_n18165), .Y(new_n18166));
  NAND2xp33_ASAP7_75t_L     g17910(.A(\a[62] ), .B(new_n18166), .Y(new_n18167));
  A2O1A1Ixp33_ASAP7_75t_L   g17911(.A1(\b[41] ), .A2(new_n10632), .B(new_n18165), .C(new_n10622), .Y(new_n18168));
  NAND4xp25_ASAP7_75t_L     g17912(.A(new_n18163), .B(new_n18167), .C(new_n18168), .D(new_n18161), .Y(new_n18169));
  NAND2xp33_ASAP7_75t_L     g17913(.A(new_n18161), .B(new_n18163), .Y(new_n18170));
  NAND2xp33_ASAP7_75t_L     g17914(.A(new_n18168), .B(new_n18167), .Y(new_n18171));
  NAND2xp33_ASAP7_75t_L     g17915(.A(new_n18171), .B(new_n18170), .Y(new_n18172));
  NAND2xp33_ASAP7_75t_L     g17916(.A(new_n18169), .B(new_n18172), .Y(new_n18173));
  AOI22xp33_ASAP7_75t_L     g17917(.A1(new_n9700), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n10027), .Y(new_n18174));
  OAI221xp5_ASAP7_75t_L     g17918(.A1(new_n10024), .A2(new_n5829), .B1(new_n9696), .B2(new_n6329), .C(new_n18174), .Y(new_n18175));
  XNOR2x2_ASAP7_75t_L       g17919(.A(\a[59] ), .B(new_n18175), .Y(new_n18176));
  INVx1_ASAP7_75t_L         g17920(.A(new_n18176), .Y(new_n18177));
  NAND2xp33_ASAP7_75t_L     g17921(.A(new_n18177), .B(new_n18173), .Y(new_n18178));
  NAND3xp33_ASAP7_75t_L     g17922(.A(new_n18172), .B(new_n18169), .C(new_n18176), .Y(new_n18179));
  AND2x2_ASAP7_75t_L        g17923(.A(new_n18179), .B(new_n18178), .Y(new_n18180));
  INVx1_ASAP7_75t_L         g17924(.A(new_n18180), .Y(new_n18181));
  NAND2xp33_ASAP7_75t_L     g17925(.A(new_n18053), .B(new_n18054), .Y(new_n18182));
  NOR2xp33_ASAP7_75t_L      g17926(.A(new_n18182), .B(new_n18181), .Y(new_n18183));
  O2A1O1Ixp33_ASAP7_75t_L   g17927(.A1(new_n18047), .A2(new_n18051), .B(new_n18054), .C(new_n18180), .Y(new_n18184));
  NOR2xp33_ASAP7_75t_L      g17928(.A(new_n18184), .B(new_n18183), .Y(new_n18185));
  XNOR2x2_ASAP7_75t_L       g17929(.A(new_n18149), .B(new_n18185), .Y(new_n18186));
  A2O1A1Ixp33_ASAP7_75t_L   g17930(.A1(new_n18061), .A2(new_n18064), .B(new_n18059), .C(new_n18186), .Y(new_n18187));
  A2O1A1Ixp33_ASAP7_75t_L   g17931(.A1(new_n17929), .A2(new_n17923), .B(new_n18058), .C(new_n18065), .Y(new_n18188));
  NOR2xp33_ASAP7_75t_L      g17932(.A(new_n18186), .B(new_n18188), .Y(new_n18189));
  INVx1_ASAP7_75t_L         g17933(.A(new_n18189), .Y(new_n18190));
  NAND2xp33_ASAP7_75t_L     g17934(.A(new_n18187), .B(new_n18190), .Y(new_n18191));
  AOI22xp33_ASAP7_75t_L     g17935(.A1(new_n7960), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n8537), .Y(new_n18192));
  OAI221xp5_ASAP7_75t_L     g17936(.A1(new_n8817), .A2(new_n7593), .B1(new_n7957), .B2(new_n7623), .C(new_n18192), .Y(new_n18193));
  XNOR2x2_ASAP7_75t_L       g17937(.A(\a[53] ), .B(new_n18193), .Y(new_n18194));
  NAND2xp33_ASAP7_75t_L     g17938(.A(new_n18194), .B(new_n18191), .Y(new_n18195));
  NOR2xp33_ASAP7_75t_L      g17939(.A(new_n18194), .B(new_n18191), .Y(new_n18196));
  INVx1_ASAP7_75t_L         g17940(.A(new_n18196), .Y(new_n18197));
  AND2x2_ASAP7_75t_L        g17941(.A(new_n18195), .B(new_n18197), .Y(new_n18198));
  INVx1_ASAP7_75t_L         g17942(.A(new_n18198), .Y(new_n18199));
  O2A1O1Ixp33_ASAP7_75t_L   g17943(.A1(new_n18067), .A2(new_n18069), .B(new_n18078), .C(new_n18199), .Y(new_n18200));
  A2O1A1Ixp33_ASAP7_75t_L   g17944(.A1(new_n18066), .A2(new_n18065), .B(new_n18069), .C(new_n18078), .Y(new_n18201));
  NOR2xp33_ASAP7_75t_L      g17945(.A(new_n18198), .B(new_n18201), .Y(new_n18202));
  NOR2xp33_ASAP7_75t_L      g17946(.A(new_n18200), .B(new_n18202), .Y(new_n18203));
  NAND2xp33_ASAP7_75t_L     g17947(.A(new_n18145), .B(new_n18203), .Y(new_n18204));
  OAI21xp33_ASAP7_75t_L     g17948(.A1(new_n18200), .A2(new_n18202), .B(new_n18144), .Y(new_n18205));
  AND2x2_ASAP7_75t_L        g17949(.A(new_n18205), .B(new_n18204), .Y(new_n18206));
  A2O1A1Ixp33_ASAP7_75t_L   g17950(.A1(new_n18084), .A2(new_n18032), .B(new_n18082), .C(new_n18206), .Y(new_n18207));
  OR3x1_ASAP7_75t_L         g17951(.A(new_n18086), .B(new_n18082), .C(new_n18206), .Y(new_n18208));
  NAND2xp33_ASAP7_75t_L     g17952(.A(new_n18207), .B(new_n18208), .Y(new_n18209));
  AOI22xp33_ASAP7_75t_L     g17953(.A1(new_n6376), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n6648), .Y(new_n18210));
  OAI221xp5_ASAP7_75t_L     g17954(.A1(new_n6646), .A2(new_n9323), .B1(new_n6636), .B2(new_n9627), .C(new_n18210), .Y(new_n18211));
  XNOR2x2_ASAP7_75t_L       g17955(.A(\a[47] ), .B(new_n18211), .Y(new_n18212));
  XNOR2x2_ASAP7_75t_L       g17956(.A(new_n18212), .B(new_n18209), .Y(new_n18213));
  INVx1_ASAP7_75t_L         g17957(.A(new_n18213), .Y(new_n18214));
  NAND2xp33_ASAP7_75t_L     g17958(.A(new_n18092), .B(new_n18095), .Y(new_n18215));
  NOR2xp33_ASAP7_75t_L      g17959(.A(new_n18214), .B(new_n18215), .Y(new_n18216));
  O2A1O1Ixp33_ASAP7_75t_L   g17960(.A1(new_n18089), .A2(new_n18090), .B(new_n18095), .C(new_n18213), .Y(new_n18217));
  NOR2xp33_ASAP7_75t_L      g17961(.A(new_n18217), .B(new_n18216), .Y(new_n18218));
  AOI22xp33_ASAP7_75t_L     g17962(.A1(new_n5624), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n5901), .Y(new_n18219));
  OAI221xp5_ASAP7_75t_L     g17963(.A1(new_n5900), .A2(new_n9947), .B1(new_n5892), .B2(new_n11446), .C(new_n18219), .Y(new_n18220));
  XNOR2x2_ASAP7_75t_L       g17964(.A(\a[44] ), .B(new_n18220), .Y(new_n18221));
  INVx1_ASAP7_75t_L         g17965(.A(new_n18221), .Y(new_n18222));
  XNOR2x2_ASAP7_75t_L       g17966(.A(new_n18222), .B(new_n18218), .Y(new_n18223));
  A2O1A1Ixp33_ASAP7_75t_L   g17967(.A1(new_n18105), .A2(new_n18098), .B(new_n18101), .C(new_n18223), .Y(new_n18224));
  A2O1A1Ixp33_ASAP7_75t_L   g17968(.A1(new_n18095), .A2(new_n18096), .B(new_n18100), .C(new_n18106), .Y(new_n18225));
  NOR2xp33_ASAP7_75t_L      g17969(.A(new_n18223), .B(new_n18225), .Y(new_n18226));
  INVx1_ASAP7_75t_L         g17970(.A(new_n18226), .Y(new_n18227));
  NAND2xp33_ASAP7_75t_L     g17971(.A(new_n18224), .B(new_n18227), .Y(new_n18228));
  AOI22xp33_ASAP7_75t_L     g17972(.A1(new_n4920), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n5167), .Y(new_n18229));
  A2O1A1Ixp33_ASAP7_75t_L   g17973(.A1(new_n11470), .A2(new_n11473), .B(new_n5158), .C(new_n18229), .Y(new_n18230));
  AOI21xp33_ASAP7_75t_L     g17974(.A1(new_n4924), .A2(\b[62] ), .B(new_n18230), .Y(new_n18231));
  NAND2xp33_ASAP7_75t_L     g17975(.A(\a[41] ), .B(new_n18231), .Y(new_n18232));
  A2O1A1Ixp33_ASAP7_75t_L   g17976(.A1(\b[62] ), .A2(new_n4924), .B(new_n18230), .C(new_n4915), .Y(new_n18233));
  NAND2xp33_ASAP7_75t_L     g17977(.A(new_n18233), .B(new_n18232), .Y(new_n18234));
  XOR2x2_ASAP7_75t_L        g17978(.A(new_n18234), .B(new_n18228), .Y(new_n18235));
  A2O1A1Ixp33_ASAP7_75t_L   g17979(.A1(new_n18113), .A2(new_n18116), .B(new_n18111), .C(new_n18235), .Y(new_n18236));
  A2O1A1Ixp33_ASAP7_75t_L   g17980(.A1(new_n17991), .A2(new_n17982), .B(new_n18110), .C(new_n18117), .Y(new_n18237));
  NOR2xp33_ASAP7_75t_L      g17981(.A(new_n18235), .B(new_n18237), .Y(new_n18238));
  INVx1_ASAP7_75t_L         g17982(.A(new_n18238), .Y(new_n18239));
  NAND2xp33_ASAP7_75t_L     g17983(.A(new_n18236), .B(new_n18239), .Y(new_n18240));
  O2A1O1Ixp33_ASAP7_75t_L   g17984(.A1(new_n18120), .A2(new_n18141), .B(new_n18126), .C(new_n18240), .Y(new_n18241));
  INVx1_ASAP7_75t_L         g17985(.A(new_n18241), .Y(new_n18242));
  OAI211xp5_ASAP7_75t_L     g17986(.A1(new_n18120), .A2(new_n18141), .B(new_n18240), .C(new_n18126), .Y(new_n18243));
  AND2x2_ASAP7_75t_L        g17987(.A(new_n18243), .B(new_n18242), .Y(new_n18244));
  INVx1_ASAP7_75t_L         g17988(.A(new_n18244), .Y(new_n18245));
  A2O1A1O1Ixp25_ASAP7_75t_L g17989(.A1(new_n18140), .A2(new_n18018), .B(new_n18137), .C(new_n18131), .D(new_n18245), .Y(new_n18246));
  A2O1A1Ixp33_ASAP7_75t_L   g17990(.A1(new_n18018), .A2(new_n18140), .B(new_n18137), .C(new_n18131), .Y(new_n18247));
  NOR2xp33_ASAP7_75t_L      g17991(.A(new_n18244), .B(new_n18247), .Y(new_n18248));
  NOR2xp33_ASAP7_75t_L      g17992(.A(new_n18246), .B(new_n18248), .Y(\f[102] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17993(.A1(new_n18232), .A2(new_n18233), .B(new_n18228), .C(new_n18239), .Y(new_n18250));
  NOR2xp33_ASAP7_75t_L      g17994(.A(new_n11172), .B(new_n5160), .Y(new_n18251));
  AOI221xp5_ASAP7_75t_L     g17995(.A1(\b[63] ), .A2(new_n4924), .B1(new_n4917), .B2(new_n12322), .C(new_n18251), .Y(new_n18252));
  XNOR2x2_ASAP7_75t_L       g17996(.A(new_n4915), .B(new_n18252), .Y(new_n18253));
  INVx1_ASAP7_75t_L         g17997(.A(new_n18253), .Y(new_n18254));
  A2O1A1Ixp33_ASAP7_75t_L   g17998(.A1(new_n18222), .A2(new_n18218), .B(new_n18226), .C(new_n18254), .Y(new_n18255));
  AOI21xp33_ASAP7_75t_L     g17999(.A1(new_n18222), .A2(new_n18218), .B(new_n18226), .Y(new_n18256));
  NAND2xp33_ASAP7_75t_L     g18000(.A(new_n18253), .B(new_n18256), .Y(new_n18257));
  AND2x2_ASAP7_75t_L        g18001(.A(new_n18255), .B(new_n18257), .Y(new_n18258));
  INVx1_ASAP7_75t_L         g18002(.A(new_n18183), .Y(new_n18259));
  NOR2xp33_ASAP7_75t_L      g18003(.A(new_n4848), .B(new_n11535), .Y(new_n18260));
  O2A1O1Ixp33_ASAP7_75t_L   g18004(.A1(new_n11247), .A2(new_n11249), .B(\b[40] ), .C(new_n18260), .Y(new_n18261));
  INVx1_ASAP7_75t_L         g18005(.A(new_n18261), .Y(new_n18262));
  A2O1A1Ixp33_ASAP7_75t_L   g18006(.A1(new_n11533), .A2(\b[37] ), .B(new_n17909), .C(new_n4268), .Y(new_n18263));
  A2O1A1O1Ixp25_ASAP7_75t_L g18007(.A1(new_n18152), .A2(new_n18154), .B(new_n18158), .C(new_n18263), .D(new_n18262), .Y(new_n18264));
  INVx1_ASAP7_75t_L         g18008(.A(new_n18264), .Y(new_n18265));
  A2O1A1O1Ixp25_ASAP7_75t_L g18009(.A1(new_n11533), .A2(\b[37] ), .B(new_n17909), .C(new_n4268), .D(new_n18157), .Y(new_n18266));
  A2O1A1Ixp33_ASAP7_75t_L   g18010(.A1(new_n11533), .A2(\b[40] ), .B(new_n18260), .C(new_n18266), .Y(new_n18267));
  NAND2xp33_ASAP7_75t_L     g18011(.A(new_n18265), .B(new_n18267), .Y(new_n18268));
  NAND2xp33_ASAP7_75t_L     g18012(.A(\b[42] ), .B(new_n10632), .Y(new_n18269));
  OAI221xp5_ASAP7_75t_L     g18013(.A1(new_n10630), .A2(new_n5805), .B1(new_n5321), .B2(new_n11257), .C(new_n18269), .Y(new_n18270));
  AOI21xp33_ASAP7_75t_L     g18014(.A1(new_n5812), .A2(new_n11256), .B(new_n18270), .Y(new_n18271));
  NAND2xp33_ASAP7_75t_L     g18015(.A(\a[62] ), .B(new_n18271), .Y(new_n18272));
  A2O1A1Ixp33_ASAP7_75t_L   g18016(.A1(new_n5812), .A2(new_n11256), .B(new_n18270), .C(new_n10622), .Y(new_n18273));
  NAND2xp33_ASAP7_75t_L     g18017(.A(new_n18273), .B(new_n18272), .Y(new_n18274));
  XNOR2x2_ASAP7_75t_L       g18018(.A(new_n18268), .B(new_n18274), .Y(new_n18275));
  NAND3xp33_ASAP7_75t_L     g18019(.A(new_n18169), .B(new_n18163), .C(new_n18275), .Y(new_n18276));
  O2A1O1Ixp33_ASAP7_75t_L   g18020(.A1(new_n18171), .A2(new_n18170), .B(new_n18163), .C(new_n18275), .Y(new_n18277));
  INVx1_ASAP7_75t_L         g18021(.A(new_n18277), .Y(new_n18278));
  AOI22xp33_ASAP7_75t_L     g18022(.A1(new_n9700), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n10027), .Y(new_n18279));
  OAI221xp5_ASAP7_75t_L     g18023(.A1(new_n10024), .A2(new_n6321), .B1(new_n9696), .B2(new_n6573), .C(new_n18279), .Y(new_n18280));
  XNOR2x2_ASAP7_75t_L       g18024(.A(\a[59] ), .B(new_n18280), .Y(new_n18281));
  NAND3xp33_ASAP7_75t_L     g18025(.A(new_n18278), .B(new_n18276), .C(new_n18281), .Y(new_n18282));
  AO21x2_ASAP7_75t_L        g18026(.A1(new_n18276), .A2(new_n18278), .B(new_n18281), .Y(new_n18283));
  AND2x2_ASAP7_75t_L        g18027(.A(new_n18282), .B(new_n18283), .Y(new_n18284));
  NAND3xp33_ASAP7_75t_L     g18028(.A(new_n18259), .B(new_n18178), .C(new_n18284), .Y(new_n18285));
  INVx1_ASAP7_75t_L         g18029(.A(new_n18284), .Y(new_n18286));
  A2O1A1Ixp33_ASAP7_75t_L   g18030(.A1(new_n18177), .A2(new_n18173), .B(new_n18183), .C(new_n18286), .Y(new_n18287));
  NAND2xp33_ASAP7_75t_L     g18031(.A(\b[47] ), .B(new_n9115), .Y(new_n18288));
  OAI221xp5_ASAP7_75t_L     g18032(.A1(new_n9113), .A2(new_n7317), .B1(new_n10016), .B2(new_n7323), .C(new_n18288), .Y(new_n18289));
  AOI21xp33_ASAP7_75t_L     g18033(.A1(new_n8835), .A2(\b[48] ), .B(new_n18289), .Y(new_n18290));
  NAND2xp33_ASAP7_75t_L     g18034(.A(\a[56] ), .B(new_n18290), .Y(new_n18291));
  A2O1A1Ixp33_ASAP7_75t_L   g18035(.A1(\b[48] ), .A2(new_n8835), .B(new_n18289), .C(new_n8826), .Y(new_n18292));
  AND2x2_ASAP7_75t_L        g18036(.A(new_n18292), .B(new_n18291), .Y(new_n18293));
  NAND3xp33_ASAP7_75t_L     g18037(.A(new_n18285), .B(new_n18287), .C(new_n18293), .Y(new_n18294));
  AO21x2_ASAP7_75t_L        g18038(.A1(new_n18287), .A2(new_n18285), .B(new_n18293), .Y(new_n18295));
  AND2x2_ASAP7_75t_L        g18039(.A(new_n18294), .B(new_n18295), .Y(new_n18296));
  INVx1_ASAP7_75t_L         g18040(.A(new_n18296), .Y(new_n18297));
  AOI21xp33_ASAP7_75t_L     g18041(.A1(new_n18185), .A2(new_n18149), .B(new_n18189), .Y(new_n18298));
  INVx1_ASAP7_75t_L         g18042(.A(new_n18298), .Y(new_n18299));
  NOR2xp33_ASAP7_75t_L      g18043(.A(new_n18297), .B(new_n18299), .Y(new_n18300));
  INVx1_ASAP7_75t_L         g18044(.A(new_n18300), .Y(new_n18301));
  A2O1A1Ixp33_ASAP7_75t_L   g18045(.A1(new_n18185), .A2(new_n18149), .B(new_n18189), .C(new_n18297), .Y(new_n18302));
  NAND2xp33_ASAP7_75t_L     g18046(.A(new_n18302), .B(new_n18301), .Y(new_n18303));
  AOI22xp33_ASAP7_75t_L     g18047(.A1(new_n7960), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n8537), .Y(new_n18304));
  OAI221xp5_ASAP7_75t_L     g18048(.A1(new_n8817), .A2(new_n7616), .B1(new_n7957), .B2(new_n7906), .C(new_n18304), .Y(new_n18305));
  XNOR2x2_ASAP7_75t_L       g18049(.A(\a[53] ), .B(new_n18305), .Y(new_n18306));
  INVx1_ASAP7_75t_L         g18050(.A(new_n18306), .Y(new_n18307));
  NOR2xp33_ASAP7_75t_L      g18051(.A(new_n18307), .B(new_n18303), .Y(new_n18308));
  INVx1_ASAP7_75t_L         g18052(.A(new_n18308), .Y(new_n18309));
  NAND2xp33_ASAP7_75t_L     g18053(.A(new_n18307), .B(new_n18303), .Y(new_n18310));
  AND2x2_ASAP7_75t_L        g18054(.A(new_n18310), .B(new_n18309), .Y(new_n18311));
  INVx1_ASAP7_75t_L         g18055(.A(new_n18311), .Y(new_n18312));
  O2A1O1Ixp33_ASAP7_75t_L   g18056(.A1(new_n18070), .A2(new_n18077), .B(new_n18195), .C(new_n18196), .Y(new_n18313));
  NAND2xp33_ASAP7_75t_L     g18057(.A(new_n18313), .B(new_n18312), .Y(new_n18314));
  A2O1A1Ixp33_ASAP7_75t_L   g18058(.A1(new_n18195), .A2(new_n18201), .B(new_n18196), .C(new_n18311), .Y(new_n18315));
  AND2x2_ASAP7_75t_L        g18059(.A(new_n18315), .B(new_n18314), .Y(new_n18316));
  NAND2xp33_ASAP7_75t_L     g18060(.A(\b[53] ), .B(new_n7391), .Y(new_n18317));
  OAI221xp5_ASAP7_75t_L     g18061(.A1(new_n7389), .A2(new_n8762), .B1(new_n8237), .B2(new_n8768), .C(new_n18317), .Y(new_n18318));
  AOI21xp33_ASAP7_75t_L     g18062(.A1(new_n7115), .A2(\b[54] ), .B(new_n18318), .Y(new_n18319));
  NAND2xp33_ASAP7_75t_L     g18063(.A(\a[50] ), .B(new_n18319), .Y(new_n18320));
  A2O1A1Ixp33_ASAP7_75t_L   g18064(.A1(\b[54] ), .A2(new_n7115), .B(new_n18318), .C(new_n7106), .Y(new_n18321));
  AND2x2_ASAP7_75t_L        g18065(.A(new_n18321), .B(new_n18320), .Y(new_n18322));
  INVx1_ASAP7_75t_L         g18066(.A(new_n18322), .Y(new_n18323));
  XNOR2x2_ASAP7_75t_L       g18067(.A(new_n18323), .B(new_n18316), .Y(new_n18324));
  INVx1_ASAP7_75t_L         g18068(.A(new_n18324), .Y(new_n18325));
  NAND3xp33_ASAP7_75t_L     g18069(.A(new_n18325), .B(new_n18207), .C(new_n18204), .Y(new_n18326));
  INVx1_ASAP7_75t_L         g18070(.A(new_n18207), .Y(new_n18327));
  A2O1A1Ixp33_ASAP7_75t_L   g18071(.A1(new_n18203), .A2(new_n18145), .B(new_n18327), .C(new_n18324), .Y(new_n18328));
  NAND2xp33_ASAP7_75t_L     g18072(.A(\b[56] ), .B(new_n6648), .Y(new_n18329));
  OAI221xp5_ASAP7_75t_L     g18073(.A1(new_n6880), .A2(new_n9920), .B1(new_n6636), .B2(new_n9925), .C(new_n18329), .Y(new_n18330));
  AOI21xp33_ASAP7_75t_L     g18074(.A1(new_n6380), .A2(\b[57] ), .B(new_n18330), .Y(new_n18331));
  NAND2xp33_ASAP7_75t_L     g18075(.A(\a[47] ), .B(new_n18331), .Y(new_n18332));
  A2O1A1Ixp33_ASAP7_75t_L   g18076(.A1(\b[57] ), .A2(new_n6380), .B(new_n18330), .C(new_n6371), .Y(new_n18333));
  AND2x2_ASAP7_75t_L        g18077(.A(new_n18333), .B(new_n18332), .Y(new_n18334));
  NAND3xp33_ASAP7_75t_L     g18078(.A(new_n18326), .B(new_n18328), .C(new_n18334), .Y(new_n18335));
  AO21x2_ASAP7_75t_L        g18079(.A1(new_n18328), .A2(new_n18326), .B(new_n18334), .Y(new_n18336));
  NAND2xp33_ASAP7_75t_L     g18080(.A(new_n18335), .B(new_n18336), .Y(new_n18337));
  NOR2xp33_ASAP7_75t_L      g18081(.A(new_n18212), .B(new_n18209), .Y(new_n18338));
  NOR3xp33_ASAP7_75t_L      g18082(.A(new_n18217), .B(new_n18337), .C(new_n18338), .Y(new_n18339));
  A2O1A1Ixp33_ASAP7_75t_L   g18083(.A1(new_n18215), .A2(new_n18214), .B(new_n18338), .C(new_n18337), .Y(new_n18340));
  INVx1_ASAP7_75t_L         g18084(.A(new_n18340), .Y(new_n18341));
  NOR2xp33_ASAP7_75t_L      g18085(.A(new_n18339), .B(new_n18341), .Y(new_n18342));
  NAND2xp33_ASAP7_75t_L     g18086(.A(\b[59] ), .B(new_n5901), .Y(new_n18343));
  OAI221xp5_ASAP7_75t_L     g18087(.A1(new_n5894), .A2(new_n10847), .B1(new_n5892), .B2(new_n10855), .C(new_n18343), .Y(new_n18344));
  AOI21xp33_ASAP7_75t_L     g18088(.A1(new_n5628), .A2(\b[60] ), .B(new_n18344), .Y(new_n18345));
  NAND2xp33_ASAP7_75t_L     g18089(.A(\a[44] ), .B(new_n18345), .Y(new_n18346));
  A2O1A1Ixp33_ASAP7_75t_L   g18090(.A1(\b[60] ), .A2(new_n5628), .B(new_n18344), .C(new_n5619), .Y(new_n18347));
  NAND2xp33_ASAP7_75t_L     g18091(.A(new_n18347), .B(new_n18346), .Y(new_n18348));
  NAND2xp33_ASAP7_75t_L     g18092(.A(new_n18348), .B(new_n18342), .Y(new_n18349));
  INVx1_ASAP7_75t_L         g18093(.A(new_n18349), .Y(new_n18350));
  NOR2xp33_ASAP7_75t_L      g18094(.A(new_n18348), .B(new_n18342), .Y(new_n18351));
  NOR2xp33_ASAP7_75t_L      g18095(.A(new_n18351), .B(new_n18350), .Y(new_n18352));
  NAND2xp33_ASAP7_75t_L     g18096(.A(new_n18352), .B(new_n18258), .Y(new_n18353));
  INVx1_ASAP7_75t_L         g18097(.A(new_n18353), .Y(new_n18354));
  NOR2xp33_ASAP7_75t_L      g18098(.A(new_n18352), .B(new_n18258), .Y(new_n18355));
  NOR2xp33_ASAP7_75t_L      g18099(.A(new_n18355), .B(new_n18354), .Y(new_n18356));
  NOR2xp33_ASAP7_75t_L      g18100(.A(new_n18356), .B(new_n18250), .Y(new_n18357));
  INVx1_ASAP7_75t_L         g18101(.A(new_n18356), .Y(new_n18358));
  A2O1A1O1Ixp25_ASAP7_75t_L g18102(.A1(new_n18232), .A2(new_n18233), .B(new_n18228), .C(new_n18239), .D(new_n18358), .Y(new_n18359));
  NOR2xp33_ASAP7_75t_L      g18103(.A(new_n18359), .B(new_n18357), .Y(new_n18360));
  A2O1A1Ixp33_ASAP7_75t_L   g18104(.A1(new_n18247), .A2(new_n18244), .B(new_n18241), .C(new_n18360), .Y(new_n18361));
  INVx1_ASAP7_75t_L         g18105(.A(new_n18361), .Y(new_n18362));
  A2O1A1Ixp33_ASAP7_75t_L   g18106(.A1(new_n18135), .A2(new_n18131), .B(new_n18245), .C(new_n18242), .Y(new_n18363));
  NOR2xp33_ASAP7_75t_L      g18107(.A(new_n18360), .B(new_n18363), .Y(new_n18364));
  NOR2xp33_ASAP7_75t_L      g18108(.A(new_n18364), .B(new_n18362), .Y(\f[103] ));
  NAND2xp33_ASAP7_75t_L     g18109(.A(new_n18204), .B(new_n18207), .Y(new_n18366));
  INVx1_ASAP7_75t_L         g18110(.A(new_n18316), .Y(new_n18367));
  A2O1A1O1Ixp25_ASAP7_75t_L g18111(.A1(new_n18078), .A2(new_n18071), .B(new_n18199), .C(new_n18197), .D(new_n18311), .Y(new_n18368));
  AOI22xp33_ASAP7_75t_L     g18112(.A1(new_n7111), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n7391), .Y(new_n18369));
  OAI221xp5_ASAP7_75t_L     g18113(.A1(new_n8558), .A2(new_n8762), .B1(new_n8237), .B2(new_n9331), .C(new_n18369), .Y(new_n18370));
  XNOR2x2_ASAP7_75t_L       g18114(.A(\a[50] ), .B(new_n18370), .Y(new_n18371));
  AOI22xp33_ASAP7_75t_L     g18115(.A1(new_n7960), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n8537), .Y(new_n18372));
  OAI221xp5_ASAP7_75t_L     g18116(.A1(new_n8817), .A2(new_n7900), .B1(new_n7957), .B2(new_n8174), .C(new_n18372), .Y(new_n18373));
  XNOR2x2_ASAP7_75t_L       g18117(.A(\a[53] ), .B(new_n18373), .Y(new_n18374));
  AOI22xp33_ASAP7_75t_L     g18118(.A1(new_n9700), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n10027), .Y(new_n18375));
  OAI221xp5_ASAP7_75t_L     g18119(.A1(new_n10024), .A2(new_n6568), .B1(new_n9696), .B2(new_n6820), .C(new_n18375), .Y(new_n18376));
  XNOR2x2_ASAP7_75t_L       g18120(.A(\a[59] ), .B(new_n18376), .Y(new_n18377));
  INVx1_ASAP7_75t_L         g18121(.A(new_n18377), .Y(new_n18378));
  NAND2xp33_ASAP7_75t_L     g18122(.A(\b[40] ), .B(new_n11534), .Y(new_n18379));
  OAI211xp5_ASAP7_75t_L     g18123(.A1(new_n11253), .A2(new_n5321), .B(new_n18261), .C(new_n18379), .Y(new_n18380));
  A2O1A1Ixp33_ASAP7_75t_L   g18124(.A1(new_n14788), .A2(new_n14789), .B(new_n5321), .C(new_n18379), .Y(new_n18381));
  A2O1A1Ixp33_ASAP7_75t_L   g18125(.A1(new_n11533), .A2(\b[40] ), .B(new_n18260), .C(new_n18381), .Y(new_n18382));
  AND2x2_ASAP7_75t_L        g18126(.A(new_n18382), .B(new_n18380), .Y(new_n18383));
  A2O1A1Ixp33_ASAP7_75t_L   g18127(.A1(new_n18274), .A2(new_n18267), .B(new_n18264), .C(new_n18383), .Y(new_n18384));
  A2O1A1Ixp33_ASAP7_75t_L   g18128(.A1(new_n18272), .A2(new_n18273), .B(new_n18268), .C(new_n18265), .Y(new_n18385));
  AO21x2_ASAP7_75t_L        g18129(.A1(new_n18382), .A2(new_n18380), .B(new_n18385), .Y(new_n18386));
  AND2x2_ASAP7_75t_L        g18130(.A(new_n18384), .B(new_n18386), .Y(new_n18387));
  AOI22xp33_ASAP7_75t_L     g18131(.A1(\b[42] ), .A2(new_n10939), .B1(\b[44] ), .B2(new_n10938), .Y(new_n18388));
  OAI221xp5_ASAP7_75t_L     g18132(.A1(new_n10937), .A2(new_n5805), .B1(new_n10629), .B2(new_n5835), .C(new_n18388), .Y(new_n18389));
  XNOR2x2_ASAP7_75t_L       g18133(.A(\a[62] ), .B(new_n18389), .Y(new_n18390));
  NOR2xp33_ASAP7_75t_L      g18134(.A(new_n18390), .B(new_n18387), .Y(new_n18391));
  INVx1_ASAP7_75t_L         g18135(.A(new_n18391), .Y(new_n18392));
  NAND2xp33_ASAP7_75t_L     g18136(.A(new_n18390), .B(new_n18387), .Y(new_n18393));
  NAND3xp33_ASAP7_75t_L     g18137(.A(new_n18378), .B(new_n18392), .C(new_n18393), .Y(new_n18394));
  AO21x2_ASAP7_75t_L        g18138(.A1(new_n18393), .A2(new_n18392), .B(new_n18378), .Y(new_n18395));
  AND2x2_ASAP7_75t_L        g18139(.A(new_n18394), .B(new_n18395), .Y(new_n18396));
  A2O1A1O1Ixp25_ASAP7_75t_L g18140(.A1(new_n18169), .A2(new_n18163), .B(new_n18275), .C(new_n18282), .D(new_n18396), .Y(new_n18397));
  INVx1_ASAP7_75t_L         g18141(.A(new_n18396), .Y(new_n18398));
  A2O1A1Ixp33_ASAP7_75t_L   g18142(.A1(new_n18169), .A2(new_n18163), .B(new_n18275), .C(new_n18282), .Y(new_n18399));
  NOR2xp33_ASAP7_75t_L      g18143(.A(new_n18399), .B(new_n18398), .Y(new_n18400));
  NOR2xp33_ASAP7_75t_L      g18144(.A(new_n18397), .B(new_n18400), .Y(new_n18401));
  INVx1_ASAP7_75t_L         g18145(.A(new_n18401), .Y(new_n18402));
  AOI22xp33_ASAP7_75t_L     g18146(.A1(new_n8831), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n9115), .Y(new_n18403));
  OAI221xp5_ASAP7_75t_L     g18147(.A1(new_n10343), .A2(new_n7317), .B1(new_n10016), .B2(new_n7602), .C(new_n18403), .Y(new_n18404));
  XNOR2x2_ASAP7_75t_L       g18148(.A(\a[56] ), .B(new_n18404), .Y(new_n18405));
  NAND2xp33_ASAP7_75t_L     g18149(.A(new_n18405), .B(new_n18402), .Y(new_n18406));
  NOR2xp33_ASAP7_75t_L      g18150(.A(new_n18405), .B(new_n18402), .Y(new_n18407));
  INVx1_ASAP7_75t_L         g18151(.A(new_n18407), .Y(new_n18408));
  AND2x2_ASAP7_75t_L        g18152(.A(new_n18406), .B(new_n18408), .Y(new_n18409));
  AND3x1_ASAP7_75t_L        g18153(.A(new_n18409), .B(new_n18294), .C(new_n18285), .Y(new_n18410));
  A2O1A1Ixp33_ASAP7_75t_L   g18154(.A1(new_n18172), .A2(new_n18169), .B(new_n18176), .C(new_n18259), .Y(new_n18411));
  O2A1O1Ixp33_ASAP7_75t_L   g18155(.A1(new_n18286), .A2(new_n18411), .B(new_n18294), .C(new_n18409), .Y(new_n18412));
  NOR3xp33_ASAP7_75t_L      g18156(.A(new_n18410), .B(new_n18412), .C(new_n18374), .Y(new_n18413));
  INVx1_ASAP7_75t_L         g18157(.A(new_n18374), .Y(new_n18414));
  NOR2xp33_ASAP7_75t_L      g18158(.A(new_n18412), .B(new_n18410), .Y(new_n18415));
  NOR2xp33_ASAP7_75t_L      g18159(.A(new_n18414), .B(new_n18415), .Y(new_n18416));
  NOR2xp33_ASAP7_75t_L      g18160(.A(new_n18413), .B(new_n18416), .Y(new_n18417));
  NOR2xp33_ASAP7_75t_L      g18161(.A(new_n18300), .B(new_n18308), .Y(new_n18418));
  NAND2xp33_ASAP7_75t_L     g18162(.A(new_n18418), .B(new_n18417), .Y(new_n18419));
  INVx1_ASAP7_75t_L         g18163(.A(new_n18419), .Y(new_n18420));
  O2A1O1Ixp33_ASAP7_75t_L   g18164(.A1(new_n18303), .A2(new_n18307), .B(new_n18301), .C(new_n18417), .Y(new_n18421));
  OR3x1_ASAP7_75t_L         g18165(.A(new_n18420), .B(new_n18371), .C(new_n18421), .Y(new_n18422));
  OAI21xp33_ASAP7_75t_L     g18166(.A1(new_n18421), .A2(new_n18420), .B(new_n18371), .Y(new_n18423));
  AND2x2_ASAP7_75t_L        g18167(.A(new_n18423), .B(new_n18422), .Y(new_n18424));
  A2O1A1Ixp33_ASAP7_75t_L   g18168(.A1(new_n18367), .A2(new_n18323), .B(new_n18368), .C(new_n18424), .Y(new_n18425));
  INVx1_ASAP7_75t_L         g18169(.A(new_n18368), .Y(new_n18426));
  A2O1A1Ixp33_ASAP7_75t_L   g18170(.A1(new_n18314), .A2(new_n18315), .B(new_n18322), .C(new_n18426), .Y(new_n18427));
  NOR2xp33_ASAP7_75t_L      g18171(.A(new_n18427), .B(new_n18424), .Y(new_n18428));
  INVx1_ASAP7_75t_L         g18172(.A(new_n18428), .Y(new_n18429));
  AOI22xp33_ASAP7_75t_L     g18173(.A1(new_n6376), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n6648), .Y(new_n18430));
  OAI221xp5_ASAP7_75t_L     g18174(.A1(new_n6646), .A2(new_n9920), .B1(new_n6636), .B2(new_n11152), .C(new_n18430), .Y(new_n18431));
  XNOR2x2_ASAP7_75t_L       g18175(.A(\a[47] ), .B(new_n18431), .Y(new_n18432));
  NAND3xp33_ASAP7_75t_L     g18176(.A(new_n18429), .B(new_n18425), .C(new_n18432), .Y(new_n18433));
  INVx1_ASAP7_75t_L         g18177(.A(new_n18433), .Y(new_n18434));
  AOI21xp33_ASAP7_75t_L     g18178(.A1(new_n18429), .A2(new_n18425), .B(new_n18432), .Y(new_n18435));
  NOR2xp33_ASAP7_75t_L      g18179(.A(new_n18435), .B(new_n18434), .Y(new_n18436));
  INVx1_ASAP7_75t_L         g18180(.A(new_n18436), .Y(new_n18437));
  O2A1O1Ixp33_ASAP7_75t_L   g18181(.A1(new_n18366), .A2(new_n18324), .B(new_n18335), .C(new_n18437), .Y(new_n18438));
  INVx1_ASAP7_75t_L         g18182(.A(new_n18438), .Y(new_n18439));
  NAND3xp33_ASAP7_75t_L     g18183(.A(new_n18437), .B(new_n18335), .C(new_n18326), .Y(new_n18440));
  AOI22xp33_ASAP7_75t_L     g18184(.A1(new_n5624), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n5901), .Y(new_n18441));
  OAI221xp5_ASAP7_75t_L     g18185(.A1(new_n5900), .A2(new_n10847), .B1(new_n5892), .B2(new_n12047), .C(new_n18441), .Y(new_n18442));
  XNOR2x2_ASAP7_75t_L       g18186(.A(\a[44] ), .B(new_n18442), .Y(new_n18443));
  NAND3xp33_ASAP7_75t_L     g18187(.A(new_n18439), .B(new_n18440), .C(new_n18443), .Y(new_n18444));
  INVx1_ASAP7_75t_L         g18188(.A(new_n18444), .Y(new_n18445));
  AOI21xp33_ASAP7_75t_L     g18189(.A1(new_n18439), .A2(new_n18440), .B(new_n18443), .Y(new_n18446));
  NOR2xp33_ASAP7_75t_L      g18190(.A(new_n18446), .B(new_n18445), .Y(new_n18447));
  A2O1A1O1Ixp25_ASAP7_75t_L g18191(.A1(new_n4917), .A2(new_n12061), .B(new_n5167), .C(\b[63] ), .D(new_n4915), .Y(new_n18448));
  A2O1A1O1Ixp25_ASAP7_75t_L g18192(.A1(\b[61] ), .A2(new_n11471), .B(\b[62] ), .C(new_n4917), .D(new_n5167), .Y(new_n18449));
  NOR3xp33_ASAP7_75t_L      g18193(.A(new_n18449), .B(new_n11468), .C(\a[41] ), .Y(new_n18450));
  NOR2xp33_ASAP7_75t_L      g18194(.A(new_n18448), .B(new_n18450), .Y(new_n18451));
  A2O1A1O1Ixp25_ASAP7_75t_L g18195(.A1(new_n18346), .A2(new_n18347), .B(new_n18339), .C(new_n18340), .D(new_n18451), .Y(new_n18452));
  INVx1_ASAP7_75t_L         g18196(.A(new_n18452), .Y(new_n18453));
  NAND3xp33_ASAP7_75t_L     g18197(.A(new_n18349), .B(new_n18340), .C(new_n18451), .Y(new_n18454));
  NAND2xp33_ASAP7_75t_L     g18198(.A(new_n18453), .B(new_n18454), .Y(new_n18455));
  XNOR2x2_ASAP7_75t_L       g18199(.A(new_n18447), .B(new_n18455), .Y(new_n18456));
  O2A1O1Ixp33_ASAP7_75t_L   g18200(.A1(new_n18256), .A2(new_n18253), .B(new_n18353), .C(new_n18456), .Y(new_n18457));
  INVx1_ASAP7_75t_L         g18201(.A(new_n18457), .Y(new_n18458));
  A2O1A1O1Ixp25_ASAP7_75t_L g18202(.A1(new_n18222), .A2(new_n18218), .B(new_n18226), .C(new_n18254), .D(new_n18354), .Y(new_n18459));
  NAND2xp33_ASAP7_75t_L     g18203(.A(new_n18456), .B(new_n18459), .Y(new_n18460));
  AND2x2_ASAP7_75t_L        g18204(.A(new_n18458), .B(new_n18460), .Y(new_n18461));
  A2O1A1Ixp33_ASAP7_75t_L   g18205(.A1(new_n18363), .A2(new_n18360), .B(new_n18359), .C(new_n18461), .Y(new_n18462));
  A2O1A1O1Ixp25_ASAP7_75t_L g18206(.A1(new_n18244), .A2(new_n18247), .B(new_n18241), .C(new_n18360), .D(new_n18359), .Y(new_n18463));
  INVx1_ASAP7_75t_L         g18207(.A(new_n18461), .Y(new_n18464));
  NAND2xp33_ASAP7_75t_L     g18208(.A(new_n18464), .B(new_n18463), .Y(new_n18465));
  AND2x2_ASAP7_75t_L        g18209(.A(new_n18462), .B(new_n18465), .Y(\f[104] ));
  INVx1_ASAP7_75t_L         g18210(.A(new_n18359), .Y(new_n18467));
  INVx1_ASAP7_75t_L         g18211(.A(new_n18454), .Y(new_n18468));
  AOI22xp33_ASAP7_75t_L     g18212(.A1(new_n7111), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n7391), .Y(new_n18469));
  OAI221xp5_ASAP7_75t_L     g18213(.A1(new_n8558), .A2(new_n9323), .B1(new_n8237), .B2(new_n9627), .C(new_n18469), .Y(new_n18470));
  XNOR2x2_ASAP7_75t_L       g18214(.A(\a[50] ), .B(new_n18470), .Y(new_n18471));
  INVx1_ASAP7_75t_L         g18215(.A(new_n18471), .Y(new_n18472));
  NOR2xp33_ASAP7_75t_L      g18216(.A(new_n18400), .B(new_n18407), .Y(new_n18473));
  AOI22xp33_ASAP7_75t_L     g18217(.A1(new_n8831), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n9115), .Y(new_n18474));
  OAI221xp5_ASAP7_75t_L     g18218(.A1(new_n10343), .A2(new_n7593), .B1(new_n10016), .B2(new_n7623), .C(new_n18474), .Y(new_n18475));
  XNOR2x2_ASAP7_75t_L       g18219(.A(\a[56] ), .B(new_n18475), .Y(new_n18476));
  INVx1_ASAP7_75t_L         g18220(.A(new_n18476), .Y(new_n18477));
  A2O1A1Ixp33_ASAP7_75t_L   g18221(.A1(new_n11533), .A2(\b[40] ), .B(new_n18260), .C(\a[41] ), .Y(new_n18478));
  NOR2xp33_ASAP7_75t_L      g18222(.A(\a[41] ), .B(new_n18262), .Y(new_n18479));
  INVx1_ASAP7_75t_L         g18223(.A(new_n18479), .Y(new_n18480));
  AND2x2_ASAP7_75t_L        g18224(.A(new_n18478), .B(new_n18480), .Y(new_n18481));
  NOR2xp33_ASAP7_75t_L      g18225(.A(new_n5321), .B(new_n11535), .Y(new_n18482));
  O2A1O1Ixp33_ASAP7_75t_L   g18226(.A1(new_n11247), .A2(new_n11249), .B(\b[42] ), .C(new_n18482), .Y(new_n18483));
  NAND2xp33_ASAP7_75t_L     g18227(.A(new_n18483), .B(new_n18481), .Y(new_n18484));
  INVx1_ASAP7_75t_L         g18228(.A(new_n18481), .Y(new_n18485));
  A2O1A1Ixp33_ASAP7_75t_L   g18229(.A1(\b[42] ), .A2(new_n11533), .B(new_n18482), .C(new_n18485), .Y(new_n18486));
  AND2x2_ASAP7_75t_L        g18230(.A(new_n18484), .B(new_n18486), .Y(new_n18487));
  INVx1_ASAP7_75t_L         g18231(.A(new_n18487), .Y(new_n18488));
  AOI22xp33_ASAP7_75t_L     g18232(.A1(\b[43] ), .A2(new_n10939), .B1(\b[45] ), .B2(new_n10938), .Y(new_n18489));
  OAI221xp5_ASAP7_75t_L     g18233(.A1(new_n10937), .A2(new_n5829), .B1(new_n10629), .B2(new_n6329), .C(new_n18489), .Y(new_n18490));
  XNOR2x2_ASAP7_75t_L       g18234(.A(\a[62] ), .B(new_n18490), .Y(new_n18491));
  XNOR2x2_ASAP7_75t_L       g18235(.A(new_n18488), .B(new_n18491), .Y(new_n18492));
  INVx1_ASAP7_75t_L         g18236(.A(new_n18383), .Y(new_n18493));
  O2A1O1Ixp33_ASAP7_75t_L   g18237(.A1(new_n11253), .A2(new_n5321), .B(new_n18379), .C(new_n18262), .Y(new_n18494));
  A2O1A1O1Ixp25_ASAP7_75t_L g18238(.A1(new_n18267), .A2(new_n18274), .B(new_n18264), .C(new_n18493), .D(new_n18494), .Y(new_n18495));
  NAND2xp33_ASAP7_75t_L     g18239(.A(new_n18495), .B(new_n18492), .Y(new_n18496));
  INVx1_ASAP7_75t_L         g18240(.A(new_n18492), .Y(new_n18497));
  A2O1A1Ixp33_ASAP7_75t_L   g18241(.A1(new_n18385), .A2(new_n18493), .B(new_n18494), .C(new_n18497), .Y(new_n18498));
  AND2x2_ASAP7_75t_L        g18242(.A(new_n18496), .B(new_n18498), .Y(new_n18499));
  AOI22xp33_ASAP7_75t_L     g18243(.A1(new_n9700), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n10027), .Y(new_n18500));
  OAI221xp5_ASAP7_75t_L     g18244(.A1(new_n10024), .A2(new_n6812), .B1(new_n9696), .B2(new_n6837), .C(new_n18500), .Y(new_n18501));
  XNOR2x2_ASAP7_75t_L       g18245(.A(\a[59] ), .B(new_n18501), .Y(new_n18502));
  INVx1_ASAP7_75t_L         g18246(.A(new_n18502), .Y(new_n18503));
  XNOR2x2_ASAP7_75t_L       g18247(.A(new_n18503), .B(new_n18499), .Y(new_n18504));
  O2A1O1Ixp33_ASAP7_75t_L   g18248(.A1(new_n18387), .A2(new_n18390), .B(new_n18394), .C(new_n18504), .Y(new_n18505));
  A2O1A1Ixp33_ASAP7_75t_L   g18249(.A1(new_n18386), .A2(new_n18384), .B(new_n18390), .C(new_n18394), .Y(new_n18506));
  INVx1_ASAP7_75t_L         g18250(.A(new_n18506), .Y(new_n18507));
  AND2x2_ASAP7_75t_L        g18251(.A(new_n18507), .B(new_n18504), .Y(new_n18508));
  NOR2xp33_ASAP7_75t_L      g18252(.A(new_n18505), .B(new_n18508), .Y(new_n18509));
  XNOR2x2_ASAP7_75t_L       g18253(.A(new_n18477), .B(new_n18509), .Y(new_n18510));
  XNOR2x2_ASAP7_75t_L       g18254(.A(new_n18473), .B(new_n18510), .Y(new_n18511));
  AOI22xp33_ASAP7_75t_L     g18255(.A1(new_n7960), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n8537), .Y(new_n18512));
  OAI221xp5_ASAP7_75t_L     g18256(.A1(new_n8817), .A2(new_n8165), .B1(new_n7957), .B2(new_n8465), .C(new_n18512), .Y(new_n18513));
  XNOR2x2_ASAP7_75t_L       g18257(.A(\a[53] ), .B(new_n18513), .Y(new_n18514));
  AND2x2_ASAP7_75t_L        g18258(.A(new_n18514), .B(new_n18511), .Y(new_n18515));
  NOR2xp33_ASAP7_75t_L      g18259(.A(new_n18514), .B(new_n18511), .Y(new_n18516));
  NOR2xp33_ASAP7_75t_L      g18260(.A(new_n18516), .B(new_n18515), .Y(new_n18517));
  A2O1A1Ixp33_ASAP7_75t_L   g18261(.A1(new_n18415), .A2(new_n18414), .B(new_n18410), .C(new_n18517), .Y(new_n18518));
  OR3x1_ASAP7_75t_L         g18262(.A(new_n18517), .B(new_n18410), .C(new_n18413), .Y(new_n18519));
  AND2x2_ASAP7_75t_L        g18263(.A(new_n18518), .B(new_n18519), .Y(new_n18520));
  NOR2xp33_ASAP7_75t_L      g18264(.A(new_n18472), .B(new_n18520), .Y(new_n18521));
  NAND2xp33_ASAP7_75t_L     g18265(.A(new_n18472), .B(new_n18520), .Y(new_n18522));
  INVx1_ASAP7_75t_L         g18266(.A(new_n18522), .Y(new_n18523));
  NOR2xp33_ASAP7_75t_L      g18267(.A(new_n18521), .B(new_n18523), .Y(new_n18524));
  INVx1_ASAP7_75t_L         g18268(.A(new_n18524), .Y(new_n18525));
  O2A1O1Ixp33_ASAP7_75t_L   g18269(.A1(new_n18371), .A2(new_n18421), .B(new_n18419), .C(new_n18525), .Y(new_n18526));
  INVx1_ASAP7_75t_L         g18270(.A(new_n18526), .Y(new_n18527));
  NAND3xp33_ASAP7_75t_L     g18271(.A(new_n18525), .B(new_n18422), .C(new_n18419), .Y(new_n18528));
  AND2x2_ASAP7_75t_L        g18272(.A(new_n18528), .B(new_n18527), .Y(new_n18529));
  AOI22xp33_ASAP7_75t_L     g18273(.A1(new_n6376), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n6648), .Y(new_n18530));
  OAI221xp5_ASAP7_75t_L     g18274(.A1(new_n6646), .A2(new_n9947), .B1(new_n6636), .B2(new_n11446), .C(new_n18530), .Y(new_n18531));
  XNOR2x2_ASAP7_75t_L       g18275(.A(\a[47] ), .B(new_n18531), .Y(new_n18532));
  XOR2x2_ASAP7_75t_L        g18276(.A(new_n18532), .B(new_n18529), .Y(new_n18533));
  A2O1A1Ixp33_ASAP7_75t_L   g18277(.A1(new_n18432), .A2(new_n18425), .B(new_n18428), .C(new_n18533), .Y(new_n18534));
  OR3x1_ASAP7_75t_L         g18278(.A(new_n18533), .B(new_n18428), .C(new_n18434), .Y(new_n18535));
  NAND2xp33_ASAP7_75t_L     g18279(.A(new_n18534), .B(new_n18535), .Y(new_n18536));
  AOI22xp33_ASAP7_75t_L     g18280(.A1(new_n5624), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n5901), .Y(new_n18537));
  A2O1A1Ixp33_ASAP7_75t_L   g18281(.A1(new_n11470), .A2(new_n11473), .B(new_n5892), .C(new_n18537), .Y(new_n18538));
  AOI21xp33_ASAP7_75t_L     g18282(.A1(new_n5628), .A2(\b[62] ), .B(new_n18538), .Y(new_n18539));
  NAND2xp33_ASAP7_75t_L     g18283(.A(\a[44] ), .B(new_n18539), .Y(new_n18540));
  A2O1A1Ixp33_ASAP7_75t_L   g18284(.A1(\b[62] ), .A2(new_n5628), .B(new_n18538), .C(new_n5619), .Y(new_n18541));
  NAND2xp33_ASAP7_75t_L     g18285(.A(new_n18541), .B(new_n18540), .Y(new_n18542));
  XOR2x2_ASAP7_75t_L        g18286(.A(new_n18542), .B(new_n18536), .Y(new_n18543));
  A2O1A1Ixp33_ASAP7_75t_L   g18287(.A1(new_n18440), .A2(new_n18443), .B(new_n18438), .C(new_n18543), .Y(new_n18544));
  A2O1A1Ixp33_ASAP7_75t_L   g18288(.A1(new_n18335), .A2(new_n18326), .B(new_n18437), .C(new_n18444), .Y(new_n18545));
  NOR2xp33_ASAP7_75t_L      g18289(.A(new_n18545), .B(new_n18543), .Y(new_n18546));
  INVx1_ASAP7_75t_L         g18290(.A(new_n18546), .Y(new_n18547));
  NAND2xp33_ASAP7_75t_L     g18291(.A(new_n18544), .B(new_n18547), .Y(new_n18548));
  O2A1O1Ixp33_ASAP7_75t_L   g18292(.A1(new_n18447), .A2(new_n18468), .B(new_n18453), .C(new_n18548), .Y(new_n18549));
  INVx1_ASAP7_75t_L         g18293(.A(new_n18549), .Y(new_n18550));
  OAI211xp5_ASAP7_75t_L     g18294(.A1(new_n18447), .A2(new_n18468), .B(new_n18548), .C(new_n18453), .Y(new_n18551));
  AND2x2_ASAP7_75t_L        g18295(.A(new_n18551), .B(new_n18550), .Y(new_n18552));
  INVx1_ASAP7_75t_L         g18296(.A(new_n18552), .Y(new_n18553));
  A2O1A1O1Ixp25_ASAP7_75t_L g18297(.A1(new_n18467), .A2(new_n18361), .B(new_n18464), .C(new_n18458), .D(new_n18553), .Y(new_n18554));
  A2O1A1Ixp33_ASAP7_75t_L   g18298(.A1(new_n18361), .A2(new_n18467), .B(new_n18464), .C(new_n18458), .Y(new_n18555));
  NOR2xp33_ASAP7_75t_L      g18299(.A(new_n18552), .B(new_n18555), .Y(new_n18556));
  NOR2xp33_ASAP7_75t_L      g18300(.A(new_n18554), .B(new_n18556), .Y(\f[105] ));
  INVx1_ASAP7_75t_L         g18301(.A(new_n18529), .Y(new_n18558));
  OAI21xp33_ASAP7_75t_L     g18302(.A1(new_n18558), .A2(new_n18532), .B(new_n18535), .Y(new_n18559));
  OAI22xp33_ASAP7_75t_L     g18303(.A1(new_n11500), .A2(new_n5892), .B1(new_n11172), .B2(new_n5895), .Y(new_n18560));
  AOI21xp33_ASAP7_75t_L     g18304(.A1(new_n5628), .A2(\b[63] ), .B(new_n18560), .Y(new_n18561));
  NAND2xp33_ASAP7_75t_L     g18305(.A(\a[44] ), .B(new_n18561), .Y(new_n18562));
  A2O1A1Ixp33_ASAP7_75t_L   g18306(.A1(\b[63] ), .A2(new_n5628), .B(new_n18560), .C(new_n5619), .Y(new_n18563));
  NAND2xp33_ASAP7_75t_L     g18307(.A(new_n18563), .B(new_n18562), .Y(new_n18564));
  XNOR2x2_ASAP7_75t_L       g18308(.A(new_n18564), .B(new_n18559), .Y(new_n18565));
  NAND2xp33_ASAP7_75t_L     g18309(.A(\b[59] ), .B(new_n6648), .Y(new_n18566));
  OAI221xp5_ASAP7_75t_L     g18310(.A1(new_n6880), .A2(new_n10847), .B1(new_n6636), .B2(new_n10855), .C(new_n18566), .Y(new_n18567));
  AOI21xp33_ASAP7_75t_L     g18311(.A1(new_n6380), .A2(\b[60] ), .B(new_n18567), .Y(new_n18568));
  NAND2xp33_ASAP7_75t_L     g18312(.A(\a[47] ), .B(new_n18568), .Y(new_n18569));
  A2O1A1Ixp33_ASAP7_75t_L   g18313(.A1(\b[60] ), .A2(new_n6380), .B(new_n18567), .C(new_n6371), .Y(new_n18570));
  AND2x2_ASAP7_75t_L        g18314(.A(new_n18570), .B(new_n18569), .Y(new_n18571));
  NOR2xp33_ASAP7_75t_L      g18315(.A(new_n5338), .B(new_n11535), .Y(new_n18572));
  O2A1O1Ixp33_ASAP7_75t_L   g18316(.A1(new_n11247), .A2(new_n11249), .B(\b[43] ), .C(new_n18572), .Y(new_n18573));
  INVx1_ASAP7_75t_L         g18317(.A(new_n18486), .Y(new_n18574));
  A2O1A1O1Ixp25_ASAP7_75t_L g18318(.A1(new_n11533), .A2(\b[40] ), .B(new_n18260), .C(new_n4915), .D(new_n18574), .Y(new_n18575));
  NAND2xp33_ASAP7_75t_L     g18319(.A(new_n18573), .B(new_n18575), .Y(new_n18576));
  INVx1_ASAP7_75t_L         g18320(.A(new_n18573), .Y(new_n18577));
  A2O1A1Ixp33_ASAP7_75t_L   g18321(.A1(new_n18262), .A2(new_n4915), .B(new_n18574), .C(new_n18577), .Y(new_n18578));
  AND2x2_ASAP7_75t_L        g18322(.A(new_n18578), .B(new_n18576), .Y(new_n18579));
  NOR2xp33_ASAP7_75t_L      g18323(.A(new_n6568), .B(new_n10630), .Y(new_n18580));
  AOI221xp5_ASAP7_75t_L     g18324(.A1(\b[44] ), .A2(new_n10939), .B1(\b[45] ), .B2(new_n10632), .C(new_n18580), .Y(new_n18581));
  OAI211xp5_ASAP7_75t_L     g18325(.A1(new_n10629), .A2(new_n6573), .B(\a[62] ), .C(new_n18581), .Y(new_n18582));
  INVx1_ASAP7_75t_L         g18326(.A(new_n18582), .Y(new_n18583));
  O2A1O1Ixp33_ASAP7_75t_L   g18327(.A1(new_n10629), .A2(new_n6573), .B(new_n18581), .C(\a[62] ), .Y(new_n18584));
  NOR2xp33_ASAP7_75t_L      g18328(.A(new_n18584), .B(new_n18583), .Y(new_n18585));
  NOR2xp33_ASAP7_75t_L      g18329(.A(new_n18579), .B(new_n18585), .Y(new_n18586));
  INVx1_ASAP7_75t_L         g18330(.A(new_n18586), .Y(new_n18587));
  NAND2xp33_ASAP7_75t_L     g18331(.A(new_n18579), .B(new_n18585), .Y(new_n18588));
  AND2x2_ASAP7_75t_L        g18332(.A(new_n18588), .B(new_n18587), .Y(new_n18589));
  INVx1_ASAP7_75t_L         g18333(.A(new_n18589), .Y(new_n18590));
  O2A1O1Ixp33_ASAP7_75t_L   g18334(.A1(new_n18488), .A2(new_n18491), .B(new_n18498), .C(new_n18590), .Y(new_n18591));
  OA211x2_ASAP7_75t_L       g18335(.A1(new_n18491), .A2(new_n18488), .B(new_n18590), .C(new_n18498), .Y(new_n18592));
  NOR2xp33_ASAP7_75t_L      g18336(.A(new_n18591), .B(new_n18592), .Y(new_n18593));
  AOI22xp33_ASAP7_75t_L     g18337(.A1(new_n9700), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n10027), .Y(new_n18594));
  OAI221xp5_ASAP7_75t_L     g18338(.A1(new_n10024), .A2(new_n6830), .B1(new_n9696), .B2(new_n7323), .C(new_n18594), .Y(new_n18595));
  XNOR2x2_ASAP7_75t_L       g18339(.A(\a[59] ), .B(new_n18595), .Y(new_n18596));
  AND2x2_ASAP7_75t_L        g18340(.A(new_n18596), .B(new_n18593), .Y(new_n18597));
  NOR2xp33_ASAP7_75t_L      g18341(.A(new_n18596), .B(new_n18593), .Y(new_n18598));
  NAND2xp33_ASAP7_75t_L     g18342(.A(new_n18503), .B(new_n18499), .Y(new_n18599));
  A2O1A1Ixp33_ASAP7_75t_L   g18343(.A1(new_n18394), .A2(new_n18392), .B(new_n18504), .C(new_n18599), .Y(new_n18600));
  OR3x1_ASAP7_75t_L         g18344(.A(new_n18597), .B(new_n18598), .C(new_n18600), .Y(new_n18601));
  NOR2xp33_ASAP7_75t_L      g18345(.A(new_n18598), .B(new_n18597), .Y(new_n18602));
  O2A1O1Ixp33_ASAP7_75t_L   g18346(.A1(new_n18507), .A2(new_n18504), .B(new_n18599), .C(new_n18602), .Y(new_n18603));
  INVx1_ASAP7_75t_L         g18347(.A(new_n18603), .Y(new_n18604));
  NAND2xp33_ASAP7_75t_L     g18348(.A(\b[50] ), .B(new_n9115), .Y(new_n18605));
  OAI221xp5_ASAP7_75t_L     g18349(.A1(new_n9113), .A2(new_n7900), .B1(new_n10016), .B2(new_n7906), .C(new_n18605), .Y(new_n18606));
  AOI21xp33_ASAP7_75t_L     g18350(.A1(new_n8835), .A2(\b[51] ), .B(new_n18606), .Y(new_n18607));
  NAND2xp33_ASAP7_75t_L     g18351(.A(\a[56] ), .B(new_n18607), .Y(new_n18608));
  A2O1A1Ixp33_ASAP7_75t_L   g18352(.A1(\b[51] ), .A2(new_n8835), .B(new_n18606), .C(new_n8826), .Y(new_n18609));
  AND2x2_ASAP7_75t_L        g18353(.A(new_n18609), .B(new_n18608), .Y(new_n18610));
  NAND3xp33_ASAP7_75t_L     g18354(.A(new_n18604), .B(new_n18601), .C(new_n18610), .Y(new_n18611));
  AO21x2_ASAP7_75t_L        g18355(.A1(new_n18601), .A2(new_n18604), .B(new_n18610), .Y(new_n18612));
  AND2x2_ASAP7_75t_L        g18356(.A(new_n18611), .B(new_n18612), .Y(new_n18613));
  INVx1_ASAP7_75t_L         g18357(.A(new_n18613), .Y(new_n18614));
  O2A1O1Ixp33_ASAP7_75t_L   g18358(.A1(new_n18398), .A2(new_n18399), .B(new_n18408), .C(new_n18510), .Y(new_n18615));
  AOI21xp33_ASAP7_75t_L     g18359(.A1(new_n18509), .A2(new_n18477), .B(new_n18615), .Y(new_n18616));
  INVx1_ASAP7_75t_L         g18360(.A(new_n18616), .Y(new_n18617));
  NOR2xp33_ASAP7_75t_L      g18361(.A(new_n18617), .B(new_n18614), .Y(new_n18618));
  INVx1_ASAP7_75t_L         g18362(.A(new_n18618), .Y(new_n18619));
  A2O1A1Ixp33_ASAP7_75t_L   g18363(.A1(new_n18477), .A2(new_n18509), .B(new_n18615), .C(new_n18614), .Y(new_n18620));
  AOI22xp33_ASAP7_75t_L     g18364(.A1(new_n7960), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n8537), .Y(new_n18621));
  OAI221xp5_ASAP7_75t_L     g18365(.A1(new_n8817), .A2(new_n8458), .B1(new_n7957), .B2(new_n8768), .C(new_n18621), .Y(new_n18622));
  XNOR2x2_ASAP7_75t_L       g18366(.A(\a[53] ), .B(new_n18622), .Y(new_n18623));
  NAND3xp33_ASAP7_75t_L     g18367(.A(new_n18619), .B(new_n18620), .C(new_n18623), .Y(new_n18624));
  AO21x2_ASAP7_75t_L        g18368(.A1(new_n18620), .A2(new_n18619), .B(new_n18623), .Y(new_n18625));
  AND2x2_ASAP7_75t_L        g18369(.A(new_n18624), .B(new_n18625), .Y(new_n18626));
  INVx1_ASAP7_75t_L         g18370(.A(new_n18626), .Y(new_n18627));
  O2A1O1Ixp33_ASAP7_75t_L   g18371(.A1(new_n18511), .A2(new_n18514), .B(new_n18518), .C(new_n18627), .Y(new_n18628));
  O2A1O1Ixp33_ASAP7_75t_L   g18372(.A1(new_n18413), .A2(new_n18410), .B(new_n18517), .C(new_n18516), .Y(new_n18629));
  AND2x2_ASAP7_75t_L        g18373(.A(new_n18629), .B(new_n18627), .Y(new_n18630));
  NOR2xp33_ASAP7_75t_L      g18374(.A(new_n18628), .B(new_n18630), .Y(new_n18631));
  AOI22xp33_ASAP7_75t_L     g18375(.A1(new_n7111), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n7391), .Y(new_n18632));
  OAI221xp5_ASAP7_75t_L     g18376(.A1(new_n8558), .A2(new_n9620), .B1(new_n8237), .B2(new_n9925), .C(new_n18632), .Y(new_n18633));
  XNOR2x2_ASAP7_75t_L       g18377(.A(\a[50] ), .B(new_n18633), .Y(new_n18634));
  INVx1_ASAP7_75t_L         g18378(.A(new_n18634), .Y(new_n18635));
  XNOR2x2_ASAP7_75t_L       g18379(.A(new_n18635), .B(new_n18631), .Y(new_n18636));
  A2O1A1Ixp33_ASAP7_75t_L   g18380(.A1(new_n18520), .A2(new_n18472), .B(new_n18526), .C(new_n18636), .Y(new_n18637));
  A2O1A1Ixp33_ASAP7_75t_L   g18381(.A1(new_n18422), .A2(new_n18419), .B(new_n18521), .C(new_n18522), .Y(new_n18638));
  NOR2xp33_ASAP7_75t_L      g18382(.A(new_n18638), .B(new_n18636), .Y(new_n18639));
  INVx1_ASAP7_75t_L         g18383(.A(new_n18639), .Y(new_n18640));
  AOI21xp33_ASAP7_75t_L     g18384(.A1(new_n18640), .A2(new_n18637), .B(new_n18571), .Y(new_n18641));
  AND3x1_ASAP7_75t_L        g18385(.A(new_n18640), .B(new_n18637), .C(new_n18571), .Y(new_n18642));
  NOR2xp33_ASAP7_75t_L      g18386(.A(new_n18641), .B(new_n18642), .Y(new_n18643));
  XNOR2x2_ASAP7_75t_L       g18387(.A(new_n18643), .B(new_n18565), .Y(new_n18644));
  A2O1A1Ixp33_ASAP7_75t_L   g18388(.A1(new_n18540), .A2(new_n18541), .B(new_n18536), .C(new_n18547), .Y(new_n18645));
  INVx1_ASAP7_75t_L         g18389(.A(new_n18645), .Y(new_n18646));
  NAND2xp33_ASAP7_75t_L     g18390(.A(new_n18644), .B(new_n18646), .Y(new_n18647));
  A2O1A1O1Ixp25_ASAP7_75t_L g18391(.A1(new_n18540), .A2(new_n18541), .B(new_n18536), .C(new_n18547), .D(new_n18644), .Y(new_n18648));
  INVx1_ASAP7_75t_L         g18392(.A(new_n18648), .Y(new_n18649));
  AND2x2_ASAP7_75t_L        g18393(.A(new_n18649), .B(new_n18647), .Y(new_n18650));
  A2O1A1Ixp33_ASAP7_75t_L   g18394(.A1(new_n18555), .A2(new_n18552), .B(new_n18549), .C(new_n18650), .Y(new_n18651));
  INVx1_ASAP7_75t_L         g18395(.A(new_n18651), .Y(new_n18652));
  A2O1A1Ixp33_ASAP7_75t_L   g18396(.A1(new_n18462), .A2(new_n18458), .B(new_n18553), .C(new_n18550), .Y(new_n18653));
  NOR2xp33_ASAP7_75t_L      g18397(.A(new_n18650), .B(new_n18653), .Y(new_n18654));
  NOR2xp33_ASAP7_75t_L      g18398(.A(new_n18654), .B(new_n18652), .Y(\f[106] ));
  INVx1_ASAP7_75t_L         g18399(.A(new_n18643), .Y(new_n18656));
  MAJIxp5_ASAP7_75t_L       g18400(.A(new_n18559), .B(new_n18564), .C(new_n18656), .Y(new_n18657));
  AOI22xp33_ASAP7_75t_L     g18401(.A1(new_n6376), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n6648), .Y(new_n18658));
  OAI221xp5_ASAP7_75t_L     g18402(.A1(new_n6646), .A2(new_n10847), .B1(new_n6636), .B2(new_n12047), .C(new_n18658), .Y(new_n18659));
  XNOR2x2_ASAP7_75t_L       g18403(.A(\a[47] ), .B(new_n18659), .Y(new_n18660));
  INVx1_ASAP7_75t_L         g18404(.A(new_n18631), .Y(new_n18661));
  AOI22xp33_ASAP7_75t_L     g18405(.A1(new_n7960), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n8537), .Y(new_n18662));
  OAI221xp5_ASAP7_75t_L     g18406(.A1(new_n8817), .A2(new_n8762), .B1(new_n7957), .B2(new_n9331), .C(new_n18662), .Y(new_n18663));
  XNOR2x2_ASAP7_75t_L       g18407(.A(\a[53] ), .B(new_n18663), .Y(new_n18664));
  AOI22xp33_ASAP7_75t_L     g18408(.A1(new_n8831), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n9115), .Y(new_n18665));
  OAI221xp5_ASAP7_75t_L     g18409(.A1(new_n10343), .A2(new_n7900), .B1(new_n10016), .B2(new_n8174), .C(new_n18665), .Y(new_n18666));
  XNOR2x2_ASAP7_75t_L       g18410(.A(\a[56] ), .B(new_n18666), .Y(new_n18667));
  INVx1_ASAP7_75t_L         g18411(.A(new_n18667), .Y(new_n18668));
  AOI22xp33_ASAP7_75t_L     g18412(.A1(new_n9700), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n10027), .Y(new_n18669));
  OAI221xp5_ASAP7_75t_L     g18413(.A1(new_n10024), .A2(new_n7317), .B1(new_n9696), .B2(new_n7602), .C(new_n18669), .Y(new_n18670));
  XNOR2x2_ASAP7_75t_L       g18414(.A(\a[59] ), .B(new_n18670), .Y(new_n18671));
  NAND2xp33_ASAP7_75t_L     g18415(.A(\b[43] ), .B(new_n11534), .Y(new_n18672));
  O2A1O1Ixp33_ASAP7_75t_L   g18416(.A1(new_n11253), .A2(new_n5829), .B(new_n18672), .C(new_n18577), .Y(new_n18673));
  INVx1_ASAP7_75t_L         g18417(.A(new_n18572), .Y(new_n18674));
  A2O1A1Ixp33_ASAP7_75t_L   g18418(.A1(new_n14788), .A2(new_n14789), .B(new_n5829), .C(new_n18672), .Y(new_n18675));
  O2A1O1Ixp33_ASAP7_75t_L   g18419(.A1(new_n5805), .A2(new_n11253), .B(new_n18674), .C(new_n18675), .Y(new_n18676));
  NOR2xp33_ASAP7_75t_L      g18420(.A(new_n6812), .B(new_n10630), .Y(new_n18677));
  AOI221xp5_ASAP7_75t_L     g18421(.A1(\b[45] ), .A2(new_n10939), .B1(\b[46] ), .B2(new_n10632), .C(new_n18677), .Y(new_n18678));
  OA21x2_ASAP7_75t_L        g18422(.A1(new_n10629), .A2(new_n6820), .B(new_n18678), .Y(new_n18679));
  NAND2xp33_ASAP7_75t_L     g18423(.A(\a[62] ), .B(new_n18679), .Y(new_n18680));
  INVx1_ASAP7_75t_L         g18424(.A(new_n18680), .Y(new_n18681));
  O2A1O1Ixp33_ASAP7_75t_L   g18425(.A1(new_n10629), .A2(new_n6820), .B(new_n18678), .C(\a[62] ), .Y(new_n18682));
  NOR2xp33_ASAP7_75t_L      g18426(.A(new_n18682), .B(new_n18681), .Y(new_n18683));
  NOR3xp33_ASAP7_75t_L      g18427(.A(new_n18683), .B(new_n18676), .C(new_n18673), .Y(new_n18684));
  NOR2xp33_ASAP7_75t_L      g18428(.A(new_n18676), .B(new_n18673), .Y(new_n18685));
  INVx1_ASAP7_75t_L         g18429(.A(new_n18683), .Y(new_n18686));
  NOR2xp33_ASAP7_75t_L      g18430(.A(new_n18685), .B(new_n18686), .Y(new_n18687));
  NOR2xp33_ASAP7_75t_L      g18431(.A(new_n18684), .B(new_n18687), .Y(new_n18688));
  INVx1_ASAP7_75t_L         g18432(.A(new_n18688), .Y(new_n18689));
  O2A1O1Ixp33_ASAP7_75t_L   g18433(.A1(new_n18577), .A2(new_n18575), .B(new_n18587), .C(new_n18689), .Y(new_n18690));
  INVx1_ASAP7_75t_L         g18434(.A(new_n18690), .Y(new_n18691));
  A2O1A1O1Ixp25_ASAP7_75t_L g18435(.A1(new_n18262), .A2(new_n4915), .B(new_n18574), .C(new_n18573), .D(new_n18586), .Y(new_n18692));
  NAND2xp33_ASAP7_75t_L     g18436(.A(new_n18692), .B(new_n18689), .Y(new_n18693));
  NAND2xp33_ASAP7_75t_L     g18437(.A(new_n18693), .B(new_n18691), .Y(new_n18694));
  NOR2xp33_ASAP7_75t_L      g18438(.A(new_n18671), .B(new_n18694), .Y(new_n18695));
  INVx1_ASAP7_75t_L         g18439(.A(new_n18695), .Y(new_n18696));
  NAND2xp33_ASAP7_75t_L     g18440(.A(new_n18671), .B(new_n18694), .Y(new_n18697));
  AND2x2_ASAP7_75t_L        g18441(.A(new_n18697), .B(new_n18696), .Y(new_n18698));
  INVx1_ASAP7_75t_L         g18442(.A(new_n18698), .Y(new_n18699));
  OR3x1_ASAP7_75t_L         g18443(.A(new_n18699), .B(new_n18592), .C(new_n18597), .Y(new_n18700));
  A2O1A1Ixp33_ASAP7_75t_L   g18444(.A1(new_n18593), .A2(new_n18596), .B(new_n18592), .C(new_n18699), .Y(new_n18701));
  NAND3xp33_ASAP7_75t_L     g18445(.A(new_n18701), .B(new_n18700), .C(new_n18668), .Y(new_n18702));
  AO21x2_ASAP7_75t_L        g18446(.A1(new_n18701), .A2(new_n18700), .B(new_n18668), .Y(new_n18703));
  AND2x2_ASAP7_75t_L        g18447(.A(new_n18702), .B(new_n18703), .Y(new_n18704));
  AND3x1_ASAP7_75t_L        g18448(.A(new_n18704), .B(new_n18611), .C(new_n18601), .Y(new_n18705));
  INVx1_ASAP7_75t_L         g18449(.A(new_n18610), .Y(new_n18706));
  O2A1O1Ixp33_ASAP7_75t_L   g18450(.A1(new_n18603), .A2(new_n18706), .B(new_n18601), .C(new_n18704), .Y(new_n18707));
  NOR2xp33_ASAP7_75t_L      g18451(.A(new_n18707), .B(new_n18705), .Y(new_n18708));
  XNOR2x2_ASAP7_75t_L       g18452(.A(new_n18664), .B(new_n18708), .Y(new_n18709));
  NAND3xp33_ASAP7_75t_L     g18453(.A(new_n18709), .B(new_n18624), .C(new_n18619), .Y(new_n18710));
  O2A1O1Ixp33_ASAP7_75t_L   g18454(.A1(new_n18614), .A2(new_n18617), .B(new_n18624), .C(new_n18709), .Y(new_n18711));
  INVx1_ASAP7_75t_L         g18455(.A(new_n18711), .Y(new_n18712));
  AOI22xp33_ASAP7_75t_L     g18456(.A1(new_n7111), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n7391), .Y(new_n18713));
  OAI221xp5_ASAP7_75t_L     g18457(.A1(new_n8558), .A2(new_n9920), .B1(new_n8237), .B2(new_n11152), .C(new_n18713), .Y(new_n18714));
  XNOR2x2_ASAP7_75t_L       g18458(.A(\a[50] ), .B(new_n18714), .Y(new_n18715));
  NAND3xp33_ASAP7_75t_L     g18459(.A(new_n18712), .B(new_n18710), .C(new_n18715), .Y(new_n18716));
  AO21x2_ASAP7_75t_L        g18460(.A1(new_n18710), .A2(new_n18712), .B(new_n18715), .Y(new_n18717));
  AND2x2_ASAP7_75t_L        g18461(.A(new_n18716), .B(new_n18717), .Y(new_n18718));
  INVx1_ASAP7_75t_L         g18462(.A(new_n18718), .Y(new_n18719));
  O2A1O1Ixp33_ASAP7_75t_L   g18463(.A1(new_n18511), .A2(new_n18514), .B(new_n18518), .C(new_n18626), .Y(new_n18720));
  A2O1A1Ixp33_ASAP7_75t_L   g18464(.A1(new_n18661), .A2(new_n18635), .B(new_n18720), .C(new_n18719), .Y(new_n18721));
  O2A1O1Ixp33_ASAP7_75t_L   g18465(.A1(new_n18628), .A2(new_n18630), .B(new_n18635), .C(new_n18720), .Y(new_n18722));
  NAND2xp33_ASAP7_75t_L     g18466(.A(new_n18722), .B(new_n18718), .Y(new_n18723));
  NAND3xp33_ASAP7_75t_L     g18467(.A(new_n18721), .B(new_n18660), .C(new_n18723), .Y(new_n18724));
  AO21x2_ASAP7_75t_L        g18468(.A1(new_n18723), .A2(new_n18721), .B(new_n18660), .Y(new_n18725));
  NAND2xp33_ASAP7_75t_L     g18469(.A(new_n18724), .B(new_n18725), .Y(new_n18726));
  A2O1A1Ixp33_ASAP7_75t_L   g18470(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n5621), .Y(new_n18727));
  A2O1A1Ixp33_ASAP7_75t_L   g18471(.A1(new_n18727), .A2(new_n5895), .B(new_n11468), .C(\a[44] ), .Y(new_n18728));
  O2A1O1Ixp33_ASAP7_75t_L   g18472(.A1(new_n5892), .A2(new_n12060), .B(new_n5895), .C(new_n11468), .Y(new_n18729));
  NAND2xp33_ASAP7_75t_L     g18473(.A(new_n5619), .B(new_n18729), .Y(new_n18730));
  NAND2xp33_ASAP7_75t_L     g18474(.A(new_n18730), .B(new_n18728), .Y(new_n18731));
  NOR2xp33_ASAP7_75t_L      g18475(.A(new_n18639), .B(new_n18642), .Y(new_n18732));
  NAND2xp33_ASAP7_75t_L     g18476(.A(new_n18731), .B(new_n18732), .Y(new_n18733));
  NOR2xp33_ASAP7_75t_L      g18477(.A(new_n18731), .B(new_n18732), .Y(new_n18734));
  INVx1_ASAP7_75t_L         g18478(.A(new_n18734), .Y(new_n18735));
  NAND2xp33_ASAP7_75t_L     g18479(.A(new_n18733), .B(new_n18735), .Y(new_n18736));
  XOR2x2_ASAP7_75t_L        g18480(.A(new_n18726), .B(new_n18736), .Y(new_n18737));
  NOR2xp33_ASAP7_75t_L      g18481(.A(new_n18657), .B(new_n18737), .Y(new_n18738));
  INVx1_ASAP7_75t_L         g18482(.A(new_n18738), .Y(new_n18739));
  NAND2xp33_ASAP7_75t_L     g18483(.A(new_n18657), .B(new_n18737), .Y(new_n18740));
  AND2x2_ASAP7_75t_L        g18484(.A(new_n18740), .B(new_n18739), .Y(new_n18741));
  A2O1A1Ixp33_ASAP7_75t_L   g18485(.A1(new_n18653), .A2(new_n18650), .B(new_n18648), .C(new_n18741), .Y(new_n18742));
  A2O1A1O1Ixp25_ASAP7_75t_L g18486(.A1(new_n18552), .A2(new_n18555), .B(new_n18549), .C(new_n18650), .D(new_n18648), .Y(new_n18743));
  INVx1_ASAP7_75t_L         g18487(.A(new_n18741), .Y(new_n18744));
  NAND2xp33_ASAP7_75t_L     g18488(.A(new_n18744), .B(new_n18743), .Y(new_n18745));
  AND2x2_ASAP7_75t_L        g18489(.A(new_n18742), .B(new_n18745), .Y(\f[107] ));
  AOI22xp33_ASAP7_75t_L     g18490(.A1(new_n7111), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n7391), .Y(new_n18747));
  OAI221xp5_ASAP7_75t_L     g18491(.A1(new_n8558), .A2(new_n9947), .B1(new_n8237), .B2(new_n11446), .C(new_n18747), .Y(new_n18748));
  XNOR2x2_ASAP7_75t_L       g18492(.A(\a[50] ), .B(new_n18748), .Y(new_n18749));
  INVx1_ASAP7_75t_L         g18493(.A(new_n18664), .Y(new_n18750));
  AOI22xp33_ASAP7_75t_L     g18494(.A1(new_n7960), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n8537), .Y(new_n18751));
  OAI221xp5_ASAP7_75t_L     g18495(.A1(new_n8817), .A2(new_n9323), .B1(new_n7957), .B2(new_n9627), .C(new_n18751), .Y(new_n18752));
  XNOR2x2_ASAP7_75t_L       g18496(.A(\a[53] ), .B(new_n18752), .Y(new_n18753));
  NOR3xp33_ASAP7_75t_L      g18497(.A(new_n18699), .B(new_n18597), .C(new_n18592), .Y(new_n18754));
  AOI22xp33_ASAP7_75t_L     g18498(.A1(new_n8831), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n9115), .Y(new_n18755));
  OAI221xp5_ASAP7_75t_L     g18499(.A1(new_n10343), .A2(new_n8165), .B1(new_n10016), .B2(new_n8465), .C(new_n18755), .Y(new_n18756));
  XNOR2x2_ASAP7_75t_L       g18500(.A(\a[56] ), .B(new_n18756), .Y(new_n18757));
  INVx1_ASAP7_75t_L         g18501(.A(new_n18757), .Y(new_n18758));
  AOI22xp33_ASAP7_75t_L     g18502(.A1(new_n9700), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n10027), .Y(new_n18759));
  OAI221xp5_ASAP7_75t_L     g18503(.A1(new_n10024), .A2(new_n7593), .B1(new_n9696), .B2(new_n7623), .C(new_n18759), .Y(new_n18760));
  XNOR2x2_ASAP7_75t_L       g18504(.A(\a[59] ), .B(new_n18760), .Y(new_n18761));
  INVx1_ASAP7_75t_L         g18505(.A(new_n18761), .Y(new_n18762));
  AOI22xp33_ASAP7_75t_L     g18506(.A1(\b[46] ), .A2(new_n10939), .B1(\b[48] ), .B2(new_n10938), .Y(new_n18763));
  OAI221xp5_ASAP7_75t_L     g18507(.A1(new_n10937), .A2(new_n6812), .B1(new_n10629), .B2(new_n6837), .C(new_n18763), .Y(new_n18764));
  XNOR2x2_ASAP7_75t_L       g18508(.A(\a[62] ), .B(new_n18764), .Y(new_n18765));
  O2A1O1Ixp33_ASAP7_75t_L   g18509(.A1(new_n18682), .A2(new_n18681), .B(new_n18685), .C(new_n18673), .Y(new_n18766));
  NOR2xp33_ASAP7_75t_L      g18510(.A(new_n5829), .B(new_n11535), .Y(new_n18767));
  A2O1A1Ixp33_ASAP7_75t_L   g18511(.A1(new_n11533), .A2(\b[45] ), .B(new_n18767), .C(new_n5619), .Y(new_n18768));
  INVx1_ASAP7_75t_L         g18512(.A(new_n18768), .Y(new_n18769));
  O2A1O1Ixp33_ASAP7_75t_L   g18513(.A1(new_n11247), .A2(new_n11249), .B(\b[45] ), .C(new_n18767), .Y(new_n18770));
  NAND2xp33_ASAP7_75t_L     g18514(.A(\a[44] ), .B(new_n18770), .Y(new_n18771));
  INVx1_ASAP7_75t_L         g18515(.A(new_n18771), .Y(new_n18772));
  OAI21xp33_ASAP7_75t_L     g18516(.A1(new_n18769), .A2(new_n18772), .B(new_n18573), .Y(new_n18773));
  NOR2xp33_ASAP7_75t_L      g18517(.A(new_n18769), .B(new_n18772), .Y(new_n18774));
  A2O1A1Ixp33_ASAP7_75t_L   g18518(.A1(new_n11533), .A2(\b[43] ), .B(new_n18572), .C(new_n18774), .Y(new_n18775));
  AND2x2_ASAP7_75t_L        g18519(.A(new_n18773), .B(new_n18775), .Y(new_n18776));
  XNOR2x2_ASAP7_75t_L       g18520(.A(new_n18776), .B(new_n18766), .Y(new_n18777));
  INVx1_ASAP7_75t_L         g18521(.A(new_n18777), .Y(new_n18778));
  NOR2xp33_ASAP7_75t_L      g18522(.A(new_n18765), .B(new_n18778), .Y(new_n18779));
  INVx1_ASAP7_75t_L         g18523(.A(new_n18779), .Y(new_n18780));
  NAND2xp33_ASAP7_75t_L     g18524(.A(new_n18765), .B(new_n18778), .Y(new_n18781));
  AND2x2_ASAP7_75t_L        g18525(.A(new_n18781), .B(new_n18780), .Y(new_n18782));
  NOR2xp33_ASAP7_75t_L      g18526(.A(new_n18762), .B(new_n18782), .Y(new_n18783));
  NAND2xp33_ASAP7_75t_L     g18527(.A(new_n18762), .B(new_n18782), .Y(new_n18784));
  INVx1_ASAP7_75t_L         g18528(.A(new_n18784), .Y(new_n18785));
  NOR2xp33_ASAP7_75t_L      g18529(.A(new_n18783), .B(new_n18785), .Y(new_n18786));
  INVx1_ASAP7_75t_L         g18530(.A(new_n18786), .Y(new_n18787));
  O2A1O1Ixp33_ASAP7_75t_L   g18531(.A1(new_n18692), .A2(new_n18689), .B(new_n18696), .C(new_n18787), .Y(new_n18788));
  INVx1_ASAP7_75t_L         g18532(.A(new_n18788), .Y(new_n18789));
  A2O1A1Ixp33_ASAP7_75t_L   g18533(.A1(new_n11533), .A2(\b[40] ), .B(new_n18260), .C(new_n4915), .Y(new_n18790));
  A2O1A1O1Ixp25_ASAP7_75t_L g18534(.A1(new_n18478), .A2(new_n18480), .B(new_n18483), .C(new_n18790), .D(new_n18577), .Y(new_n18791));
  O2A1O1Ixp33_ASAP7_75t_L   g18535(.A1(new_n18586), .A2(new_n18791), .B(new_n18688), .C(new_n18695), .Y(new_n18792));
  NAND2xp33_ASAP7_75t_L     g18536(.A(new_n18792), .B(new_n18787), .Y(new_n18793));
  AO21x2_ASAP7_75t_L        g18537(.A1(new_n18793), .A2(new_n18789), .B(new_n18758), .Y(new_n18794));
  NAND3xp33_ASAP7_75t_L     g18538(.A(new_n18789), .B(new_n18758), .C(new_n18793), .Y(new_n18795));
  AND2x2_ASAP7_75t_L        g18539(.A(new_n18795), .B(new_n18794), .Y(new_n18796));
  A2O1A1Ixp33_ASAP7_75t_L   g18540(.A1(new_n18701), .A2(new_n18668), .B(new_n18754), .C(new_n18796), .Y(new_n18797));
  INVx1_ASAP7_75t_L         g18541(.A(new_n18796), .Y(new_n18798));
  NAND3xp33_ASAP7_75t_L     g18542(.A(new_n18798), .B(new_n18702), .C(new_n18700), .Y(new_n18799));
  AND2x2_ASAP7_75t_L        g18543(.A(new_n18797), .B(new_n18799), .Y(new_n18800));
  INVx1_ASAP7_75t_L         g18544(.A(new_n18800), .Y(new_n18801));
  NAND2xp33_ASAP7_75t_L     g18545(.A(new_n18753), .B(new_n18801), .Y(new_n18802));
  INVx1_ASAP7_75t_L         g18546(.A(new_n18753), .Y(new_n18803));
  NAND2xp33_ASAP7_75t_L     g18547(.A(new_n18803), .B(new_n18800), .Y(new_n18804));
  AND2x2_ASAP7_75t_L        g18548(.A(new_n18804), .B(new_n18802), .Y(new_n18805));
  A2O1A1Ixp33_ASAP7_75t_L   g18549(.A1(new_n18708), .A2(new_n18750), .B(new_n18705), .C(new_n18805), .Y(new_n18806));
  INVx1_ASAP7_75t_L         g18550(.A(new_n18806), .Y(new_n18807));
  AOI211xp5_ASAP7_75t_L     g18551(.A1(new_n18708), .A2(new_n18750), .B(new_n18705), .C(new_n18805), .Y(new_n18808));
  OAI21xp33_ASAP7_75t_L     g18552(.A1(new_n18808), .A2(new_n18807), .B(new_n18749), .Y(new_n18809));
  OR3x1_ASAP7_75t_L         g18553(.A(new_n18807), .B(new_n18749), .C(new_n18808), .Y(new_n18810));
  AND2x2_ASAP7_75t_L        g18554(.A(new_n18809), .B(new_n18810), .Y(new_n18811));
  NAND3xp33_ASAP7_75t_L     g18555(.A(new_n18811), .B(new_n18716), .C(new_n18712), .Y(new_n18812));
  INVx1_ASAP7_75t_L         g18556(.A(new_n18811), .Y(new_n18813));
  A2O1A1Ixp33_ASAP7_75t_L   g18557(.A1(new_n18715), .A2(new_n18710), .B(new_n18711), .C(new_n18813), .Y(new_n18814));
  NAND2xp33_ASAP7_75t_L     g18558(.A(new_n18812), .B(new_n18814), .Y(new_n18815));
  AOI22xp33_ASAP7_75t_L     g18559(.A1(new_n6376), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n6648), .Y(new_n18816));
  A2O1A1Ixp33_ASAP7_75t_L   g18560(.A1(new_n11470), .A2(new_n11473), .B(new_n6636), .C(new_n18816), .Y(new_n18817));
  AOI21xp33_ASAP7_75t_L     g18561(.A1(new_n6380), .A2(\b[62] ), .B(new_n18817), .Y(new_n18818));
  NAND2xp33_ASAP7_75t_L     g18562(.A(\a[47] ), .B(new_n18818), .Y(new_n18819));
  A2O1A1Ixp33_ASAP7_75t_L   g18563(.A1(\b[62] ), .A2(new_n6380), .B(new_n18817), .C(new_n6371), .Y(new_n18820));
  NAND2xp33_ASAP7_75t_L     g18564(.A(new_n18820), .B(new_n18819), .Y(new_n18821));
  XNOR2x2_ASAP7_75t_L       g18565(.A(new_n18821), .B(new_n18815), .Y(new_n18822));
  AO21x2_ASAP7_75t_L        g18566(.A1(new_n18723), .A2(new_n18724), .B(new_n18822), .Y(new_n18823));
  NAND3xp33_ASAP7_75t_L     g18567(.A(new_n18822), .B(new_n18724), .C(new_n18723), .Y(new_n18824));
  AND2x2_ASAP7_75t_L        g18568(.A(new_n18824), .B(new_n18823), .Y(new_n18825));
  INVx1_ASAP7_75t_L         g18569(.A(new_n18825), .Y(new_n18826));
  A2O1A1O1Ixp25_ASAP7_75t_L g18570(.A1(new_n18725), .A2(new_n18724), .B(new_n18734), .C(new_n18733), .D(new_n18826), .Y(new_n18827));
  INVx1_ASAP7_75t_L         g18571(.A(new_n18827), .Y(new_n18828));
  A2O1A1Ixp33_ASAP7_75t_L   g18572(.A1(new_n18725), .A2(new_n18724), .B(new_n18734), .C(new_n18733), .Y(new_n18829));
  AO21x2_ASAP7_75t_L        g18573(.A1(new_n18824), .A2(new_n18823), .B(new_n18829), .Y(new_n18830));
  AND2x2_ASAP7_75t_L        g18574(.A(new_n18830), .B(new_n18828), .Y(new_n18831));
  INVx1_ASAP7_75t_L         g18575(.A(new_n18831), .Y(new_n18832));
  A2O1A1O1Ixp25_ASAP7_75t_L g18576(.A1(new_n18649), .A2(new_n18651), .B(new_n18744), .C(new_n18739), .D(new_n18832), .Y(new_n18833));
  A2O1A1Ixp33_ASAP7_75t_L   g18577(.A1(new_n18651), .A2(new_n18649), .B(new_n18744), .C(new_n18739), .Y(new_n18834));
  NOR2xp33_ASAP7_75t_L      g18578(.A(new_n18831), .B(new_n18834), .Y(new_n18835));
  NOR2xp33_ASAP7_75t_L      g18579(.A(new_n18833), .B(new_n18835), .Y(\f[108] ));
  NAND2xp33_ASAP7_75t_L     g18580(.A(new_n18810), .B(new_n18812), .Y(new_n18837));
  OAI22xp33_ASAP7_75t_L     g18581(.A1(new_n11500), .A2(new_n6636), .B1(new_n11172), .B2(new_n6638), .Y(new_n18838));
  AOI21xp33_ASAP7_75t_L     g18582(.A1(new_n6380), .A2(\b[63] ), .B(new_n18838), .Y(new_n18839));
  NAND2xp33_ASAP7_75t_L     g18583(.A(\a[47] ), .B(new_n18839), .Y(new_n18840));
  A2O1A1Ixp33_ASAP7_75t_L   g18584(.A1(\b[63] ), .A2(new_n6380), .B(new_n18838), .C(new_n6371), .Y(new_n18841));
  NAND2xp33_ASAP7_75t_L     g18585(.A(new_n18841), .B(new_n18840), .Y(new_n18842));
  XNOR2x2_ASAP7_75t_L       g18586(.A(new_n18842), .B(new_n18837), .Y(new_n18843));
  AOI22xp33_ASAP7_75t_L     g18587(.A1(new_n7111), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n7391), .Y(new_n18844));
  OAI221xp5_ASAP7_75t_L     g18588(.A1(new_n8558), .A2(new_n10250), .B1(new_n8237), .B2(new_n10855), .C(new_n18844), .Y(new_n18845));
  XNOR2x2_ASAP7_75t_L       g18589(.A(\a[50] ), .B(new_n18845), .Y(new_n18846));
  AOI22xp33_ASAP7_75t_L     g18590(.A1(new_n7960), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n8537), .Y(new_n18847));
  OAI221xp5_ASAP7_75t_L     g18591(.A1(new_n8817), .A2(new_n9620), .B1(new_n7957), .B2(new_n9925), .C(new_n18847), .Y(new_n18848));
  XNOR2x2_ASAP7_75t_L       g18592(.A(\a[53] ), .B(new_n18848), .Y(new_n18849));
  INVx1_ASAP7_75t_L         g18593(.A(new_n18849), .Y(new_n18850));
  AOI22xp33_ASAP7_75t_L     g18594(.A1(new_n9700), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n10027), .Y(new_n18851));
  OAI221xp5_ASAP7_75t_L     g18595(.A1(new_n10024), .A2(new_n7616), .B1(new_n9696), .B2(new_n7906), .C(new_n18851), .Y(new_n18852));
  XNOR2x2_ASAP7_75t_L       g18596(.A(\a[59] ), .B(new_n18852), .Y(new_n18853));
  INVx1_ASAP7_75t_L         g18597(.A(new_n18853), .Y(new_n18854));
  A2O1A1Ixp33_ASAP7_75t_L   g18598(.A1(new_n18686), .A2(new_n18685), .B(new_n18673), .C(new_n18776), .Y(new_n18855));
  NOR2xp33_ASAP7_75t_L      g18599(.A(new_n6321), .B(new_n11535), .Y(new_n18856));
  A2O1A1O1Ixp25_ASAP7_75t_L g18600(.A1(new_n11533), .A2(\b[43] ), .B(new_n18572), .C(new_n18771), .D(new_n18769), .Y(new_n18857));
  A2O1A1Ixp33_ASAP7_75t_L   g18601(.A1(new_n11533), .A2(\b[46] ), .B(new_n18856), .C(new_n18857), .Y(new_n18858));
  O2A1O1Ixp33_ASAP7_75t_L   g18602(.A1(new_n11247), .A2(new_n11249), .B(\b[46] ), .C(new_n18856), .Y(new_n18859));
  INVx1_ASAP7_75t_L         g18603(.A(new_n18859), .Y(new_n18860));
  O2A1O1Ixp33_ASAP7_75t_L   g18604(.A1(new_n18573), .A2(new_n18772), .B(new_n18768), .C(new_n18860), .Y(new_n18861));
  INVx1_ASAP7_75t_L         g18605(.A(new_n18861), .Y(new_n18862));
  NAND2xp33_ASAP7_75t_L     g18606(.A(new_n18858), .B(new_n18862), .Y(new_n18863));
  NAND2xp33_ASAP7_75t_L     g18607(.A(\b[47] ), .B(new_n10939), .Y(new_n18864));
  OAI221xp5_ASAP7_75t_L     g18608(.A1(new_n10630), .A2(new_n7317), .B1(new_n10629), .B2(new_n7323), .C(new_n18864), .Y(new_n18865));
  AOI21xp33_ASAP7_75t_L     g18609(.A1(new_n10632), .A2(\b[48] ), .B(new_n18865), .Y(new_n18866));
  NAND2xp33_ASAP7_75t_L     g18610(.A(\a[62] ), .B(new_n18866), .Y(new_n18867));
  A2O1A1Ixp33_ASAP7_75t_L   g18611(.A1(\b[48] ), .A2(new_n10632), .B(new_n18865), .C(new_n10622), .Y(new_n18868));
  AND3x1_ASAP7_75t_L        g18612(.A(new_n18867), .B(new_n18868), .C(new_n18863), .Y(new_n18869));
  AND2x2_ASAP7_75t_L        g18613(.A(new_n18868), .B(new_n18867), .Y(new_n18870));
  NOR2xp33_ASAP7_75t_L      g18614(.A(new_n18863), .B(new_n18870), .Y(new_n18871));
  NOR2xp33_ASAP7_75t_L      g18615(.A(new_n18869), .B(new_n18871), .Y(new_n18872));
  INVx1_ASAP7_75t_L         g18616(.A(new_n18872), .Y(new_n18873));
  O2A1O1Ixp33_ASAP7_75t_L   g18617(.A1(new_n18765), .A2(new_n18778), .B(new_n18855), .C(new_n18873), .Y(new_n18874));
  INVx1_ASAP7_75t_L         g18618(.A(new_n18874), .Y(new_n18875));
  O2A1O1Ixp33_ASAP7_75t_L   g18619(.A1(new_n18673), .A2(new_n18684), .B(new_n18776), .C(new_n18779), .Y(new_n18876));
  NAND2xp33_ASAP7_75t_L     g18620(.A(new_n18873), .B(new_n18876), .Y(new_n18877));
  NAND3xp33_ASAP7_75t_L     g18621(.A(new_n18875), .B(new_n18854), .C(new_n18877), .Y(new_n18878));
  AO21x2_ASAP7_75t_L        g18622(.A1(new_n18877), .A2(new_n18875), .B(new_n18854), .Y(new_n18879));
  AND2x2_ASAP7_75t_L        g18623(.A(new_n18878), .B(new_n18879), .Y(new_n18880));
  A2O1A1Ixp33_ASAP7_75t_L   g18624(.A1(new_n18782), .A2(new_n18762), .B(new_n18788), .C(new_n18880), .Y(new_n18881));
  A2O1A1Ixp33_ASAP7_75t_L   g18625(.A1(new_n18696), .A2(new_n18691), .B(new_n18783), .C(new_n18784), .Y(new_n18882));
  NOR2xp33_ASAP7_75t_L      g18626(.A(new_n18882), .B(new_n18880), .Y(new_n18883));
  INVx1_ASAP7_75t_L         g18627(.A(new_n18883), .Y(new_n18884));
  AOI22xp33_ASAP7_75t_L     g18628(.A1(new_n8831), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n9115), .Y(new_n18885));
  OAI221xp5_ASAP7_75t_L     g18629(.A1(new_n10343), .A2(new_n8458), .B1(new_n10016), .B2(new_n8768), .C(new_n18885), .Y(new_n18886));
  XNOR2x2_ASAP7_75t_L       g18630(.A(\a[56] ), .B(new_n18886), .Y(new_n18887));
  NAND3xp33_ASAP7_75t_L     g18631(.A(new_n18881), .B(new_n18884), .C(new_n18887), .Y(new_n18888));
  INVx1_ASAP7_75t_L         g18632(.A(new_n18888), .Y(new_n18889));
  AOI21xp33_ASAP7_75t_L     g18633(.A1(new_n18881), .A2(new_n18884), .B(new_n18887), .Y(new_n18890));
  NOR2xp33_ASAP7_75t_L      g18634(.A(new_n18890), .B(new_n18889), .Y(new_n18891));
  A2O1A1O1Ixp25_ASAP7_75t_L g18635(.A1(new_n18702), .A2(new_n18700), .B(new_n18798), .C(new_n18795), .D(new_n18891), .Y(new_n18892));
  INVx1_ASAP7_75t_L         g18636(.A(new_n18892), .Y(new_n18893));
  NAND3xp33_ASAP7_75t_L     g18637(.A(new_n18797), .B(new_n18795), .C(new_n18891), .Y(new_n18894));
  AO21x2_ASAP7_75t_L        g18638(.A1(new_n18894), .A2(new_n18893), .B(new_n18850), .Y(new_n18895));
  NAND3xp33_ASAP7_75t_L     g18639(.A(new_n18893), .B(new_n18850), .C(new_n18894), .Y(new_n18896));
  AND2x2_ASAP7_75t_L        g18640(.A(new_n18896), .B(new_n18895), .Y(new_n18897));
  INVx1_ASAP7_75t_L         g18641(.A(new_n18897), .Y(new_n18898));
  O2A1O1Ixp33_ASAP7_75t_L   g18642(.A1(new_n18753), .A2(new_n18801), .B(new_n18806), .C(new_n18898), .Y(new_n18899));
  INVx1_ASAP7_75t_L         g18643(.A(new_n18804), .Y(new_n18900));
  A2O1A1O1Ixp25_ASAP7_75t_L g18644(.A1(new_n18750), .A2(new_n18708), .B(new_n18705), .C(new_n18802), .D(new_n18900), .Y(new_n18901));
  NAND2xp33_ASAP7_75t_L     g18645(.A(new_n18901), .B(new_n18898), .Y(new_n18902));
  INVx1_ASAP7_75t_L         g18646(.A(new_n18902), .Y(new_n18903));
  NOR2xp33_ASAP7_75t_L      g18647(.A(new_n18903), .B(new_n18899), .Y(new_n18904));
  XNOR2x2_ASAP7_75t_L       g18648(.A(new_n18846), .B(new_n18904), .Y(new_n18905));
  XNOR2x2_ASAP7_75t_L       g18649(.A(new_n18905), .B(new_n18843), .Y(new_n18906));
  A2O1A1Ixp33_ASAP7_75t_L   g18650(.A1(new_n18819), .A2(new_n18820), .B(new_n18815), .C(new_n18824), .Y(new_n18907));
  NOR2xp33_ASAP7_75t_L      g18651(.A(new_n18906), .B(new_n18907), .Y(new_n18908));
  NAND2xp33_ASAP7_75t_L     g18652(.A(new_n18906), .B(new_n18907), .Y(new_n18909));
  INVx1_ASAP7_75t_L         g18653(.A(new_n18909), .Y(new_n18910));
  NOR2xp33_ASAP7_75t_L      g18654(.A(new_n18908), .B(new_n18910), .Y(new_n18911));
  A2O1A1Ixp33_ASAP7_75t_L   g18655(.A1(new_n18742), .A2(new_n18739), .B(new_n18832), .C(new_n18828), .Y(new_n18912));
  XOR2x2_ASAP7_75t_L        g18656(.A(new_n18911), .B(new_n18912), .Y(\f[109] ));
  AOI22xp33_ASAP7_75t_L     g18657(.A1(new_n7111), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n7391), .Y(new_n18914));
  OAI221xp5_ASAP7_75t_L     g18658(.A1(new_n8558), .A2(new_n10847), .B1(new_n8237), .B2(new_n12047), .C(new_n18914), .Y(new_n18915));
  XNOR2x2_ASAP7_75t_L       g18659(.A(\a[50] ), .B(new_n18915), .Y(new_n18916));
  AOI22xp33_ASAP7_75t_L     g18660(.A1(new_n8831), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n9115), .Y(new_n18917));
  OAI221xp5_ASAP7_75t_L     g18661(.A1(new_n10343), .A2(new_n8762), .B1(new_n10016), .B2(new_n9331), .C(new_n18917), .Y(new_n18918));
  XNOR2x2_ASAP7_75t_L       g18662(.A(\a[56] ), .B(new_n18918), .Y(new_n18919));
  INVx1_ASAP7_75t_L         g18663(.A(new_n18919), .Y(new_n18920));
  AOI22xp33_ASAP7_75t_L     g18664(.A1(new_n9700), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n10027), .Y(new_n18921));
  OAI221xp5_ASAP7_75t_L     g18665(.A1(new_n10024), .A2(new_n7900), .B1(new_n9696), .B2(new_n8174), .C(new_n18921), .Y(new_n18922));
  XNOR2x2_ASAP7_75t_L       g18666(.A(\a[59] ), .B(new_n18922), .Y(new_n18923));
  INVx1_ASAP7_75t_L         g18667(.A(new_n18923), .Y(new_n18924));
  AOI22xp33_ASAP7_75t_L     g18668(.A1(\b[48] ), .A2(new_n10939), .B1(\b[50] ), .B2(new_n10938), .Y(new_n18925));
  OAI221xp5_ASAP7_75t_L     g18669(.A1(new_n10937), .A2(new_n7317), .B1(new_n10629), .B2(new_n7602), .C(new_n18925), .Y(new_n18926));
  XNOR2x2_ASAP7_75t_L       g18670(.A(\a[62] ), .B(new_n18926), .Y(new_n18927));
  O2A1O1Ixp33_ASAP7_75t_L   g18671(.A1(new_n5805), .A2(new_n11253), .B(new_n18674), .C(new_n18772), .Y(new_n18928));
  O2A1O1Ixp33_ASAP7_75t_L   g18672(.A1(new_n18769), .A2(new_n18928), .B(new_n18859), .C(new_n18871), .Y(new_n18929));
  NOR2xp33_ASAP7_75t_L      g18673(.A(new_n6568), .B(new_n11535), .Y(new_n18930));
  A2O1A1Ixp33_ASAP7_75t_L   g18674(.A1(\b[47] ), .A2(new_n11533), .B(new_n18930), .C(new_n18859), .Y(new_n18931));
  O2A1O1Ixp33_ASAP7_75t_L   g18675(.A1(new_n11247), .A2(new_n11249), .B(\b[47] ), .C(new_n18930), .Y(new_n18932));
  A2O1A1Ixp33_ASAP7_75t_L   g18676(.A1(new_n11533), .A2(\b[46] ), .B(new_n18856), .C(new_n18932), .Y(new_n18933));
  AND2x2_ASAP7_75t_L        g18677(.A(new_n18931), .B(new_n18933), .Y(new_n18934));
  AND2x2_ASAP7_75t_L        g18678(.A(new_n18934), .B(new_n18929), .Y(new_n18935));
  A2O1A1O1Ixp25_ASAP7_75t_L g18679(.A1(new_n18868), .A2(new_n18867), .B(new_n18863), .C(new_n18862), .D(new_n18934), .Y(new_n18936));
  NOR2xp33_ASAP7_75t_L      g18680(.A(new_n18936), .B(new_n18935), .Y(new_n18937));
  NOR2xp33_ASAP7_75t_L      g18681(.A(new_n18927), .B(new_n18937), .Y(new_n18938));
  INVx1_ASAP7_75t_L         g18682(.A(new_n18938), .Y(new_n18939));
  NAND2xp33_ASAP7_75t_L     g18683(.A(new_n18927), .B(new_n18937), .Y(new_n18940));
  NAND3xp33_ASAP7_75t_L     g18684(.A(new_n18939), .B(new_n18924), .C(new_n18940), .Y(new_n18941));
  INVx1_ASAP7_75t_L         g18685(.A(new_n18941), .Y(new_n18942));
  AOI21xp33_ASAP7_75t_L     g18686(.A1(new_n18939), .A2(new_n18940), .B(new_n18924), .Y(new_n18943));
  NOR2xp33_ASAP7_75t_L      g18687(.A(new_n18943), .B(new_n18942), .Y(new_n18944));
  INVx1_ASAP7_75t_L         g18688(.A(new_n18944), .Y(new_n18945));
  O2A1O1Ixp33_ASAP7_75t_L   g18689(.A1(new_n18876), .A2(new_n18873), .B(new_n18878), .C(new_n18945), .Y(new_n18946));
  INVx1_ASAP7_75t_L         g18690(.A(new_n18946), .Y(new_n18947));
  NAND3xp33_ASAP7_75t_L     g18691(.A(new_n18945), .B(new_n18878), .C(new_n18875), .Y(new_n18948));
  AND2x2_ASAP7_75t_L        g18692(.A(new_n18948), .B(new_n18947), .Y(new_n18949));
  NAND2xp33_ASAP7_75t_L     g18693(.A(new_n18920), .B(new_n18949), .Y(new_n18950));
  INVx1_ASAP7_75t_L         g18694(.A(new_n18950), .Y(new_n18951));
  NOR2xp33_ASAP7_75t_L      g18695(.A(new_n18920), .B(new_n18949), .Y(new_n18952));
  NOR2xp33_ASAP7_75t_L      g18696(.A(new_n18952), .B(new_n18951), .Y(new_n18953));
  NAND3xp33_ASAP7_75t_L     g18697(.A(new_n18953), .B(new_n18888), .C(new_n18884), .Y(new_n18954));
  O2A1O1Ixp33_ASAP7_75t_L   g18698(.A1(new_n18882), .A2(new_n18880), .B(new_n18888), .C(new_n18953), .Y(new_n18955));
  INVx1_ASAP7_75t_L         g18699(.A(new_n18955), .Y(new_n18956));
  AOI22xp33_ASAP7_75t_L     g18700(.A1(new_n7960), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n8537), .Y(new_n18957));
  OAI221xp5_ASAP7_75t_L     g18701(.A1(new_n8817), .A2(new_n9920), .B1(new_n7957), .B2(new_n11152), .C(new_n18957), .Y(new_n18958));
  XNOR2x2_ASAP7_75t_L       g18702(.A(\a[53] ), .B(new_n18958), .Y(new_n18959));
  NAND3xp33_ASAP7_75t_L     g18703(.A(new_n18956), .B(new_n18954), .C(new_n18959), .Y(new_n18960));
  AO21x2_ASAP7_75t_L        g18704(.A1(new_n18954), .A2(new_n18956), .B(new_n18959), .Y(new_n18961));
  AND2x2_ASAP7_75t_L        g18705(.A(new_n18960), .B(new_n18961), .Y(new_n18962));
  INVx1_ASAP7_75t_L         g18706(.A(new_n18962), .Y(new_n18963));
  A2O1A1Ixp33_ASAP7_75t_L   g18707(.A1(new_n18894), .A2(new_n18850), .B(new_n18892), .C(new_n18963), .Y(new_n18964));
  NAND3xp33_ASAP7_75t_L     g18708(.A(new_n18962), .B(new_n18896), .C(new_n18893), .Y(new_n18965));
  NAND3xp33_ASAP7_75t_L     g18709(.A(new_n18964), .B(new_n18916), .C(new_n18965), .Y(new_n18966));
  AO21x2_ASAP7_75t_L        g18710(.A1(new_n18965), .A2(new_n18964), .B(new_n18916), .Y(new_n18967));
  NAND2xp33_ASAP7_75t_L     g18711(.A(new_n18966), .B(new_n18967), .Y(new_n18968));
  INVx1_ASAP7_75t_L         g18712(.A(new_n18846), .Y(new_n18969));
  A2O1A1O1Ixp25_ASAP7_75t_L g18713(.A1(new_n6373), .A2(new_n12061), .B(new_n6648), .C(\b[63] ), .D(new_n6371), .Y(new_n18970));
  A2O1A1Ixp33_ASAP7_75t_L   g18714(.A1(new_n12061), .A2(new_n6373), .B(new_n6648), .C(\b[63] ), .Y(new_n18971));
  NOR2xp33_ASAP7_75t_L      g18715(.A(\a[47] ), .B(new_n18971), .Y(new_n18972));
  OAI221xp5_ASAP7_75t_L     g18716(.A1(new_n18972), .A2(new_n18970), .B1(new_n18969), .B2(new_n18899), .C(new_n18902), .Y(new_n18973));
  NOR2xp33_ASAP7_75t_L      g18717(.A(new_n18970), .B(new_n18972), .Y(new_n18974));
  A2O1A1Ixp33_ASAP7_75t_L   g18718(.A1(new_n18904), .A2(new_n18846), .B(new_n18903), .C(new_n18974), .Y(new_n18975));
  NAND2xp33_ASAP7_75t_L     g18719(.A(new_n18973), .B(new_n18975), .Y(new_n18976));
  NAND2xp33_ASAP7_75t_L     g18720(.A(new_n18976), .B(new_n18968), .Y(new_n18977));
  NOR2xp33_ASAP7_75t_L      g18721(.A(new_n18976), .B(new_n18968), .Y(new_n18978));
  INVx1_ASAP7_75t_L         g18722(.A(new_n18978), .Y(new_n18979));
  NAND2xp33_ASAP7_75t_L     g18723(.A(new_n18977), .B(new_n18979), .Y(new_n18980));
  MAJx2_ASAP7_75t_L         g18724(.A(new_n18837), .B(new_n18842), .C(new_n18905), .Y(new_n18981));
  NOR2xp33_ASAP7_75t_L      g18725(.A(new_n18981), .B(new_n18980), .Y(new_n18982));
  NAND2xp33_ASAP7_75t_L     g18726(.A(new_n18981), .B(new_n18980), .Y(new_n18983));
  INVx1_ASAP7_75t_L         g18727(.A(new_n18983), .Y(new_n18984));
  NOR2xp33_ASAP7_75t_L      g18728(.A(new_n18982), .B(new_n18984), .Y(new_n18985));
  A2O1A1Ixp33_ASAP7_75t_L   g18729(.A1(new_n18912), .A2(new_n18911), .B(new_n18910), .C(new_n18985), .Y(new_n18986));
  INVx1_ASAP7_75t_L         g18730(.A(new_n18986), .Y(new_n18987));
  INVx1_ASAP7_75t_L         g18731(.A(new_n18833), .Y(new_n18988));
  A2O1A1Ixp33_ASAP7_75t_L   g18732(.A1(new_n18988), .A2(new_n18828), .B(new_n18908), .C(new_n18909), .Y(new_n18989));
  NOR2xp33_ASAP7_75t_L      g18733(.A(new_n18985), .B(new_n18989), .Y(new_n18990));
  NOR2xp33_ASAP7_75t_L      g18734(.A(new_n18987), .B(new_n18990), .Y(\f[110] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18735(.A1(new_n18834), .A2(new_n18831), .B(new_n18827), .C(new_n18911), .Y(new_n18992));
  AOI22xp33_ASAP7_75t_L     g18736(.A1(new_n7960), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n8537), .Y(new_n18993));
  OAI221xp5_ASAP7_75t_L     g18737(.A1(new_n8817), .A2(new_n9947), .B1(new_n7957), .B2(new_n11446), .C(new_n18993), .Y(new_n18994));
  XNOR2x2_ASAP7_75t_L       g18738(.A(\a[53] ), .B(new_n18994), .Y(new_n18995));
  AOI22xp33_ASAP7_75t_L     g18739(.A1(new_n8831), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n9115), .Y(new_n18996));
  OAI221xp5_ASAP7_75t_L     g18740(.A1(new_n10343), .A2(new_n9323), .B1(new_n10016), .B2(new_n9627), .C(new_n18996), .Y(new_n18997));
  XNOR2x2_ASAP7_75t_L       g18741(.A(\a[56] ), .B(new_n18997), .Y(new_n18998));
  INVx1_ASAP7_75t_L         g18742(.A(new_n18998), .Y(new_n18999));
  AOI22xp33_ASAP7_75t_L     g18743(.A1(\b[49] ), .A2(new_n10939), .B1(\b[51] ), .B2(new_n10938), .Y(new_n19000));
  OAI221xp5_ASAP7_75t_L     g18744(.A1(new_n10937), .A2(new_n7593), .B1(new_n10629), .B2(new_n7623), .C(new_n19000), .Y(new_n19001));
  XNOR2x2_ASAP7_75t_L       g18745(.A(\a[62] ), .B(new_n19001), .Y(new_n19002));
  NOR2xp33_ASAP7_75t_L      g18746(.A(new_n6812), .B(new_n11535), .Y(new_n19003));
  INVx1_ASAP7_75t_L         g18747(.A(new_n19003), .Y(new_n19004));
  A2O1A1Ixp33_ASAP7_75t_L   g18748(.A1(new_n11533), .A2(\b[47] ), .B(new_n18930), .C(\a[47] ), .Y(new_n19005));
  INVx1_ASAP7_75t_L         g18749(.A(new_n18932), .Y(new_n19006));
  NOR2xp33_ASAP7_75t_L      g18750(.A(\a[47] ), .B(new_n19006), .Y(new_n19007));
  INVx1_ASAP7_75t_L         g18751(.A(new_n19007), .Y(new_n19008));
  AND2x2_ASAP7_75t_L        g18752(.A(new_n19005), .B(new_n19008), .Y(new_n19009));
  O2A1O1Ixp33_ASAP7_75t_L   g18753(.A1(new_n6830), .A2(new_n11253), .B(new_n19004), .C(new_n19009), .Y(new_n19010));
  O2A1O1Ixp33_ASAP7_75t_L   g18754(.A1(new_n11247), .A2(new_n11249), .B(\b[48] ), .C(new_n19003), .Y(new_n19011));
  AND3x1_ASAP7_75t_L        g18755(.A(new_n19008), .B(new_n19005), .C(new_n19011), .Y(new_n19012));
  NOR2xp33_ASAP7_75t_L      g18756(.A(new_n19012), .B(new_n19010), .Y(new_n19013));
  INVx1_ASAP7_75t_L         g18757(.A(new_n19013), .Y(new_n19014));
  XNOR2x2_ASAP7_75t_L       g18758(.A(new_n19014), .B(new_n19002), .Y(new_n19015));
  A2O1A1O1Ixp25_ASAP7_75t_L g18759(.A1(\b[47] ), .A2(new_n11533), .B(new_n18930), .C(new_n18859), .D(new_n18929), .Y(new_n19016));
  A2O1A1Ixp33_ASAP7_75t_L   g18760(.A1(new_n18860), .A2(new_n18932), .B(new_n19016), .C(new_n19015), .Y(new_n19017));
  INVx1_ASAP7_75t_L         g18761(.A(new_n19015), .Y(new_n19018));
  A2O1A1O1Ixp25_ASAP7_75t_L g18762(.A1(new_n11533), .A2(\b[46] ), .B(new_n18856), .C(new_n18932), .D(new_n19016), .Y(new_n19019));
  NAND2xp33_ASAP7_75t_L     g18763(.A(new_n19018), .B(new_n19019), .Y(new_n19020));
  AND2x2_ASAP7_75t_L        g18764(.A(new_n19017), .B(new_n19020), .Y(new_n19021));
  AOI22xp33_ASAP7_75t_L     g18765(.A1(new_n9700), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n10027), .Y(new_n19022));
  OAI221xp5_ASAP7_75t_L     g18766(.A1(new_n10024), .A2(new_n8165), .B1(new_n9696), .B2(new_n8465), .C(new_n19022), .Y(new_n19023));
  XNOR2x2_ASAP7_75t_L       g18767(.A(\a[59] ), .B(new_n19023), .Y(new_n19024));
  NAND2xp33_ASAP7_75t_L     g18768(.A(new_n19024), .B(new_n19021), .Y(new_n19025));
  NOR2xp33_ASAP7_75t_L      g18769(.A(new_n19024), .B(new_n19021), .Y(new_n19026));
  INVx1_ASAP7_75t_L         g18770(.A(new_n19026), .Y(new_n19027));
  AND2x2_ASAP7_75t_L        g18771(.A(new_n19025), .B(new_n19027), .Y(new_n19028));
  INVx1_ASAP7_75t_L         g18772(.A(new_n19028), .Y(new_n19029));
  O2A1O1Ixp33_ASAP7_75t_L   g18773(.A1(new_n18927), .A2(new_n18937), .B(new_n18941), .C(new_n19029), .Y(new_n19030));
  INVx1_ASAP7_75t_L         g18774(.A(new_n19030), .Y(new_n19031));
  NAND3xp33_ASAP7_75t_L     g18775(.A(new_n19029), .B(new_n18941), .C(new_n18939), .Y(new_n19032));
  AO21x2_ASAP7_75t_L        g18776(.A1(new_n19032), .A2(new_n19031), .B(new_n18999), .Y(new_n19033));
  AND2x2_ASAP7_75t_L        g18777(.A(new_n19032), .B(new_n19031), .Y(new_n19034));
  NAND2xp33_ASAP7_75t_L     g18778(.A(new_n18999), .B(new_n19034), .Y(new_n19035));
  AND2x2_ASAP7_75t_L        g18779(.A(new_n19033), .B(new_n19035), .Y(new_n19036));
  A2O1A1Ixp33_ASAP7_75t_L   g18780(.A1(new_n18948), .A2(new_n18920), .B(new_n18946), .C(new_n19036), .Y(new_n19037));
  INVx1_ASAP7_75t_L         g18781(.A(new_n19037), .Y(new_n19038));
  A2O1A1Ixp33_ASAP7_75t_L   g18782(.A1(new_n18878), .A2(new_n18875), .B(new_n18945), .C(new_n18950), .Y(new_n19039));
  NOR2xp33_ASAP7_75t_L      g18783(.A(new_n19039), .B(new_n19036), .Y(new_n19040));
  OAI21xp33_ASAP7_75t_L     g18784(.A1(new_n19040), .A2(new_n19038), .B(new_n18995), .Y(new_n19041));
  INVx1_ASAP7_75t_L         g18785(.A(new_n18995), .Y(new_n19042));
  NOR2xp33_ASAP7_75t_L      g18786(.A(new_n19040), .B(new_n19038), .Y(new_n19043));
  NAND2xp33_ASAP7_75t_L     g18787(.A(new_n19042), .B(new_n19043), .Y(new_n19044));
  AND2x2_ASAP7_75t_L        g18788(.A(new_n19041), .B(new_n19044), .Y(new_n19045));
  INVx1_ASAP7_75t_L         g18789(.A(new_n19045), .Y(new_n19046));
  A2O1A1Ixp33_ASAP7_75t_L   g18790(.A1(new_n18888), .A2(new_n18884), .B(new_n18953), .C(new_n18960), .Y(new_n19047));
  NOR2xp33_ASAP7_75t_L      g18791(.A(new_n19047), .B(new_n19046), .Y(new_n19048));
  INVx1_ASAP7_75t_L         g18792(.A(new_n19048), .Y(new_n19049));
  A2O1A1Ixp33_ASAP7_75t_L   g18793(.A1(new_n18959), .A2(new_n18954), .B(new_n18955), .C(new_n19046), .Y(new_n19050));
  NAND2xp33_ASAP7_75t_L     g18794(.A(new_n19050), .B(new_n19049), .Y(new_n19051));
  AOI22xp33_ASAP7_75t_L     g18795(.A1(new_n7111), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n7391), .Y(new_n19052));
  A2O1A1Ixp33_ASAP7_75t_L   g18796(.A1(new_n11470), .A2(new_n11473), .B(new_n8237), .C(new_n19052), .Y(new_n19053));
  AOI21xp33_ASAP7_75t_L     g18797(.A1(new_n7115), .A2(\b[62] ), .B(new_n19053), .Y(new_n19054));
  NAND2xp33_ASAP7_75t_L     g18798(.A(\a[50] ), .B(new_n19054), .Y(new_n19055));
  A2O1A1Ixp33_ASAP7_75t_L   g18799(.A1(\b[62] ), .A2(new_n7115), .B(new_n19053), .C(new_n7106), .Y(new_n19056));
  NAND2xp33_ASAP7_75t_L     g18800(.A(new_n19056), .B(new_n19055), .Y(new_n19057));
  XNOR2x2_ASAP7_75t_L       g18801(.A(new_n19057), .B(new_n19051), .Y(new_n19058));
  AO21x2_ASAP7_75t_L        g18802(.A1(new_n18965), .A2(new_n18966), .B(new_n19058), .Y(new_n19059));
  NAND3xp33_ASAP7_75t_L     g18803(.A(new_n19058), .B(new_n18966), .C(new_n18965), .Y(new_n19060));
  AND2x2_ASAP7_75t_L        g18804(.A(new_n19060), .B(new_n19059), .Y(new_n19061));
  O2A1O1Ixp33_ASAP7_75t_L   g18805(.A1(new_n18968), .A2(new_n18976), .B(new_n18975), .C(new_n19061), .Y(new_n19062));
  INVx1_ASAP7_75t_L         g18806(.A(new_n19061), .Y(new_n19063));
  A2O1A1O1Ixp25_ASAP7_75t_L g18807(.A1(new_n18846), .A2(new_n18904), .B(new_n18903), .C(new_n18974), .D(new_n18978), .Y(new_n19064));
  INVx1_ASAP7_75t_L         g18808(.A(new_n19064), .Y(new_n19065));
  NOR2xp33_ASAP7_75t_L      g18809(.A(new_n19065), .B(new_n19063), .Y(new_n19066));
  NOR2xp33_ASAP7_75t_L      g18810(.A(new_n19062), .B(new_n19066), .Y(new_n19067));
  INVx1_ASAP7_75t_L         g18811(.A(new_n19067), .Y(new_n19068));
  A2O1A1O1Ixp25_ASAP7_75t_L g18812(.A1(new_n18909), .A2(new_n18992), .B(new_n18982), .C(new_n18983), .D(new_n19068), .Y(new_n19069));
  A2O1A1Ixp33_ASAP7_75t_L   g18813(.A1(new_n18992), .A2(new_n18909), .B(new_n18982), .C(new_n18983), .Y(new_n19070));
  NOR2xp33_ASAP7_75t_L      g18814(.A(new_n19067), .B(new_n19070), .Y(new_n19071));
  NOR2xp33_ASAP7_75t_L      g18815(.A(new_n19069), .B(new_n19071), .Y(\f[111] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18816(.A1(new_n19055), .A2(new_n19056), .B(new_n19051), .C(new_n19060), .Y(new_n19073));
  AOI22xp33_ASAP7_75t_L     g18817(.A1(new_n7960), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n8537), .Y(new_n19074));
  OAI221xp5_ASAP7_75t_L     g18818(.A1(new_n8817), .A2(new_n10250), .B1(new_n7957), .B2(new_n10855), .C(new_n19074), .Y(new_n19075));
  NOR2xp33_ASAP7_75t_L      g18819(.A(new_n7954), .B(new_n19075), .Y(new_n19076));
  AND2x2_ASAP7_75t_L        g18820(.A(new_n7954), .B(new_n19075), .Y(new_n19077));
  INVx1_ASAP7_75t_L         g18821(.A(new_n19035), .Y(new_n19078));
  AOI22xp33_ASAP7_75t_L     g18822(.A1(new_n8831), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n9115), .Y(new_n19079));
  OAI221xp5_ASAP7_75t_L     g18823(.A1(new_n10343), .A2(new_n9620), .B1(new_n10016), .B2(new_n9925), .C(new_n19079), .Y(new_n19080));
  XNOR2x2_ASAP7_75t_L       g18824(.A(\a[56] ), .B(new_n19080), .Y(new_n19081));
  AOI22xp33_ASAP7_75t_L     g18825(.A1(new_n9700), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n10027), .Y(new_n19082));
  OAI221xp5_ASAP7_75t_L     g18826(.A1(new_n10024), .A2(new_n8458), .B1(new_n9696), .B2(new_n8768), .C(new_n19082), .Y(new_n19083));
  XNOR2x2_ASAP7_75t_L       g18827(.A(\a[59] ), .B(new_n19083), .Y(new_n19084));
  INVx1_ASAP7_75t_L         g18828(.A(new_n19084), .Y(new_n19085));
  A2O1A1Ixp33_ASAP7_75t_L   g18829(.A1(new_n18860), .A2(new_n18932), .B(new_n19016), .C(new_n19018), .Y(new_n19086));
  NOR2xp33_ASAP7_75t_L      g18830(.A(new_n6830), .B(new_n11535), .Y(new_n19087));
  O2A1O1Ixp33_ASAP7_75t_L   g18831(.A1(new_n11247), .A2(new_n11249), .B(\b[49] ), .C(new_n19087), .Y(new_n19088));
  INVx1_ASAP7_75t_L         g18832(.A(new_n19088), .Y(new_n19089));
  A2O1A1Ixp33_ASAP7_75t_L   g18833(.A1(new_n11533), .A2(\b[47] ), .B(new_n18930), .C(new_n6371), .Y(new_n19090));
  A2O1A1O1Ixp25_ASAP7_75t_L g18834(.A1(new_n19005), .A2(new_n19008), .B(new_n19011), .C(new_n19090), .D(new_n19089), .Y(new_n19091));
  INVx1_ASAP7_75t_L         g18835(.A(new_n19087), .Y(new_n19092));
  A2O1A1Ixp33_ASAP7_75t_L   g18836(.A1(new_n19008), .A2(new_n19005), .B(new_n19011), .C(new_n19090), .Y(new_n19093));
  O2A1O1Ixp33_ASAP7_75t_L   g18837(.A1(new_n7317), .A2(new_n11253), .B(new_n19092), .C(new_n19093), .Y(new_n19094));
  NOR2xp33_ASAP7_75t_L      g18838(.A(new_n19091), .B(new_n19094), .Y(new_n19095));
  INVx1_ASAP7_75t_L         g18839(.A(new_n19095), .Y(new_n19096));
  NOR2xp33_ASAP7_75t_L      g18840(.A(new_n7900), .B(new_n10630), .Y(new_n19097));
  AOI221xp5_ASAP7_75t_L     g18841(.A1(\b[50] ), .A2(new_n10939), .B1(\b[51] ), .B2(new_n10632), .C(new_n19097), .Y(new_n19098));
  OAI211xp5_ASAP7_75t_L     g18842(.A1(new_n10629), .A2(new_n7906), .B(\a[62] ), .C(new_n19098), .Y(new_n19099));
  INVx1_ASAP7_75t_L         g18843(.A(new_n19099), .Y(new_n19100));
  O2A1O1Ixp33_ASAP7_75t_L   g18844(.A1(new_n10629), .A2(new_n7906), .B(new_n19098), .C(\a[62] ), .Y(new_n19101));
  NOR2xp33_ASAP7_75t_L      g18845(.A(new_n19101), .B(new_n19100), .Y(new_n19102));
  NOR2xp33_ASAP7_75t_L      g18846(.A(new_n19096), .B(new_n19102), .Y(new_n19103));
  INVx1_ASAP7_75t_L         g18847(.A(new_n19103), .Y(new_n19104));
  NAND2xp33_ASAP7_75t_L     g18848(.A(new_n19096), .B(new_n19102), .Y(new_n19105));
  NAND2xp33_ASAP7_75t_L     g18849(.A(new_n19105), .B(new_n19104), .Y(new_n19106));
  INVx1_ASAP7_75t_L         g18850(.A(new_n19106), .Y(new_n19107));
  O2A1O1Ixp33_ASAP7_75t_L   g18851(.A1(new_n19002), .A2(new_n19014), .B(new_n19086), .C(new_n19107), .Y(new_n19108));
  OA211x2_ASAP7_75t_L       g18852(.A1(new_n19002), .A2(new_n19014), .B(new_n19086), .C(new_n19107), .Y(new_n19109));
  NOR2xp33_ASAP7_75t_L      g18853(.A(new_n19108), .B(new_n19109), .Y(new_n19110));
  XNOR2x2_ASAP7_75t_L       g18854(.A(new_n19085), .B(new_n19110), .Y(new_n19111));
  INVx1_ASAP7_75t_L         g18855(.A(new_n19111), .Y(new_n19112));
  A2O1A1O1Ixp25_ASAP7_75t_L g18856(.A1(new_n18941), .A2(new_n18939), .B(new_n19029), .C(new_n19027), .D(new_n19112), .Y(new_n19113));
  A2O1A1O1Ixp25_ASAP7_75t_L g18857(.A1(new_n18924), .A2(new_n18940), .B(new_n18938), .C(new_n19025), .D(new_n19026), .Y(new_n19114));
  INVx1_ASAP7_75t_L         g18858(.A(new_n19114), .Y(new_n19115));
  NOR2xp33_ASAP7_75t_L      g18859(.A(new_n19111), .B(new_n19115), .Y(new_n19116));
  NOR3xp33_ASAP7_75t_L      g18860(.A(new_n19113), .B(new_n19116), .C(new_n19081), .Y(new_n19117));
  OA21x2_ASAP7_75t_L        g18861(.A1(new_n19116), .A2(new_n19113), .B(new_n19081), .Y(new_n19118));
  NOR2xp33_ASAP7_75t_L      g18862(.A(new_n19117), .B(new_n19118), .Y(new_n19119));
  A2O1A1Ixp33_ASAP7_75t_L   g18863(.A1(new_n19033), .A2(new_n19039), .B(new_n19078), .C(new_n19119), .Y(new_n19120));
  O2A1O1Ixp33_ASAP7_75t_L   g18864(.A1(new_n18946), .A2(new_n18951), .B(new_n19033), .C(new_n19078), .Y(new_n19121));
  INVx1_ASAP7_75t_L         g18865(.A(new_n19119), .Y(new_n19122));
  NAND2xp33_ASAP7_75t_L     g18866(.A(new_n19122), .B(new_n19121), .Y(new_n19123));
  AND2x2_ASAP7_75t_L        g18867(.A(new_n19120), .B(new_n19123), .Y(new_n19124));
  OAI21xp33_ASAP7_75t_L     g18868(.A1(new_n19076), .A2(new_n19077), .B(new_n19124), .Y(new_n19125));
  OR3x1_ASAP7_75t_L         g18869(.A(new_n19124), .B(new_n19076), .C(new_n19077), .Y(new_n19126));
  AND2x2_ASAP7_75t_L        g18870(.A(new_n19125), .B(new_n19126), .Y(new_n19127));
  A2O1A1Ixp33_ASAP7_75t_L   g18871(.A1(new_n19043), .A2(new_n19042), .B(new_n19048), .C(new_n19127), .Y(new_n19128));
  NAND2xp33_ASAP7_75t_L     g18872(.A(new_n19044), .B(new_n19049), .Y(new_n19129));
  NOR2xp33_ASAP7_75t_L      g18873(.A(new_n19127), .B(new_n19129), .Y(new_n19130));
  INVx1_ASAP7_75t_L         g18874(.A(new_n19130), .Y(new_n19131));
  NAND2xp33_ASAP7_75t_L     g18875(.A(new_n19128), .B(new_n19131), .Y(new_n19132));
  NAND2xp33_ASAP7_75t_L     g18876(.A(\b[63] ), .B(new_n7115), .Y(new_n19133));
  OAI221xp5_ASAP7_75t_L     g18877(.A1(new_n7676), .A2(new_n11172), .B1(new_n8237), .B2(new_n11500), .C(new_n19133), .Y(new_n19134));
  XNOR2x2_ASAP7_75t_L       g18878(.A(\a[50] ), .B(new_n19134), .Y(new_n19135));
  XOR2x2_ASAP7_75t_L        g18879(.A(new_n19135), .B(new_n19132), .Y(new_n19136));
  NOR2xp33_ASAP7_75t_L      g18880(.A(new_n19073), .B(new_n19136), .Y(new_n19137));
  NAND2xp33_ASAP7_75t_L     g18881(.A(new_n19073), .B(new_n19136), .Y(new_n19138));
  INVx1_ASAP7_75t_L         g18882(.A(new_n19138), .Y(new_n19139));
  NOR2xp33_ASAP7_75t_L      g18883(.A(new_n19137), .B(new_n19139), .Y(new_n19140));
  A2O1A1Ixp33_ASAP7_75t_L   g18884(.A1(new_n19070), .A2(new_n19067), .B(new_n19066), .C(new_n19140), .Y(new_n19141));
  INVx1_ASAP7_75t_L         g18885(.A(new_n19141), .Y(new_n19142));
  INVx1_ASAP7_75t_L         g18886(.A(new_n19066), .Y(new_n19143));
  A2O1A1Ixp33_ASAP7_75t_L   g18887(.A1(new_n18986), .A2(new_n18983), .B(new_n19068), .C(new_n19143), .Y(new_n19144));
  NOR2xp33_ASAP7_75t_L      g18888(.A(new_n19140), .B(new_n19144), .Y(new_n19145));
  NOR2xp33_ASAP7_75t_L      g18889(.A(new_n19145), .B(new_n19142), .Y(\f[112] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18890(.A1(new_n19002), .A2(new_n19014), .B(new_n19086), .C(new_n19106), .Y(new_n19147));
  O2A1O1Ixp33_ASAP7_75t_L   g18891(.A1(new_n19108), .A2(new_n19109), .B(new_n19085), .C(new_n19147), .Y(new_n19148));
  INVx1_ASAP7_75t_L         g18892(.A(new_n19148), .Y(new_n19149));
  NAND2xp33_ASAP7_75t_L     g18893(.A(\b[51] ), .B(new_n10939), .Y(new_n19150));
  OAI221xp5_ASAP7_75t_L     g18894(.A1(new_n10630), .A2(new_n8165), .B1(new_n10629), .B2(new_n8174), .C(new_n19150), .Y(new_n19151));
  AOI21xp33_ASAP7_75t_L     g18895(.A1(new_n10632), .A2(\b[52] ), .B(new_n19151), .Y(new_n19152));
  NAND2xp33_ASAP7_75t_L     g18896(.A(\a[62] ), .B(new_n19152), .Y(new_n19153));
  A2O1A1Ixp33_ASAP7_75t_L   g18897(.A1(\b[52] ), .A2(new_n10632), .B(new_n19151), .C(new_n10622), .Y(new_n19154));
  NAND2xp33_ASAP7_75t_L     g18898(.A(new_n19154), .B(new_n19153), .Y(new_n19155));
  NOR2xp33_ASAP7_75t_L      g18899(.A(new_n7317), .B(new_n11535), .Y(new_n19156));
  O2A1O1Ixp33_ASAP7_75t_L   g18900(.A1(new_n11247), .A2(new_n11249), .B(\b[50] ), .C(new_n19156), .Y(new_n19157));
  AND2x2_ASAP7_75t_L        g18901(.A(new_n19088), .B(new_n19157), .Y(new_n19158));
  O2A1O1Ixp33_ASAP7_75t_L   g18902(.A1(new_n7317), .A2(new_n11253), .B(new_n19092), .C(new_n19157), .Y(new_n19159));
  NOR2xp33_ASAP7_75t_L      g18903(.A(new_n19159), .B(new_n19158), .Y(new_n19160));
  XOR2x2_ASAP7_75t_L        g18904(.A(new_n19160), .B(new_n19155), .Y(new_n19161));
  A2O1A1O1Ixp25_ASAP7_75t_L g18905(.A1(new_n11533), .A2(\b[47] ), .B(new_n18930), .C(new_n6371), .D(new_n19010), .Y(new_n19162));
  A2O1A1Ixp33_ASAP7_75t_L   g18906(.A1(new_n11533), .A2(\b[49] ), .B(new_n19087), .C(new_n19162), .Y(new_n19163));
  O2A1O1Ixp33_ASAP7_75t_L   g18907(.A1(new_n19101), .A2(new_n19100), .B(new_n19163), .C(new_n19091), .Y(new_n19164));
  NAND2xp33_ASAP7_75t_L     g18908(.A(new_n19164), .B(new_n19161), .Y(new_n19165));
  INVx1_ASAP7_75t_L         g18909(.A(new_n19091), .Y(new_n19166));
  O2A1O1Ixp33_ASAP7_75t_L   g18910(.A1(new_n19096), .A2(new_n19102), .B(new_n19166), .C(new_n19161), .Y(new_n19167));
  INVx1_ASAP7_75t_L         g18911(.A(new_n19167), .Y(new_n19168));
  AOI22xp33_ASAP7_75t_L     g18912(.A1(new_n9700), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n10027), .Y(new_n19169));
  OAI221xp5_ASAP7_75t_L     g18913(.A1(new_n10024), .A2(new_n8762), .B1(new_n9696), .B2(new_n9331), .C(new_n19169), .Y(new_n19170));
  XNOR2x2_ASAP7_75t_L       g18914(.A(\a[59] ), .B(new_n19170), .Y(new_n19171));
  INVx1_ASAP7_75t_L         g18915(.A(new_n19171), .Y(new_n19172));
  AO21x2_ASAP7_75t_L        g18916(.A1(new_n19165), .A2(new_n19168), .B(new_n19172), .Y(new_n19173));
  NAND3xp33_ASAP7_75t_L     g18917(.A(new_n19168), .B(new_n19165), .C(new_n19172), .Y(new_n19174));
  AND2x2_ASAP7_75t_L        g18918(.A(new_n19174), .B(new_n19173), .Y(new_n19175));
  NAND2xp33_ASAP7_75t_L     g18919(.A(new_n19149), .B(new_n19175), .Y(new_n19176));
  NOR2xp33_ASAP7_75t_L      g18920(.A(new_n19149), .B(new_n19175), .Y(new_n19177));
  INVx1_ASAP7_75t_L         g18921(.A(new_n19177), .Y(new_n19178));
  AOI22xp33_ASAP7_75t_L     g18922(.A1(new_n8831), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n9115), .Y(new_n19179));
  OAI221xp5_ASAP7_75t_L     g18923(.A1(new_n10343), .A2(new_n9920), .B1(new_n10016), .B2(new_n11152), .C(new_n19179), .Y(new_n19180));
  XNOR2x2_ASAP7_75t_L       g18924(.A(\a[56] ), .B(new_n19180), .Y(new_n19181));
  NAND3xp33_ASAP7_75t_L     g18925(.A(new_n19178), .B(new_n19176), .C(new_n19181), .Y(new_n19182));
  AO21x2_ASAP7_75t_L        g18926(.A1(new_n19176), .A2(new_n19178), .B(new_n19181), .Y(new_n19183));
  AND2x2_ASAP7_75t_L        g18927(.A(new_n19182), .B(new_n19183), .Y(new_n19184));
  O2A1O1Ixp33_ASAP7_75t_L   g18928(.A1(new_n19026), .A2(new_n19030), .B(new_n19111), .C(new_n19117), .Y(new_n19185));
  NAND2xp33_ASAP7_75t_L     g18929(.A(new_n19185), .B(new_n19184), .Y(new_n19186));
  INVx1_ASAP7_75t_L         g18930(.A(new_n19184), .Y(new_n19187));
  A2O1A1Ixp33_ASAP7_75t_L   g18931(.A1(new_n19111), .A2(new_n19115), .B(new_n19117), .C(new_n19187), .Y(new_n19188));
  AOI22xp33_ASAP7_75t_L     g18932(.A1(new_n7960), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n8537), .Y(new_n19189));
  OAI221xp5_ASAP7_75t_L     g18933(.A1(new_n8817), .A2(new_n10847), .B1(new_n7957), .B2(new_n12047), .C(new_n19189), .Y(new_n19190));
  XNOR2x2_ASAP7_75t_L       g18934(.A(\a[53] ), .B(new_n19190), .Y(new_n19191));
  NAND3xp33_ASAP7_75t_L     g18935(.A(new_n19188), .B(new_n19186), .C(new_n19191), .Y(new_n19192));
  AO21x2_ASAP7_75t_L        g18936(.A1(new_n19186), .A2(new_n19188), .B(new_n19191), .Y(new_n19193));
  NAND2xp33_ASAP7_75t_L     g18937(.A(new_n19192), .B(new_n19193), .Y(new_n19194));
  A2O1A1Ixp33_ASAP7_75t_L   g18938(.A1(new_n19037), .A2(new_n19035), .B(new_n19122), .C(new_n19125), .Y(new_n19195));
  A2O1A1Ixp33_ASAP7_75t_L   g18939(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n7108), .Y(new_n19196));
  A2O1A1Ixp33_ASAP7_75t_L   g18940(.A1(new_n19196), .A2(new_n7676), .B(new_n11468), .C(\a[50] ), .Y(new_n19197));
  O2A1O1Ixp33_ASAP7_75t_L   g18941(.A1(new_n8237), .A2(new_n12060), .B(new_n7676), .C(new_n11468), .Y(new_n19198));
  NAND2xp33_ASAP7_75t_L     g18942(.A(new_n7106), .B(new_n19198), .Y(new_n19199));
  NAND2xp33_ASAP7_75t_L     g18943(.A(new_n19199), .B(new_n19197), .Y(new_n19200));
  NAND2xp33_ASAP7_75t_L     g18944(.A(new_n19200), .B(new_n19195), .Y(new_n19201));
  NOR2xp33_ASAP7_75t_L      g18945(.A(new_n19200), .B(new_n19195), .Y(new_n19202));
  INVx1_ASAP7_75t_L         g18946(.A(new_n19202), .Y(new_n19203));
  NAND2xp33_ASAP7_75t_L     g18947(.A(new_n19201), .B(new_n19203), .Y(new_n19204));
  NAND2xp33_ASAP7_75t_L     g18948(.A(new_n19194), .B(new_n19204), .Y(new_n19205));
  NOR2xp33_ASAP7_75t_L      g18949(.A(new_n19194), .B(new_n19204), .Y(new_n19206));
  INVx1_ASAP7_75t_L         g18950(.A(new_n19206), .Y(new_n19207));
  NAND2xp33_ASAP7_75t_L     g18951(.A(new_n19205), .B(new_n19207), .Y(new_n19208));
  OAI21xp33_ASAP7_75t_L     g18952(.A1(new_n19135), .A2(new_n19130), .B(new_n19128), .Y(new_n19209));
  NOR2xp33_ASAP7_75t_L      g18953(.A(new_n19208), .B(new_n19209), .Y(new_n19210));
  NAND2xp33_ASAP7_75t_L     g18954(.A(new_n19208), .B(new_n19209), .Y(new_n19211));
  INVx1_ASAP7_75t_L         g18955(.A(new_n19211), .Y(new_n19212));
  NOR2xp33_ASAP7_75t_L      g18956(.A(new_n19210), .B(new_n19212), .Y(new_n19213));
  A2O1A1Ixp33_ASAP7_75t_L   g18957(.A1(new_n19144), .A2(new_n19140), .B(new_n19139), .C(new_n19213), .Y(new_n19214));
  INVx1_ASAP7_75t_L         g18958(.A(new_n19214), .Y(new_n19215));
  INVx1_ASAP7_75t_L         g18959(.A(new_n19069), .Y(new_n19216));
  A2O1A1Ixp33_ASAP7_75t_L   g18960(.A1(new_n19216), .A2(new_n19143), .B(new_n19137), .C(new_n19138), .Y(new_n19217));
  NOR2xp33_ASAP7_75t_L      g18961(.A(new_n19213), .B(new_n19217), .Y(new_n19218));
  NOR2xp33_ASAP7_75t_L      g18962(.A(new_n19215), .B(new_n19218), .Y(\f[113] ));
  AOI22xp33_ASAP7_75t_L     g18963(.A1(new_n8831), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n9115), .Y(new_n19220));
  OAI221xp5_ASAP7_75t_L     g18964(.A1(new_n10343), .A2(new_n9947), .B1(new_n10016), .B2(new_n11446), .C(new_n19220), .Y(new_n19221));
  XNOR2x2_ASAP7_75t_L       g18965(.A(\a[56] ), .B(new_n19221), .Y(new_n19222));
  AOI22xp33_ASAP7_75t_L     g18966(.A1(new_n9700), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n10027), .Y(new_n19223));
  OAI221xp5_ASAP7_75t_L     g18967(.A1(new_n10024), .A2(new_n9323), .B1(new_n9696), .B2(new_n9627), .C(new_n19223), .Y(new_n19224));
  XNOR2x2_ASAP7_75t_L       g18968(.A(\a[59] ), .B(new_n19224), .Y(new_n19225));
  INVx1_ASAP7_75t_L         g18969(.A(new_n19225), .Y(new_n19226));
  AOI22xp33_ASAP7_75t_L     g18970(.A1(\b[52] ), .A2(new_n10939), .B1(\b[54] ), .B2(new_n10938), .Y(new_n19227));
  OAI221xp5_ASAP7_75t_L     g18971(.A1(new_n10937), .A2(new_n8165), .B1(new_n10629), .B2(new_n8465), .C(new_n19227), .Y(new_n19228));
  XNOR2x2_ASAP7_75t_L       g18972(.A(\a[62] ), .B(new_n19228), .Y(new_n19229));
  A2O1A1Ixp33_ASAP7_75t_L   g18973(.A1(\b[50] ), .A2(new_n11533), .B(new_n19156), .C(new_n19088), .Y(new_n19230));
  NOR2xp33_ASAP7_75t_L      g18974(.A(new_n7593), .B(new_n11535), .Y(new_n19231));
  A2O1A1Ixp33_ASAP7_75t_L   g18975(.A1(new_n11533), .A2(\b[51] ), .B(new_n19231), .C(new_n7106), .Y(new_n19232));
  INVx1_ASAP7_75t_L         g18976(.A(new_n19232), .Y(new_n19233));
  O2A1O1Ixp33_ASAP7_75t_L   g18977(.A1(new_n11247), .A2(new_n11249), .B(\b[51] ), .C(new_n19231), .Y(new_n19234));
  NAND2xp33_ASAP7_75t_L     g18978(.A(\a[50] ), .B(new_n19234), .Y(new_n19235));
  INVx1_ASAP7_75t_L         g18979(.A(new_n19235), .Y(new_n19236));
  NOR2xp33_ASAP7_75t_L      g18980(.A(new_n19233), .B(new_n19236), .Y(new_n19237));
  INVx1_ASAP7_75t_L         g18981(.A(new_n19237), .Y(new_n19238));
  O2A1O1Ixp33_ASAP7_75t_L   g18982(.A1(new_n7317), .A2(new_n11253), .B(new_n19092), .C(new_n19238), .Y(new_n19239));
  INVx1_ASAP7_75t_L         g18983(.A(new_n19239), .Y(new_n19240));
  NAND2xp33_ASAP7_75t_L     g18984(.A(new_n19088), .B(new_n19238), .Y(new_n19241));
  AND2x2_ASAP7_75t_L        g18985(.A(new_n19241), .B(new_n19240), .Y(new_n19242));
  A2O1A1O1Ixp25_ASAP7_75t_L g18986(.A1(new_n19154), .A2(new_n19153), .B(new_n19160), .C(new_n19230), .D(new_n19242), .Y(new_n19243));
  A2O1A1Ixp33_ASAP7_75t_L   g18987(.A1(new_n19153), .A2(new_n19154), .B(new_n19160), .C(new_n19230), .Y(new_n19244));
  INVx1_ASAP7_75t_L         g18988(.A(new_n19242), .Y(new_n19245));
  NOR2xp33_ASAP7_75t_L      g18989(.A(new_n19245), .B(new_n19244), .Y(new_n19246));
  NOR2xp33_ASAP7_75t_L      g18990(.A(new_n19243), .B(new_n19246), .Y(new_n19247));
  NOR2xp33_ASAP7_75t_L      g18991(.A(new_n19229), .B(new_n19247), .Y(new_n19248));
  INVx1_ASAP7_75t_L         g18992(.A(new_n19229), .Y(new_n19249));
  NOR3xp33_ASAP7_75t_L      g18993(.A(new_n19246), .B(new_n19249), .C(new_n19243), .Y(new_n19250));
  NOR2xp33_ASAP7_75t_L      g18994(.A(new_n19250), .B(new_n19248), .Y(new_n19251));
  XNOR2x2_ASAP7_75t_L       g18995(.A(new_n19226), .B(new_n19251), .Y(new_n19252));
  O2A1O1Ixp33_ASAP7_75t_L   g18996(.A1(new_n19161), .A2(new_n19164), .B(new_n19174), .C(new_n19252), .Y(new_n19253));
  AND3x1_ASAP7_75t_L        g18997(.A(new_n19252), .B(new_n19174), .C(new_n19168), .Y(new_n19254));
  OR3x1_ASAP7_75t_L         g18998(.A(new_n19254), .B(new_n19222), .C(new_n19253), .Y(new_n19255));
  OAI21xp33_ASAP7_75t_L     g18999(.A1(new_n19253), .A2(new_n19254), .B(new_n19222), .Y(new_n19256));
  AND2x2_ASAP7_75t_L        g19000(.A(new_n19256), .B(new_n19255), .Y(new_n19257));
  NAND3xp33_ASAP7_75t_L     g19001(.A(new_n19257), .B(new_n19182), .C(new_n19178), .Y(new_n19258));
  INVx1_ASAP7_75t_L         g19002(.A(new_n19257), .Y(new_n19259));
  A2O1A1Ixp33_ASAP7_75t_L   g19003(.A1(new_n19181), .A2(new_n19176), .B(new_n19177), .C(new_n19259), .Y(new_n19260));
  NAND2xp33_ASAP7_75t_L     g19004(.A(new_n19258), .B(new_n19260), .Y(new_n19261));
  AOI22xp33_ASAP7_75t_L     g19005(.A1(new_n7960), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n8537), .Y(new_n19262));
  A2O1A1Ixp33_ASAP7_75t_L   g19006(.A1(new_n11470), .A2(new_n11473), .B(new_n7957), .C(new_n19262), .Y(new_n19263));
  AOI21xp33_ASAP7_75t_L     g19007(.A1(new_n7963), .A2(\b[62] ), .B(new_n19263), .Y(new_n19264));
  NAND2xp33_ASAP7_75t_L     g19008(.A(\a[53] ), .B(new_n19264), .Y(new_n19265));
  A2O1A1Ixp33_ASAP7_75t_L   g19009(.A1(\b[62] ), .A2(new_n7963), .B(new_n19263), .C(new_n7954), .Y(new_n19266));
  NAND2xp33_ASAP7_75t_L     g19010(.A(new_n19266), .B(new_n19265), .Y(new_n19267));
  XNOR2x2_ASAP7_75t_L       g19011(.A(new_n19267), .B(new_n19261), .Y(new_n19268));
  AO21x2_ASAP7_75t_L        g19012(.A1(new_n19186), .A2(new_n19192), .B(new_n19268), .Y(new_n19269));
  NAND3xp33_ASAP7_75t_L     g19013(.A(new_n19268), .B(new_n19192), .C(new_n19186), .Y(new_n19270));
  AND2x2_ASAP7_75t_L        g19014(.A(new_n19270), .B(new_n19269), .Y(new_n19271));
  O2A1O1Ixp33_ASAP7_75t_L   g19015(.A1(new_n19194), .A2(new_n19204), .B(new_n19203), .C(new_n19271), .Y(new_n19272));
  INVx1_ASAP7_75t_L         g19016(.A(new_n19271), .Y(new_n19273));
  NOR2xp33_ASAP7_75t_L      g19017(.A(new_n19202), .B(new_n19206), .Y(new_n19274));
  INVx1_ASAP7_75t_L         g19018(.A(new_n19274), .Y(new_n19275));
  NOR2xp33_ASAP7_75t_L      g19019(.A(new_n19273), .B(new_n19275), .Y(new_n19276));
  NOR2xp33_ASAP7_75t_L      g19020(.A(new_n19272), .B(new_n19276), .Y(new_n19277));
  INVx1_ASAP7_75t_L         g19021(.A(new_n19277), .Y(new_n19278));
  A2O1A1O1Ixp25_ASAP7_75t_L g19022(.A1(new_n19138), .A2(new_n19141), .B(new_n19210), .C(new_n19211), .D(new_n19278), .Y(new_n19279));
  A2O1A1Ixp33_ASAP7_75t_L   g19023(.A1(new_n19141), .A2(new_n19138), .B(new_n19210), .C(new_n19211), .Y(new_n19280));
  NOR2xp33_ASAP7_75t_L      g19024(.A(new_n19277), .B(new_n19280), .Y(new_n19281));
  NOR2xp33_ASAP7_75t_L      g19025(.A(new_n19279), .B(new_n19281), .Y(\f[114] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19026(.A1(new_n19265), .A2(new_n19266), .B(new_n19261), .C(new_n19270), .Y(new_n19283));
  NAND2xp33_ASAP7_75t_L     g19027(.A(new_n19255), .B(new_n19258), .Y(new_n19284));
  AOI22xp33_ASAP7_75t_L     g19028(.A1(new_n8831), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n9115), .Y(new_n19285));
  OAI221xp5_ASAP7_75t_L     g19029(.A1(new_n10343), .A2(new_n10250), .B1(new_n10016), .B2(new_n10855), .C(new_n19285), .Y(new_n19286));
  NOR2xp33_ASAP7_75t_L      g19030(.A(new_n8826), .B(new_n19286), .Y(new_n19287));
  AND2x2_ASAP7_75t_L        g19031(.A(new_n8826), .B(new_n19286), .Y(new_n19288));
  NOR2xp33_ASAP7_75t_L      g19032(.A(new_n19287), .B(new_n19288), .Y(new_n19289));
  NAND2xp33_ASAP7_75t_L     g19033(.A(new_n19226), .B(new_n19251), .Y(new_n19290));
  AOI22xp33_ASAP7_75t_L     g19034(.A1(new_n9700), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n10027), .Y(new_n19291));
  OAI221xp5_ASAP7_75t_L     g19035(.A1(new_n10024), .A2(new_n9620), .B1(new_n9696), .B2(new_n9925), .C(new_n19291), .Y(new_n19292));
  XNOR2x2_ASAP7_75t_L       g19036(.A(\a[59] ), .B(new_n19292), .Y(new_n19293));
  NOR2xp33_ASAP7_75t_L      g19037(.A(new_n7616), .B(new_n11535), .Y(new_n19294));
  A2O1A1O1Ixp25_ASAP7_75t_L g19038(.A1(new_n11533), .A2(\b[49] ), .B(new_n19087), .C(new_n19235), .D(new_n19233), .Y(new_n19295));
  A2O1A1Ixp33_ASAP7_75t_L   g19039(.A1(new_n11533), .A2(\b[52] ), .B(new_n19294), .C(new_n19295), .Y(new_n19296));
  O2A1O1Ixp33_ASAP7_75t_L   g19040(.A1(new_n11247), .A2(new_n11249), .B(\b[52] ), .C(new_n19294), .Y(new_n19297));
  INVx1_ASAP7_75t_L         g19041(.A(new_n19297), .Y(new_n19298));
  O2A1O1Ixp33_ASAP7_75t_L   g19042(.A1(new_n19088), .A2(new_n19236), .B(new_n19232), .C(new_n19298), .Y(new_n19299));
  INVx1_ASAP7_75t_L         g19043(.A(new_n19299), .Y(new_n19300));
  NAND2xp33_ASAP7_75t_L     g19044(.A(new_n19296), .B(new_n19300), .Y(new_n19301));
  NAND2xp33_ASAP7_75t_L     g19045(.A(\b[53] ), .B(new_n10939), .Y(new_n19302));
  OAI221xp5_ASAP7_75t_L     g19046(.A1(new_n10630), .A2(new_n8762), .B1(new_n10629), .B2(new_n8768), .C(new_n19302), .Y(new_n19303));
  AOI21xp33_ASAP7_75t_L     g19047(.A1(new_n10632), .A2(\b[54] ), .B(new_n19303), .Y(new_n19304));
  NAND2xp33_ASAP7_75t_L     g19048(.A(\a[62] ), .B(new_n19304), .Y(new_n19305));
  A2O1A1Ixp33_ASAP7_75t_L   g19049(.A1(\b[54] ), .A2(new_n10632), .B(new_n19303), .C(new_n10622), .Y(new_n19306));
  AND2x2_ASAP7_75t_L        g19050(.A(new_n19306), .B(new_n19305), .Y(new_n19307));
  NAND2xp33_ASAP7_75t_L     g19051(.A(new_n19301), .B(new_n19307), .Y(new_n19308));
  NOR2xp33_ASAP7_75t_L      g19052(.A(new_n19301), .B(new_n19307), .Y(new_n19309));
  INVx1_ASAP7_75t_L         g19053(.A(new_n19309), .Y(new_n19310));
  AND2x2_ASAP7_75t_L        g19054(.A(new_n19308), .B(new_n19310), .Y(new_n19311));
  A2O1A1Ixp33_ASAP7_75t_L   g19055(.A1(new_n19242), .A2(new_n19244), .B(new_n19248), .C(new_n19311), .Y(new_n19312));
  INVx1_ASAP7_75t_L         g19056(.A(new_n19312), .Y(new_n19313));
  A2O1A1O1Ixp25_ASAP7_75t_L g19057(.A1(new_n19154), .A2(new_n19153), .B(new_n19160), .C(new_n19230), .D(new_n19245), .Y(new_n19314));
  O2A1O1Ixp33_ASAP7_75t_L   g19058(.A1(new_n19243), .A2(new_n19246), .B(new_n19249), .C(new_n19314), .Y(new_n19315));
  INVx1_ASAP7_75t_L         g19059(.A(new_n19315), .Y(new_n19316));
  NOR2xp33_ASAP7_75t_L      g19060(.A(new_n19316), .B(new_n19311), .Y(new_n19317));
  NOR2xp33_ASAP7_75t_L      g19061(.A(new_n19317), .B(new_n19313), .Y(new_n19318));
  INVx1_ASAP7_75t_L         g19062(.A(new_n19318), .Y(new_n19319));
  NOR2xp33_ASAP7_75t_L      g19063(.A(new_n19293), .B(new_n19319), .Y(new_n19320));
  INVx1_ASAP7_75t_L         g19064(.A(new_n19320), .Y(new_n19321));
  NAND2xp33_ASAP7_75t_L     g19065(.A(new_n19293), .B(new_n19319), .Y(new_n19322));
  AND2x2_ASAP7_75t_L        g19066(.A(new_n19322), .B(new_n19321), .Y(new_n19323));
  INVx1_ASAP7_75t_L         g19067(.A(new_n19323), .Y(new_n19324));
  A2O1A1O1Ixp25_ASAP7_75t_L g19068(.A1(new_n19174), .A2(new_n19168), .B(new_n19252), .C(new_n19290), .D(new_n19324), .Y(new_n19325));
  A2O1A1Ixp33_ASAP7_75t_L   g19069(.A1(new_n19174), .A2(new_n19168), .B(new_n19252), .C(new_n19290), .Y(new_n19326));
  NOR2xp33_ASAP7_75t_L      g19070(.A(new_n19326), .B(new_n19323), .Y(new_n19327));
  NOR2xp33_ASAP7_75t_L      g19071(.A(new_n19327), .B(new_n19325), .Y(new_n19328));
  XNOR2x2_ASAP7_75t_L       g19072(.A(new_n19289), .B(new_n19328), .Y(new_n19329));
  NAND2xp33_ASAP7_75t_L     g19073(.A(new_n19284), .B(new_n19329), .Y(new_n19330));
  NOR2xp33_ASAP7_75t_L      g19074(.A(new_n19284), .B(new_n19329), .Y(new_n19331));
  INVx1_ASAP7_75t_L         g19075(.A(new_n19331), .Y(new_n19332));
  NAND2xp33_ASAP7_75t_L     g19076(.A(new_n19330), .B(new_n19332), .Y(new_n19333));
  NAND2xp33_ASAP7_75t_L     g19077(.A(\b[63] ), .B(new_n7963), .Y(new_n19334));
  OAI221xp5_ASAP7_75t_L     g19078(.A1(new_n8247), .A2(new_n11172), .B1(new_n7957), .B2(new_n11500), .C(new_n19334), .Y(new_n19335));
  XNOR2x2_ASAP7_75t_L       g19079(.A(\a[53] ), .B(new_n19335), .Y(new_n19336));
  XOR2x2_ASAP7_75t_L        g19080(.A(new_n19336), .B(new_n19333), .Y(new_n19337));
  NOR2xp33_ASAP7_75t_L      g19081(.A(new_n19283), .B(new_n19337), .Y(new_n19338));
  NAND2xp33_ASAP7_75t_L     g19082(.A(new_n19283), .B(new_n19337), .Y(new_n19339));
  INVx1_ASAP7_75t_L         g19083(.A(new_n19339), .Y(new_n19340));
  NOR2xp33_ASAP7_75t_L      g19084(.A(new_n19338), .B(new_n19340), .Y(new_n19341));
  A2O1A1Ixp33_ASAP7_75t_L   g19085(.A1(new_n19280), .A2(new_n19277), .B(new_n19276), .C(new_n19341), .Y(new_n19342));
  INVx1_ASAP7_75t_L         g19086(.A(new_n19342), .Y(new_n19343));
  INVx1_ASAP7_75t_L         g19087(.A(new_n19276), .Y(new_n19344));
  A2O1A1Ixp33_ASAP7_75t_L   g19088(.A1(new_n19214), .A2(new_n19211), .B(new_n19278), .C(new_n19344), .Y(new_n19345));
  NOR2xp33_ASAP7_75t_L      g19089(.A(new_n19341), .B(new_n19345), .Y(new_n19346));
  NOR2xp33_ASAP7_75t_L      g19090(.A(new_n19346), .B(new_n19343), .Y(\f[115] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19091(.A1(new_n19248), .A2(new_n19314), .B(new_n19311), .C(new_n19320), .Y(new_n19348));
  AOI22xp33_ASAP7_75t_L     g19092(.A1(new_n9700), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n10027), .Y(new_n19349));
  OAI221xp5_ASAP7_75t_L     g19093(.A1(new_n10024), .A2(new_n9920), .B1(new_n9696), .B2(new_n11152), .C(new_n19349), .Y(new_n19350));
  XNOR2x2_ASAP7_75t_L       g19094(.A(\a[59] ), .B(new_n19350), .Y(new_n19351));
  INVx1_ASAP7_75t_L         g19095(.A(new_n19351), .Y(new_n19352));
  AOI22xp33_ASAP7_75t_L     g19096(.A1(\b[54] ), .A2(new_n10939), .B1(\b[56] ), .B2(new_n10938), .Y(new_n19353));
  OAI221xp5_ASAP7_75t_L     g19097(.A1(new_n10937), .A2(new_n8762), .B1(new_n10629), .B2(new_n9331), .C(new_n19353), .Y(new_n19354));
  XNOR2x2_ASAP7_75t_L       g19098(.A(\a[62] ), .B(new_n19354), .Y(new_n19355));
  NOR2xp33_ASAP7_75t_L      g19099(.A(new_n7900), .B(new_n11535), .Y(new_n19356));
  A2O1A1Ixp33_ASAP7_75t_L   g19100(.A1(\b[53] ), .A2(new_n11533), .B(new_n19356), .C(new_n19297), .Y(new_n19357));
  O2A1O1Ixp33_ASAP7_75t_L   g19101(.A1(new_n11247), .A2(new_n11249), .B(\b[53] ), .C(new_n19356), .Y(new_n19358));
  A2O1A1Ixp33_ASAP7_75t_L   g19102(.A1(new_n11533), .A2(\b[52] ), .B(new_n19294), .C(new_n19358), .Y(new_n19359));
  AND2x2_ASAP7_75t_L        g19103(.A(new_n19357), .B(new_n19359), .Y(new_n19360));
  AND3x1_ASAP7_75t_L        g19104(.A(new_n19310), .B(new_n19360), .C(new_n19300), .Y(new_n19361));
  A2O1A1O1Ixp25_ASAP7_75t_L g19105(.A1(new_n19306), .A2(new_n19305), .B(new_n19301), .C(new_n19300), .D(new_n19360), .Y(new_n19362));
  NOR2xp33_ASAP7_75t_L      g19106(.A(new_n19362), .B(new_n19361), .Y(new_n19363));
  NOR2xp33_ASAP7_75t_L      g19107(.A(new_n19355), .B(new_n19363), .Y(new_n19364));
  INVx1_ASAP7_75t_L         g19108(.A(new_n19364), .Y(new_n19365));
  NAND2xp33_ASAP7_75t_L     g19109(.A(new_n19355), .B(new_n19363), .Y(new_n19366));
  NAND3xp33_ASAP7_75t_L     g19110(.A(new_n19365), .B(new_n19352), .C(new_n19366), .Y(new_n19367));
  AO21x2_ASAP7_75t_L        g19111(.A1(new_n19366), .A2(new_n19365), .B(new_n19352), .Y(new_n19368));
  AND2x2_ASAP7_75t_L        g19112(.A(new_n19367), .B(new_n19368), .Y(new_n19369));
  INVx1_ASAP7_75t_L         g19113(.A(new_n19369), .Y(new_n19370));
  NAND2xp33_ASAP7_75t_L     g19114(.A(new_n19348), .B(new_n19370), .Y(new_n19371));
  A2O1A1Ixp33_ASAP7_75t_L   g19115(.A1(new_n19311), .A2(new_n19316), .B(new_n19320), .C(new_n19369), .Y(new_n19372));
  AOI22xp33_ASAP7_75t_L     g19116(.A1(new_n8831), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n9115), .Y(new_n19373));
  OAI221xp5_ASAP7_75t_L     g19117(.A1(new_n10343), .A2(new_n10847), .B1(new_n10016), .B2(new_n12047), .C(new_n19373), .Y(new_n19374));
  XNOR2x2_ASAP7_75t_L       g19118(.A(\a[56] ), .B(new_n19374), .Y(new_n19375));
  NAND3xp33_ASAP7_75t_L     g19119(.A(new_n19371), .B(new_n19372), .C(new_n19375), .Y(new_n19376));
  AO21x2_ASAP7_75t_L        g19120(.A1(new_n19372), .A2(new_n19371), .B(new_n19375), .Y(new_n19377));
  INVx1_ASAP7_75t_L         g19121(.A(new_n19289), .Y(new_n19378));
  A2O1A1Ixp33_ASAP7_75t_L   g19122(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n7958), .Y(new_n19379));
  A2O1A1Ixp33_ASAP7_75t_L   g19123(.A1(new_n19379), .A2(new_n8247), .B(new_n11468), .C(\a[53] ), .Y(new_n19380));
  O2A1O1Ixp33_ASAP7_75t_L   g19124(.A1(new_n7957), .A2(new_n12060), .B(new_n8247), .C(new_n11468), .Y(new_n19381));
  NAND2xp33_ASAP7_75t_L     g19125(.A(new_n7954), .B(new_n19381), .Y(new_n19382));
  NAND2xp33_ASAP7_75t_L     g19126(.A(new_n19382), .B(new_n19380), .Y(new_n19383));
  A2O1A1Ixp33_ASAP7_75t_L   g19127(.A1(new_n19328), .A2(new_n19378), .B(new_n19325), .C(new_n19383), .Y(new_n19384));
  O2A1O1Ixp33_ASAP7_75t_L   g19128(.A1(new_n19288), .A2(new_n19287), .B(new_n19328), .C(new_n19325), .Y(new_n19385));
  NAND3xp33_ASAP7_75t_L     g19129(.A(new_n19385), .B(new_n19380), .C(new_n19382), .Y(new_n19386));
  AOI22xp33_ASAP7_75t_L     g19130(.A1(new_n19376), .A2(new_n19377), .B1(new_n19384), .B2(new_n19386), .Y(new_n19387));
  NAND2xp33_ASAP7_75t_L     g19131(.A(new_n19376), .B(new_n19377), .Y(new_n19388));
  NAND2xp33_ASAP7_75t_L     g19132(.A(new_n19384), .B(new_n19386), .Y(new_n19389));
  NOR2xp33_ASAP7_75t_L      g19133(.A(new_n19388), .B(new_n19389), .Y(new_n19390));
  NOR2xp33_ASAP7_75t_L      g19134(.A(new_n19387), .B(new_n19390), .Y(new_n19391));
  OAI211xp5_ASAP7_75t_L     g19135(.A1(new_n19331), .A2(new_n19336), .B(new_n19391), .C(new_n19330), .Y(new_n19392));
  O2A1O1Ixp33_ASAP7_75t_L   g19136(.A1(new_n19331), .A2(new_n19336), .B(new_n19330), .C(new_n19391), .Y(new_n19393));
  INVx1_ASAP7_75t_L         g19137(.A(new_n19393), .Y(new_n19394));
  AND2x2_ASAP7_75t_L        g19138(.A(new_n19392), .B(new_n19394), .Y(new_n19395));
  A2O1A1Ixp33_ASAP7_75t_L   g19139(.A1(new_n19345), .A2(new_n19341), .B(new_n19340), .C(new_n19395), .Y(new_n19396));
  INVx1_ASAP7_75t_L         g19140(.A(new_n19395), .Y(new_n19397));
  A2O1A1O1Ixp25_ASAP7_75t_L g19141(.A1(new_n19277), .A2(new_n19280), .B(new_n19276), .C(new_n19341), .D(new_n19340), .Y(new_n19398));
  NAND2xp33_ASAP7_75t_L     g19142(.A(new_n19397), .B(new_n19398), .Y(new_n19399));
  AND2x2_ASAP7_75t_L        g19143(.A(new_n19396), .B(new_n19399), .Y(\f[116] ));
  AOI22xp33_ASAP7_75t_L     g19144(.A1(new_n8831), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n9115), .Y(new_n19401));
  A2O1A1Ixp33_ASAP7_75t_L   g19145(.A1(new_n11470), .A2(new_n11473), .B(new_n10016), .C(new_n19401), .Y(new_n19402));
  AOI21xp33_ASAP7_75t_L     g19146(.A1(new_n8835), .A2(\b[62] ), .B(new_n19402), .Y(new_n19403));
  NAND2xp33_ASAP7_75t_L     g19147(.A(\a[56] ), .B(new_n19403), .Y(new_n19404));
  A2O1A1Ixp33_ASAP7_75t_L   g19148(.A1(\b[62] ), .A2(new_n8835), .B(new_n19402), .C(new_n8826), .Y(new_n19405));
  INVx1_ASAP7_75t_L         g19149(.A(new_n19348), .Y(new_n19406));
  A2O1A1Ixp33_ASAP7_75t_L   g19150(.A1(new_n19367), .A2(new_n19368), .B(new_n19406), .C(new_n19376), .Y(new_n19407));
  AOI21xp33_ASAP7_75t_L     g19151(.A1(new_n19405), .A2(new_n19404), .B(new_n19407), .Y(new_n19408));
  NAND2xp33_ASAP7_75t_L     g19152(.A(new_n19405), .B(new_n19404), .Y(new_n19409));
  O2A1O1Ixp33_ASAP7_75t_L   g19153(.A1(new_n19406), .A2(new_n19369), .B(new_n19376), .C(new_n19409), .Y(new_n19410));
  AOI22xp33_ASAP7_75t_L     g19154(.A1(new_n9700), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n10027), .Y(new_n19411));
  OAI221xp5_ASAP7_75t_L     g19155(.A1(new_n10024), .A2(new_n9947), .B1(new_n9696), .B2(new_n11446), .C(new_n19411), .Y(new_n19412));
  XNOR2x2_ASAP7_75t_L       g19156(.A(\a[59] ), .B(new_n19412), .Y(new_n19413));
  INVx1_ASAP7_75t_L         g19157(.A(new_n19413), .Y(new_n19414));
  A2O1A1Ixp33_ASAP7_75t_L   g19158(.A1(new_n11533), .A2(\b[53] ), .B(new_n19356), .C(\a[53] ), .Y(new_n19415));
  INVx1_ASAP7_75t_L         g19159(.A(new_n19358), .Y(new_n19416));
  NOR2xp33_ASAP7_75t_L      g19160(.A(\a[53] ), .B(new_n19416), .Y(new_n19417));
  INVx1_ASAP7_75t_L         g19161(.A(new_n19417), .Y(new_n19418));
  AND2x2_ASAP7_75t_L        g19162(.A(new_n19415), .B(new_n19418), .Y(new_n19419));
  INVx1_ASAP7_75t_L         g19163(.A(new_n19419), .Y(new_n19420));
  NOR2xp33_ASAP7_75t_L      g19164(.A(new_n8165), .B(new_n11535), .Y(new_n19421));
  INVx1_ASAP7_75t_L         g19165(.A(new_n19421), .Y(new_n19422));
  A2O1A1Ixp33_ASAP7_75t_L   g19166(.A1(new_n14788), .A2(new_n14789), .B(new_n8458), .C(new_n19422), .Y(new_n19423));
  NOR2xp33_ASAP7_75t_L      g19167(.A(new_n19423), .B(new_n19420), .Y(new_n19424));
  O2A1O1Ixp33_ASAP7_75t_L   g19168(.A1(new_n11253), .A2(new_n8458), .B(new_n19422), .C(new_n19419), .Y(new_n19425));
  NOR2xp33_ASAP7_75t_L      g19169(.A(new_n19425), .B(new_n19424), .Y(new_n19426));
  INVx1_ASAP7_75t_L         g19170(.A(new_n19426), .Y(new_n19427));
  AOI22xp33_ASAP7_75t_L     g19171(.A1(\b[55] ), .A2(new_n10939), .B1(\b[57] ), .B2(new_n10938), .Y(new_n19428));
  OAI221xp5_ASAP7_75t_L     g19172(.A1(new_n10937), .A2(new_n9323), .B1(new_n10629), .B2(new_n9627), .C(new_n19428), .Y(new_n19429));
  XNOR2x2_ASAP7_75t_L       g19173(.A(\a[62] ), .B(new_n19429), .Y(new_n19430));
  XNOR2x2_ASAP7_75t_L       g19174(.A(new_n19427), .B(new_n19430), .Y(new_n19431));
  INVx1_ASAP7_75t_L         g19175(.A(new_n19431), .Y(new_n19432));
  O2A1O1Ixp33_ASAP7_75t_L   g19176(.A1(new_n19233), .A2(new_n19239), .B(new_n19297), .C(new_n19309), .Y(new_n19433));
  A2O1A1O1Ixp25_ASAP7_75t_L g19177(.A1(\b[53] ), .A2(new_n11533), .B(new_n19356), .C(new_n19297), .D(new_n19433), .Y(new_n19434));
  A2O1A1Ixp33_ASAP7_75t_L   g19178(.A1(new_n19298), .A2(new_n19358), .B(new_n19434), .C(new_n19432), .Y(new_n19435));
  A2O1A1O1Ixp25_ASAP7_75t_L g19179(.A1(new_n11533), .A2(\b[52] ), .B(new_n19294), .C(new_n19358), .D(new_n19434), .Y(new_n19436));
  NAND2xp33_ASAP7_75t_L     g19180(.A(new_n19431), .B(new_n19436), .Y(new_n19437));
  AND2x2_ASAP7_75t_L        g19181(.A(new_n19435), .B(new_n19437), .Y(new_n19438));
  XNOR2x2_ASAP7_75t_L       g19182(.A(new_n19414), .B(new_n19438), .Y(new_n19439));
  O2A1O1Ixp33_ASAP7_75t_L   g19183(.A1(new_n19355), .A2(new_n19363), .B(new_n19367), .C(new_n19439), .Y(new_n19440));
  AND3x1_ASAP7_75t_L        g19184(.A(new_n19439), .B(new_n19367), .C(new_n19365), .Y(new_n19441));
  NOR2xp33_ASAP7_75t_L      g19185(.A(new_n19440), .B(new_n19441), .Y(new_n19442));
  INVx1_ASAP7_75t_L         g19186(.A(new_n19442), .Y(new_n19443));
  OR3x1_ASAP7_75t_L         g19187(.A(new_n19408), .B(new_n19410), .C(new_n19443), .Y(new_n19444));
  OAI21xp33_ASAP7_75t_L     g19188(.A1(new_n19410), .A2(new_n19408), .B(new_n19443), .Y(new_n19445));
  AND2x2_ASAP7_75t_L        g19189(.A(new_n19445), .B(new_n19444), .Y(new_n19446));
  INVx1_ASAP7_75t_L         g19190(.A(new_n19446), .Y(new_n19447));
  OAI21xp33_ASAP7_75t_L     g19191(.A1(new_n19388), .A2(new_n19389), .B(new_n19386), .Y(new_n19448));
  NOR2xp33_ASAP7_75t_L      g19192(.A(new_n19448), .B(new_n19447), .Y(new_n19449));
  O2A1O1Ixp33_ASAP7_75t_L   g19193(.A1(new_n19388), .A2(new_n19389), .B(new_n19386), .C(new_n19446), .Y(new_n19450));
  NOR2xp33_ASAP7_75t_L      g19194(.A(new_n19450), .B(new_n19449), .Y(new_n19451));
  INVx1_ASAP7_75t_L         g19195(.A(new_n19451), .Y(new_n19452));
  A2O1A1O1Ixp25_ASAP7_75t_L g19196(.A1(new_n19339), .A2(new_n19342), .B(new_n19397), .C(new_n19394), .D(new_n19452), .Y(new_n19453));
  A2O1A1Ixp33_ASAP7_75t_L   g19197(.A1(new_n19342), .A2(new_n19339), .B(new_n19397), .C(new_n19394), .Y(new_n19454));
  NOR2xp33_ASAP7_75t_L      g19198(.A(new_n19451), .B(new_n19454), .Y(new_n19455));
  NOR2xp33_ASAP7_75t_L      g19199(.A(new_n19453), .B(new_n19455), .Y(\f[117] ));
  AOI22xp33_ASAP7_75t_L     g19200(.A1(new_n9700), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n10027), .Y(new_n19457));
  OAI221xp5_ASAP7_75t_L     g19201(.A1(new_n10024), .A2(new_n10250), .B1(new_n9696), .B2(new_n10855), .C(new_n19457), .Y(new_n19458));
  XNOR2x2_ASAP7_75t_L       g19202(.A(\a[59] ), .B(new_n19458), .Y(new_n19459));
  O2A1O1Ixp33_ASAP7_75t_L   g19203(.A1(new_n11247), .A2(new_n11249), .B(\b[54] ), .C(new_n19421), .Y(new_n19460));
  NOR2xp33_ASAP7_75t_L      g19204(.A(new_n8458), .B(new_n11535), .Y(new_n19461));
  O2A1O1Ixp33_ASAP7_75t_L   g19205(.A1(new_n11247), .A2(new_n11249), .B(\b[55] ), .C(new_n19461), .Y(new_n19462));
  INVx1_ASAP7_75t_L         g19206(.A(new_n19462), .Y(new_n19463));
  A2O1A1Ixp33_ASAP7_75t_L   g19207(.A1(new_n11533), .A2(\b[53] ), .B(new_n19356), .C(new_n7954), .Y(new_n19464));
  A2O1A1O1Ixp25_ASAP7_75t_L g19208(.A1(new_n19415), .A2(new_n19418), .B(new_n19460), .C(new_n19464), .D(new_n19463), .Y(new_n19465));
  INVx1_ASAP7_75t_L         g19209(.A(new_n19465), .Y(new_n19466));
  A2O1A1O1Ixp25_ASAP7_75t_L g19210(.A1(new_n11533), .A2(\b[53] ), .B(new_n19356), .C(new_n7954), .D(new_n19425), .Y(new_n19467));
  A2O1A1Ixp33_ASAP7_75t_L   g19211(.A1(new_n11533), .A2(\b[55] ), .B(new_n19461), .C(new_n19467), .Y(new_n19468));
  NOR2xp33_ASAP7_75t_L      g19212(.A(new_n9920), .B(new_n10630), .Y(new_n19469));
  AOI221xp5_ASAP7_75t_L     g19213(.A1(\b[56] ), .A2(new_n10939), .B1(\b[57] ), .B2(new_n10632), .C(new_n19469), .Y(new_n19470));
  OA211x2_ASAP7_75t_L       g19214(.A1(new_n10629), .A2(new_n9925), .B(\a[62] ), .C(new_n19470), .Y(new_n19471));
  O2A1O1Ixp33_ASAP7_75t_L   g19215(.A1(new_n10629), .A2(new_n9925), .B(new_n19470), .C(\a[62] ), .Y(new_n19472));
  OA211x2_ASAP7_75t_L       g19216(.A1(new_n19472), .A2(new_n19471), .B(new_n19466), .C(new_n19468), .Y(new_n19473));
  AOI211xp5_ASAP7_75t_L     g19217(.A1(new_n19468), .A2(new_n19466), .B(new_n19472), .C(new_n19471), .Y(new_n19474));
  NOR2xp33_ASAP7_75t_L      g19218(.A(new_n19474), .B(new_n19473), .Y(new_n19475));
  INVx1_ASAP7_75t_L         g19219(.A(new_n19475), .Y(new_n19476));
  O2A1O1Ixp33_ASAP7_75t_L   g19220(.A1(new_n19427), .A2(new_n19430), .B(new_n19435), .C(new_n19476), .Y(new_n19477));
  INVx1_ASAP7_75t_L         g19221(.A(new_n19477), .Y(new_n19478));
  OAI211xp5_ASAP7_75t_L     g19222(.A1(new_n19430), .A2(new_n19427), .B(new_n19435), .C(new_n19476), .Y(new_n19479));
  NAND2xp33_ASAP7_75t_L     g19223(.A(new_n19479), .B(new_n19478), .Y(new_n19480));
  NOR2xp33_ASAP7_75t_L      g19224(.A(new_n19459), .B(new_n19480), .Y(new_n19481));
  AND2x2_ASAP7_75t_L        g19225(.A(new_n19459), .B(new_n19480), .Y(new_n19482));
  NOR2xp33_ASAP7_75t_L      g19226(.A(new_n19481), .B(new_n19482), .Y(new_n19483));
  A2O1A1Ixp33_ASAP7_75t_L   g19227(.A1(new_n19438), .A2(new_n19414), .B(new_n19440), .C(new_n19483), .Y(new_n19484));
  NAND2xp33_ASAP7_75t_L     g19228(.A(new_n19414), .B(new_n19438), .Y(new_n19485));
  A2O1A1Ixp33_ASAP7_75t_L   g19229(.A1(new_n19367), .A2(new_n19365), .B(new_n19439), .C(new_n19485), .Y(new_n19486));
  NOR2xp33_ASAP7_75t_L      g19230(.A(new_n19483), .B(new_n19486), .Y(new_n19487));
  INVx1_ASAP7_75t_L         g19231(.A(new_n19487), .Y(new_n19488));
  NAND2xp33_ASAP7_75t_L     g19232(.A(\b[63] ), .B(new_n8835), .Y(new_n19489));
  OAI221xp5_ASAP7_75t_L     g19233(.A1(new_n9418), .A2(new_n11172), .B1(new_n10016), .B2(new_n11500), .C(new_n19489), .Y(new_n19490));
  XNOR2x2_ASAP7_75t_L       g19234(.A(\a[56] ), .B(new_n19490), .Y(new_n19491));
  AND3x1_ASAP7_75t_L        g19235(.A(new_n19488), .B(new_n19491), .C(new_n19484), .Y(new_n19492));
  AOI21xp33_ASAP7_75t_L     g19236(.A1(new_n19488), .A2(new_n19484), .B(new_n19491), .Y(new_n19493));
  NOR2xp33_ASAP7_75t_L      g19237(.A(new_n19493), .B(new_n19492), .Y(new_n19494));
  A2O1A1O1Ixp25_ASAP7_75t_L g19238(.A1(new_n19405), .A2(new_n19404), .B(new_n19407), .C(new_n19444), .D(new_n19494), .Y(new_n19495));
  INVx1_ASAP7_75t_L         g19239(.A(new_n19495), .Y(new_n19496));
  A2O1A1Ixp33_ASAP7_75t_L   g19240(.A1(new_n19405), .A2(new_n19404), .B(new_n19407), .C(new_n19444), .Y(new_n19497));
  OR3x1_ASAP7_75t_L         g19241(.A(new_n19497), .B(new_n19492), .C(new_n19493), .Y(new_n19498));
  AND2x2_ASAP7_75t_L        g19242(.A(new_n19496), .B(new_n19498), .Y(new_n19499));
  A2O1A1Ixp33_ASAP7_75t_L   g19243(.A1(new_n19454), .A2(new_n19451), .B(new_n19449), .C(new_n19499), .Y(new_n19500));
  INVx1_ASAP7_75t_L         g19244(.A(new_n19500), .Y(new_n19501));
  INVx1_ASAP7_75t_L         g19245(.A(new_n19449), .Y(new_n19502));
  A2O1A1Ixp33_ASAP7_75t_L   g19246(.A1(new_n19396), .A2(new_n19394), .B(new_n19452), .C(new_n19502), .Y(new_n19503));
  NOR2xp33_ASAP7_75t_L      g19247(.A(new_n19499), .B(new_n19503), .Y(new_n19504));
  NOR2xp33_ASAP7_75t_L      g19248(.A(new_n19504), .B(new_n19501), .Y(\f[118] ));
  NAND2xp33_ASAP7_75t_L     g19249(.A(\b[57] ), .B(new_n10939), .Y(new_n19506));
  OAI221xp5_ASAP7_75t_L     g19250(.A1(new_n10630), .A2(new_n9947), .B1(new_n10629), .B2(new_n11152), .C(new_n19506), .Y(new_n19507));
  AOI21xp33_ASAP7_75t_L     g19251(.A1(new_n10632), .A2(\b[58] ), .B(new_n19507), .Y(new_n19508));
  NAND2xp33_ASAP7_75t_L     g19252(.A(\a[62] ), .B(new_n19508), .Y(new_n19509));
  A2O1A1Ixp33_ASAP7_75t_L   g19253(.A1(\b[58] ), .A2(new_n10632), .B(new_n19507), .C(new_n10622), .Y(new_n19510));
  NAND2xp33_ASAP7_75t_L     g19254(.A(new_n19510), .B(new_n19509), .Y(new_n19511));
  NOR2xp33_ASAP7_75t_L      g19255(.A(new_n8762), .B(new_n11535), .Y(new_n19512));
  O2A1O1Ixp33_ASAP7_75t_L   g19256(.A1(new_n11247), .A2(new_n11249), .B(\b[56] ), .C(new_n19512), .Y(new_n19513));
  NAND2xp33_ASAP7_75t_L     g19257(.A(new_n19513), .B(new_n19462), .Y(new_n19514));
  A2O1A1Ixp33_ASAP7_75t_L   g19258(.A1(\b[56] ), .A2(new_n11533), .B(new_n19512), .C(new_n19463), .Y(new_n19515));
  AND2x2_ASAP7_75t_L        g19259(.A(new_n19514), .B(new_n19515), .Y(new_n19516));
  INVx1_ASAP7_75t_L         g19260(.A(new_n19516), .Y(new_n19517));
  XNOR2x2_ASAP7_75t_L       g19261(.A(new_n19517), .B(new_n19511), .Y(new_n19518));
  O2A1O1Ixp33_ASAP7_75t_L   g19262(.A1(new_n19472), .A2(new_n19471), .B(new_n19468), .C(new_n19465), .Y(new_n19519));
  NAND2xp33_ASAP7_75t_L     g19263(.A(new_n19519), .B(new_n19518), .Y(new_n19520));
  INVx1_ASAP7_75t_L         g19264(.A(new_n19467), .Y(new_n19521));
  INVx1_ASAP7_75t_L         g19265(.A(new_n19518), .Y(new_n19522));
  A2O1A1Ixp33_ASAP7_75t_L   g19266(.A1(new_n19521), .A2(new_n19462), .B(new_n19473), .C(new_n19522), .Y(new_n19523));
  AOI22xp33_ASAP7_75t_L     g19267(.A1(new_n9700), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n10027), .Y(new_n19524));
  OAI221xp5_ASAP7_75t_L     g19268(.A1(new_n10024), .A2(new_n10847), .B1(new_n9696), .B2(new_n12047), .C(new_n19524), .Y(new_n19525));
  XNOR2x2_ASAP7_75t_L       g19269(.A(\a[59] ), .B(new_n19525), .Y(new_n19526));
  NAND3xp33_ASAP7_75t_L     g19270(.A(new_n19523), .B(new_n19520), .C(new_n19526), .Y(new_n19527));
  AO21x2_ASAP7_75t_L        g19271(.A1(new_n19520), .A2(new_n19523), .B(new_n19526), .Y(new_n19528));
  NAND2xp33_ASAP7_75t_L     g19272(.A(new_n19527), .B(new_n19528), .Y(new_n19529));
  A2O1A1Ixp33_ASAP7_75t_L   g19273(.A1(new_n11471), .A2(\b[61] ), .B(\b[62] ), .C(new_n8828), .Y(new_n19530));
  A2O1A1Ixp33_ASAP7_75t_L   g19274(.A1(new_n19530), .A2(new_n9418), .B(new_n11468), .C(\a[56] ), .Y(new_n19531));
  O2A1O1Ixp33_ASAP7_75t_L   g19275(.A1(new_n10016), .A2(new_n12060), .B(new_n9418), .C(new_n11468), .Y(new_n19532));
  NAND2xp33_ASAP7_75t_L     g19276(.A(new_n8826), .B(new_n19532), .Y(new_n19533));
  AND2x2_ASAP7_75t_L        g19277(.A(new_n19533), .B(new_n19531), .Y(new_n19534));
  O2A1O1Ixp33_ASAP7_75t_L   g19278(.A1(new_n19459), .A2(new_n19480), .B(new_n19478), .C(new_n19534), .Y(new_n19535));
  NOR2xp33_ASAP7_75t_L      g19279(.A(new_n19477), .B(new_n19481), .Y(new_n19536));
  INVx1_ASAP7_75t_L         g19280(.A(new_n19536), .Y(new_n19537));
  INVx1_ASAP7_75t_L         g19281(.A(new_n19534), .Y(new_n19538));
  NOR2xp33_ASAP7_75t_L      g19282(.A(new_n19538), .B(new_n19537), .Y(new_n19539));
  NOR2xp33_ASAP7_75t_L      g19283(.A(new_n19535), .B(new_n19539), .Y(new_n19540));
  INVx1_ASAP7_75t_L         g19284(.A(new_n19540), .Y(new_n19541));
  NAND2xp33_ASAP7_75t_L     g19285(.A(new_n19529), .B(new_n19541), .Y(new_n19542));
  NOR2xp33_ASAP7_75t_L      g19286(.A(new_n19529), .B(new_n19541), .Y(new_n19543));
  INVx1_ASAP7_75t_L         g19287(.A(new_n19543), .Y(new_n19544));
  NAND2xp33_ASAP7_75t_L     g19288(.A(new_n19542), .B(new_n19544), .Y(new_n19545));
  OAI21xp33_ASAP7_75t_L     g19289(.A1(new_n19491), .A2(new_n19487), .B(new_n19484), .Y(new_n19546));
  NOR2xp33_ASAP7_75t_L      g19290(.A(new_n19546), .B(new_n19545), .Y(new_n19547));
  NAND2xp33_ASAP7_75t_L     g19291(.A(new_n19546), .B(new_n19545), .Y(new_n19548));
  INVx1_ASAP7_75t_L         g19292(.A(new_n19548), .Y(new_n19549));
  NOR2xp33_ASAP7_75t_L      g19293(.A(new_n19547), .B(new_n19549), .Y(new_n19550));
  A2O1A1Ixp33_ASAP7_75t_L   g19294(.A1(new_n19503), .A2(new_n19499), .B(new_n19495), .C(new_n19550), .Y(new_n19551));
  INVx1_ASAP7_75t_L         g19295(.A(new_n19551), .Y(new_n19552));
  INVx1_ASAP7_75t_L         g19296(.A(new_n19408), .Y(new_n19553));
  A2O1A1Ixp33_ASAP7_75t_L   g19297(.A1(new_n19444), .A2(new_n19553), .B(new_n19494), .C(new_n19500), .Y(new_n19554));
  NOR2xp33_ASAP7_75t_L      g19298(.A(new_n19550), .B(new_n19554), .Y(new_n19555));
  NOR2xp33_ASAP7_75t_L      g19299(.A(new_n19552), .B(new_n19555), .Y(\f[119] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19300(.A1(\b[56] ), .A2(new_n11533), .B(new_n19512), .C(new_n19462), .Y(new_n19557));
  A2O1A1Ixp33_ASAP7_75t_L   g19301(.A1(new_n19509), .A2(new_n19510), .B(new_n19516), .C(new_n19557), .Y(new_n19558));
  NOR2xp33_ASAP7_75t_L      g19302(.A(new_n9323), .B(new_n11535), .Y(new_n19559));
  O2A1O1Ixp33_ASAP7_75t_L   g19303(.A1(new_n11247), .A2(new_n11249), .B(\b[57] ), .C(new_n19559), .Y(new_n19560));
  INVx1_ASAP7_75t_L         g19304(.A(new_n19560), .Y(new_n19561));
  NOR2xp33_ASAP7_75t_L      g19305(.A(\a[56] ), .B(new_n19561), .Y(new_n19562));
  INVx1_ASAP7_75t_L         g19306(.A(new_n19562), .Y(new_n19563));
  A2O1A1Ixp33_ASAP7_75t_L   g19307(.A1(new_n11533), .A2(\b[57] ), .B(new_n19559), .C(\a[56] ), .Y(new_n19564));
  NAND2xp33_ASAP7_75t_L     g19308(.A(new_n19564), .B(new_n19563), .Y(new_n19565));
  A2O1A1Ixp33_ASAP7_75t_L   g19309(.A1(new_n11533), .A2(\b[55] ), .B(new_n19461), .C(new_n19565), .Y(new_n19566));
  NAND3xp33_ASAP7_75t_L     g19310(.A(new_n19563), .B(new_n19462), .C(new_n19564), .Y(new_n19567));
  AND2x2_ASAP7_75t_L        g19311(.A(new_n19567), .B(new_n19566), .Y(new_n19568));
  NOR2xp33_ASAP7_75t_L      g19312(.A(new_n19568), .B(new_n19558), .Y(new_n19569));
  INVx1_ASAP7_75t_L         g19313(.A(new_n19568), .Y(new_n19570));
  A2O1A1O1Ixp25_ASAP7_75t_L g19314(.A1(new_n19510), .A2(new_n19509), .B(new_n19516), .C(new_n19557), .D(new_n19570), .Y(new_n19571));
  NOR2xp33_ASAP7_75t_L      g19315(.A(new_n19571), .B(new_n19569), .Y(new_n19572));
  AOI22xp33_ASAP7_75t_L     g19316(.A1(\b[58] ), .A2(new_n10939), .B1(\b[60] ), .B2(new_n10938), .Y(new_n19573));
  OAI221xp5_ASAP7_75t_L     g19317(.A1(new_n10937), .A2(new_n9947), .B1(new_n10629), .B2(new_n11446), .C(new_n19573), .Y(new_n19574));
  XNOR2x2_ASAP7_75t_L       g19318(.A(\a[62] ), .B(new_n19574), .Y(new_n19575));
  XNOR2x2_ASAP7_75t_L       g19319(.A(new_n19575), .B(new_n19572), .Y(new_n19576));
  AOI22xp33_ASAP7_75t_L     g19320(.A1(new_n9700), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n10027), .Y(new_n19577));
  A2O1A1Ixp33_ASAP7_75t_L   g19321(.A1(new_n11470), .A2(new_n11473), .B(new_n9696), .C(new_n19577), .Y(new_n19578));
  AOI21xp33_ASAP7_75t_L     g19322(.A1(new_n9703), .A2(\b[62] ), .B(new_n19578), .Y(new_n19579));
  NAND2xp33_ASAP7_75t_L     g19323(.A(\a[59] ), .B(new_n19579), .Y(new_n19580));
  A2O1A1Ixp33_ASAP7_75t_L   g19324(.A1(\b[62] ), .A2(new_n9703), .B(new_n19578), .C(new_n9693), .Y(new_n19581));
  NAND2xp33_ASAP7_75t_L     g19325(.A(new_n19520), .B(new_n19527), .Y(new_n19582));
  AOI21xp33_ASAP7_75t_L     g19326(.A1(new_n19581), .A2(new_n19580), .B(new_n19582), .Y(new_n19583));
  INVx1_ASAP7_75t_L         g19327(.A(new_n19583), .Y(new_n19584));
  NAND3xp33_ASAP7_75t_L     g19328(.A(new_n19582), .B(new_n19581), .C(new_n19580), .Y(new_n19585));
  NAND3xp33_ASAP7_75t_L     g19329(.A(new_n19584), .B(new_n19576), .C(new_n19585), .Y(new_n19586));
  AO21x2_ASAP7_75t_L        g19330(.A1(new_n19585), .A2(new_n19584), .B(new_n19576), .Y(new_n19587));
  AND2x2_ASAP7_75t_L        g19331(.A(new_n19586), .B(new_n19587), .Y(new_n19588));
  O2A1O1Ixp33_ASAP7_75t_L   g19332(.A1(new_n19537), .A2(new_n19538), .B(new_n19544), .C(new_n19588), .Y(new_n19589));
  INVx1_ASAP7_75t_L         g19333(.A(new_n19588), .Y(new_n19590));
  NOR2xp33_ASAP7_75t_L      g19334(.A(new_n19539), .B(new_n19543), .Y(new_n19591));
  INVx1_ASAP7_75t_L         g19335(.A(new_n19591), .Y(new_n19592));
  NOR2xp33_ASAP7_75t_L      g19336(.A(new_n19590), .B(new_n19592), .Y(new_n19593));
  NOR2xp33_ASAP7_75t_L      g19337(.A(new_n19589), .B(new_n19593), .Y(new_n19594));
  INVx1_ASAP7_75t_L         g19338(.A(new_n19594), .Y(new_n19595));
  A2O1A1O1Ixp25_ASAP7_75t_L g19339(.A1(new_n19496), .A2(new_n19500), .B(new_n19547), .C(new_n19548), .D(new_n19595), .Y(new_n19596));
  A2O1A1Ixp33_ASAP7_75t_L   g19340(.A1(new_n19500), .A2(new_n19496), .B(new_n19547), .C(new_n19548), .Y(new_n19597));
  NOR2xp33_ASAP7_75t_L      g19341(.A(new_n19594), .B(new_n19597), .Y(new_n19598));
  NOR2xp33_ASAP7_75t_L      g19342(.A(new_n19596), .B(new_n19598), .Y(\f[120] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19343(.A1(new_n19581), .A2(new_n19580), .B(new_n19582), .C(new_n19586), .Y(new_n19600));
  INVx1_ASAP7_75t_L         g19344(.A(new_n19600), .Y(new_n19601));
  INVx1_ASAP7_75t_L         g19345(.A(new_n19575), .Y(new_n19602));
  NOR2xp33_ASAP7_75t_L      g19346(.A(new_n9620), .B(new_n11535), .Y(new_n19603));
  INVx1_ASAP7_75t_L         g19347(.A(new_n19566), .Y(new_n19604));
  A2O1A1O1Ixp25_ASAP7_75t_L g19348(.A1(new_n11533), .A2(\b[57] ), .B(new_n19559), .C(new_n8826), .D(new_n19604), .Y(new_n19605));
  A2O1A1Ixp33_ASAP7_75t_L   g19349(.A1(new_n11533), .A2(\b[58] ), .B(new_n19603), .C(new_n19605), .Y(new_n19606));
  O2A1O1Ixp33_ASAP7_75t_L   g19350(.A1(new_n11247), .A2(new_n11249), .B(\b[58] ), .C(new_n19603), .Y(new_n19607));
  INVx1_ASAP7_75t_L         g19351(.A(new_n19607), .Y(new_n19608));
  A2O1A1Ixp33_ASAP7_75t_L   g19352(.A1(new_n11533), .A2(\b[57] ), .B(new_n19559), .C(new_n8826), .Y(new_n19609));
  A2O1A1O1Ixp25_ASAP7_75t_L g19353(.A1(new_n19564), .A2(new_n19563), .B(new_n19462), .C(new_n19609), .D(new_n19608), .Y(new_n19610));
  INVx1_ASAP7_75t_L         g19354(.A(new_n19610), .Y(new_n19611));
  NAND2xp33_ASAP7_75t_L     g19355(.A(new_n19611), .B(new_n19606), .Y(new_n19612));
  INVx1_ASAP7_75t_L         g19356(.A(new_n19612), .Y(new_n19613));
  NAND2xp33_ASAP7_75t_L     g19357(.A(\b[60] ), .B(new_n10632), .Y(new_n19614));
  OAI221xp5_ASAP7_75t_L     g19358(.A1(new_n10630), .A2(new_n10847), .B1(new_n9947), .B2(new_n11257), .C(new_n19614), .Y(new_n19615));
  AOI21xp33_ASAP7_75t_L     g19359(.A1(new_n11759), .A2(new_n11256), .B(new_n19615), .Y(new_n19616));
  NAND2xp33_ASAP7_75t_L     g19360(.A(\a[62] ), .B(new_n19616), .Y(new_n19617));
  A2O1A1Ixp33_ASAP7_75t_L   g19361(.A1(new_n11759), .A2(new_n11256), .B(new_n19615), .C(new_n10622), .Y(new_n19618));
  NAND2xp33_ASAP7_75t_L     g19362(.A(new_n19618), .B(new_n19617), .Y(new_n19619));
  NAND2xp33_ASAP7_75t_L     g19363(.A(new_n19613), .B(new_n19619), .Y(new_n19620));
  INVx1_ASAP7_75t_L         g19364(.A(new_n19620), .Y(new_n19621));
  NOR2xp33_ASAP7_75t_L      g19365(.A(new_n19613), .B(new_n19619), .Y(new_n19622));
  NOR2xp33_ASAP7_75t_L      g19366(.A(new_n19622), .B(new_n19621), .Y(new_n19623));
  A2O1A1Ixp33_ASAP7_75t_L   g19367(.A1(new_n19572), .A2(new_n19602), .B(new_n19571), .C(new_n19623), .Y(new_n19624));
  AO21x2_ASAP7_75t_L        g19368(.A1(new_n19602), .A2(new_n19572), .B(new_n19571), .Y(new_n19625));
  NOR2xp33_ASAP7_75t_L      g19369(.A(new_n19623), .B(new_n19625), .Y(new_n19626));
  INVx1_ASAP7_75t_L         g19370(.A(new_n19626), .Y(new_n19627));
  NAND2xp33_ASAP7_75t_L     g19371(.A(new_n19624), .B(new_n19627), .Y(new_n19628));
  AOI22xp33_ASAP7_75t_L     g19372(.A1(new_n9703), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n10027), .Y(new_n19629));
  OAI211xp5_ASAP7_75t_L     g19373(.A1(new_n9696), .A2(new_n11500), .B(\a[59] ), .C(new_n19629), .Y(new_n19630));
  INVx1_ASAP7_75t_L         g19374(.A(new_n19630), .Y(new_n19631));
  O2A1O1Ixp33_ASAP7_75t_L   g19375(.A1(new_n9696), .A2(new_n11500), .B(new_n19629), .C(\a[59] ), .Y(new_n19632));
  NOR2xp33_ASAP7_75t_L      g19376(.A(new_n19632), .B(new_n19631), .Y(new_n19633));
  XNOR2x2_ASAP7_75t_L       g19377(.A(new_n19633), .B(new_n19628), .Y(new_n19634));
  NAND2xp33_ASAP7_75t_L     g19378(.A(new_n19634), .B(new_n19601), .Y(new_n19635));
  A2O1A1O1Ixp25_ASAP7_75t_L g19379(.A1(new_n19581), .A2(new_n19580), .B(new_n19582), .C(new_n19586), .D(new_n19634), .Y(new_n19636));
  INVx1_ASAP7_75t_L         g19380(.A(new_n19636), .Y(new_n19637));
  AND2x2_ASAP7_75t_L        g19381(.A(new_n19637), .B(new_n19635), .Y(new_n19638));
  A2O1A1Ixp33_ASAP7_75t_L   g19382(.A1(new_n19597), .A2(new_n19594), .B(new_n19593), .C(new_n19638), .Y(new_n19639));
  INVx1_ASAP7_75t_L         g19383(.A(new_n19639), .Y(new_n19640));
  INVx1_ASAP7_75t_L         g19384(.A(new_n19593), .Y(new_n19641));
  A2O1A1Ixp33_ASAP7_75t_L   g19385(.A1(new_n19551), .A2(new_n19548), .B(new_n19595), .C(new_n19641), .Y(new_n19642));
  NOR2xp33_ASAP7_75t_L      g19386(.A(new_n19638), .B(new_n19642), .Y(new_n19643));
  NOR2xp33_ASAP7_75t_L      g19387(.A(new_n19643), .B(new_n19640), .Y(\f[121] ));
  AOI22xp33_ASAP7_75t_L     g19388(.A1(\b[60] ), .A2(new_n10939), .B1(\b[62] ), .B2(new_n10938), .Y(new_n19645));
  OAI221xp5_ASAP7_75t_L     g19389(.A1(new_n10937), .A2(new_n10847), .B1(new_n10629), .B2(new_n12047), .C(new_n19645), .Y(new_n19646));
  XNOR2x2_ASAP7_75t_L       g19390(.A(\a[62] ), .B(new_n19646), .Y(new_n19647));
  A2O1A1O1Ixp25_ASAP7_75t_L g19391(.A1(new_n9697), .A2(new_n12061), .B(new_n10027), .C(\b[63] ), .D(new_n9693), .Y(new_n19648));
  A2O1A1Ixp33_ASAP7_75t_L   g19392(.A1(new_n12061), .A2(new_n9697), .B(new_n10027), .C(\b[63] ), .Y(new_n19649));
  NOR2xp33_ASAP7_75t_L      g19393(.A(\a[59] ), .B(new_n19649), .Y(new_n19650));
  NOR2xp33_ASAP7_75t_L      g19394(.A(new_n19648), .B(new_n19650), .Y(new_n19651));
  NOR2xp33_ASAP7_75t_L      g19395(.A(new_n19651), .B(new_n19647), .Y(new_n19652));
  NAND2xp33_ASAP7_75t_L     g19396(.A(new_n19651), .B(new_n19647), .Y(new_n19653));
  INVx1_ASAP7_75t_L         g19397(.A(new_n19653), .Y(new_n19654));
  NOR2xp33_ASAP7_75t_L      g19398(.A(new_n19652), .B(new_n19654), .Y(new_n19655));
  NOR2xp33_ASAP7_75t_L      g19399(.A(new_n9920), .B(new_n11535), .Y(new_n19656));
  A2O1A1Ixp33_ASAP7_75t_L   g19400(.A1(\b[59] ), .A2(new_n11533), .B(new_n19656), .C(new_n19607), .Y(new_n19657));
  O2A1O1Ixp33_ASAP7_75t_L   g19401(.A1(new_n11247), .A2(new_n11249), .B(\b[59] ), .C(new_n19656), .Y(new_n19658));
  A2O1A1Ixp33_ASAP7_75t_L   g19402(.A1(new_n11533), .A2(\b[58] ), .B(new_n19603), .C(new_n19658), .Y(new_n19659));
  AND2x2_ASAP7_75t_L        g19403(.A(new_n19657), .B(new_n19659), .Y(new_n19660));
  AND3x1_ASAP7_75t_L        g19404(.A(new_n19620), .B(new_n19660), .C(new_n19611), .Y(new_n19661));
  A2O1A1O1Ixp25_ASAP7_75t_L g19405(.A1(new_n19618), .A2(new_n19617), .B(new_n19612), .C(new_n19611), .D(new_n19660), .Y(new_n19662));
  NOR2xp33_ASAP7_75t_L      g19406(.A(new_n19662), .B(new_n19661), .Y(new_n19663));
  XOR2x2_ASAP7_75t_L        g19407(.A(new_n19663), .B(new_n19655), .Y(new_n19664));
  O2A1O1Ixp33_ASAP7_75t_L   g19408(.A1(new_n19626), .A2(new_n19633), .B(new_n19624), .C(new_n19664), .Y(new_n19665));
  INVx1_ASAP7_75t_L         g19409(.A(new_n19665), .Y(new_n19666));
  OAI211xp5_ASAP7_75t_L     g19410(.A1(new_n19626), .A2(new_n19633), .B(new_n19664), .C(new_n19624), .Y(new_n19667));
  AND2x2_ASAP7_75t_L        g19411(.A(new_n19667), .B(new_n19666), .Y(new_n19668));
  A2O1A1Ixp33_ASAP7_75t_L   g19412(.A1(new_n19642), .A2(new_n19638), .B(new_n19636), .C(new_n19668), .Y(new_n19669));
  A2O1A1O1Ixp25_ASAP7_75t_L g19413(.A1(new_n19594), .A2(new_n19597), .B(new_n19593), .C(new_n19638), .D(new_n19636), .Y(new_n19670));
  INVx1_ASAP7_75t_L         g19414(.A(new_n19668), .Y(new_n19671));
  NAND2xp33_ASAP7_75t_L     g19415(.A(new_n19671), .B(new_n19670), .Y(new_n19672));
  AND2x2_ASAP7_75t_L        g19416(.A(new_n19669), .B(new_n19672), .Y(\f[122] ));
  INVx1_ASAP7_75t_L         g19417(.A(new_n19652), .Y(new_n19674));
  INVx1_ASAP7_75t_L         g19418(.A(new_n19658), .Y(new_n19675));
  A2O1A1Ixp33_ASAP7_75t_L   g19419(.A1(new_n11533), .A2(\b[59] ), .B(new_n19656), .C(\a[59] ), .Y(new_n19676));
  NOR2xp33_ASAP7_75t_L      g19420(.A(\a[59] ), .B(new_n19675), .Y(new_n19677));
  INVx1_ASAP7_75t_L         g19421(.A(new_n19677), .Y(new_n19678));
  NOR2xp33_ASAP7_75t_L      g19422(.A(new_n9947), .B(new_n11535), .Y(new_n19679));
  O2A1O1Ixp33_ASAP7_75t_L   g19423(.A1(new_n11247), .A2(new_n11249), .B(\b[60] ), .C(new_n19679), .Y(new_n19680));
  NAND3xp33_ASAP7_75t_L     g19424(.A(new_n19678), .B(new_n19676), .C(new_n19680), .Y(new_n19681));
  NAND2xp33_ASAP7_75t_L     g19425(.A(new_n19676), .B(new_n19678), .Y(new_n19682));
  A2O1A1Ixp33_ASAP7_75t_L   g19426(.A1(\b[60] ), .A2(new_n11533), .B(new_n19679), .C(new_n19682), .Y(new_n19683));
  AND2x2_ASAP7_75t_L        g19427(.A(new_n19681), .B(new_n19683), .Y(new_n19684));
  AOI22xp33_ASAP7_75t_L     g19428(.A1(\b[61] ), .A2(new_n10939), .B1(\b[63] ), .B2(new_n10938), .Y(new_n19685));
  A2O1A1Ixp33_ASAP7_75t_L   g19429(.A1(new_n11470), .A2(new_n11473), .B(new_n10629), .C(new_n19685), .Y(new_n19686));
  AOI21xp33_ASAP7_75t_L     g19430(.A1(new_n10632), .A2(\b[62] ), .B(new_n19686), .Y(new_n19687));
  NAND2xp33_ASAP7_75t_L     g19431(.A(\a[62] ), .B(new_n19687), .Y(new_n19688));
  A2O1A1Ixp33_ASAP7_75t_L   g19432(.A1(\b[62] ), .A2(new_n10632), .B(new_n19686), .C(new_n10622), .Y(new_n19689));
  NAND2xp33_ASAP7_75t_L     g19433(.A(new_n19689), .B(new_n19688), .Y(new_n19690));
  XNOR2x2_ASAP7_75t_L       g19434(.A(new_n19684), .B(new_n19690), .Y(new_n19691));
  A2O1A1Ixp33_ASAP7_75t_L   g19435(.A1(new_n19619), .A2(new_n19613), .B(new_n19610), .C(new_n19657), .Y(new_n19692));
  O2A1O1Ixp33_ASAP7_75t_L   g19436(.A1(new_n19675), .A2(new_n19607), .B(new_n19692), .C(new_n19691), .Y(new_n19693));
  AND3x1_ASAP7_75t_L        g19437(.A(new_n19691), .B(new_n19692), .C(new_n19659), .Y(new_n19694));
  NOR2xp33_ASAP7_75t_L      g19438(.A(new_n19693), .B(new_n19694), .Y(new_n19695));
  INVx1_ASAP7_75t_L         g19439(.A(new_n19695), .Y(new_n19696));
  O2A1O1Ixp33_ASAP7_75t_L   g19440(.A1(new_n19654), .A2(new_n19663), .B(new_n19674), .C(new_n19696), .Y(new_n19697));
  INVx1_ASAP7_75t_L         g19441(.A(new_n19697), .Y(new_n19698));
  O2A1O1Ixp33_ASAP7_75t_L   g19442(.A1(new_n19662), .A2(new_n19661), .B(new_n19653), .C(new_n19652), .Y(new_n19699));
  NAND2xp33_ASAP7_75t_L     g19443(.A(new_n19699), .B(new_n19696), .Y(new_n19700));
  AND2x2_ASAP7_75t_L        g19444(.A(new_n19700), .B(new_n19698), .Y(new_n19701));
  INVx1_ASAP7_75t_L         g19445(.A(new_n19701), .Y(new_n19702));
  A2O1A1O1Ixp25_ASAP7_75t_L g19446(.A1(new_n19637), .A2(new_n19639), .B(new_n19671), .C(new_n19666), .D(new_n19702), .Y(new_n19703));
  A2O1A1Ixp33_ASAP7_75t_L   g19447(.A1(new_n19639), .A2(new_n19637), .B(new_n19671), .C(new_n19666), .Y(new_n19704));
  NOR2xp33_ASAP7_75t_L      g19448(.A(new_n19701), .B(new_n19704), .Y(new_n19705));
  NOR2xp33_ASAP7_75t_L      g19449(.A(new_n19703), .B(new_n19705), .Y(\f[123] ));
  INVx1_ASAP7_75t_L         g19450(.A(new_n19684), .Y(new_n19707));
  INVx1_ASAP7_75t_L         g19451(.A(new_n19691), .Y(new_n19708));
  A2O1A1O1Ixp25_ASAP7_75t_L g19452(.A1(new_n19561), .A2(new_n8826), .B(new_n19604), .C(new_n19607), .D(new_n19621), .Y(new_n19709));
  A2O1A1O1Ixp25_ASAP7_75t_L g19453(.A1(\b[59] ), .A2(new_n11533), .B(new_n19656), .C(new_n19607), .D(new_n19709), .Y(new_n19710));
  A2O1A1Ixp33_ASAP7_75t_L   g19454(.A1(new_n19608), .A2(new_n19658), .B(new_n19710), .C(new_n19708), .Y(new_n19711));
  NOR2xp33_ASAP7_75t_L      g19455(.A(new_n10250), .B(new_n11535), .Y(new_n19712));
  O2A1O1Ixp33_ASAP7_75t_L   g19456(.A1(new_n11247), .A2(new_n11249), .B(\b[61] ), .C(new_n19712), .Y(new_n19713));
  INVx1_ASAP7_75t_L         g19457(.A(new_n19713), .Y(new_n19714));
  A2O1A1Ixp33_ASAP7_75t_L   g19458(.A1(new_n11533), .A2(\b[59] ), .B(new_n19656), .C(new_n9693), .Y(new_n19715));
  A2O1A1O1Ixp25_ASAP7_75t_L g19459(.A1(new_n19676), .A2(new_n19678), .B(new_n19680), .C(new_n19715), .D(new_n19714), .Y(new_n19716));
  INVx1_ASAP7_75t_L         g19460(.A(new_n19716), .Y(new_n19717));
  INVx1_ASAP7_75t_L         g19461(.A(new_n19683), .Y(new_n19718));
  A2O1A1O1Ixp25_ASAP7_75t_L g19462(.A1(new_n11533), .A2(\b[59] ), .B(new_n19656), .C(new_n9693), .D(new_n19718), .Y(new_n19719));
  A2O1A1Ixp33_ASAP7_75t_L   g19463(.A1(new_n11533), .A2(\b[61] ), .B(new_n19712), .C(new_n19719), .Y(new_n19720));
  NAND2xp33_ASAP7_75t_L     g19464(.A(new_n19717), .B(new_n19720), .Y(new_n19721));
  OAI22xp33_ASAP7_75t_L     g19465(.A1(new_n11500), .A2(new_n10629), .B1(new_n11172), .B2(new_n11257), .Y(new_n19722));
  AOI21xp33_ASAP7_75t_L     g19466(.A1(new_n10632), .A2(\b[63] ), .B(new_n19722), .Y(new_n19723));
  NAND2xp33_ASAP7_75t_L     g19467(.A(\a[62] ), .B(new_n19723), .Y(new_n19724));
  A2O1A1Ixp33_ASAP7_75t_L   g19468(.A1(\b[63] ), .A2(new_n10632), .B(new_n19722), .C(new_n10622), .Y(new_n19725));
  AND2x2_ASAP7_75t_L        g19469(.A(new_n19725), .B(new_n19724), .Y(new_n19726));
  NOR2xp33_ASAP7_75t_L      g19470(.A(new_n19721), .B(new_n19726), .Y(new_n19727));
  AND3x1_ASAP7_75t_L        g19471(.A(new_n19724), .B(new_n19725), .C(new_n19721), .Y(new_n19728));
  NOR2xp33_ASAP7_75t_L      g19472(.A(new_n19728), .B(new_n19727), .Y(new_n19729));
  INVx1_ASAP7_75t_L         g19473(.A(new_n19729), .Y(new_n19730));
  A2O1A1O1Ixp25_ASAP7_75t_L g19474(.A1(new_n19688), .A2(new_n19689), .B(new_n19707), .C(new_n19711), .D(new_n19730), .Y(new_n19731));
  INVx1_ASAP7_75t_L         g19475(.A(new_n19731), .Y(new_n19732));
  A2O1A1Ixp33_ASAP7_75t_L   g19476(.A1(new_n19688), .A2(new_n19689), .B(new_n19707), .C(new_n19711), .Y(new_n19733));
  INVx1_ASAP7_75t_L         g19477(.A(new_n19733), .Y(new_n19734));
  NAND2xp33_ASAP7_75t_L     g19478(.A(new_n19730), .B(new_n19734), .Y(new_n19735));
  AND2x2_ASAP7_75t_L        g19479(.A(new_n19732), .B(new_n19735), .Y(new_n19736));
  A2O1A1Ixp33_ASAP7_75t_L   g19480(.A1(new_n19704), .A2(new_n19701), .B(new_n19697), .C(new_n19736), .Y(new_n19737));
  A2O1A1Ixp33_ASAP7_75t_L   g19481(.A1(new_n19586), .A2(new_n19584), .B(new_n19634), .C(new_n19639), .Y(new_n19738));
  A2O1A1O1Ixp25_ASAP7_75t_L g19482(.A1(new_n19667), .A2(new_n19738), .B(new_n19665), .C(new_n19701), .D(new_n19697), .Y(new_n19739));
  INVx1_ASAP7_75t_L         g19483(.A(new_n19736), .Y(new_n19740));
  NAND2xp33_ASAP7_75t_L     g19484(.A(new_n19740), .B(new_n19739), .Y(new_n19741));
  AND2x2_ASAP7_75t_L        g19485(.A(new_n19737), .B(new_n19741), .Y(\f[124] ));
  NAND2xp33_ASAP7_75t_L     g19486(.A(\b[61] ), .B(new_n11534), .Y(new_n19743));
  O2A1O1Ixp33_ASAP7_75t_L   g19487(.A1(new_n11253), .A2(new_n11172), .B(new_n19743), .C(new_n19714), .Y(new_n19744));
  INVx1_ASAP7_75t_L         g19488(.A(new_n19712), .Y(new_n19745));
  A2O1A1Ixp33_ASAP7_75t_L   g19489(.A1(new_n14788), .A2(new_n14789), .B(new_n11172), .C(new_n19743), .Y(new_n19746));
  O2A1O1Ixp33_ASAP7_75t_L   g19490(.A1(new_n10847), .A2(new_n11253), .B(new_n19745), .C(new_n19746), .Y(new_n19747));
  NOR2xp33_ASAP7_75t_L      g19491(.A(new_n19747), .B(new_n19744), .Y(new_n19748));
  A2O1A1O1Ixp25_ASAP7_75t_L g19492(.A1(new_n11256), .A2(new_n12061), .B(new_n10939), .C(\b[63] ), .D(new_n10622), .Y(new_n19749));
  A2O1A1Ixp33_ASAP7_75t_L   g19493(.A1(new_n12061), .A2(new_n11256), .B(new_n10939), .C(\b[63] ), .Y(new_n19750));
  NOR2xp33_ASAP7_75t_L      g19494(.A(\a[62] ), .B(new_n19750), .Y(new_n19751));
  OA21x2_ASAP7_75t_L        g19495(.A1(new_n19749), .A2(new_n19751), .B(new_n19748), .Y(new_n19752));
  NOR3xp33_ASAP7_75t_L      g19496(.A(new_n19751), .B(new_n19749), .C(new_n19748), .Y(new_n19753));
  NOR2xp33_ASAP7_75t_L      g19497(.A(new_n19753), .B(new_n19752), .Y(new_n19754));
  INVx1_ASAP7_75t_L         g19498(.A(new_n19754), .Y(new_n19755));
  A2O1A1O1Ixp25_ASAP7_75t_L g19499(.A1(new_n19725), .A2(new_n19724), .B(new_n19721), .C(new_n19717), .D(new_n19755), .Y(new_n19756));
  INVx1_ASAP7_75t_L         g19500(.A(new_n19756), .Y(new_n19757));
  A2O1A1O1Ixp25_ASAP7_75t_L g19501(.A1(new_n19675), .A2(new_n9693), .B(new_n19718), .C(new_n19713), .D(new_n19727), .Y(new_n19758));
  NAND2xp33_ASAP7_75t_L     g19502(.A(new_n19755), .B(new_n19758), .Y(new_n19759));
  AND2x2_ASAP7_75t_L        g19503(.A(new_n19757), .B(new_n19759), .Y(new_n19760));
  INVx1_ASAP7_75t_L         g19504(.A(new_n19760), .Y(new_n19761));
  O2A1O1Ixp33_ASAP7_75t_L   g19505(.A1(new_n19734), .A2(new_n19730), .B(new_n19737), .C(new_n19761), .Y(new_n19762));
  A2O1A1Ixp33_ASAP7_75t_L   g19506(.A1(new_n19669), .A2(new_n19666), .B(new_n19702), .C(new_n19698), .Y(new_n19763));
  AOI211xp5_ASAP7_75t_L     g19507(.A1(new_n19763), .A2(new_n19736), .B(new_n19760), .C(new_n19731), .Y(new_n19764));
  NOR2xp33_ASAP7_75t_L      g19508(.A(new_n19764), .B(new_n19762), .Y(\f[125] ));
  NOR2xp33_ASAP7_75t_L      g19509(.A(new_n11248), .B(new_n11468), .Y(new_n19766));
  INVx1_ASAP7_75t_L         g19510(.A(new_n19766), .Y(new_n19767));
  NOR3xp33_ASAP7_75t_L      g19511(.A(new_n10622), .B(new_n11248), .C(new_n11172), .Y(new_n19768));
  O2A1O1Ixp33_ASAP7_75t_L   g19512(.A1(new_n10622), .A2(\b[63] ), .B(new_n19767), .C(new_n19768), .Y(new_n19769));
  O2A1O1Ixp33_ASAP7_75t_L   g19513(.A1(new_n10847), .A2(new_n11253), .B(new_n19745), .C(new_n19769), .Y(new_n19770));
  INVx1_ASAP7_75t_L         g19514(.A(new_n19770), .Y(new_n19771));
  NAND2xp33_ASAP7_75t_L     g19515(.A(new_n19769), .B(new_n19713), .Y(new_n19772));
  NAND2xp33_ASAP7_75t_L     g19516(.A(new_n19772), .B(new_n19771), .Y(new_n19773));
  INVx1_ASAP7_75t_L         g19517(.A(new_n19773), .Y(new_n19774));
  A2O1A1Ixp33_ASAP7_75t_L   g19518(.A1(new_n19746), .A2(new_n19713), .B(new_n19752), .C(new_n19774), .Y(new_n19775));
  O2A1O1Ixp33_ASAP7_75t_L   g19519(.A1(new_n19749), .A2(new_n19751), .B(new_n19748), .C(new_n19744), .Y(new_n19776));
  NAND2xp33_ASAP7_75t_L     g19520(.A(new_n19773), .B(new_n19776), .Y(new_n19777));
  AND2x2_ASAP7_75t_L        g19521(.A(new_n19777), .B(new_n19775), .Y(new_n19778));
  INVx1_ASAP7_75t_L         g19522(.A(new_n19778), .Y(new_n19779));
  A2O1A1O1Ixp25_ASAP7_75t_L g19523(.A1(new_n19732), .A2(new_n19737), .B(new_n19761), .C(new_n19757), .D(new_n19779), .Y(new_n19780));
  A2O1A1Ixp33_ASAP7_75t_L   g19524(.A1(new_n19737), .A2(new_n19732), .B(new_n19761), .C(new_n19757), .Y(new_n19781));
  NOR2xp33_ASAP7_75t_L      g19525(.A(new_n19778), .B(new_n19781), .Y(new_n19782));
  NOR2xp33_ASAP7_75t_L      g19526(.A(new_n19780), .B(new_n19782), .Y(\f[126] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g19527(.A1(new_n19736), .A2(new_n19763), .B(new_n19731), .C(new_n19760), .D(new_n19756), .Y(new_n19784));
  INVx1_ASAP7_75t_L         g19528(.A(new_n19769), .Y(new_n19785));
  A2O1A1O1Ixp25_ASAP7_75t_L g19529(.A1(\b[61] ), .A2(new_n11533), .B(new_n19712), .C(new_n19785), .D(new_n19767), .Y(new_n19786));
  NOR2xp33_ASAP7_75t_L      g19530(.A(new_n19766), .B(new_n19771), .Y(new_n19787));
  NOR2xp33_ASAP7_75t_L      g19531(.A(new_n19786), .B(new_n19787), .Y(new_n19788));
  OAI211xp5_ASAP7_75t_L     g19532(.A1(new_n19779), .A2(new_n19784), .B(new_n19775), .C(new_n19788), .Y(new_n19789));
  INVx1_ASAP7_75t_L         g19533(.A(new_n19775), .Y(new_n19790));
  INVx1_ASAP7_75t_L         g19534(.A(new_n19788), .Y(new_n19791));
  A2O1A1Ixp33_ASAP7_75t_L   g19535(.A1(new_n19781), .A2(new_n19778), .B(new_n19790), .C(new_n19791), .Y(new_n19792));
  NAND2xp33_ASAP7_75t_L     g19536(.A(new_n19789), .B(new_n19792), .Y(\f[127] ));
endmodule


