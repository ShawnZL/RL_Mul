// Benchmark "top" written by ABC on Mon Dec 25 16:58:19 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386, new_n387, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1398, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1452, new_n1453, new_n1454, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1480;
  AND2x2_ASAP7_75t_L        g0000(.A(\a[0] ), .B(\b[0] ), .Y(new_n386));
  NOR2xp33_ASAP7_75t_L      g0001(.A(\a[0] ), .B(\b[0] ), .Y(new_n387));
  NOR2xp33_ASAP7_75t_L      g0002(.A(new_n387), .B(new_n386), .Y(\f[0] ));
  INVx1_ASAP7_75t_L         g0003(.A(\a[1] ), .Y(new_n389));
  INVx1_ASAP7_75t_L         g0004(.A(\b[1] ), .Y(new_n390));
  NAND2xp33_ASAP7_75t_L     g0005(.A(new_n390), .B(new_n389), .Y(new_n391));
  INVx1_ASAP7_75t_L         g0006(.A(new_n391), .Y(new_n392));
  NOR2xp33_ASAP7_75t_L      g0007(.A(new_n389), .B(new_n390), .Y(new_n393));
  NOR2xp33_ASAP7_75t_L      g0008(.A(new_n393), .B(new_n392), .Y(new_n394));
  XOR2x2_ASAP7_75t_L        g0009(.A(new_n386), .B(new_n394), .Y(\f[1] ));
  NOR2xp33_ASAP7_75t_L      g0010(.A(\a[2] ), .B(\b[2] ), .Y(new_n396));
  INVx1_ASAP7_75t_L         g0011(.A(\a[2] ), .Y(new_n397));
  INVx1_ASAP7_75t_L         g0012(.A(\b[2] ), .Y(new_n398));
  NOR2xp33_ASAP7_75t_L      g0013(.A(new_n397), .B(new_n398), .Y(new_n399));
  NOR2xp33_ASAP7_75t_L      g0014(.A(new_n396), .B(new_n399), .Y(new_n400));
  O2A1O1Ixp33_ASAP7_75t_L   g0015(.A1(new_n386), .A2(new_n393), .B(new_n391), .C(new_n400), .Y(new_n401));
  A2O1A1Ixp33_ASAP7_75t_L   g0016(.A1(\a[0] ), .A2(\b[0] ), .B(new_n393), .C(new_n391), .Y(new_n402));
  NOR3xp33_ASAP7_75t_L      g0017(.A(new_n402), .B(new_n399), .C(new_n396), .Y(new_n403));
  NOR2xp33_ASAP7_75t_L      g0018(.A(new_n401), .B(new_n403), .Y(\f[2] ));
  NOR2xp33_ASAP7_75t_L      g0019(.A(\a[3] ), .B(\b[3] ), .Y(new_n405));
  INVx1_ASAP7_75t_L         g0020(.A(\a[3] ), .Y(new_n406));
  INVx1_ASAP7_75t_L         g0021(.A(\b[3] ), .Y(new_n407));
  NOR2xp33_ASAP7_75t_L      g0022(.A(new_n406), .B(new_n407), .Y(new_n408));
  NOR2xp33_ASAP7_75t_L      g0023(.A(new_n405), .B(new_n408), .Y(new_n409));
  MAJIxp5_ASAP7_75t_L       g0024(.A(new_n402), .B(new_n397), .C(new_n398), .Y(new_n410));
  NOR2xp33_ASAP7_75t_L      g0025(.A(new_n409), .B(new_n410), .Y(new_n411));
  A2O1A1Ixp33_ASAP7_75t_L   g0026(.A1(\b[2] ), .A2(\a[2] ), .B(new_n403), .C(new_n409), .Y(new_n412));
  INVx1_ASAP7_75t_L         g0027(.A(new_n412), .Y(new_n413));
  NOR2xp33_ASAP7_75t_L      g0028(.A(new_n411), .B(new_n413), .Y(\f[3] ));
  NOR2xp33_ASAP7_75t_L      g0029(.A(\a[4] ), .B(\b[4] ), .Y(new_n415));
  INVx1_ASAP7_75t_L         g0030(.A(new_n415), .Y(new_n416));
  NAND2xp33_ASAP7_75t_L     g0031(.A(\b[4] ), .B(\a[4] ), .Y(new_n417));
  NAND2xp33_ASAP7_75t_L     g0032(.A(new_n417), .B(new_n416), .Y(new_n418));
  O2A1O1Ixp33_ASAP7_75t_L   g0033(.A1(new_n399), .A2(new_n403), .B(new_n409), .C(new_n408), .Y(new_n419));
  AND2x2_ASAP7_75t_L        g0034(.A(new_n418), .B(new_n419), .Y(new_n420));
  O2A1O1Ixp33_ASAP7_75t_L   g0035(.A1(new_n406), .A2(new_n407), .B(new_n412), .C(new_n418), .Y(new_n421));
  NOR2xp33_ASAP7_75t_L      g0036(.A(new_n421), .B(new_n420), .Y(\f[4] ));
  INVx1_ASAP7_75t_L         g0037(.A(new_n417), .Y(new_n423));
  NOR2xp33_ASAP7_75t_L      g0038(.A(\a[5] ), .B(\b[5] ), .Y(new_n424));
  INVx1_ASAP7_75t_L         g0039(.A(\a[5] ), .Y(new_n425));
  INVx1_ASAP7_75t_L         g0040(.A(\b[5] ), .Y(new_n426));
  NOR2xp33_ASAP7_75t_L      g0041(.A(new_n425), .B(new_n426), .Y(new_n427));
  NOR2xp33_ASAP7_75t_L      g0042(.A(new_n424), .B(new_n427), .Y(new_n428));
  NOR3xp33_ASAP7_75t_L      g0043(.A(new_n421), .B(new_n428), .C(new_n423), .Y(new_n429));
  A2O1A1Ixp33_ASAP7_75t_L   g0044(.A1(\b[4] ), .A2(\a[4] ), .B(new_n421), .C(new_n428), .Y(new_n430));
  INVx1_ASAP7_75t_L         g0045(.A(new_n430), .Y(new_n431));
  NOR2xp33_ASAP7_75t_L      g0046(.A(new_n429), .B(new_n431), .Y(\f[5] ));
  NOR2xp33_ASAP7_75t_L      g0047(.A(\a[6] ), .B(\b[6] ), .Y(new_n433));
  AND2x2_ASAP7_75t_L        g0048(.A(\a[6] ), .B(\b[6] ), .Y(new_n434));
  NOR2xp33_ASAP7_75t_L      g0049(.A(new_n433), .B(new_n434), .Y(new_n435));
  INVx1_ASAP7_75t_L         g0050(.A(new_n421), .Y(new_n436));
  INVx1_ASAP7_75t_L         g0051(.A(new_n427), .Y(new_n437));
  A2O1A1Ixp33_ASAP7_75t_L   g0052(.A1(new_n436), .A2(new_n417), .B(new_n424), .C(new_n437), .Y(new_n438));
  NOR2xp33_ASAP7_75t_L      g0053(.A(new_n435), .B(new_n438), .Y(new_n439));
  A2O1A1O1Ixp25_ASAP7_75t_L g0054(.A1(new_n409), .A2(new_n410), .B(new_n408), .C(new_n416), .D(new_n423), .Y(new_n440));
  INVx1_ASAP7_75t_L         g0055(.A(new_n435), .Y(new_n441));
  O2A1O1Ixp33_ASAP7_75t_L   g0056(.A1(new_n424), .A2(new_n440), .B(new_n437), .C(new_n441), .Y(new_n442));
  NOR2xp33_ASAP7_75t_L      g0057(.A(new_n442), .B(new_n439), .Y(\f[6] ));
  INVx1_ASAP7_75t_L         g0058(.A(\a[7] ), .Y(new_n444));
  INVx1_ASAP7_75t_L         g0059(.A(\b[7] ), .Y(new_n445));
  NAND2xp33_ASAP7_75t_L     g0060(.A(new_n445), .B(new_n444), .Y(new_n446));
  NOR2xp33_ASAP7_75t_L      g0061(.A(new_n444), .B(new_n445), .Y(new_n447));
  INVx1_ASAP7_75t_L         g0062(.A(new_n447), .Y(new_n448));
  AND2x2_ASAP7_75t_L        g0063(.A(new_n446), .B(new_n448), .Y(new_n449));
  O2A1O1Ixp33_ASAP7_75t_L   g0064(.A1(new_n427), .A2(new_n431), .B(new_n435), .C(new_n434), .Y(new_n450));
  XNOR2x2_ASAP7_75t_L       g0065(.A(new_n449), .B(new_n450), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g0066(.A(\a[8] ), .B(\b[8] ), .Y(new_n452));
  INVx1_ASAP7_75t_L         g0067(.A(\a[8] ), .Y(new_n453));
  INVx1_ASAP7_75t_L         g0068(.A(\b[8] ), .Y(new_n454));
  NOR2xp33_ASAP7_75t_L      g0069(.A(new_n453), .B(new_n454), .Y(new_n455));
  NOR2xp33_ASAP7_75t_L      g0070(.A(new_n452), .B(new_n455), .Y(new_n456));
  INVx1_ASAP7_75t_L         g0071(.A(new_n456), .Y(new_n457));
  O2A1O1Ixp33_ASAP7_75t_L   g0072(.A1(new_n434), .A2(new_n442), .B(new_n446), .C(new_n447), .Y(new_n458));
  AND2x2_ASAP7_75t_L        g0073(.A(new_n457), .B(new_n458), .Y(new_n459));
  A2O1A1Ixp33_ASAP7_75t_L   g0074(.A1(\b[6] ), .A2(\a[6] ), .B(new_n442), .C(new_n449), .Y(new_n460));
  O2A1O1Ixp33_ASAP7_75t_L   g0075(.A1(new_n444), .A2(new_n445), .B(new_n460), .C(new_n457), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g0076(.A(new_n461), .B(new_n459), .Y(\f[8] ));
  NOR2xp33_ASAP7_75t_L      g0077(.A(\a[9] ), .B(\b[9] ), .Y(new_n463));
  INVx1_ASAP7_75t_L         g0078(.A(\a[9] ), .Y(new_n464));
  INVx1_ASAP7_75t_L         g0079(.A(\b[9] ), .Y(new_n465));
  NOR2xp33_ASAP7_75t_L      g0080(.A(new_n464), .B(new_n465), .Y(new_n466));
  NOR2xp33_ASAP7_75t_L      g0081(.A(new_n463), .B(new_n466), .Y(new_n467));
  INVx1_ASAP7_75t_L         g0082(.A(new_n455), .Y(new_n468));
  A2O1A1Ixp33_ASAP7_75t_L   g0083(.A1(new_n460), .A2(new_n448), .B(new_n452), .C(new_n468), .Y(new_n469));
  NOR2xp33_ASAP7_75t_L      g0084(.A(new_n467), .B(new_n469), .Y(new_n470));
  A2O1A1Ixp33_ASAP7_75t_L   g0085(.A1(\b[8] ), .A2(\a[8] ), .B(new_n461), .C(new_n467), .Y(new_n471));
  INVx1_ASAP7_75t_L         g0086(.A(new_n471), .Y(new_n472));
  NOR2xp33_ASAP7_75t_L      g0087(.A(new_n470), .B(new_n472), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g0088(.A(\a[10] ), .B(\b[10] ), .Y(new_n474));
  INVx1_ASAP7_75t_L         g0089(.A(\a[10] ), .Y(new_n475));
  INVx1_ASAP7_75t_L         g0090(.A(\b[10] ), .Y(new_n476));
  NOR2xp33_ASAP7_75t_L      g0091(.A(new_n475), .B(new_n476), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g0092(.A(new_n474), .B(new_n477), .Y(new_n478));
  INVx1_ASAP7_75t_L         g0093(.A(new_n461), .Y(new_n479));
  INVx1_ASAP7_75t_L         g0094(.A(new_n466), .Y(new_n480));
  A2O1A1Ixp33_ASAP7_75t_L   g0095(.A1(new_n479), .A2(new_n468), .B(new_n463), .C(new_n480), .Y(new_n481));
  NOR2xp33_ASAP7_75t_L      g0096(.A(new_n478), .B(new_n481), .Y(new_n482));
  INVx1_ASAP7_75t_L         g0097(.A(new_n478), .Y(new_n483));
  A2O1A1O1Ixp25_ASAP7_75t_L g0098(.A1(new_n468), .A2(new_n479), .B(new_n463), .C(new_n480), .D(new_n483), .Y(new_n484));
  NOR2xp33_ASAP7_75t_L      g0099(.A(new_n484), .B(new_n482), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g0100(.A(\a[11] ), .B(\b[11] ), .Y(new_n486));
  INVx1_ASAP7_75t_L         g0101(.A(\a[11] ), .Y(new_n487));
  INVx1_ASAP7_75t_L         g0102(.A(\b[11] ), .Y(new_n488));
  NOR2xp33_ASAP7_75t_L      g0103(.A(new_n487), .B(new_n488), .Y(new_n489));
  NOR2xp33_ASAP7_75t_L      g0104(.A(new_n486), .B(new_n489), .Y(new_n490));
  INVx1_ASAP7_75t_L         g0105(.A(new_n477), .Y(new_n491));
  A2O1A1Ixp33_ASAP7_75t_L   g0106(.A1(new_n471), .A2(new_n480), .B(new_n474), .C(new_n491), .Y(new_n492));
  NOR2xp33_ASAP7_75t_L      g0107(.A(new_n490), .B(new_n492), .Y(new_n493));
  A2O1A1Ixp33_ASAP7_75t_L   g0108(.A1(new_n481), .A2(new_n478), .B(new_n477), .C(new_n490), .Y(new_n494));
  INVx1_ASAP7_75t_L         g0109(.A(new_n494), .Y(new_n495));
  NOR2xp33_ASAP7_75t_L      g0110(.A(new_n493), .B(new_n495), .Y(\f[11] ));
  NOR2xp33_ASAP7_75t_L      g0111(.A(\a[12] ), .B(\b[12] ), .Y(new_n497));
  AND2x2_ASAP7_75t_L        g0112(.A(\a[12] ), .B(\b[12] ), .Y(new_n498));
  NOR2xp33_ASAP7_75t_L      g0113(.A(new_n497), .B(new_n498), .Y(new_n499));
  NOR3xp33_ASAP7_75t_L      g0114(.A(new_n495), .B(new_n499), .C(new_n489), .Y(new_n500));
  INVx1_ASAP7_75t_L         g0115(.A(new_n499), .Y(new_n501));
  O2A1O1Ixp33_ASAP7_75t_L   g0116(.A1(new_n487), .A2(new_n488), .B(new_n494), .C(new_n501), .Y(new_n502));
  NOR2xp33_ASAP7_75t_L      g0117(.A(new_n502), .B(new_n500), .Y(\f[12] ));
  NOR2xp33_ASAP7_75t_L      g0118(.A(\a[13] ), .B(\b[13] ), .Y(new_n504));
  INVx1_ASAP7_75t_L         g0119(.A(\a[13] ), .Y(new_n505));
  INVx1_ASAP7_75t_L         g0120(.A(\b[13] ), .Y(new_n506));
  NOR2xp33_ASAP7_75t_L      g0121(.A(new_n505), .B(new_n506), .Y(new_n507));
  NOR2xp33_ASAP7_75t_L      g0122(.A(new_n504), .B(new_n507), .Y(new_n508));
  A2O1A1O1Ixp25_ASAP7_75t_L g0123(.A1(new_n490), .A2(new_n492), .B(new_n489), .C(new_n499), .D(new_n498), .Y(new_n509));
  XNOR2x2_ASAP7_75t_L       g0124(.A(new_n508), .B(new_n509), .Y(\f[13] ));
  NOR2xp33_ASAP7_75t_L      g0125(.A(\a[14] ), .B(\b[14] ), .Y(new_n511));
  AND2x2_ASAP7_75t_L        g0126(.A(\a[14] ), .B(\b[14] ), .Y(new_n512));
  NOR2xp33_ASAP7_75t_L      g0127(.A(new_n511), .B(new_n512), .Y(new_n513));
  INVx1_ASAP7_75t_L         g0128(.A(new_n513), .Y(new_n514));
  O2A1O1Ixp33_ASAP7_75t_L   g0129(.A1(new_n498), .A2(new_n502), .B(new_n508), .C(new_n507), .Y(new_n515));
  AND2x2_ASAP7_75t_L        g0130(.A(new_n514), .B(new_n515), .Y(new_n516));
  A2O1A1Ixp33_ASAP7_75t_L   g0131(.A1(\b[12] ), .A2(\a[12] ), .B(new_n502), .C(new_n508), .Y(new_n517));
  O2A1O1Ixp33_ASAP7_75t_L   g0132(.A1(new_n505), .A2(new_n506), .B(new_n517), .C(new_n514), .Y(new_n518));
  NOR2xp33_ASAP7_75t_L      g0133(.A(new_n518), .B(new_n516), .Y(\f[14] ));
  NOR2xp33_ASAP7_75t_L      g0134(.A(\a[15] ), .B(\b[15] ), .Y(new_n520));
  INVx1_ASAP7_75t_L         g0135(.A(\a[15] ), .Y(new_n521));
  INVx1_ASAP7_75t_L         g0136(.A(\b[15] ), .Y(new_n522));
  NOR2xp33_ASAP7_75t_L      g0137(.A(new_n521), .B(new_n522), .Y(new_n523));
  NOR2xp33_ASAP7_75t_L      g0138(.A(new_n520), .B(new_n523), .Y(new_n524));
  OR3x1_ASAP7_75t_L         g0139(.A(new_n518), .B(new_n512), .C(new_n524), .Y(new_n525));
  A2O1A1Ixp33_ASAP7_75t_L   g0140(.A1(\b[14] ), .A2(\a[14] ), .B(new_n518), .C(new_n524), .Y(new_n526));
  AND2x2_ASAP7_75t_L        g0141(.A(new_n526), .B(new_n525), .Y(\f[15] ));
  NOR2xp33_ASAP7_75t_L      g0142(.A(\a[16] ), .B(\b[16] ), .Y(new_n528));
  AND2x2_ASAP7_75t_L        g0143(.A(\a[16] ), .B(\b[16] ), .Y(new_n529));
  NOR2xp33_ASAP7_75t_L      g0144(.A(new_n528), .B(new_n529), .Y(new_n530));
  INVx1_ASAP7_75t_L         g0145(.A(new_n530), .Y(new_n531));
  O2A1O1Ixp33_ASAP7_75t_L   g0146(.A1(new_n512), .A2(new_n518), .B(new_n524), .C(new_n523), .Y(new_n532));
  AND2x2_ASAP7_75t_L        g0147(.A(new_n531), .B(new_n532), .Y(new_n533));
  O2A1O1Ixp33_ASAP7_75t_L   g0148(.A1(new_n521), .A2(new_n522), .B(new_n526), .C(new_n531), .Y(new_n534));
  NOR2xp33_ASAP7_75t_L      g0149(.A(new_n534), .B(new_n533), .Y(\f[16] ));
  NOR2xp33_ASAP7_75t_L      g0150(.A(\a[17] ), .B(\b[17] ), .Y(new_n536));
  INVx1_ASAP7_75t_L         g0151(.A(\a[17] ), .Y(new_n537));
  INVx1_ASAP7_75t_L         g0152(.A(\b[17] ), .Y(new_n538));
  NOR2xp33_ASAP7_75t_L      g0153(.A(new_n537), .B(new_n538), .Y(new_n539));
  NOR2xp33_ASAP7_75t_L      g0154(.A(new_n536), .B(new_n539), .Y(new_n540));
  OR3x1_ASAP7_75t_L         g0155(.A(new_n534), .B(new_n529), .C(new_n540), .Y(new_n541));
  A2O1A1Ixp33_ASAP7_75t_L   g0156(.A1(\b[16] ), .A2(\a[16] ), .B(new_n534), .C(new_n540), .Y(new_n542));
  AND2x2_ASAP7_75t_L        g0157(.A(new_n542), .B(new_n541), .Y(\f[17] ));
  NOR2xp33_ASAP7_75t_L      g0158(.A(\a[18] ), .B(\b[18] ), .Y(new_n544));
  AND2x2_ASAP7_75t_L        g0159(.A(\a[18] ), .B(\b[18] ), .Y(new_n545));
  NOR2xp33_ASAP7_75t_L      g0160(.A(new_n544), .B(new_n545), .Y(new_n546));
  INVx1_ASAP7_75t_L         g0161(.A(new_n546), .Y(new_n547));
  O2A1O1Ixp33_ASAP7_75t_L   g0162(.A1(new_n529), .A2(new_n534), .B(new_n540), .C(new_n539), .Y(new_n548));
  AND2x2_ASAP7_75t_L        g0163(.A(new_n547), .B(new_n548), .Y(new_n549));
  O2A1O1Ixp33_ASAP7_75t_L   g0164(.A1(new_n537), .A2(new_n538), .B(new_n542), .C(new_n547), .Y(new_n550));
  NOR2xp33_ASAP7_75t_L      g0165(.A(new_n550), .B(new_n549), .Y(\f[18] ));
  NOR2xp33_ASAP7_75t_L      g0166(.A(\a[19] ), .B(\b[19] ), .Y(new_n552));
  INVx1_ASAP7_75t_L         g0167(.A(\a[19] ), .Y(new_n553));
  INVx1_ASAP7_75t_L         g0168(.A(\b[19] ), .Y(new_n554));
  NOR2xp33_ASAP7_75t_L      g0169(.A(new_n553), .B(new_n554), .Y(new_n555));
  NOR2xp33_ASAP7_75t_L      g0170(.A(new_n552), .B(new_n555), .Y(new_n556));
  OR3x1_ASAP7_75t_L         g0171(.A(new_n550), .B(new_n545), .C(new_n556), .Y(new_n557));
  A2O1A1Ixp33_ASAP7_75t_L   g0172(.A1(\b[18] ), .A2(\a[18] ), .B(new_n550), .C(new_n556), .Y(new_n558));
  AND2x2_ASAP7_75t_L        g0173(.A(new_n558), .B(new_n557), .Y(\f[19] ));
  NOR2xp33_ASAP7_75t_L      g0174(.A(\a[20] ), .B(\b[20] ), .Y(new_n560));
  AND2x2_ASAP7_75t_L        g0175(.A(\a[20] ), .B(\b[20] ), .Y(new_n561));
  NOR2xp33_ASAP7_75t_L      g0176(.A(new_n560), .B(new_n561), .Y(new_n562));
  INVx1_ASAP7_75t_L         g0177(.A(new_n562), .Y(new_n563));
  O2A1O1Ixp33_ASAP7_75t_L   g0178(.A1(new_n545), .A2(new_n550), .B(new_n556), .C(new_n555), .Y(new_n564));
  AND2x2_ASAP7_75t_L        g0179(.A(new_n563), .B(new_n564), .Y(new_n565));
  O2A1O1Ixp33_ASAP7_75t_L   g0180(.A1(new_n553), .A2(new_n554), .B(new_n558), .C(new_n563), .Y(new_n566));
  NOR2xp33_ASAP7_75t_L      g0181(.A(new_n566), .B(new_n565), .Y(\f[20] ));
  NOR2xp33_ASAP7_75t_L      g0182(.A(\a[21] ), .B(\b[21] ), .Y(new_n568));
  INVx1_ASAP7_75t_L         g0183(.A(\a[21] ), .Y(new_n569));
  INVx1_ASAP7_75t_L         g0184(.A(\b[21] ), .Y(new_n570));
  NOR2xp33_ASAP7_75t_L      g0185(.A(new_n569), .B(new_n570), .Y(new_n571));
  NOR2xp33_ASAP7_75t_L      g0186(.A(new_n568), .B(new_n571), .Y(new_n572));
  OR3x1_ASAP7_75t_L         g0187(.A(new_n566), .B(new_n561), .C(new_n572), .Y(new_n573));
  A2O1A1Ixp33_ASAP7_75t_L   g0188(.A1(\b[20] ), .A2(\a[20] ), .B(new_n566), .C(new_n572), .Y(new_n574));
  AND2x2_ASAP7_75t_L        g0189(.A(new_n574), .B(new_n573), .Y(\f[21] ));
  NOR2xp33_ASAP7_75t_L      g0190(.A(\a[22] ), .B(\b[22] ), .Y(new_n576));
  AND2x2_ASAP7_75t_L        g0191(.A(\a[22] ), .B(\b[22] ), .Y(new_n577));
  NOR2xp33_ASAP7_75t_L      g0192(.A(new_n576), .B(new_n577), .Y(new_n578));
  INVx1_ASAP7_75t_L         g0193(.A(new_n578), .Y(new_n579));
  O2A1O1Ixp33_ASAP7_75t_L   g0194(.A1(new_n561), .A2(new_n566), .B(new_n572), .C(new_n571), .Y(new_n580));
  AND2x2_ASAP7_75t_L        g0195(.A(new_n579), .B(new_n580), .Y(new_n581));
  O2A1O1Ixp33_ASAP7_75t_L   g0196(.A1(new_n569), .A2(new_n570), .B(new_n574), .C(new_n579), .Y(new_n582));
  NOR2xp33_ASAP7_75t_L      g0197(.A(new_n582), .B(new_n581), .Y(\f[22] ));
  NOR2xp33_ASAP7_75t_L      g0198(.A(\a[23] ), .B(\b[23] ), .Y(new_n584));
  INVx1_ASAP7_75t_L         g0199(.A(\a[23] ), .Y(new_n585));
  INVx1_ASAP7_75t_L         g0200(.A(\b[23] ), .Y(new_n586));
  NOR2xp33_ASAP7_75t_L      g0201(.A(new_n585), .B(new_n586), .Y(new_n587));
  NOR2xp33_ASAP7_75t_L      g0202(.A(new_n584), .B(new_n587), .Y(new_n588));
  OR3x1_ASAP7_75t_L         g0203(.A(new_n582), .B(new_n577), .C(new_n588), .Y(new_n589));
  A2O1A1Ixp33_ASAP7_75t_L   g0204(.A1(\b[22] ), .A2(\a[22] ), .B(new_n582), .C(new_n588), .Y(new_n590));
  AND2x2_ASAP7_75t_L        g0205(.A(new_n590), .B(new_n589), .Y(\f[23] ));
  NOR2xp33_ASAP7_75t_L      g0206(.A(\a[24] ), .B(\b[24] ), .Y(new_n592));
  AND2x2_ASAP7_75t_L        g0207(.A(\a[24] ), .B(\b[24] ), .Y(new_n593));
  NOR2xp33_ASAP7_75t_L      g0208(.A(new_n592), .B(new_n593), .Y(new_n594));
  INVx1_ASAP7_75t_L         g0209(.A(new_n594), .Y(new_n595));
  O2A1O1Ixp33_ASAP7_75t_L   g0210(.A1(new_n577), .A2(new_n582), .B(new_n588), .C(new_n587), .Y(new_n596));
  AND2x2_ASAP7_75t_L        g0211(.A(new_n595), .B(new_n596), .Y(new_n597));
  O2A1O1Ixp33_ASAP7_75t_L   g0212(.A1(new_n585), .A2(new_n586), .B(new_n590), .C(new_n595), .Y(new_n598));
  NOR2xp33_ASAP7_75t_L      g0213(.A(new_n598), .B(new_n597), .Y(\f[24] ));
  NOR2xp33_ASAP7_75t_L      g0214(.A(\a[25] ), .B(\b[25] ), .Y(new_n600));
  INVx1_ASAP7_75t_L         g0215(.A(\a[25] ), .Y(new_n601));
  INVx1_ASAP7_75t_L         g0216(.A(\b[25] ), .Y(new_n602));
  NOR2xp33_ASAP7_75t_L      g0217(.A(new_n601), .B(new_n602), .Y(new_n603));
  NOR2xp33_ASAP7_75t_L      g0218(.A(new_n600), .B(new_n603), .Y(new_n604));
  OR3x1_ASAP7_75t_L         g0219(.A(new_n598), .B(new_n593), .C(new_n604), .Y(new_n605));
  A2O1A1Ixp33_ASAP7_75t_L   g0220(.A1(\b[24] ), .A2(\a[24] ), .B(new_n598), .C(new_n604), .Y(new_n606));
  AND2x2_ASAP7_75t_L        g0221(.A(new_n606), .B(new_n605), .Y(\f[25] ));
  NOR2xp33_ASAP7_75t_L      g0222(.A(\a[26] ), .B(\b[26] ), .Y(new_n608));
  AND2x2_ASAP7_75t_L        g0223(.A(\a[26] ), .B(\b[26] ), .Y(new_n609));
  NOR2xp33_ASAP7_75t_L      g0224(.A(new_n608), .B(new_n609), .Y(new_n610));
  INVx1_ASAP7_75t_L         g0225(.A(new_n610), .Y(new_n611));
  O2A1O1Ixp33_ASAP7_75t_L   g0226(.A1(new_n593), .A2(new_n598), .B(new_n604), .C(new_n603), .Y(new_n612));
  AND2x2_ASAP7_75t_L        g0227(.A(new_n611), .B(new_n612), .Y(new_n613));
  O2A1O1Ixp33_ASAP7_75t_L   g0228(.A1(new_n601), .A2(new_n602), .B(new_n606), .C(new_n611), .Y(new_n614));
  NOR2xp33_ASAP7_75t_L      g0229(.A(new_n614), .B(new_n613), .Y(\f[26] ));
  NOR2xp33_ASAP7_75t_L      g0230(.A(\a[27] ), .B(\b[27] ), .Y(new_n616));
  INVx1_ASAP7_75t_L         g0231(.A(\a[27] ), .Y(new_n617));
  INVx1_ASAP7_75t_L         g0232(.A(\b[27] ), .Y(new_n618));
  NOR2xp33_ASAP7_75t_L      g0233(.A(new_n617), .B(new_n618), .Y(new_n619));
  NOR2xp33_ASAP7_75t_L      g0234(.A(new_n616), .B(new_n619), .Y(new_n620));
  OR3x1_ASAP7_75t_L         g0235(.A(new_n614), .B(new_n609), .C(new_n620), .Y(new_n621));
  A2O1A1Ixp33_ASAP7_75t_L   g0236(.A1(\b[26] ), .A2(\a[26] ), .B(new_n614), .C(new_n620), .Y(new_n622));
  AND2x2_ASAP7_75t_L        g0237(.A(new_n622), .B(new_n621), .Y(\f[27] ));
  NOR2xp33_ASAP7_75t_L      g0238(.A(\a[28] ), .B(\b[28] ), .Y(new_n624));
  AND2x2_ASAP7_75t_L        g0239(.A(\a[28] ), .B(\b[28] ), .Y(new_n625));
  NOR2xp33_ASAP7_75t_L      g0240(.A(new_n624), .B(new_n625), .Y(new_n626));
  INVx1_ASAP7_75t_L         g0241(.A(new_n626), .Y(new_n627));
  O2A1O1Ixp33_ASAP7_75t_L   g0242(.A1(new_n609), .A2(new_n614), .B(new_n620), .C(new_n619), .Y(new_n628));
  AND2x2_ASAP7_75t_L        g0243(.A(new_n627), .B(new_n628), .Y(new_n629));
  O2A1O1Ixp33_ASAP7_75t_L   g0244(.A1(new_n617), .A2(new_n618), .B(new_n622), .C(new_n627), .Y(new_n630));
  NOR2xp33_ASAP7_75t_L      g0245(.A(new_n630), .B(new_n629), .Y(\f[28] ));
  NOR2xp33_ASAP7_75t_L      g0246(.A(\a[29] ), .B(\b[29] ), .Y(new_n632));
  INVx1_ASAP7_75t_L         g0247(.A(\a[29] ), .Y(new_n633));
  INVx1_ASAP7_75t_L         g0248(.A(\b[29] ), .Y(new_n634));
  NOR2xp33_ASAP7_75t_L      g0249(.A(new_n633), .B(new_n634), .Y(new_n635));
  NOR2xp33_ASAP7_75t_L      g0250(.A(new_n632), .B(new_n635), .Y(new_n636));
  OR3x1_ASAP7_75t_L         g0251(.A(new_n630), .B(new_n625), .C(new_n636), .Y(new_n637));
  A2O1A1Ixp33_ASAP7_75t_L   g0252(.A1(\b[28] ), .A2(\a[28] ), .B(new_n630), .C(new_n636), .Y(new_n638));
  AND2x2_ASAP7_75t_L        g0253(.A(new_n638), .B(new_n637), .Y(\f[29] ));
  NOR2xp33_ASAP7_75t_L      g0254(.A(\a[30] ), .B(\b[30] ), .Y(new_n640));
  AND2x2_ASAP7_75t_L        g0255(.A(\a[30] ), .B(\b[30] ), .Y(new_n641));
  NOR2xp33_ASAP7_75t_L      g0256(.A(new_n640), .B(new_n641), .Y(new_n642));
  INVx1_ASAP7_75t_L         g0257(.A(new_n642), .Y(new_n643));
  O2A1O1Ixp33_ASAP7_75t_L   g0258(.A1(new_n625), .A2(new_n630), .B(new_n636), .C(new_n635), .Y(new_n644));
  AND2x2_ASAP7_75t_L        g0259(.A(new_n643), .B(new_n644), .Y(new_n645));
  O2A1O1Ixp33_ASAP7_75t_L   g0260(.A1(new_n633), .A2(new_n634), .B(new_n638), .C(new_n643), .Y(new_n646));
  NOR2xp33_ASAP7_75t_L      g0261(.A(new_n646), .B(new_n645), .Y(\f[30] ));
  NOR2xp33_ASAP7_75t_L      g0262(.A(\a[31] ), .B(\b[31] ), .Y(new_n648));
  INVx1_ASAP7_75t_L         g0263(.A(\a[31] ), .Y(new_n649));
  INVx1_ASAP7_75t_L         g0264(.A(\b[31] ), .Y(new_n650));
  NOR2xp33_ASAP7_75t_L      g0265(.A(new_n649), .B(new_n650), .Y(new_n651));
  NOR2xp33_ASAP7_75t_L      g0266(.A(new_n648), .B(new_n651), .Y(new_n652));
  OR3x1_ASAP7_75t_L         g0267(.A(new_n646), .B(new_n641), .C(new_n652), .Y(new_n653));
  A2O1A1Ixp33_ASAP7_75t_L   g0268(.A1(\b[30] ), .A2(\a[30] ), .B(new_n646), .C(new_n652), .Y(new_n654));
  AND2x2_ASAP7_75t_L        g0269(.A(new_n654), .B(new_n653), .Y(\f[31] ));
  NOR2xp33_ASAP7_75t_L      g0270(.A(\a[32] ), .B(\b[32] ), .Y(new_n656));
  AND2x2_ASAP7_75t_L        g0271(.A(\a[32] ), .B(\b[32] ), .Y(new_n657));
  NOR2xp33_ASAP7_75t_L      g0272(.A(new_n656), .B(new_n657), .Y(new_n658));
  INVx1_ASAP7_75t_L         g0273(.A(new_n658), .Y(new_n659));
  O2A1O1Ixp33_ASAP7_75t_L   g0274(.A1(new_n641), .A2(new_n646), .B(new_n652), .C(new_n651), .Y(new_n660));
  AND2x2_ASAP7_75t_L        g0275(.A(new_n659), .B(new_n660), .Y(new_n661));
  O2A1O1Ixp33_ASAP7_75t_L   g0276(.A1(new_n649), .A2(new_n650), .B(new_n654), .C(new_n659), .Y(new_n662));
  NOR2xp33_ASAP7_75t_L      g0277(.A(new_n662), .B(new_n661), .Y(\f[32] ));
  NOR2xp33_ASAP7_75t_L      g0278(.A(\a[33] ), .B(\b[33] ), .Y(new_n664));
  INVx1_ASAP7_75t_L         g0279(.A(\a[33] ), .Y(new_n665));
  INVx1_ASAP7_75t_L         g0280(.A(\b[33] ), .Y(new_n666));
  NOR2xp33_ASAP7_75t_L      g0281(.A(new_n665), .B(new_n666), .Y(new_n667));
  NOR2xp33_ASAP7_75t_L      g0282(.A(new_n664), .B(new_n667), .Y(new_n668));
  OR3x1_ASAP7_75t_L         g0283(.A(new_n662), .B(new_n657), .C(new_n668), .Y(new_n669));
  A2O1A1Ixp33_ASAP7_75t_L   g0284(.A1(\b[32] ), .A2(\a[32] ), .B(new_n662), .C(new_n668), .Y(new_n670));
  AND2x2_ASAP7_75t_L        g0285(.A(new_n670), .B(new_n669), .Y(\f[33] ));
  NOR2xp33_ASAP7_75t_L      g0286(.A(\a[34] ), .B(\b[34] ), .Y(new_n672));
  AND2x2_ASAP7_75t_L        g0287(.A(\a[34] ), .B(\b[34] ), .Y(new_n673));
  NOR2xp33_ASAP7_75t_L      g0288(.A(new_n672), .B(new_n673), .Y(new_n674));
  INVx1_ASAP7_75t_L         g0289(.A(new_n674), .Y(new_n675));
  O2A1O1Ixp33_ASAP7_75t_L   g0290(.A1(new_n657), .A2(new_n662), .B(new_n668), .C(new_n667), .Y(new_n676));
  AND2x2_ASAP7_75t_L        g0291(.A(new_n675), .B(new_n676), .Y(new_n677));
  O2A1O1Ixp33_ASAP7_75t_L   g0292(.A1(new_n665), .A2(new_n666), .B(new_n670), .C(new_n675), .Y(new_n678));
  NOR2xp33_ASAP7_75t_L      g0293(.A(new_n678), .B(new_n677), .Y(\f[34] ));
  NOR2xp33_ASAP7_75t_L      g0294(.A(\a[35] ), .B(\b[35] ), .Y(new_n680));
  INVx1_ASAP7_75t_L         g0295(.A(\a[35] ), .Y(new_n681));
  INVx1_ASAP7_75t_L         g0296(.A(\b[35] ), .Y(new_n682));
  NOR2xp33_ASAP7_75t_L      g0297(.A(new_n681), .B(new_n682), .Y(new_n683));
  NOR2xp33_ASAP7_75t_L      g0298(.A(new_n680), .B(new_n683), .Y(new_n684));
  OR3x1_ASAP7_75t_L         g0299(.A(new_n678), .B(new_n673), .C(new_n684), .Y(new_n685));
  A2O1A1Ixp33_ASAP7_75t_L   g0300(.A1(\b[34] ), .A2(\a[34] ), .B(new_n678), .C(new_n684), .Y(new_n686));
  AND2x2_ASAP7_75t_L        g0301(.A(new_n686), .B(new_n685), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g0302(.A(\a[36] ), .B(\b[36] ), .Y(new_n688));
  AND2x2_ASAP7_75t_L        g0303(.A(\a[36] ), .B(\b[36] ), .Y(new_n689));
  NOR2xp33_ASAP7_75t_L      g0304(.A(new_n688), .B(new_n689), .Y(new_n690));
  INVx1_ASAP7_75t_L         g0305(.A(new_n690), .Y(new_n691));
  O2A1O1Ixp33_ASAP7_75t_L   g0306(.A1(new_n673), .A2(new_n678), .B(new_n684), .C(new_n683), .Y(new_n692));
  AND2x2_ASAP7_75t_L        g0307(.A(new_n691), .B(new_n692), .Y(new_n693));
  O2A1O1Ixp33_ASAP7_75t_L   g0308(.A1(new_n681), .A2(new_n682), .B(new_n686), .C(new_n691), .Y(new_n694));
  NOR2xp33_ASAP7_75t_L      g0309(.A(new_n694), .B(new_n693), .Y(\f[36] ));
  INVx1_ASAP7_75t_L         g0310(.A(\a[37] ), .Y(new_n696));
  INVx1_ASAP7_75t_L         g0311(.A(\b[37] ), .Y(new_n697));
  NAND2xp33_ASAP7_75t_L     g0312(.A(new_n697), .B(new_n696), .Y(new_n698));
  NOR2xp33_ASAP7_75t_L      g0313(.A(new_n696), .B(new_n697), .Y(new_n699));
  INVx1_ASAP7_75t_L         g0314(.A(new_n699), .Y(new_n700));
  AND2x2_ASAP7_75t_L        g0315(.A(new_n698), .B(new_n700), .Y(new_n701));
  OR3x1_ASAP7_75t_L         g0316(.A(new_n694), .B(new_n689), .C(new_n701), .Y(new_n702));
  A2O1A1Ixp33_ASAP7_75t_L   g0317(.A1(\b[36] ), .A2(\a[36] ), .B(new_n694), .C(new_n701), .Y(new_n703));
  AND2x2_ASAP7_75t_L        g0318(.A(new_n703), .B(new_n702), .Y(\f[37] ));
  NOR2xp33_ASAP7_75t_L      g0319(.A(\a[38] ), .B(\b[38] ), .Y(new_n705));
  INVx1_ASAP7_75t_L         g0320(.A(\a[38] ), .Y(new_n706));
  INVx1_ASAP7_75t_L         g0321(.A(\b[38] ), .Y(new_n707));
  NOR2xp33_ASAP7_75t_L      g0322(.A(new_n706), .B(new_n707), .Y(new_n708));
  NOR2xp33_ASAP7_75t_L      g0323(.A(new_n705), .B(new_n708), .Y(new_n709));
  INVx1_ASAP7_75t_L         g0324(.A(new_n709), .Y(new_n710));
  O2A1O1Ixp33_ASAP7_75t_L   g0325(.A1(new_n689), .A2(new_n694), .B(new_n698), .C(new_n699), .Y(new_n711));
  AND2x2_ASAP7_75t_L        g0326(.A(new_n710), .B(new_n711), .Y(new_n712));
  O2A1O1Ixp33_ASAP7_75t_L   g0327(.A1(new_n696), .A2(new_n697), .B(new_n703), .C(new_n710), .Y(new_n713));
  NOR2xp33_ASAP7_75t_L      g0328(.A(new_n713), .B(new_n712), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g0329(.A(\a[39] ), .B(\b[39] ), .Y(new_n715));
  AND2x2_ASAP7_75t_L        g0330(.A(\a[39] ), .B(\b[39] ), .Y(new_n716));
  NOR2xp33_ASAP7_75t_L      g0331(.A(new_n715), .B(new_n716), .Y(new_n717));
  INVx1_ASAP7_75t_L         g0332(.A(new_n708), .Y(new_n718));
  A2O1A1Ixp33_ASAP7_75t_L   g0333(.A1(new_n703), .A2(new_n700), .B(new_n705), .C(new_n718), .Y(new_n719));
  NOR2xp33_ASAP7_75t_L      g0334(.A(new_n717), .B(new_n719), .Y(new_n720));
  A2O1A1Ixp33_ASAP7_75t_L   g0335(.A1(\b[38] ), .A2(\a[38] ), .B(new_n713), .C(new_n717), .Y(new_n721));
  INVx1_ASAP7_75t_L         g0336(.A(new_n721), .Y(new_n722));
  NOR2xp33_ASAP7_75t_L      g0337(.A(new_n720), .B(new_n722), .Y(\f[39] ));
  INVx1_ASAP7_75t_L         g0338(.A(\a[40] ), .Y(new_n724));
  INVx1_ASAP7_75t_L         g0339(.A(\b[40] ), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g0340(.A(new_n725), .B(new_n724), .Y(new_n726));
  NOR2xp33_ASAP7_75t_L      g0341(.A(new_n724), .B(new_n725), .Y(new_n727));
  INVx1_ASAP7_75t_L         g0342(.A(new_n727), .Y(new_n728));
  AND2x2_ASAP7_75t_L        g0343(.A(new_n726), .B(new_n728), .Y(new_n729));
  O2A1O1Ixp33_ASAP7_75t_L   g0344(.A1(new_n708), .A2(new_n713), .B(new_n717), .C(new_n716), .Y(new_n730));
  XNOR2x2_ASAP7_75t_L       g0345(.A(new_n729), .B(new_n730), .Y(\f[40] ));
  A2O1A1Ixp33_ASAP7_75t_L   g0346(.A1(new_n719), .A2(new_n717), .B(new_n716), .C(new_n729), .Y(new_n732));
  NOR2xp33_ASAP7_75t_L      g0347(.A(\a[41] ), .B(\b[41] ), .Y(new_n733));
  INVx1_ASAP7_75t_L         g0348(.A(\a[41] ), .Y(new_n734));
  INVx1_ASAP7_75t_L         g0349(.A(\b[41] ), .Y(new_n735));
  NOR2xp33_ASAP7_75t_L      g0350(.A(new_n734), .B(new_n735), .Y(new_n736));
  NOR2xp33_ASAP7_75t_L      g0351(.A(new_n733), .B(new_n736), .Y(new_n737));
  INVx1_ASAP7_75t_L         g0352(.A(new_n737), .Y(new_n738));
  AND3x1_ASAP7_75t_L        g0353(.A(new_n732), .B(new_n738), .C(new_n728), .Y(new_n739));
  O2A1O1Ixp33_ASAP7_75t_L   g0354(.A1(new_n724), .A2(new_n725), .B(new_n732), .C(new_n738), .Y(new_n740));
  NOR2xp33_ASAP7_75t_L      g0355(.A(new_n740), .B(new_n739), .Y(\f[41] ));
  NOR2xp33_ASAP7_75t_L      g0356(.A(\a[42] ), .B(\b[42] ), .Y(new_n742));
  AND2x2_ASAP7_75t_L        g0357(.A(\a[42] ), .B(\b[42] ), .Y(new_n743));
  NOR2xp33_ASAP7_75t_L      g0358(.A(new_n742), .B(new_n743), .Y(new_n744));
  INVx1_ASAP7_75t_L         g0359(.A(new_n736), .Y(new_n745));
  A2O1A1Ixp33_ASAP7_75t_L   g0360(.A1(new_n732), .A2(new_n728), .B(new_n733), .C(new_n745), .Y(new_n746));
  NOR2xp33_ASAP7_75t_L      g0361(.A(new_n744), .B(new_n746), .Y(new_n747));
  A2O1A1Ixp33_ASAP7_75t_L   g0362(.A1(\b[41] ), .A2(\a[41] ), .B(new_n740), .C(new_n744), .Y(new_n748));
  INVx1_ASAP7_75t_L         g0363(.A(new_n748), .Y(new_n749));
  NOR2xp33_ASAP7_75t_L      g0364(.A(new_n747), .B(new_n749), .Y(\f[42] ));
  NOR2xp33_ASAP7_75t_L      g0365(.A(\a[43] ), .B(\b[43] ), .Y(new_n751));
  INVx1_ASAP7_75t_L         g0366(.A(\a[43] ), .Y(new_n752));
  INVx1_ASAP7_75t_L         g0367(.A(\b[43] ), .Y(new_n753));
  NOR2xp33_ASAP7_75t_L      g0368(.A(new_n752), .B(new_n753), .Y(new_n754));
  NOR2xp33_ASAP7_75t_L      g0369(.A(new_n751), .B(new_n754), .Y(new_n755));
  NOR3xp33_ASAP7_75t_L      g0370(.A(new_n749), .B(new_n755), .C(new_n743), .Y(new_n756));
  A2O1A1Ixp33_ASAP7_75t_L   g0371(.A1(new_n746), .A2(new_n744), .B(new_n743), .C(new_n755), .Y(new_n757));
  INVx1_ASAP7_75t_L         g0372(.A(new_n757), .Y(new_n758));
  NOR2xp33_ASAP7_75t_L      g0373(.A(new_n758), .B(new_n756), .Y(\f[43] ));
  NOR2xp33_ASAP7_75t_L      g0374(.A(\a[44] ), .B(\b[44] ), .Y(new_n760));
  NAND2xp33_ASAP7_75t_L     g0375(.A(\b[44] ), .B(\a[44] ), .Y(new_n761));
  INVx1_ASAP7_75t_L         g0376(.A(new_n761), .Y(new_n762));
  NOR2xp33_ASAP7_75t_L      g0377(.A(new_n760), .B(new_n762), .Y(new_n763));
  A2O1A1O1Ixp25_ASAP7_75t_L g0378(.A1(new_n744), .A2(new_n746), .B(new_n743), .C(new_n755), .D(new_n754), .Y(new_n764));
  XNOR2x2_ASAP7_75t_L       g0379(.A(new_n763), .B(new_n764), .Y(\f[44] ));
  NOR2xp33_ASAP7_75t_L      g0380(.A(\a[45] ), .B(\b[45] ), .Y(new_n766));
  INVx1_ASAP7_75t_L         g0381(.A(\a[45] ), .Y(new_n767));
  INVx1_ASAP7_75t_L         g0382(.A(\b[45] ), .Y(new_n768));
  NOR2xp33_ASAP7_75t_L      g0383(.A(new_n767), .B(new_n768), .Y(new_n769));
  NOR2xp33_ASAP7_75t_L      g0384(.A(new_n766), .B(new_n769), .Y(new_n770));
  INVx1_ASAP7_75t_L         g0385(.A(new_n754), .Y(new_n771));
  A2O1A1Ixp33_ASAP7_75t_L   g0386(.A1(new_n757), .A2(new_n771), .B(new_n760), .C(new_n761), .Y(new_n772));
  XOR2x2_ASAP7_75t_L        g0387(.A(new_n770), .B(new_n772), .Y(\f[45] ));
  NOR2xp33_ASAP7_75t_L      g0388(.A(\a[46] ), .B(\b[46] ), .Y(new_n774));
  INVx1_ASAP7_75t_L         g0389(.A(\a[46] ), .Y(new_n775));
  INVx1_ASAP7_75t_L         g0390(.A(\b[46] ), .Y(new_n776));
  NOR2xp33_ASAP7_75t_L      g0391(.A(new_n775), .B(new_n776), .Y(new_n777));
  NOR2xp33_ASAP7_75t_L      g0392(.A(new_n774), .B(new_n777), .Y(new_n778));
  A2O1A1Ixp33_ASAP7_75t_L   g0393(.A1(\b[43] ), .A2(\a[43] ), .B(new_n758), .C(new_n763), .Y(new_n779));
  INVx1_ASAP7_75t_L         g0394(.A(new_n769), .Y(new_n780));
  A2O1A1Ixp33_ASAP7_75t_L   g0395(.A1(new_n779), .A2(new_n761), .B(new_n766), .C(new_n780), .Y(new_n781));
  NOR2xp33_ASAP7_75t_L      g0396(.A(new_n778), .B(new_n781), .Y(new_n782));
  A2O1A1Ixp33_ASAP7_75t_L   g0397(.A1(new_n772), .A2(new_n770), .B(new_n769), .C(new_n778), .Y(new_n783));
  INVx1_ASAP7_75t_L         g0398(.A(new_n783), .Y(new_n784));
  NOR2xp33_ASAP7_75t_L      g0399(.A(new_n784), .B(new_n782), .Y(\f[46] ));
  NOR2xp33_ASAP7_75t_L      g0400(.A(\a[47] ), .B(\b[47] ), .Y(new_n786));
  NAND2xp33_ASAP7_75t_L     g0401(.A(\b[47] ), .B(\a[47] ), .Y(new_n787));
  INVx1_ASAP7_75t_L         g0402(.A(new_n787), .Y(new_n788));
  NOR2xp33_ASAP7_75t_L      g0403(.A(new_n786), .B(new_n788), .Y(new_n789));
  A2O1A1O1Ixp25_ASAP7_75t_L g0404(.A1(new_n770), .A2(new_n772), .B(new_n769), .C(new_n778), .D(new_n777), .Y(new_n790));
  XNOR2x2_ASAP7_75t_L       g0405(.A(new_n789), .B(new_n790), .Y(\f[47] ));
  NOR2xp33_ASAP7_75t_L      g0406(.A(\a[48] ), .B(\b[48] ), .Y(new_n792));
  INVx1_ASAP7_75t_L         g0407(.A(\a[48] ), .Y(new_n793));
  INVx1_ASAP7_75t_L         g0408(.A(\b[48] ), .Y(new_n794));
  NOR2xp33_ASAP7_75t_L      g0409(.A(new_n793), .B(new_n794), .Y(new_n795));
  NOR2xp33_ASAP7_75t_L      g0410(.A(new_n792), .B(new_n795), .Y(new_n796));
  INVx1_ASAP7_75t_L         g0411(.A(new_n777), .Y(new_n797));
  A2O1A1Ixp33_ASAP7_75t_L   g0412(.A1(new_n783), .A2(new_n797), .B(new_n786), .C(new_n787), .Y(new_n798));
  XOR2x2_ASAP7_75t_L        g0413(.A(new_n796), .B(new_n798), .Y(\f[48] ));
  NOR2xp33_ASAP7_75t_L      g0414(.A(\a[49] ), .B(\b[49] ), .Y(new_n800));
  INVx1_ASAP7_75t_L         g0415(.A(\a[49] ), .Y(new_n801));
  INVx1_ASAP7_75t_L         g0416(.A(\b[49] ), .Y(new_n802));
  NOR2xp33_ASAP7_75t_L      g0417(.A(new_n801), .B(new_n802), .Y(new_n803));
  NOR2xp33_ASAP7_75t_L      g0418(.A(new_n800), .B(new_n803), .Y(new_n804));
  A2O1A1Ixp33_ASAP7_75t_L   g0419(.A1(new_n781), .A2(new_n778), .B(new_n777), .C(new_n789), .Y(new_n805));
  INVx1_ASAP7_75t_L         g0420(.A(new_n795), .Y(new_n806));
  A2O1A1Ixp33_ASAP7_75t_L   g0421(.A1(new_n805), .A2(new_n787), .B(new_n792), .C(new_n806), .Y(new_n807));
  NOR2xp33_ASAP7_75t_L      g0422(.A(new_n804), .B(new_n807), .Y(new_n808));
  A2O1A1Ixp33_ASAP7_75t_L   g0423(.A1(new_n798), .A2(new_n796), .B(new_n795), .C(new_n804), .Y(new_n809));
  INVx1_ASAP7_75t_L         g0424(.A(new_n809), .Y(new_n810));
  NOR2xp33_ASAP7_75t_L      g0425(.A(new_n810), .B(new_n808), .Y(\f[49] ));
  NOR2xp33_ASAP7_75t_L      g0426(.A(\a[50] ), .B(\b[50] ), .Y(new_n812));
  NAND2xp33_ASAP7_75t_L     g0427(.A(\b[50] ), .B(\a[50] ), .Y(new_n813));
  INVx1_ASAP7_75t_L         g0428(.A(new_n813), .Y(new_n814));
  NOR2xp33_ASAP7_75t_L      g0429(.A(new_n812), .B(new_n814), .Y(new_n815));
  A2O1A1O1Ixp25_ASAP7_75t_L g0430(.A1(new_n796), .A2(new_n798), .B(new_n795), .C(new_n804), .D(new_n803), .Y(new_n816));
  XNOR2x2_ASAP7_75t_L       g0431(.A(new_n815), .B(new_n816), .Y(\f[50] ));
  NOR2xp33_ASAP7_75t_L      g0432(.A(\a[51] ), .B(\b[51] ), .Y(new_n818));
  INVx1_ASAP7_75t_L         g0433(.A(\a[51] ), .Y(new_n819));
  INVx1_ASAP7_75t_L         g0434(.A(\b[51] ), .Y(new_n820));
  NOR2xp33_ASAP7_75t_L      g0435(.A(new_n819), .B(new_n820), .Y(new_n821));
  NOR2xp33_ASAP7_75t_L      g0436(.A(new_n818), .B(new_n821), .Y(new_n822));
  INVx1_ASAP7_75t_L         g0437(.A(new_n803), .Y(new_n823));
  A2O1A1Ixp33_ASAP7_75t_L   g0438(.A1(new_n809), .A2(new_n823), .B(new_n812), .C(new_n813), .Y(new_n824));
  XOR2x2_ASAP7_75t_L        g0439(.A(new_n822), .B(new_n824), .Y(\f[51] ));
  NOR2xp33_ASAP7_75t_L      g0440(.A(\a[52] ), .B(\b[52] ), .Y(new_n826));
  INVx1_ASAP7_75t_L         g0441(.A(\a[52] ), .Y(new_n827));
  INVx1_ASAP7_75t_L         g0442(.A(\b[52] ), .Y(new_n828));
  NOR2xp33_ASAP7_75t_L      g0443(.A(new_n827), .B(new_n828), .Y(new_n829));
  NOR2xp33_ASAP7_75t_L      g0444(.A(new_n826), .B(new_n829), .Y(new_n830));
  A2O1A1Ixp33_ASAP7_75t_L   g0445(.A1(new_n807), .A2(new_n804), .B(new_n803), .C(new_n815), .Y(new_n831));
  INVx1_ASAP7_75t_L         g0446(.A(new_n821), .Y(new_n832));
  A2O1A1Ixp33_ASAP7_75t_L   g0447(.A1(new_n831), .A2(new_n813), .B(new_n818), .C(new_n832), .Y(new_n833));
  NOR2xp33_ASAP7_75t_L      g0448(.A(new_n830), .B(new_n833), .Y(new_n834));
  A2O1A1Ixp33_ASAP7_75t_L   g0449(.A1(new_n824), .A2(new_n822), .B(new_n821), .C(new_n830), .Y(new_n835));
  INVx1_ASAP7_75t_L         g0450(.A(new_n835), .Y(new_n836));
  NOR2xp33_ASAP7_75t_L      g0451(.A(new_n836), .B(new_n834), .Y(\f[52] ));
  NOR2xp33_ASAP7_75t_L      g0452(.A(\a[53] ), .B(\b[53] ), .Y(new_n838));
  NAND2xp33_ASAP7_75t_L     g0453(.A(\b[53] ), .B(\a[53] ), .Y(new_n839));
  INVx1_ASAP7_75t_L         g0454(.A(new_n839), .Y(new_n840));
  NOR2xp33_ASAP7_75t_L      g0455(.A(new_n838), .B(new_n840), .Y(new_n841));
  A2O1A1O1Ixp25_ASAP7_75t_L g0456(.A1(new_n822), .A2(new_n824), .B(new_n821), .C(new_n830), .D(new_n829), .Y(new_n842));
  XNOR2x2_ASAP7_75t_L       g0457(.A(new_n841), .B(new_n842), .Y(\f[53] ));
  NOR2xp33_ASAP7_75t_L      g0458(.A(\a[54] ), .B(\b[54] ), .Y(new_n844));
  INVx1_ASAP7_75t_L         g0459(.A(\a[54] ), .Y(new_n845));
  INVx1_ASAP7_75t_L         g0460(.A(\b[54] ), .Y(new_n846));
  NOR2xp33_ASAP7_75t_L      g0461(.A(new_n845), .B(new_n846), .Y(new_n847));
  NOR2xp33_ASAP7_75t_L      g0462(.A(new_n844), .B(new_n847), .Y(new_n848));
  INVx1_ASAP7_75t_L         g0463(.A(new_n829), .Y(new_n849));
  A2O1A1Ixp33_ASAP7_75t_L   g0464(.A1(new_n835), .A2(new_n849), .B(new_n838), .C(new_n839), .Y(new_n850));
  XOR2x2_ASAP7_75t_L        g0465(.A(new_n848), .B(new_n850), .Y(\f[54] ));
  NOR2xp33_ASAP7_75t_L      g0466(.A(\a[55] ), .B(\b[55] ), .Y(new_n852));
  INVx1_ASAP7_75t_L         g0467(.A(\a[55] ), .Y(new_n853));
  INVx1_ASAP7_75t_L         g0468(.A(\b[55] ), .Y(new_n854));
  NOR2xp33_ASAP7_75t_L      g0469(.A(new_n853), .B(new_n854), .Y(new_n855));
  NOR2xp33_ASAP7_75t_L      g0470(.A(new_n852), .B(new_n855), .Y(new_n856));
  A2O1A1Ixp33_ASAP7_75t_L   g0471(.A1(new_n833), .A2(new_n830), .B(new_n829), .C(new_n841), .Y(new_n857));
  INVx1_ASAP7_75t_L         g0472(.A(new_n847), .Y(new_n858));
  A2O1A1Ixp33_ASAP7_75t_L   g0473(.A1(new_n857), .A2(new_n839), .B(new_n844), .C(new_n858), .Y(new_n859));
  NOR2xp33_ASAP7_75t_L      g0474(.A(new_n856), .B(new_n859), .Y(new_n860));
  A2O1A1Ixp33_ASAP7_75t_L   g0475(.A1(new_n850), .A2(new_n848), .B(new_n847), .C(new_n856), .Y(new_n861));
  INVx1_ASAP7_75t_L         g0476(.A(new_n861), .Y(new_n862));
  NOR2xp33_ASAP7_75t_L      g0477(.A(new_n862), .B(new_n860), .Y(\f[55] ));
  NOR2xp33_ASAP7_75t_L      g0478(.A(\a[56] ), .B(\b[56] ), .Y(new_n864));
  NAND2xp33_ASAP7_75t_L     g0479(.A(\b[56] ), .B(\a[56] ), .Y(new_n865));
  INVx1_ASAP7_75t_L         g0480(.A(new_n865), .Y(new_n866));
  NOR2xp33_ASAP7_75t_L      g0481(.A(new_n864), .B(new_n866), .Y(new_n867));
  A2O1A1O1Ixp25_ASAP7_75t_L g0482(.A1(new_n848), .A2(new_n850), .B(new_n847), .C(new_n856), .D(new_n855), .Y(new_n868));
  XNOR2x2_ASAP7_75t_L       g0483(.A(new_n867), .B(new_n868), .Y(\f[56] ));
  NOR2xp33_ASAP7_75t_L      g0484(.A(\a[57] ), .B(\b[57] ), .Y(new_n870));
  INVx1_ASAP7_75t_L         g0485(.A(\a[57] ), .Y(new_n871));
  INVx1_ASAP7_75t_L         g0486(.A(\b[57] ), .Y(new_n872));
  NOR2xp33_ASAP7_75t_L      g0487(.A(new_n871), .B(new_n872), .Y(new_n873));
  NOR2xp33_ASAP7_75t_L      g0488(.A(new_n870), .B(new_n873), .Y(new_n874));
  INVx1_ASAP7_75t_L         g0489(.A(new_n855), .Y(new_n875));
  A2O1A1Ixp33_ASAP7_75t_L   g0490(.A1(new_n861), .A2(new_n875), .B(new_n864), .C(new_n865), .Y(new_n876));
  XOR2x2_ASAP7_75t_L        g0491(.A(new_n874), .B(new_n876), .Y(\f[57] ));
  NOR2xp33_ASAP7_75t_L      g0492(.A(\a[58] ), .B(\b[58] ), .Y(new_n878));
  INVx1_ASAP7_75t_L         g0493(.A(\a[58] ), .Y(new_n879));
  INVx1_ASAP7_75t_L         g0494(.A(\b[58] ), .Y(new_n880));
  NOR2xp33_ASAP7_75t_L      g0495(.A(new_n879), .B(new_n880), .Y(new_n881));
  NOR2xp33_ASAP7_75t_L      g0496(.A(new_n878), .B(new_n881), .Y(new_n882));
  A2O1A1Ixp33_ASAP7_75t_L   g0497(.A1(new_n859), .A2(new_n856), .B(new_n855), .C(new_n867), .Y(new_n883));
  INVx1_ASAP7_75t_L         g0498(.A(new_n873), .Y(new_n884));
  A2O1A1Ixp33_ASAP7_75t_L   g0499(.A1(new_n883), .A2(new_n865), .B(new_n870), .C(new_n884), .Y(new_n885));
  NOR2xp33_ASAP7_75t_L      g0500(.A(new_n882), .B(new_n885), .Y(new_n886));
  A2O1A1Ixp33_ASAP7_75t_L   g0501(.A1(new_n876), .A2(new_n874), .B(new_n873), .C(new_n882), .Y(new_n887));
  INVx1_ASAP7_75t_L         g0502(.A(new_n887), .Y(new_n888));
  NOR2xp33_ASAP7_75t_L      g0503(.A(new_n888), .B(new_n886), .Y(\f[58] ));
  NOR2xp33_ASAP7_75t_L      g0504(.A(\a[59] ), .B(\b[59] ), .Y(new_n890));
  NAND2xp33_ASAP7_75t_L     g0505(.A(\b[59] ), .B(\a[59] ), .Y(new_n891));
  INVx1_ASAP7_75t_L         g0506(.A(new_n891), .Y(new_n892));
  NOR2xp33_ASAP7_75t_L      g0507(.A(new_n890), .B(new_n892), .Y(new_n893));
  A2O1A1O1Ixp25_ASAP7_75t_L g0508(.A1(new_n874), .A2(new_n876), .B(new_n873), .C(new_n882), .D(new_n881), .Y(new_n894));
  XNOR2x2_ASAP7_75t_L       g0509(.A(new_n893), .B(new_n894), .Y(\f[59] ));
  NOR2xp33_ASAP7_75t_L      g0510(.A(\a[60] ), .B(\b[60] ), .Y(new_n896));
  INVx1_ASAP7_75t_L         g0511(.A(\a[60] ), .Y(new_n897));
  INVx1_ASAP7_75t_L         g0512(.A(\b[60] ), .Y(new_n898));
  NOR2xp33_ASAP7_75t_L      g0513(.A(new_n897), .B(new_n898), .Y(new_n899));
  NOR2xp33_ASAP7_75t_L      g0514(.A(new_n896), .B(new_n899), .Y(new_n900));
  INVx1_ASAP7_75t_L         g0515(.A(new_n881), .Y(new_n901));
  A2O1A1Ixp33_ASAP7_75t_L   g0516(.A1(new_n887), .A2(new_n901), .B(new_n890), .C(new_n891), .Y(new_n902));
  XOR2x2_ASAP7_75t_L        g0517(.A(new_n900), .B(new_n902), .Y(\f[60] ));
  NOR2xp33_ASAP7_75t_L      g0518(.A(\a[61] ), .B(\b[61] ), .Y(new_n904));
  INVx1_ASAP7_75t_L         g0519(.A(\a[61] ), .Y(new_n905));
  INVx1_ASAP7_75t_L         g0520(.A(\b[61] ), .Y(new_n906));
  NOR2xp33_ASAP7_75t_L      g0521(.A(new_n905), .B(new_n906), .Y(new_n907));
  NOR2xp33_ASAP7_75t_L      g0522(.A(new_n904), .B(new_n907), .Y(new_n908));
  A2O1A1Ixp33_ASAP7_75t_L   g0523(.A1(new_n885), .A2(new_n882), .B(new_n881), .C(new_n893), .Y(new_n909));
  INVx1_ASAP7_75t_L         g0524(.A(new_n899), .Y(new_n910));
  A2O1A1Ixp33_ASAP7_75t_L   g0525(.A1(new_n909), .A2(new_n891), .B(new_n896), .C(new_n910), .Y(new_n911));
  NOR2xp33_ASAP7_75t_L      g0526(.A(new_n908), .B(new_n911), .Y(new_n912));
  A2O1A1Ixp33_ASAP7_75t_L   g0527(.A1(new_n902), .A2(new_n900), .B(new_n899), .C(new_n908), .Y(new_n913));
  INVx1_ASAP7_75t_L         g0528(.A(new_n913), .Y(new_n914));
  NOR2xp33_ASAP7_75t_L      g0529(.A(new_n914), .B(new_n912), .Y(\f[61] ));
  NOR2xp33_ASAP7_75t_L      g0530(.A(\a[62] ), .B(\b[62] ), .Y(new_n916));
  NAND2xp33_ASAP7_75t_L     g0531(.A(\b[62] ), .B(\a[62] ), .Y(new_n917));
  INVx1_ASAP7_75t_L         g0532(.A(new_n917), .Y(new_n918));
  NOR2xp33_ASAP7_75t_L      g0533(.A(new_n916), .B(new_n918), .Y(new_n919));
  A2O1A1O1Ixp25_ASAP7_75t_L g0534(.A1(new_n900), .A2(new_n902), .B(new_n899), .C(new_n908), .D(new_n907), .Y(new_n920));
  XNOR2x2_ASAP7_75t_L       g0535(.A(new_n919), .B(new_n920), .Y(\f[62] ));
  NOR2xp33_ASAP7_75t_L      g0536(.A(\a[63] ), .B(\b[63] ), .Y(new_n922));
  INVx1_ASAP7_75t_L         g0537(.A(\a[63] ), .Y(new_n923));
  INVx1_ASAP7_75t_L         g0538(.A(\b[63] ), .Y(new_n924));
  NOR2xp33_ASAP7_75t_L      g0539(.A(new_n923), .B(new_n924), .Y(new_n925));
  NOR2xp33_ASAP7_75t_L      g0540(.A(new_n922), .B(new_n925), .Y(new_n926));
  INVx1_ASAP7_75t_L         g0541(.A(new_n907), .Y(new_n927));
  A2O1A1Ixp33_ASAP7_75t_L   g0542(.A1(new_n913), .A2(new_n927), .B(new_n916), .C(new_n917), .Y(new_n928));
  XOR2x2_ASAP7_75t_L        g0543(.A(new_n926), .B(new_n928), .Y(\f[63] ));
  NOR2xp33_ASAP7_75t_L      g0544(.A(\a[64] ), .B(\b[64] ), .Y(new_n930));
  INVx1_ASAP7_75t_L         g0545(.A(\a[64] ), .Y(new_n931));
  INVx1_ASAP7_75t_L         g0546(.A(\b[64] ), .Y(new_n932));
  NOR2xp33_ASAP7_75t_L      g0547(.A(new_n931), .B(new_n932), .Y(new_n933));
  NOR2xp33_ASAP7_75t_L      g0548(.A(new_n930), .B(new_n933), .Y(new_n934));
  A2O1A1Ixp33_ASAP7_75t_L   g0549(.A1(new_n911), .A2(new_n908), .B(new_n907), .C(new_n919), .Y(new_n935));
  INVx1_ASAP7_75t_L         g0550(.A(new_n925), .Y(new_n936));
  A2O1A1Ixp33_ASAP7_75t_L   g0551(.A1(new_n935), .A2(new_n917), .B(new_n922), .C(new_n936), .Y(new_n937));
  NOR2xp33_ASAP7_75t_L      g0552(.A(new_n934), .B(new_n937), .Y(new_n938));
  A2O1A1Ixp33_ASAP7_75t_L   g0553(.A1(new_n928), .A2(new_n926), .B(new_n925), .C(new_n934), .Y(new_n939));
  INVx1_ASAP7_75t_L         g0554(.A(new_n939), .Y(new_n940));
  NOR2xp33_ASAP7_75t_L      g0555(.A(new_n940), .B(new_n938), .Y(\f[64] ));
  NOR2xp33_ASAP7_75t_L      g0556(.A(\a[65] ), .B(\b[65] ), .Y(new_n942));
  NAND2xp33_ASAP7_75t_L     g0557(.A(\b[65] ), .B(\a[65] ), .Y(new_n943));
  INVx1_ASAP7_75t_L         g0558(.A(new_n943), .Y(new_n944));
  NOR2xp33_ASAP7_75t_L      g0559(.A(new_n942), .B(new_n944), .Y(new_n945));
  A2O1A1O1Ixp25_ASAP7_75t_L g0560(.A1(new_n926), .A2(new_n928), .B(new_n925), .C(new_n934), .D(new_n933), .Y(new_n946));
  XNOR2x2_ASAP7_75t_L       g0561(.A(new_n945), .B(new_n946), .Y(\f[65] ));
  NOR2xp33_ASAP7_75t_L      g0562(.A(\a[66] ), .B(\b[66] ), .Y(new_n948));
  INVx1_ASAP7_75t_L         g0563(.A(\a[66] ), .Y(new_n949));
  INVx1_ASAP7_75t_L         g0564(.A(\b[66] ), .Y(new_n950));
  NOR2xp33_ASAP7_75t_L      g0565(.A(new_n949), .B(new_n950), .Y(new_n951));
  NOR2xp33_ASAP7_75t_L      g0566(.A(new_n948), .B(new_n951), .Y(new_n952));
  INVx1_ASAP7_75t_L         g0567(.A(new_n933), .Y(new_n953));
  A2O1A1Ixp33_ASAP7_75t_L   g0568(.A1(new_n939), .A2(new_n953), .B(new_n942), .C(new_n943), .Y(new_n954));
  XOR2x2_ASAP7_75t_L        g0569(.A(new_n952), .B(new_n954), .Y(\f[66] ));
  NOR2xp33_ASAP7_75t_L      g0570(.A(\a[67] ), .B(\b[67] ), .Y(new_n956));
  INVx1_ASAP7_75t_L         g0571(.A(\a[67] ), .Y(new_n957));
  INVx1_ASAP7_75t_L         g0572(.A(\b[67] ), .Y(new_n958));
  NOR2xp33_ASAP7_75t_L      g0573(.A(new_n957), .B(new_n958), .Y(new_n959));
  NOR2xp33_ASAP7_75t_L      g0574(.A(new_n956), .B(new_n959), .Y(new_n960));
  A2O1A1Ixp33_ASAP7_75t_L   g0575(.A1(new_n937), .A2(new_n934), .B(new_n933), .C(new_n945), .Y(new_n961));
  INVx1_ASAP7_75t_L         g0576(.A(new_n951), .Y(new_n962));
  A2O1A1Ixp33_ASAP7_75t_L   g0577(.A1(new_n961), .A2(new_n943), .B(new_n948), .C(new_n962), .Y(new_n963));
  NOR2xp33_ASAP7_75t_L      g0578(.A(new_n960), .B(new_n963), .Y(new_n964));
  A2O1A1Ixp33_ASAP7_75t_L   g0579(.A1(new_n954), .A2(new_n952), .B(new_n951), .C(new_n960), .Y(new_n965));
  INVx1_ASAP7_75t_L         g0580(.A(new_n965), .Y(new_n966));
  NOR2xp33_ASAP7_75t_L      g0581(.A(new_n966), .B(new_n964), .Y(\f[67] ));
  NOR2xp33_ASAP7_75t_L      g0582(.A(\a[68] ), .B(\b[68] ), .Y(new_n968));
  NAND2xp33_ASAP7_75t_L     g0583(.A(\b[68] ), .B(\a[68] ), .Y(new_n969));
  INVx1_ASAP7_75t_L         g0584(.A(new_n969), .Y(new_n970));
  NOR2xp33_ASAP7_75t_L      g0585(.A(new_n968), .B(new_n970), .Y(new_n971));
  A2O1A1O1Ixp25_ASAP7_75t_L g0586(.A1(new_n952), .A2(new_n954), .B(new_n951), .C(new_n960), .D(new_n959), .Y(new_n972));
  XNOR2x2_ASAP7_75t_L       g0587(.A(new_n971), .B(new_n972), .Y(\f[68] ));
  NOR2xp33_ASAP7_75t_L      g0588(.A(\a[69] ), .B(\b[69] ), .Y(new_n974));
  INVx1_ASAP7_75t_L         g0589(.A(\a[69] ), .Y(new_n975));
  INVx1_ASAP7_75t_L         g0590(.A(\b[69] ), .Y(new_n976));
  NOR2xp33_ASAP7_75t_L      g0591(.A(new_n975), .B(new_n976), .Y(new_n977));
  NOR2xp33_ASAP7_75t_L      g0592(.A(new_n974), .B(new_n977), .Y(new_n978));
  INVx1_ASAP7_75t_L         g0593(.A(new_n959), .Y(new_n979));
  A2O1A1Ixp33_ASAP7_75t_L   g0594(.A1(new_n965), .A2(new_n979), .B(new_n968), .C(new_n969), .Y(new_n980));
  XOR2x2_ASAP7_75t_L        g0595(.A(new_n978), .B(new_n980), .Y(\f[69] ));
  NOR2xp33_ASAP7_75t_L      g0596(.A(\a[70] ), .B(\b[70] ), .Y(new_n982));
  INVx1_ASAP7_75t_L         g0597(.A(\a[70] ), .Y(new_n983));
  INVx1_ASAP7_75t_L         g0598(.A(\b[70] ), .Y(new_n984));
  NOR2xp33_ASAP7_75t_L      g0599(.A(new_n983), .B(new_n984), .Y(new_n985));
  NOR2xp33_ASAP7_75t_L      g0600(.A(new_n982), .B(new_n985), .Y(new_n986));
  A2O1A1Ixp33_ASAP7_75t_L   g0601(.A1(new_n963), .A2(new_n960), .B(new_n959), .C(new_n971), .Y(new_n987));
  INVx1_ASAP7_75t_L         g0602(.A(new_n977), .Y(new_n988));
  A2O1A1Ixp33_ASAP7_75t_L   g0603(.A1(new_n987), .A2(new_n969), .B(new_n974), .C(new_n988), .Y(new_n989));
  NOR2xp33_ASAP7_75t_L      g0604(.A(new_n986), .B(new_n989), .Y(new_n990));
  A2O1A1Ixp33_ASAP7_75t_L   g0605(.A1(new_n980), .A2(new_n978), .B(new_n977), .C(new_n986), .Y(new_n991));
  INVx1_ASAP7_75t_L         g0606(.A(new_n991), .Y(new_n992));
  NOR2xp33_ASAP7_75t_L      g0607(.A(new_n992), .B(new_n990), .Y(\f[70] ));
  NOR2xp33_ASAP7_75t_L      g0608(.A(\a[71] ), .B(\b[71] ), .Y(new_n994));
  NAND2xp33_ASAP7_75t_L     g0609(.A(\b[71] ), .B(\a[71] ), .Y(new_n995));
  INVx1_ASAP7_75t_L         g0610(.A(new_n995), .Y(new_n996));
  NOR2xp33_ASAP7_75t_L      g0611(.A(new_n994), .B(new_n996), .Y(new_n997));
  A2O1A1O1Ixp25_ASAP7_75t_L g0612(.A1(new_n978), .A2(new_n980), .B(new_n977), .C(new_n986), .D(new_n985), .Y(new_n998));
  XNOR2x2_ASAP7_75t_L       g0613(.A(new_n997), .B(new_n998), .Y(\f[71] ));
  NOR2xp33_ASAP7_75t_L      g0614(.A(\a[72] ), .B(\b[72] ), .Y(new_n1000));
  INVx1_ASAP7_75t_L         g0615(.A(\a[72] ), .Y(new_n1001));
  INVx1_ASAP7_75t_L         g0616(.A(\b[72] ), .Y(new_n1002));
  NOR2xp33_ASAP7_75t_L      g0617(.A(new_n1001), .B(new_n1002), .Y(new_n1003));
  NOR2xp33_ASAP7_75t_L      g0618(.A(new_n1000), .B(new_n1003), .Y(new_n1004));
  INVx1_ASAP7_75t_L         g0619(.A(new_n985), .Y(new_n1005));
  A2O1A1Ixp33_ASAP7_75t_L   g0620(.A1(new_n991), .A2(new_n1005), .B(new_n994), .C(new_n995), .Y(new_n1006));
  XOR2x2_ASAP7_75t_L        g0621(.A(new_n1004), .B(new_n1006), .Y(\f[72] ));
  NOR2xp33_ASAP7_75t_L      g0622(.A(\a[73] ), .B(\b[73] ), .Y(new_n1008));
  INVx1_ASAP7_75t_L         g0623(.A(\a[73] ), .Y(new_n1009));
  INVx1_ASAP7_75t_L         g0624(.A(\b[73] ), .Y(new_n1010));
  NOR2xp33_ASAP7_75t_L      g0625(.A(new_n1009), .B(new_n1010), .Y(new_n1011));
  NOR2xp33_ASAP7_75t_L      g0626(.A(new_n1008), .B(new_n1011), .Y(new_n1012));
  A2O1A1Ixp33_ASAP7_75t_L   g0627(.A1(new_n989), .A2(new_n986), .B(new_n985), .C(new_n997), .Y(new_n1013));
  INVx1_ASAP7_75t_L         g0628(.A(new_n1003), .Y(new_n1014));
  A2O1A1Ixp33_ASAP7_75t_L   g0629(.A1(new_n1013), .A2(new_n995), .B(new_n1000), .C(new_n1014), .Y(new_n1015));
  NOR2xp33_ASAP7_75t_L      g0630(.A(new_n1012), .B(new_n1015), .Y(new_n1016));
  A2O1A1Ixp33_ASAP7_75t_L   g0631(.A1(new_n1006), .A2(new_n1004), .B(new_n1003), .C(new_n1012), .Y(new_n1017));
  INVx1_ASAP7_75t_L         g0632(.A(new_n1017), .Y(new_n1018));
  NOR2xp33_ASAP7_75t_L      g0633(.A(new_n1018), .B(new_n1016), .Y(\f[73] ));
  NOR2xp33_ASAP7_75t_L      g0634(.A(\a[74] ), .B(\b[74] ), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g0635(.A(\b[74] ), .B(\a[74] ), .Y(new_n1021));
  INVx1_ASAP7_75t_L         g0636(.A(new_n1021), .Y(new_n1022));
  NOR2xp33_ASAP7_75t_L      g0637(.A(new_n1020), .B(new_n1022), .Y(new_n1023));
  A2O1A1O1Ixp25_ASAP7_75t_L g0638(.A1(new_n1004), .A2(new_n1006), .B(new_n1003), .C(new_n1012), .D(new_n1011), .Y(new_n1024));
  XNOR2x2_ASAP7_75t_L       g0639(.A(new_n1023), .B(new_n1024), .Y(\f[74] ));
  NOR2xp33_ASAP7_75t_L      g0640(.A(\a[75] ), .B(\b[75] ), .Y(new_n1026));
  INVx1_ASAP7_75t_L         g0641(.A(\a[75] ), .Y(new_n1027));
  INVx1_ASAP7_75t_L         g0642(.A(\b[75] ), .Y(new_n1028));
  NOR2xp33_ASAP7_75t_L      g0643(.A(new_n1027), .B(new_n1028), .Y(new_n1029));
  NOR2xp33_ASAP7_75t_L      g0644(.A(new_n1026), .B(new_n1029), .Y(new_n1030));
  INVx1_ASAP7_75t_L         g0645(.A(new_n1011), .Y(new_n1031));
  A2O1A1Ixp33_ASAP7_75t_L   g0646(.A1(new_n1017), .A2(new_n1031), .B(new_n1020), .C(new_n1021), .Y(new_n1032));
  XOR2x2_ASAP7_75t_L        g0647(.A(new_n1030), .B(new_n1032), .Y(\f[75] ));
  NOR2xp33_ASAP7_75t_L      g0648(.A(\a[76] ), .B(\b[76] ), .Y(new_n1034));
  INVx1_ASAP7_75t_L         g0649(.A(\a[76] ), .Y(new_n1035));
  INVx1_ASAP7_75t_L         g0650(.A(\b[76] ), .Y(new_n1036));
  NOR2xp33_ASAP7_75t_L      g0651(.A(new_n1035), .B(new_n1036), .Y(new_n1037));
  NOR2xp33_ASAP7_75t_L      g0652(.A(new_n1034), .B(new_n1037), .Y(new_n1038));
  A2O1A1Ixp33_ASAP7_75t_L   g0653(.A1(new_n1015), .A2(new_n1012), .B(new_n1011), .C(new_n1023), .Y(new_n1039));
  INVx1_ASAP7_75t_L         g0654(.A(new_n1029), .Y(new_n1040));
  A2O1A1Ixp33_ASAP7_75t_L   g0655(.A1(new_n1039), .A2(new_n1021), .B(new_n1026), .C(new_n1040), .Y(new_n1041));
  NOR2xp33_ASAP7_75t_L      g0656(.A(new_n1038), .B(new_n1041), .Y(new_n1042));
  A2O1A1Ixp33_ASAP7_75t_L   g0657(.A1(new_n1032), .A2(new_n1030), .B(new_n1029), .C(new_n1038), .Y(new_n1043));
  INVx1_ASAP7_75t_L         g0658(.A(new_n1043), .Y(new_n1044));
  NOR2xp33_ASAP7_75t_L      g0659(.A(new_n1044), .B(new_n1042), .Y(\f[76] ));
  NOR2xp33_ASAP7_75t_L      g0660(.A(\a[77] ), .B(\b[77] ), .Y(new_n1046));
  NAND2xp33_ASAP7_75t_L     g0661(.A(\b[77] ), .B(\a[77] ), .Y(new_n1047));
  INVx1_ASAP7_75t_L         g0662(.A(new_n1047), .Y(new_n1048));
  NOR2xp33_ASAP7_75t_L      g0663(.A(new_n1046), .B(new_n1048), .Y(new_n1049));
  A2O1A1O1Ixp25_ASAP7_75t_L g0664(.A1(new_n1030), .A2(new_n1032), .B(new_n1029), .C(new_n1038), .D(new_n1037), .Y(new_n1050));
  XNOR2x2_ASAP7_75t_L       g0665(.A(new_n1049), .B(new_n1050), .Y(\f[77] ));
  NOR2xp33_ASAP7_75t_L      g0666(.A(\a[78] ), .B(\b[78] ), .Y(new_n1052));
  INVx1_ASAP7_75t_L         g0667(.A(\a[78] ), .Y(new_n1053));
  INVx1_ASAP7_75t_L         g0668(.A(\b[78] ), .Y(new_n1054));
  NOR2xp33_ASAP7_75t_L      g0669(.A(new_n1053), .B(new_n1054), .Y(new_n1055));
  NOR2xp33_ASAP7_75t_L      g0670(.A(new_n1052), .B(new_n1055), .Y(new_n1056));
  INVx1_ASAP7_75t_L         g0671(.A(new_n1037), .Y(new_n1057));
  A2O1A1Ixp33_ASAP7_75t_L   g0672(.A1(new_n1043), .A2(new_n1057), .B(new_n1046), .C(new_n1047), .Y(new_n1058));
  XOR2x2_ASAP7_75t_L        g0673(.A(new_n1056), .B(new_n1058), .Y(\f[78] ));
  NOR2xp33_ASAP7_75t_L      g0674(.A(\a[79] ), .B(\b[79] ), .Y(new_n1060));
  INVx1_ASAP7_75t_L         g0675(.A(\a[79] ), .Y(new_n1061));
  INVx1_ASAP7_75t_L         g0676(.A(\b[79] ), .Y(new_n1062));
  NOR2xp33_ASAP7_75t_L      g0677(.A(new_n1061), .B(new_n1062), .Y(new_n1063));
  NOR2xp33_ASAP7_75t_L      g0678(.A(new_n1060), .B(new_n1063), .Y(new_n1064));
  A2O1A1Ixp33_ASAP7_75t_L   g0679(.A1(new_n1041), .A2(new_n1038), .B(new_n1037), .C(new_n1049), .Y(new_n1065));
  INVx1_ASAP7_75t_L         g0680(.A(new_n1055), .Y(new_n1066));
  A2O1A1Ixp33_ASAP7_75t_L   g0681(.A1(new_n1065), .A2(new_n1047), .B(new_n1052), .C(new_n1066), .Y(new_n1067));
  NOR2xp33_ASAP7_75t_L      g0682(.A(new_n1064), .B(new_n1067), .Y(new_n1068));
  A2O1A1Ixp33_ASAP7_75t_L   g0683(.A1(new_n1058), .A2(new_n1056), .B(new_n1055), .C(new_n1064), .Y(new_n1069));
  INVx1_ASAP7_75t_L         g0684(.A(new_n1069), .Y(new_n1070));
  NOR2xp33_ASAP7_75t_L      g0685(.A(new_n1070), .B(new_n1068), .Y(\f[79] ));
  NOR2xp33_ASAP7_75t_L      g0686(.A(\a[80] ), .B(\b[80] ), .Y(new_n1072));
  NAND2xp33_ASAP7_75t_L     g0687(.A(\b[80] ), .B(\a[80] ), .Y(new_n1073));
  INVx1_ASAP7_75t_L         g0688(.A(new_n1073), .Y(new_n1074));
  NOR2xp33_ASAP7_75t_L      g0689(.A(new_n1072), .B(new_n1074), .Y(new_n1075));
  A2O1A1O1Ixp25_ASAP7_75t_L g0690(.A1(new_n1056), .A2(new_n1058), .B(new_n1055), .C(new_n1064), .D(new_n1063), .Y(new_n1076));
  XNOR2x2_ASAP7_75t_L       g0691(.A(new_n1075), .B(new_n1076), .Y(\f[80] ));
  NOR2xp33_ASAP7_75t_L      g0692(.A(\a[81] ), .B(\b[81] ), .Y(new_n1078));
  INVx1_ASAP7_75t_L         g0693(.A(\a[81] ), .Y(new_n1079));
  INVx1_ASAP7_75t_L         g0694(.A(\b[81] ), .Y(new_n1080));
  NOR2xp33_ASAP7_75t_L      g0695(.A(new_n1079), .B(new_n1080), .Y(new_n1081));
  NOR2xp33_ASAP7_75t_L      g0696(.A(new_n1078), .B(new_n1081), .Y(new_n1082));
  INVx1_ASAP7_75t_L         g0697(.A(new_n1063), .Y(new_n1083));
  A2O1A1Ixp33_ASAP7_75t_L   g0698(.A1(new_n1069), .A2(new_n1083), .B(new_n1072), .C(new_n1073), .Y(new_n1084));
  XOR2x2_ASAP7_75t_L        g0699(.A(new_n1082), .B(new_n1084), .Y(\f[81] ));
  NOR2xp33_ASAP7_75t_L      g0700(.A(\a[82] ), .B(\b[82] ), .Y(new_n1086));
  INVx1_ASAP7_75t_L         g0701(.A(\a[82] ), .Y(new_n1087));
  INVx1_ASAP7_75t_L         g0702(.A(\b[82] ), .Y(new_n1088));
  NOR2xp33_ASAP7_75t_L      g0703(.A(new_n1087), .B(new_n1088), .Y(new_n1089));
  NOR2xp33_ASAP7_75t_L      g0704(.A(new_n1086), .B(new_n1089), .Y(new_n1090));
  A2O1A1Ixp33_ASAP7_75t_L   g0705(.A1(new_n1067), .A2(new_n1064), .B(new_n1063), .C(new_n1075), .Y(new_n1091));
  INVx1_ASAP7_75t_L         g0706(.A(new_n1081), .Y(new_n1092));
  A2O1A1Ixp33_ASAP7_75t_L   g0707(.A1(new_n1091), .A2(new_n1073), .B(new_n1078), .C(new_n1092), .Y(new_n1093));
  NOR2xp33_ASAP7_75t_L      g0708(.A(new_n1090), .B(new_n1093), .Y(new_n1094));
  A2O1A1Ixp33_ASAP7_75t_L   g0709(.A1(new_n1084), .A2(new_n1082), .B(new_n1081), .C(new_n1090), .Y(new_n1095));
  INVx1_ASAP7_75t_L         g0710(.A(new_n1095), .Y(new_n1096));
  NOR2xp33_ASAP7_75t_L      g0711(.A(new_n1096), .B(new_n1094), .Y(\f[82] ));
  NOR2xp33_ASAP7_75t_L      g0712(.A(\a[83] ), .B(\b[83] ), .Y(new_n1098));
  NAND2xp33_ASAP7_75t_L     g0713(.A(\b[83] ), .B(\a[83] ), .Y(new_n1099));
  INVx1_ASAP7_75t_L         g0714(.A(new_n1099), .Y(new_n1100));
  NOR2xp33_ASAP7_75t_L      g0715(.A(new_n1098), .B(new_n1100), .Y(new_n1101));
  A2O1A1O1Ixp25_ASAP7_75t_L g0716(.A1(new_n1082), .A2(new_n1084), .B(new_n1081), .C(new_n1090), .D(new_n1089), .Y(new_n1102));
  XNOR2x2_ASAP7_75t_L       g0717(.A(new_n1101), .B(new_n1102), .Y(\f[83] ));
  NOR2xp33_ASAP7_75t_L      g0718(.A(\a[84] ), .B(\b[84] ), .Y(new_n1104));
  INVx1_ASAP7_75t_L         g0719(.A(\a[84] ), .Y(new_n1105));
  INVx1_ASAP7_75t_L         g0720(.A(\b[84] ), .Y(new_n1106));
  NOR2xp33_ASAP7_75t_L      g0721(.A(new_n1105), .B(new_n1106), .Y(new_n1107));
  NOR2xp33_ASAP7_75t_L      g0722(.A(new_n1104), .B(new_n1107), .Y(new_n1108));
  INVx1_ASAP7_75t_L         g0723(.A(new_n1089), .Y(new_n1109));
  A2O1A1Ixp33_ASAP7_75t_L   g0724(.A1(new_n1095), .A2(new_n1109), .B(new_n1098), .C(new_n1099), .Y(new_n1110));
  XOR2x2_ASAP7_75t_L        g0725(.A(new_n1108), .B(new_n1110), .Y(\f[84] ));
  NOR2xp33_ASAP7_75t_L      g0726(.A(\a[85] ), .B(\b[85] ), .Y(new_n1112));
  INVx1_ASAP7_75t_L         g0727(.A(\a[85] ), .Y(new_n1113));
  INVx1_ASAP7_75t_L         g0728(.A(\b[85] ), .Y(new_n1114));
  NOR2xp33_ASAP7_75t_L      g0729(.A(new_n1113), .B(new_n1114), .Y(new_n1115));
  NOR2xp33_ASAP7_75t_L      g0730(.A(new_n1112), .B(new_n1115), .Y(new_n1116));
  A2O1A1Ixp33_ASAP7_75t_L   g0731(.A1(new_n1093), .A2(new_n1090), .B(new_n1089), .C(new_n1101), .Y(new_n1117));
  INVx1_ASAP7_75t_L         g0732(.A(new_n1107), .Y(new_n1118));
  A2O1A1Ixp33_ASAP7_75t_L   g0733(.A1(new_n1117), .A2(new_n1099), .B(new_n1104), .C(new_n1118), .Y(new_n1119));
  NOR2xp33_ASAP7_75t_L      g0734(.A(new_n1116), .B(new_n1119), .Y(new_n1120));
  A2O1A1Ixp33_ASAP7_75t_L   g0735(.A1(new_n1110), .A2(new_n1108), .B(new_n1107), .C(new_n1116), .Y(new_n1121));
  INVx1_ASAP7_75t_L         g0736(.A(new_n1121), .Y(new_n1122));
  NOR2xp33_ASAP7_75t_L      g0737(.A(new_n1122), .B(new_n1120), .Y(\f[85] ));
  NOR2xp33_ASAP7_75t_L      g0738(.A(\a[86] ), .B(\b[86] ), .Y(new_n1124));
  NAND2xp33_ASAP7_75t_L     g0739(.A(\b[86] ), .B(\a[86] ), .Y(new_n1125));
  INVx1_ASAP7_75t_L         g0740(.A(new_n1125), .Y(new_n1126));
  NOR2xp33_ASAP7_75t_L      g0741(.A(new_n1124), .B(new_n1126), .Y(new_n1127));
  A2O1A1O1Ixp25_ASAP7_75t_L g0742(.A1(new_n1108), .A2(new_n1110), .B(new_n1107), .C(new_n1116), .D(new_n1115), .Y(new_n1128));
  XNOR2x2_ASAP7_75t_L       g0743(.A(new_n1127), .B(new_n1128), .Y(\f[86] ));
  NOR2xp33_ASAP7_75t_L      g0744(.A(\a[87] ), .B(\b[87] ), .Y(new_n1130));
  INVx1_ASAP7_75t_L         g0745(.A(\a[87] ), .Y(new_n1131));
  INVx1_ASAP7_75t_L         g0746(.A(\b[87] ), .Y(new_n1132));
  NOR2xp33_ASAP7_75t_L      g0747(.A(new_n1131), .B(new_n1132), .Y(new_n1133));
  NOR2xp33_ASAP7_75t_L      g0748(.A(new_n1130), .B(new_n1133), .Y(new_n1134));
  INVx1_ASAP7_75t_L         g0749(.A(new_n1115), .Y(new_n1135));
  A2O1A1Ixp33_ASAP7_75t_L   g0750(.A1(new_n1121), .A2(new_n1135), .B(new_n1124), .C(new_n1125), .Y(new_n1136));
  XOR2x2_ASAP7_75t_L        g0751(.A(new_n1134), .B(new_n1136), .Y(\f[87] ));
  NOR2xp33_ASAP7_75t_L      g0752(.A(\a[88] ), .B(\b[88] ), .Y(new_n1138));
  INVx1_ASAP7_75t_L         g0753(.A(\a[88] ), .Y(new_n1139));
  INVx1_ASAP7_75t_L         g0754(.A(\b[88] ), .Y(new_n1140));
  NOR2xp33_ASAP7_75t_L      g0755(.A(new_n1139), .B(new_n1140), .Y(new_n1141));
  NOR2xp33_ASAP7_75t_L      g0756(.A(new_n1138), .B(new_n1141), .Y(new_n1142));
  A2O1A1Ixp33_ASAP7_75t_L   g0757(.A1(new_n1119), .A2(new_n1116), .B(new_n1115), .C(new_n1127), .Y(new_n1143));
  INVx1_ASAP7_75t_L         g0758(.A(new_n1133), .Y(new_n1144));
  A2O1A1Ixp33_ASAP7_75t_L   g0759(.A1(new_n1143), .A2(new_n1125), .B(new_n1130), .C(new_n1144), .Y(new_n1145));
  NOR2xp33_ASAP7_75t_L      g0760(.A(new_n1142), .B(new_n1145), .Y(new_n1146));
  A2O1A1Ixp33_ASAP7_75t_L   g0761(.A1(new_n1136), .A2(new_n1134), .B(new_n1133), .C(new_n1142), .Y(new_n1147));
  INVx1_ASAP7_75t_L         g0762(.A(new_n1147), .Y(new_n1148));
  NOR2xp33_ASAP7_75t_L      g0763(.A(new_n1148), .B(new_n1146), .Y(\f[88] ));
  NOR2xp33_ASAP7_75t_L      g0764(.A(\a[89] ), .B(\b[89] ), .Y(new_n1150));
  NAND2xp33_ASAP7_75t_L     g0765(.A(\b[89] ), .B(\a[89] ), .Y(new_n1151));
  INVx1_ASAP7_75t_L         g0766(.A(new_n1151), .Y(new_n1152));
  NOR2xp33_ASAP7_75t_L      g0767(.A(new_n1150), .B(new_n1152), .Y(new_n1153));
  A2O1A1O1Ixp25_ASAP7_75t_L g0768(.A1(new_n1134), .A2(new_n1136), .B(new_n1133), .C(new_n1142), .D(new_n1141), .Y(new_n1154));
  XNOR2x2_ASAP7_75t_L       g0769(.A(new_n1153), .B(new_n1154), .Y(\f[89] ));
  NOR2xp33_ASAP7_75t_L      g0770(.A(\a[90] ), .B(\b[90] ), .Y(new_n1156));
  INVx1_ASAP7_75t_L         g0771(.A(\a[90] ), .Y(new_n1157));
  INVx1_ASAP7_75t_L         g0772(.A(\b[90] ), .Y(new_n1158));
  NOR2xp33_ASAP7_75t_L      g0773(.A(new_n1157), .B(new_n1158), .Y(new_n1159));
  NOR2xp33_ASAP7_75t_L      g0774(.A(new_n1156), .B(new_n1159), .Y(new_n1160));
  INVx1_ASAP7_75t_L         g0775(.A(new_n1141), .Y(new_n1161));
  A2O1A1Ixp33_ASAP7_75t_L   g0776(.A1(new_n1147), .A2(new_n1161), .B(new_n1150), .C(new_n1151), .Y(new_n1162));
  XOR2x2_ASAP7_75t_L        g0777(.A(new_n1160), .B(new_n1162), .Y(\f[90] ));
  NOR2xp33_ASAP7_75t_L      g0778(.A(\a[91] ), .B(\b[91] ), .Y(new_n1164));
  INVx1_ASAP7_75t_L         g0779(.A(\a[91] ), .Y(new_n1165));
  INVx1_ASAP7_75t_L         g0780(.A(\b[91] ), .Y(new_n1166));
  NOR2xp33_ASAP7_75t_L      g0781(.A(new_n1165), .B(new_n1166), .Y(new_n1167));
  NOR2xp33_ASAP7_75t_L      g0782(.A(new_n1164), .B(new_n1167), .Y(new_n1168));
  A2O1A1Ixp33_ASAP7_75t_L   g0783(.A1(new_n1145), .A2(new_n1142), .B(new_n1141), .C(new_n1153), .Y(new_n1169));
  INVx1_ASAP7_75t_L         g0784(.A(new_n1159), .Y(new_n1170));
  A2O1A1Ixp33_ASAP7_75t_L   g0785(.A1(new_n1169), .A2(new_n1151), .B(new_n1156), .C(new_n1170), .Y(new_n1171));
  NOR2xp33_ASAP7_75t_L      g0786(.A(new_n1168), .B(new_n1171), .Y(new_n1172));
  A2O1A1Ixp33_ASAP7_75t_L   g0787(.A1(new_n1162), .A2(new_n1160), .B(new_n1159), .C(new_n1168), .Y(new_n1173));
  INVx1_ASAP7_75t_L         g0788(.A(new_n1173), .Y(new_n1174));
  NOR2xp33_ASAP7_75t_L      g0789(.A(new_n1174), .B(new_n1172), .Y(\f[91] ));
  NOR2xp33_ASAP7_75t_L      g0790(.A(\a[92] ), .B(\b[92] ), .Y(new_n1176));
  NAND2xp33_ASAP7_75t_L     g0791(.A(\b[92] ), .B(\a[92] ), .Y(new_n1177));
  INVx1_ASAP7_75t_L         g0792(.A(new_n1177), .Y(new_n1178));
  NOR2xp33_ASAP7_75t_L      g0793(.A(new_n1176), .B(new_n1178), .Y(new_n1179));
  A2O1A1O1Ixp25_ASAP7_75t_L g0794(.A1(new_n1160), .A2(new_n1162), .B(new_n1159), .C(new_n1168), .D(new_n1167), .Y(new_n1180));
  XNOR2x2_ASAP7_75t_L       g0795(.A(new_n1179), .B(new_n1180), .Y(\f[92] ));
  NOR2xp33_ASAP7_75t_L      g0796(.A(\a[93] ), .B(\b[93] ), .Y(new_n1182));
  INVx1_ASAP7_75t_L         g0797(.A(\a[93] ), .Y(new_n1183));
  INVx1_ASAP7_75t_L         g0798(.A(\b[93] ), .Y(new_n1184));
  NOR2xp33_ASAP7_75t_L      g0799(.A(new_n1183), .B(new_n1184), .Y(new_n1185));
  NOR2xp33_ASAP7_75t_L      g0800(.A(new_n1182), .B(new_n1185), .Y(new_n1186));
  INVx1_ASAP7_75t_L         g0801(.A(new_n1167), .Y(new_n1187));
  A2O1A1Ixp33_ASAP7_75t_L   g0802(.A1(new_n1173), .A2(new_n1187), .B(new_n1176), .C(new_n1177), .Y(new_n1188));
  XOR2x2_ASAP7_75t_L        g0803(.A(new_n1186), .B(new_n1188), .Y(\f[93] ));
  NOR2xp33_ASAP7_75t_L      g0804(.A(\a[94] ), .B(\b[94] ), .Y(new_n1190));
  INVx1_ASAP7_75t_L         g0805(.A(\a[94] ), .Y(new_n1191));
  INVx1_ASAP7_75t_L         g0806(.A(\b[94] ), .Y(new_n1192));
  NOR2xp33_ASAP7_75t_L      g0807(.A(new_n1191), .B(new_n1192), .Y(new_n1193));
  NOR2xp33_ASAP7_75t_L      g0808(.A(new_n1190), .B(new_n1193), .Y(new_n1194));
  A2O1A1Ixp33_ASAP7_75t_L   g0809(.A1(new_n1171), .A2(new_n1168), .B(new_n1167), .C(new_n1179), .Y(new_n1195));
  INVx1_ASAP7_75t_L         g0810(.A(new_n1185), .Y(new_n1196));
  A2O1A1Ixp33_ASAP7_75t_L   g0811(.A1(new_n1195), .A2(new_n1177), .B(new_n1182), .C(new_n1196), .Y(new_n1197));
  NOR2xp33_ASAP7_75t_L      g0812(.A(new_n1194), .B(new_n1197), .Y(new_n1198));
  A2O1A1Ixp33_ASAP7_75t_L   g0813(.A1(new_n1188), .A2(new_n1186), .B(new_n1185), .C(new_n1194), .Y(new_n1199));
  INVx1_ASAP7_75t_L         g0814(.A(new_n1199), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g0815(.A(new_n1200), .B(new_n1198), .Y(\f[94] ));
  NOR2xp33_ASAP7_75t_L      g0816(.A(\a[95] ), .B(\b[95] ), .Y(new_n1202));
  NAND2xp33_ASAP7_75t_L     g0817(.A(\b[95] ), .B(\a[95] ), .Y(new_n1203));
  INVx1_ASAP7_75t_L         g0818(.A(new_n1203), .Y(new_n1204));
  NOR2xp33_ASAP7_75t_L      g0819(.A(new_n1202), .B(new_n1204), .Y(new_n1205));
  A2O1A1O1Ixp25_ASAP7_75t_L g0820(.A1(new_n1186), .A2(new_n1188), .B(new_n1185), .C(new_n1194), .D(new_n1193), .Y(new_n1206));
  XNOR2x2_ASAP7_75t_L       g0821(.A(new_n1205), .B(new_n1206), .Y(\f[95] ));
  NOR2xp33_ASAP7_75t_L      g0822(.A(\a[96] ), .B(\b[96] ), .Y(new_n1208));
  INVx1_ASAP7_75t_L         g0823(.A(\a[96] ), .Y(new_n1209));
  INVx1_ASAP7_75t_L         g0824(.A(\b[96] ), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g0825(.A(new_n1209), .B(new_n1210), .Y(new_n1211));
  NOR2xp33_ASAP7_75t_L      g0826(.A(new_n1208), .B(new_n1211), .Y(new_n1212));
  INVx1_ASAP7_75t_L         g0827(.A(new_n1193), .Y(new_n1213));
  A2O1A1Ixp33_ASAP7_75t_L   g0828(.A1(new_n1199), .A2(new_n1213), .B(new_n1202), .C(new_n1203), .Y(new_n1214));
  XOR2x2_ASAP7_75t_L        g0829(.A(new_n1212), .B(new_n1214), .Y(\f[96] ));
  NOR2xp33_ASAP7_75t_L      g0830(.A(\a[97] ), .B(\b[97] ), .Y(new_n1216));
  INVx1_ASAP7_75t_L         g0831(.A(\a[97] ), .Y(new_n1217));
  INVx1_ASAP7_75t_L         g0832(.A(\b[97] ), .Y(new_n1218));
  NOR2xp33_ASAP7_75t_L      g0833(.A(new_n1217), .B(new_n1218), .Y(new_n1219));
  NOR2xp33_ASAP7_75t_L      g0834(.A(new_n1216), .B(new_n1219), .Y(new_n1220));
  A2O1A1Ixp33_ASAP7_75t_L   g0835(.A1(new_n1197), .A2(new_n1194), .B(new_n1193), .C(new_n1205), .Y(new_n1221));
  INVx1_ASAP7_75t_L         g0836(.A(new_n1211), .Y(new_n1222));
  A2O1A1Ixp33_ASAP7_75t_L   g0837(.A1(new_n1221), .A2(new_n1203), .B(new_n1208), .C(new_n1222), .Y(new_n1223));
  NOR2xp33_ASAP7_75t_L      g0838(.A(new_n1220), .B(new_n1223), .Y(new_n1224));
  A2O1A1Ixp33_ASAP7_75t_L   g0839(.A1(new_n1214), .A2(new_n1212), .B(new_n1211), .C(new_n1220), .Y(new_n1225));
  INVx1_ASAP7_75t_L         g0840(.A(new_n1225), .Y(new_n1226));
  NOR2xp33_ASAP7_75t_L      g0841(.A(new_n1226), .B(new_n1224), .Y(\f[97] ));
  NOR2xp33_ASAP7_75t_L      g0842(.A(\a[98] ), .B(\b[98] ), .Y(new_n1228));
  NAND2xp33_ASAP7_75t_L     g0843(.A(\b[98] ), .B(\a[98] ), .Y(new_n1229));
  INVx1_ASAP7_75t_L         g0844(.A(new_n1229), .Y(new_n1230));
  NOR2xp33_ASAP7_75t_L      g0845(.A(new_n1228), .B(new_n1230), .Y(new_n1231));
  A2O1A1O1Ixp25_ASAP7_75t_L g0846(.A1(new_n1212), .A2(new_n1214), .B(new_n1211), .C(new_n1220), .D(new_n1219), .Y(new_n1232));
  XNOR2x2_ASAP7_75t_L       g0847(.A(new_n1231), .B(new_n1232), .Y(\f[98] ));
  NOR2xp33_ASAP7_75t_L      g0848(.A(\a[99] ), .B(\b[99] ), .Y(new_n1234));
  INVx1_ASAP7_75t_L         g0849(.A(\a[99] ), .Y(new_n1235));
  INVx1_ASAP7_75t_L         g0850(.A(\b[99] ), .Y(new_n1236));
  NOR2xp33_ASAP7_75t_L      g0851(.A(new_n1235), .B(new_n1236), .Y(new_n1237));
  NOR2xp33_ASAP7_75t_L      g0852(.A(new_n1234), .B(new_n1237), .Y(new_n1238));
  INVx1_ASAP7_75t_L         g0853(.A(new_n1219), .Y(new_n1239));
  A2O1A1Ixp33_ASAP7_75t_L   g0854(.A1(new_n1225), .A2(new_n1239), .B(new_n1228), .C(new_n1229), .Y(new_n1240));
  XOR2x2_ASAP7_75t_L        g0855(.A(new_n1238), .B(new_n1240), .Y(\f[99] ));
  NOR2xp33_ASAP7_75t_L      g0856(.A(\a[100] ), .B(\b[100] ), .Y(new_n1242));
  INVx1_ASAP7_75t_L         g0857(.A(\a[100] ), .Y(new_n1243));
  INVx1_ASAP7_75t_L         g0858(.A(\b[100] ), .Y(new_n1244));
  NOR2xp33_ASAP7_75t_L      g0859(.A(new_n1243), .B(new_n1244), .Y(new_n1245));
  NOR2xp33_ASAP7_75t_L      g0860(.A(new_n1242), .B(new_n1245), .Y(new_n1246));
  A2O1A1Ixp33_ASAP7_75t_L   g0861(.A1(new_n1223), .A2(new_n1220), .B(new_n1219), .C(new_n1231), .Y(new_n1247));
  INVx1_ASAP7_75t_L         g0862(.A(new_n1237), .Y(new_n1248));
  A2O1A1Ixp33_ASAP7_75t_L   g0863(.A1(new_n1247), .A2(new_n1229), .B(new_n1234), .C(new_n1248), .Y(new_n1249));
  NOR2xp33_ASAP7_75t_L      g0864(.A(new_n1246), .B(new_n1249), .Y(new_n1250));
  A2O1A1Ixp33_ASAP7_75t_L   g0865(.A1(new_n1240), .A2(new_n1238), .B(new_n1237), .C(new_n1246), .Y(new_n1251));
  INVx1_ASAP7_75t_L         g0866(.A(new_n1251), .Y(new_n1252));
  NOR2xp33_ASAP7_75t_L      g0867(.A(new_n1252), .B(new_n1250), .Y(\f[100] ));
  NOR2xp33_ASAP7_75t_L      g0868(.A(\a[101] ), .B(\b[101] ), .Y(new_n1254));
  NAND2xp33_ASAP7_75t_L     g0869(.A(\b[101] ), .B(\a[101] ), .Y(new_n1255));
  INVx1_ASAP7_75t_L         g0870(.A(new_n1255), .Y(new_n1256));
  NOR2xp33_ASAP7_75t_L      g0871(.A(new_n1254), .B(new_n1256), .Y(new_n1257));
  A2O1A1O1Ixp25_ASAP7_75t_L g0872(.A1(new_n1238), .A2(new_n1240), .B(new_n1237), .C(new_n1246), .D(new_n1245), .Y(new_n1258));
  XNOR2x2_ASAP7_75t_L       g0873(.A(new_n1257), .B(new_n1258), .Y(\f[101] ));
  NOR2xp33_ASAP7_75t_L      g0874(.A(\a[102] ), .B(\b[102] ), .Y(new_n1260));
  INVx1_ASAP7_75t_L         g0875(.A(\a[102] ), .Y(new_n1261));
  INVx1_ASAP7_75t_L         g0876(.A(\b[102] ), .Y(new_n1262));
  NOR2xp33_ASAP7_75t_L      g0877(.A(new_n1261), .B(new_n1262), .Y(new_n1263));
  NOR2xp33_ASAP7_75t_L      g0878(.A(new_n1260), .B(new_n1263), .Y(new_n1264));
  INVx1_ASAP7_75t_L         g0879(.A(new_n1245), .Y(new_n1265));
  A2O1A1Ixp33_ASAP7_75t_L   g0880(.A1(new_n1251), .A2(new_n1265), .B(new_n1254), .C(new_n1255), .Y(new_n1266));
  XOR2x2_ASAP7_75t_L        g0881(.A(new_n1264), .B(new_n1266), .Y(\f[102] ));
  NOR2xp33_ASAP7_75t_L      g0882(.A(\a[103] ), .B(\b[103] ), .Y(new_n1268));
  INVx1_ASAP7_75t_L         g0883(.A(\a[103] ), .Y(new_n1269));
  INVx1_ASAP7_75t_L         g0884(.A(\b[103] ), .Y(new_n1270));
  NOR2xp33_ASAP7_75t_L      g0885(.A(new_n1269), .B(new_n1270), .Y(new_n1271));
  NOR2xp33_ASAP7_75t_L      g0886(.A(new_n1268), .B(new_n1271), .Y(new_n1272));
  A2O1A1Ixp33_ASAP7_75t_L   g0887(.A1(new_n1249), .A2(new_n1246), .B(new_n1245), .C(new_n1257), .Y(new_n1273));
  INVx1_ASAP7_75t_L         g0888(.A(new_n1263), .Y(new_n1274));
  A2O1A1Ixp33_ASAP7_75t_L   g0889(.A1(new_n1273), .A2(new_n1255), .B(new_n1260), .C(new_n1274), .Y(new_n1275));
  NOR2xp33_ASAP7_75t_L      g0890(.A(new_n1272), .B(new_n1275), .Y(new_n1276));
  A2O1A1Ixp33_ASAP7_75t_L   g0891(.A1(new_n1266), .A2(new_n1264), .B(new_n1263), .C(new_n1272), .Y(new_n1277));
  INVx1_ASAP7_75t_L         g0892(.A(new_n1277), .Y(new_n1278));
  NOR2xp33_ASAP7_75t_L      g0893(.A(new_n1278), .B(new_n1276), .Y(\f[103] ));
  NOR2xp33_ASAP7_75t_L      g0894(.A(\a[104] ), .B(\b[104] ), .Y(new_n1280));
  NAND2xp33_ASAP7_75t_L     g0895(.A(\b[104] ), .B(\a[104] ), .Y(new_n1281));
  INVx1_ASAP7_75t_L         g0896(.A(new_n1281), .Y(new_n1282));
  NOR2xp33_ASAP7_75t_L      g0897(.A(new_n1280), .B(new_n1282), .Y(new_n1283));
  A2O1A1O1Ixp25_ASAP7_75t_L g0898(.A1(new_n1264), .A2(new_n1266), .B(new_n1263), .C(new_n1272), .D(new_n1271), .Y(new_n1284));
  XNOR2x2_ASAP7_75t_L       g0899(.A(new_n1283), .B(new_n1284), .Y(\f[104] ));
  NOR2xp33_ASAP7_75t_L      g0900(.A(\a[105] ), .B(\b[105] ), .Y(new_n1286));
  INVx1_ASAP7_75t_L         g0901(.A(\a[105] ), .Y(new_n1287));
  INVx1_ASAP7_75t_L         g0902(.A(\b[105] ), .Y(new_n1288));
  NOR2xp33_ASAP7_75t_L      g0903(.A(new_n1287), .B(new_n1288), .Y(new_n1289));
  NOR2xp33_ASAP7_75t_L      g0904(.A(new_n1286), .B(new_n1289), .Y(new_n1290));
  INVx1_ASAP7_75t_L         g0905(.A(new_n1271), .Y(new_n1291));
  A2O1A1Ixp33_ASAP7_75t_L   g0906(.A1(new_n1277), .A2(new_n1291), .B(new_n1280), .C(new_n1281), .Y(new_n1292));
  XOR2x2_ASAP7_75t_L        g0907(.A(new_n1290), .B(new_n1292), .Y(\f[105] ));
  NOR2xp33_ASAP7_75t_L      g0908(.A(\a[106] ), .B(\b[106] ), .Y(new_n1294));
  INVx1_ASAP7_75t_L         g0909(.A(\a[106] ), .Y(new_n1295));
  INVx1_ASAP7_75t_L         g0910(.A(\b[106] ), .Y(new_n1296));
  NOR2xp33_ASAP7_75t_L      g0911(.A(new_n1295), .B(new_n1296), .Y(new_n1297));
  NOR2xp33_ASAP7_75t_L      g0912(.A(new_n1294), .B(new_n1297), .Y(new_n1298));
  A2O1A1Ixp33_ASAP7_75t_L   g0913(.A1(new_n1275), .A2(new_n1272), .B(new_n1271), .C(new_n1283), .Y(new_n1299));
  INVx1_ASAP7_75t_L         g0914(.A(new_n1289), .Y(new_n1300));
  A2O1A1Ixp33_ASAP7_75t_L   g0915(.A1(new_n1299), .A2(new_n1281), .B(new_n1286), .C(new_n1300), .Y(new_n1301));
  NOR2xp33_ASAP7_75t_L      g0916(.A(new_n1298), .B(new_n1301), .Y(new_n1302));
  A2O1A1Ixp33_ASAP7_75t_L   g0917(.A1(new_n1292), .A2(new_n1290), .B(new_n1289), .C(new_n1298), .Y(new_n1303));
  INVx1_ASAP7_75t_L         g0918(.A(new_n1303), .Y(new_n1304));
  NOR2xp33_ASAP7_75t_L      g0919(.A(new_n1304), .B(new_n1302), .Y(\f[106] ));
  NOR2xp33_ASAP7_75t_L      g0920(.A(\a[107] ), .B(\b[107] ), .Y(new_n1306));
  NAND2xp33_ASAP7_75t_L     g0921(.A(\b[107] ), .B(\a[107] ), .Y(new_n1307));
  INVx1_ASAP7_75t_L         g0922(.A(new_n1307), .Y(new_n1308));
  NOR2xp33_ASAP7_75t_L      g0923(.A(new_n1306), .B(new_n1308), .Y(new_n1309));
  A2O1A1O1Ixp25_ASAP7_75t_L g0924(.A1(new_n1290), .A2(new_n1292), .B(new_n1289), .C(new_n1298), .D(new_n1297), .Y(new_n1310));
  XNOR2x2_ASAP7_75t_L       g0925(.A(new_n1309), .B(new_n1310), .Y(\f[107] ));
  NOR2xp33_ASAP7_75t_L      g0926(.A(\a[108] ), .B(\b[108] ), .Y(new_n1312));
  INVx1_ASAP7_75t_L         g0927(.A(\a[108] ), .Y(new_n1313));
  INVx1_ASAP7_75t_L         g0928(.A(\b[108] ), .Y(new_n1314));
  NOR2xp33_ASAP7_75t_L      g0929(.A(new_n1313), .B(new_n1314), .Y(new_n1315));
  NOR2xp33_ASAP7_75t_L      g0930(.A(new_n1312), .B(new_n1315), .Y(new_n1316));
  INVx1_ASAP7_75t_L         g0931(.A(new_n1297), .Y(new_n1317));
  A2O1A1Ixp33_ASAP7_75t_L   g0932(.A1(new_n1303), .A2(new_n1317), .B(new_n1306), .C(new_n1307), .Y(new_n1318));
  XOR2x2_ASAP7_75t_L        g0933(.A(new_n1316), .B(new_n1318), .Y(\f[108] ));
  NOR2xp33_ASAP7_75t_L      g0934(.A(\a[109] ), .B(\b[109] ), .Y(new_n1320));
  INVx1_ASAP7_75t_L         g0935(.A(\a[109] ), .Y(new_n1321));
  INVx1_ASAP7_75t_L         g0936(.A(\b[109] ), .Y(new_n1322));
  NOR2xp33_ASAP7_75t_L      g0937(.A(new_n1321), .B(new_n1322), .Y(new_n1323));
  NOR2xp33_ASAP7_75t_L      g0938(.A(new_n1320), .B(new_n1323), .Y(new_n1324));
  A2O1A1Ixp33_ASAP7_75t_L   g0939(.A1(new_n1301), .A2(new_n1298), .B(new_n1297), .C(new_n1309), .Y(new_n1325));
  INVx1_ASAP7_75t_L         g0940(.A(new_n1315), .Y(new_n1326));
  A2O1A1Ixp33_ASAP7_75t_L   g0941(.A1(new_n1325), .A2(new_n1307), .B(new_n1312), .C(new_n1326), .Y(new_n1327));
  NOR2xp33_ASAP7_75t_L      g0942(.A(new_n1324), .B(new_n1327), .Y(new_n1328));
  A2O1A1Ixp33_ASAP7_75t_L   g0943(.A1(new_n1318), .A2(new_n1316), .B(new_n1315), .C(new_n1324), .Y(new_n1329));
  INVx1_ASAP7_75t_L         g0944(.A(new_n1329), .Y(new_n1330));
  NOR2xp33_ASAP7_75t_L      g0945(.A(new_n1330), .B(new_n1328), .Y(\f[109] ));
  NOR2xp33_ASAP7_75t_L      g0946(.A(\a[110] ), .B(\b[110] ), .Y(new_n1332));
  NAND2xp33_ASAP7_75t_L     g0947(.A(\b[110] ), .B(\a[110] ), .Y(new_n1333));
  INVx1_ASAP7_75t_L         g0948(.A(new_n1333), .Y(new_n1334));
  NOR2xp33_ASAP7_75t_L      g0949(.A(new_n1332), .B(new_n1334), .Y(new_n1335));
  A2O1A1O1Ixp25_ASAP7_75t_L g0950(.A1(new_n1316), .A2(new_n1318), .B(new_n1315), .C(new_n1324), .D(new_n1323), .Y(new_n1336));
  XNOR2x2_ASAP7_75t_L       g0951(.A(new_n1335), .B(new_n1336), .Y(\f[110] ));
  NOR2xp33_ASAP7_75t_L      g0952(.A(\a[111] ), .B(\b[111] ), .Y(new_n1338));
  INVx1_ASAP7_75t_L         g0953(.A(\a[111] ), .Y(new_n1339));
  INVx1_ASAP7_75t_L         g0954(.A(\b[111] ), .Y(new_n1340));
  NOR2xp33_ASAP7_75t_L      g0955(.A(new_n1339), .B(new_n1340), .Y(new_n1341));
  NOR2xp33_ASAP7_75t_L      g0956(.A(new_n1338), .B(new_n1341), .Y(new_n1342));
  INVx1_ASAP7_75t_L         g0957(.A(new_n1323), .Y(new_n1343));
  A2O1A1Ixp33_ASAP7_75t_L   g0958(.A1(new_n1329), .A2(new_n1343), .B(new_n1332), .C(new_n1333), .Y(new_n1344));
  XOR2x2_ASAP7_75t_L        g0959(.A(new_n1342), .B(new_n1344), .Y(\f[111] ));
  NOR2xp33_ASAP7_75t_L      g0960(.A(\a[112] ), .B(\b[112] ), .Y(new_n1346));
  INVx1_ASAP7_75t_L         g0961(.A(\a[112] ), .Y(new_n1347));
  INVx1_ASAP7_75t_L         g0962(.A(\b[112] ), .Y(new_n1348));
  NOR2xp33_ASAP7_75t_L      g0963(.A(new_n1347), .B(new_n1348), .Y(new_n1349));
  NOR2xp33_ASAP7_75t_L      g0964(.A(new_n1346), .B(new_n1349), .Y(new_n1350));
  A2O1A1Ixp33_ASAP7_75t_L   g0965(.A1(new_n1327), .A2(new_n1324), .B(new_n1323), .C(new_n1335), .Y(new_n1351));
  INVx1_ASAP7_75t_L         g0966(.A(new_n1341), .Y(new_n1352));
  A2O1A1Ixp33_ASAP7_75t_L   g0967(.A1(new_n1351), .A2(new_n1333), .B(new_n1338), .C(new_n1352), .Y(new_n1353));
  NOR2xp33_ASAP7_75t_L      g0968(.A(new_n1350), .B(new_n1353), .Y(new_n1354));
  A2O1A1Ixp33_ASAP7_75t_L   g0969(.A1(new_n1344), .A2(new_n1342), .B(new_n1341), .C(new_n1350), .Y(new_n1355));
  INVx1_ASAP7_75t_L         g0970(.A(new_n1355), .Y(new_n1356));
  NOR2xp33_ASAP7_75t_L      g0971(.A(new_n1356), .B(new_n1354), .Y(\f[112] ));
  NOR2xp33_ASAP7_75t_L      g0972(.A(\a[113] ), .B(\b[113] ), .Y(new_n1358));
  NAND2xp33_ASAP7_75t_L     g0973(.A(\b[113] ), .B(\a[113] ), .Y(new_n1359));
  INVx1_ASAP7_75t_L         g0974(.A(new_n1359), .Y(new_n1360));
  NOR2xp33_ASAP7_75t_L      g0975(.A(new_n1358), .B(new_n1360), .Y(new_n1361));
  A2O1A1O1Ixp25_ASAP7_75t_L g0976(.A1(new_n1342), .A2(new_n1344), .B(new_n1341), .C(new_n1350), .D(new_n1349), .Y(new_n1362));
  XNOR2x2_ASAP7_75t_L       g0977(.A(new_n1361), .B(new_n1362), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g0978(.A(\a[114] ), .B(\b[114] ), .Y(new_n1364));
  INVx1_ASAP7_75t_L         g0979(.A(\a[114] ), .Y(new_n1365));
  INVx1_ASAP7_75t_L         g0980(.A(\b[114] ), .Y(new_n1366));
  NOR2xp33_ASAP7_75t_L      g0981(.A(new_n1365), .B(new_n1366), .Y(new_n1367));
  NOR2xp33_ASAP7_75t_L      g0982(.A(new_n1364), .B(new_n1367), .Y(new_n1368));
  INVx1_ASAP7_75t_L         g0983(.A(new_n1349), .Y(new_n1369));
  A2O1A1Ixp33_ASAP7_75t_L   g0984(.A1(new_n1355), .A2(new_n1369), .B(new_n1358), .C(new_n1359), .Y(new_n1370));
  XOR2x2_ASAP7_75t_L        g0985(.A(new_n1368), .B(new_n1370), .Y(\f[114] ));
  NOR2xp33_ASAP7_75t_L      g0986(.A(\a[115] ), .B(\b[115] ), .Y(new_n1372));
  INVx1_ASAP7_75t_L         g0987(.A(\a[115] ), .Y(new_n1373));
  INVx1_ASAP7_75t_L         g0988(.A(\b[115] ), .Y(new_n1374));
  NOR2xp33_ASAP7_75t_L      g0989(.A(new_n1373), .B(new_n1374), .Y(new_n1375));
  NOR2xp33_ASAP7_75t_L      g0990(.A(new_n1372), .B(new_n1375), .Y(new_n1376));
  A2O1A1Ixp33_ASAP7_75t_L   g0991(.A1(new_n1353), .A2(new_n1350), .B(new_n1349), .C(new_n1361), .Y(new_n1377));
  INVx1_ASAP7_75t_L         g0992(.A(new_n1367), .Y(new_n1378));
  A2O1A1Ixp33_ASAP7_75t_L   g0993(.A1(new_n1377), .A2(new_n1359), .B(new_n1364), .C(new_n1378), .Y(new_n1379));
  NOR2xp33_ASAP7_75t_L      g0994(.A(new_n1376), .B(new_n1379), .Y(new_n1380));
  A2O1A1Ixp33_ASAP7_75t_L   g0995(.A1(new_n1370), .A2(new_n1368), .B(new_n1367), .C(new_n1376), .Y(new_n1381));
  INVx1_ASAP7_75t_L         g0996(.A(new_n1381), .Y(new_n1382));
  NOR2xp33_ASAP7_75t_L      g0997(.A(new_n1382), .B(new_n1380), .Y(\f[115] ));
  NOR2xp33_ASAP7_75t_L      g0998(.A(\a[116] ), .B(\b[116] ), .Y(new_n1384));
  NAND2xp33_ASAP7_75t_L     g0999(.A(\b[116] ), .B(\a[116] ), .Y(new_n1385));
  INVx1_ASAP7_75t_L         g1000(.A(new_n1385), .Y(new_n1386));
  NOR2xp33_ASAP7_75t_L      g1001(.A(new_n1384), .B(new_n1386), .Y(new_n1387));
  A2O1A1O1Ixp25_ASAP7_75t_L g1002(.A1(new_n1368), .A2(new_n1370), .B(new_n1367), .C(new_n1376), .D(new_n1375), .Y(new_n1388));
  XNOR2x2_ASAP7_75t_L       g1003(.A(new_n1387), .B(new_n1388), .Y(\f[116] ));
  NOR2xp33_ASAP7_75t_L      g1004(.A(\a[117] ), .B(\b[117] ), .Y(new_n1390));
  INVx1_ASAP7_75t_L         g1005(.A(\a[117] ), .Y(new_n1391));
  INVx1_ASAP7_75t_L         g1006(.A(\b[117] ), .Y(new_n1392));
  NOR2xp33_ASAP7_75t_L      g1007(.A(new_n1391), .B(new_n1392), .Y(new_n1393));
  NOR2xp33_ASAP7_75t_L      g1008(.A(new_n1390), .B(new_n1393), .Y(new_n1394));
  INVx1_ASAP7_75t_L         g1009(.A(new_n1375), .Y(new_n1395));
  A2O1A1Ixp33_ASAP7_75t_L   g1010(.A1(new_n1381), .A2(new_n1395), .B(new_n1384), .C(new_n1385), .Y(new_n1396));
  XOR2x2_ASAP7_75t_L        g1011(.A(new_n1394), .B(new_n1396), .Y(\f[117] ));
  NOR2xp33_ASAP7_75t_L      g1012(.A(\a[118] ), .B(\b[118] ), .Y(new_n1398));
  INVx1_ASAP7_75t_L         g1013(.A(\a[118] ), .Y(new_n1399));
  INVx1_ASAP7_75t_L         g1014(.A(\b[118] ), .Y(new_n1400));
  NOR2xp33_ASAP7_75t_L      g1015(.A(new_n1399), .B(new_n1400), .Y(new_n1401));
  NOR2xp33_ASAP7_75t_L      g1016(.A(new_n1398), .B(new_n1401), .Y(new_n1402));
  A2O1A1Ixp33_ASAP7_75t_L   g1017(.A1(new_n1379), .A2(new_n1376), .B(new_n1375), .C(new_n1387), .Y(new_n1403));
  INVx1_ASAP7_75t_L         g1018(.A(new_n1393), .Y(new_n1404));
  A2O1A1Ixp33_ASAP7_75t_L   g1019(.A1(new_n1403), .A2(new_n1385), .B(new_n1390), .C(new_n1404), .Y(new_n1405));
  NOR2xp33_ASAP7_75t_L      g1020(.A(new_n1402), .B(new_n1405), .Y(new_n1406));
  A2O1A1Ixp33_ASAP7_75t_L   g1021(.A1(new_n1396), .A2(new_n1394), .B(new_n1393), .C(new_n1402), .Y(new_n1407));
  INVx1_ASAP7_75t_L         g1022(.A(new_n1407), .Y(new_n1408));
  NOR2xp33_ASAP7_75t_L      g1023(.A(new_n1408), .B(new_n1406), .Y(\f[118] ));
  NOR2xp33_ASAP7_75t_L      g1024(.A(\a[119] ), .B(\b[119] ), .Y(new_n1410));
  INVx1_ASAP7_75t_L         g1025(.A(new_n1410), .Y(new_n1411));
  NAND2xp33_ASAP7_75t_L     g1026(.A(\b[119] ), .B(\a[119] ), .Y(new_n1412));
  AND2x2_ASAP7_75t_L        g1027(.A(new_n1412), .B(new_n1411), .Y(new_n1413));
  NOR3xp33_ASAP7_75t_L      g1028(.A(new_n1408), .B(new_n1413), .C(new_n1401), .Y(new_n1414));
  A2O1A1Ixp33_ASAP7_75t_L   g1029(.A1(new_n1405), .A2(new_n1402), .B(new_n1401), .C(new_n1413), .Y(new_n1415));
  INVx1_ASAP7_75t_L         g1030(.A(new_n1415), .Y(new_n1416));
  NOR2xp33_ASAP7_75t_L      g1031(.A(new_n1414), .B(new_n1416), .Y(\f[119] ));
  NOR2xp33_ASAP7_75t_L      g1032(.A(\a[120] ), .B(\b[120] ), .Y(new_n1418));
  INVx1_ASAP7_75t_L         g1033(.A(\a[120] ), .Y(new_n1419));
  INVx1_ASAP7_75t_L         g1034(.A(\b[120] ), .Y(new_n1420));
  NOR2xp33_ASAP7_75t_L      g1035(.A(new_n1419), .B(new_n1420), .Y(new_n1421));
  NOR2xp33_ASAP7_75t_L      g1036(.A(new_n1418), .B(new_n1421), .Y(new_n1422));
  INVx1_ASAP7_75t_L         g1037(.A(new_n1401), .Y(new_n1423));
  A2O1A1Ixp33_ASAP7_75t_L   g1038(.A1(new_n1407), .A2(new_n1423), .B(new_n1410), .C(new_n1412), .Y(new_n1424));
  XOR2x2_ASAP7_75t_L        g1039(.A(new_n1422), .B(new_n1424), .Y(\f[120] ));
  NOR2xp33_ASAP7_75t_L      g1040(.A(\a[121] ), .B(\b[121] ), .Y(new_n1426));
  NAND2xp33_ASAP7_75t_L     g1041(.A(\b[121] ), .B(\a[121] ), .Y(new_n1427));
  INVx1_ASAP7_75t_L         g1042(.A(new_n1427), .Y(new_n1428));
  NOR2xp33_ASAP7_75t_L      g1043(.A(new_n1426), .B(new_n1428), .Y(new_n1429));
  INVx1_ASAP7_75t_L         g1044(.A(new_n1421), .Y(new_n1430));
  A2O1A1Ixp33_ASAP7_75t_L   g1045(.A1(new_n1415), .A2(new_n1412), .B(new_n1418), .C(new_n1430), .Y(new_n1431));
  NOR2xp33_ASAP7_75t_L      g1046(.A(new_n1429), .B(new_n1431), .Y(new_n1432));
  A2O1A1Ixp33_ASAP7_75t_L   g1047(.A1(new_n1424), .A2(new_n1422), .B(new_n1421), .C(new_n1429), .Y(new_n1433));
  INVx1_ASAP7_75t_L         g1048(.A(new_n1433), .Y(new_n1434));
  NOR2xp33_ASAP7_75t_L      g1049(.A(new_n1434), .B(new_n1432), .Y(\f[121] ));
  NOR2xp33_ASAP7_75t_L      g1050(.A(\a[122] ), .B(\b[122] ), .Y(new_n1436));
  NAND2xp33_ASAP7_75t_L     g1051(.A(\b[122] ), .B(\a[122] ), .Y(new_n1437));
  INVx1_ASAP7_75t_L         g1052(.A(new_n1437), .Y(new_n1438));
  NOR2xp33_ASAP7_75t_L      g1053(.A(new_n1436), .B(new_n1438), .Y(new_n1439));
  A2O1A1O1Ixp25_ASAP7_75t_L g1054(.A1(new_n1422), .A2(new_n1424), .B(new_n1421), .C(new_n1429), .D(new_n1428), .Y(new_n1440));
  XNOR2x2_ASAP7_75t_L       g1055(.A(new_n1439), .B(new_n1440), .Y(\f[122] ));
  NOR2xp33_ASAP7_75t_L      g1056(.A(\a[123] ), .B(\b[123] ), .Y(new_n1442));
  NAND2xp33_ASAP7_75t_L     g1057(.A(\b[123] ), .B(\a[123] ), .Y(new_n1443));
  INVx1_ASAP7_75t_L         g1058(.A(new_n1443), .Y(new_n1444));
  NOR2xp33_ASAP7_75t_L      g1059(.A(new_n1442), .B(new_n1444), .Y(new_n1445));
  A2O1A1Ixp33_ASAP7_75t_L   g1060(.A1(new_n1433), .A2(new_n1427), .B(new_n1436), .C(new_n1437), .Y(new_n1446));
  XOR2x2_ASAP7_75t_L        g1061(.A(new_n1445), .B(new_n1446), .Y(\f[123] ));
  NOR2xp33_ASAP7_75t_L      g1062(.A(\a[124] ), .B(\b[124] ), .Y(new_n1448));
  INVx1_ASAP7_75t_L         g1063(.A(\a[124] ), .Y(new_n1449));
  INVx1_ASAP7_75t_L         g1064(.A(\b[124] ), .Y(new_n1450));
  NOR2xp33_ASAP7_75t_L      g1065(.A(new_n1449), .B(new_n1450), .Y(new_n1451));
  NOR2xp33_ASAP7_75t_L      g1066(.A(new_n1448), .B(new_n1451), .Y(new_n1452));
  INVx1_ASAP7_75t_L         g1067(.A(new_n1440), .Y(new_n1453));
  A2O1A1O1Ixp25_ASAP7_75t_L g1068(.A1(new_n1439), .A2(new_n1453), .B(new_n1438), .C(new_n1445), .D(new_n1444), .Y(new_n1454));
  XNOR2x2_ASAP7_75t_L       g1069(.A(new_n1452), .B(new_n1454), .Y(\f[124] ));
  NOR2xp33_ASAP7_75t_L      g1070(.A(\a[125] ), .B(\b[125] ), .Y(new_n1456));
  INVx1_ASAP7_75t_L         g1071(.A(new_n1456), .Y(new_n1457));
  NAND2xp33_ASAP7_75t_L     g1072(.A(\b[125] ), .B(\a[125] ), .Y(new_n1458));
  AND2x2_ASAP7_75t_L        g1073(.A(new_n1458), .B(new_n1457), .Y(new_n1459));
  A2O1A1Ixp33_ASAP7_75t_L   g1074(.A1(new_n1453), .A2(new_n1439), .B(new_n1438), .C(new_n1445), .Y(new_n1460));
  INVx1_ASAP7_75t_L         g1075(.A(new_n1451), .Y(new_n1461));
  A2O1A1Ixp33_ASAP7_75t_L   g1076(.A1(new_n1460), .A2(new_n1443), .B(new_n1448), .C(new_n1461), .Y(new_n1462));
  NOR2xp33_ASAP7_75t_L      g1077(.A(new_n1459), .B(new_n1462), .Y(new_n1463));
  A2O1A1Ixp33_ASAP7_75t_L   g1078(.A1(new_n1446), .A2(new_n1445), .B(new_n1444), .C(new_n1452), .Y(new_n1464));
  INVx1_ASAP7_75t_L         g1079(.A(new_n1459), .Y(new_n1465));
  O2A1O1Ixp33_ASAP7_75t_L   g1080(.A1(new_n1449), .A2(new_n1450), .B(new_n1464), .C(new_n1465), .Y(new_n1466));
  NOR2xp33_ASAP7_75t_L      g1081(.A(new_n1466), .B(new_n1463), .Y(\f[125] ));
  NOR2xp33_ASAP7_75t_L      g1082(.A(\a[126] ), .B(\b[126] ), .Y(new_n1468));
  NAND2xp33_ASAP7_75t_L     g1083(.A(\b[126] ), .B(\a[126] ), .Y(new_n1469));
  INVx1_ASAP7_75t_L         g1084(.A(new_n1469), .Y(new_n1470));
  NOR2xp33_ASAP7_75t_L      g1085(.A(new_n1468), .B(new_n1470), .Y(new_n1471));
  A2O1A1Ixp33_ASAP7_75t_L   g1086(.A1(new_n1464), .A2(new_n1461), .B(new_n1456), .C(new_n1458), .Y(new_n1472));
  XOR2x2_ASAP7_75t_L        g1087(.A(new_n1471), .B(new_n1472), .Y(\f[126] ));
  NOR2xp33_ASAP7_75t_L      g1088(.A(\a[127] ), .B(\b[127] ), .Y(new_n1474));
  NAND2xp33_ASAP7_75t_L     g1089(.A(\b[127] ), .B(\a[127] ), .Y(new_n1475));
  INVx1_ASAP7_75t_L         g1090(.A(new_n1475), .Y(new_n1476));
  NOR2xp33_ASAP7_75t_L      g1091(.A(new_n1474), .B(new_n1476), .Y(new_n1477));
  A2O1A1O1Ixp25_ASAP7_75t_L g1092(.A1(\b[125] ), .A2(\a[125] ), .B(new_n1466), .C(new_n1471), .D(new_n1470), .Y(new_n1478));
  XNOR2x2_ASAP7_75t_L       g1093(.A(new_n1477), .B(new_n1478), .Y(\f[127] ));
  A2O1A1Ixp33_ASAP7_75t_L   g1094(.A1(\b[125] ), .A2(\a[125] ), .B(new_n1466), .C(new_n1471), .Y(new_n1480));
  A2O1A1Ixp33_ASAP7_75t_L   g1095(.A1(new_n1480), .A2(new_n1469), .B(new_n1474), .C(new_n1475), .Y(cOut));
endmodule


